`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CncNK4FCRbhq2wSizbRTVHnAqJdmJyFM0zrTZFM0xviq/ReMLSj8w/pC7qbGHLMIvnDYxIw45VEB
xdL+zJ5MGw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VLYwsd3GMIG1D2lwWLTQPYLgGoiE1QUQSpt3aY4lzm9d4Lqv45EZwCa670pueNnM+Z7PwB3aitXo
MiH4t4uRN3hDn1QhJ2ClBmI2tsNgPALuYc0J5qU9JN9IKy4uaQ3zjakv5TqVIC2xNUxXGrl2pfeB
dSA5/YnpeYKjqC4w3M8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
EZn5uWxHY0yseLdi5uzrVV8wyQUJ/G2NN5dEQiVOWEBDJDGqkeu1QG7PdyFoWY2RzkUL8+6w+9eF
/B1G1Y+RSfeQzkYBeU05tvDWMuRmYH1Ukl+elkmapPCfkKn7H4lO+I5C8xhpYnfH6tQi+kgcqTBs
sDwu06UnFZ0Xq7DSyKWpLJvtvV8nDJyD1p8DbCzywf8K0uDGcEJ9O1L0vkw/pyd65tElbEY2VOtd
XaXCqk0xcHEZdxLyJoNgRTlskmenwbhh+nNA88ngjm+W+YP+RpJ+//V96HCjJdLtubVQ9XTJqCNx
Ki/q30UOMuiU3L+jjTmO16ZY5jjRi35gkYlk6A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eNZ6hQq/cQZkIPHHXOfpixt9YG3Yx/ggZQD/py6rjiuOMQPoqCLax/NXs1d47RPQHg9KnYsgYsvC
jvNIVkgutfS2qiFh4lVqW09Chym3fVnvg/4bx4WkTkU4r2SP3B+4KT+/yaO5QQ423rNP8gdK4FJj
wR4E8ckzvzPRNIMM8oc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mtNNcvnOs8KnjkG0lm7b5bmphqS20d2JbyEKm+vqPAFGe9wC4v45yZtoTwl6QtdJiWZXPUIR9rWn
EvyLAhZHQV9rNJ5q+JaoTRlyUiMbjWeGA97jBjmAIKa/tBlww43vfIaM/GtlOJ7uIbqTCuvp/WP9
HZo3KniAVlqFzuLNANuvkOWahTSI75Zp1roegn6wfolUm0OiI/FcauvC0Fc8PmQmFqAlOIw45IyR
Vdomk/OQaUKPRJW/72/nn8SaH/epsM1CKt6O3k1MB10FbQS/OGhwDEzy3lzWQhv2xu/9WXN7MTR4
/x/mgSkZN+mjpeHJq9xsmEUTh086k2HuODuOHw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38784)
`protect data_block
4w/5u/NHk659yEsUlY65gCE68R9PPldq3x68LXy63h+qYTfY3WAs8IKwHl7AEqmUIkG+844zDHqj
NXGs9cXmDIrjO99j0p4LgoY29bHCnQKGbC3RH85hLX5VWKhZ1r3zmkaakhKrRYLFWFpuXvDgS1F3
sFM74giLeZ25P8PqfNzv7m6vbNkiBaCT3goT7L+4UXEU8nrfjBzNUTlf6f4CgjLMOyUK/1H/74Zl
4iO6tsewjXiH1AtR9z0bSYLTob4w3HEhuHgsI0z4MZz8+/Jn/aTWLIgYm2ni/ymMWwQ5toyZS9eK
qUGpJzorfvv31Ij4cRIEp0oTK90tYpZ0UOwejqBMgYrAIox0HLc55NdS3Zvh5nrZDNJ8qEmZYvIX
b3ytxZCcsQ2UMerb7XkZvgBhzROXFoyvD6o9Gho2bqjettFH6B14mV/CrXiV/FTXWA9fiJ0oJ9IQ
6v7fkr8iemTENZyVJ6z0cayWmlKnW56gMHDfafuTIUIApYa+rM/CbCPv4XJ1jsV/7wlTnJSARDYb
4wNmwZVzuwyvFit97frLI/+I4/VtNDggroTVeypxxUrSMp/Db0+oDyM4YBbFEyqcITqlsTuhbXXg
s0flggBsHG7XVx2+pAOE2hTlJ4Kf4Luut6eRhGM7VEd1dStlGMVD0q0nhutMSrXwuqvedRE/Tf2i
SKwQ012ckkI1YsXed8bMxSmjfVpi6jLYcXYqco6DK0wj9nMD2B5HL6s8k7BfQIOLlXQI37Ug5/Z7
GoLqp1GXxpsJJezA8GvWtgdTjvuUXZYe7arelC5jjjxLTcpDUI8m+62qfajvMiE4kANP5auoiqmx
e83YD/NL4AOhkHdbbZiNCVjDJ9yRfg7Kl0RjGZEnuv+RZNyjz4v3HHM4duPhQc2JthRImenL7Lz3
+FiqwlRt1EFMpn6sRXwBVkh7zSBKf/akm7oS1kiyPXq8g07K9qKWB2Dy2UuS8QCu6RRtOWHNct9h
cD/OjrrT+v7FYGL7WWUEEW/yaOdEYaU4QXFrncWV4lqYF8KvXO7nnlinI/GKGzBtcnZRe2LqbmeD
egYUxdbWn14UacC8H72d9wZENrT6l5Q8a7bTSYpuSzwq4LlNMN4hdnSMs6FlTy3RXCL5dmfA/o6s
z5fhBW55z4zFKHuScJWAtds7R0+DEs3Y9rNr8oaF0HPON/J36cp72RQKffiNMNb8limVmcLPoKuM
vs0Rz+imaUif6y9JqMmhcZ74J/pHpoT//Y1G6YkUntQawELs+7VYcvDJJHgLvT1SI2BBdR4d/N3N
ftiv1zmAyKL7q6WHNa2z/2RchSLIhaY1lXTXenSeLHdu+tDTtLm0QmVXg1i9KwSVVPCaD6CU93jE
lipgYvtpMkqil1fxUveUT7QqnKYHcraAiI4OAXOtpyC2EIfI1RbXiwcavm/AcSvdqkm3r/F9GqGu
8xyxlis1UgIqkyWy2ly/spb5YwEtbn2Ls7+qn4ioeFC7k2IbeVVoltqlwM+k9R0Q9dnBiOmB/5LX
WQGeqPvAIobE5hRxogI6nOLgwSyl7teg17tF8vmPSvvkqmaokz9Lb24op7ggPMOWdvKOtz7FPO/g
OZTP61C1v1rHEsMZSi2zWa+8feluTbs/OmsZ6fcEgUhzzih9WRWsX6oOJ0mKEHKvGri13J0yYY1T
9ycFZIkmuDbmTpnWjT9vm1BoyBfLTKDGTD07JFJBlbQPXK8DIN8oH/3q1W8SrbVtAGuA0pYV9z5N
GI50xkNmbVl+QfoiuVSTz5VbNNWQpWjO1Nu3a2CXT38EL6iHO5mYuT6DcJVmtHuQ8v3qLNUua2cr
JvQtmHzzLc0lQn53SEELSWgvLSUn+pNAlxhJPybrkLPWWvlJRKXLfYRDBCUhv1unL2T8/Tlqkxsr
lgxpesY6jgEORsgFl+whAuIbKIdDRef21M2Aai7SLoR1BxfjjiIJvLIsEl26Ww7V2I7mvCHw5RUP
BZTJ4qBxfwgfRVEUijt54lmufPQ+Za45GGrYIRUt7xM3+x6IEAKQc9xE2iOISUsAZF714GQt7Fd8
+i4corHlLwsAUmfV8Pw+pP2s9KJcAKE+F/AXn21trSLICO3J5SrY6knbLX1LWZOmjlTjcnA+EF/J
etRYbqVSpvD9IIECuXVNW8GdU84daFX/MNz4Gey1NL6IHTC+hRrc6Lj1fEWCxShOC6J7ZFVloW4R
fAc2x5pBZuVs9m7UsDBt6is8flYzV627+Uja8l2qWIbQHFMBjp3+nA/Utkwy2Ih3EzdqDnmT9Vbc
BkjIdO5CrK878SUjS1DkCyDMbmZ/ZuFmN7XwAdgqL+gSEVGuOLfwin0inzy9lZdFota0zfY+E3EA
PDuE/T3bW43CvlYxFU0FAChQGhbIlGksB0w54TyiHg9ECFHb8Zxzny0pQ0UHvDd5JKBoRpW7unZk
ZL6m3RLLeuzQi7MM2AOVJE5d1De/ksPGPRyoj7QH15i9lspjKg1h8JmrwbGTtMuLIZKWbHiyEk0+
cuUHgCyAgORufB0dgbAjZvtjEx5jaDJzhAbtBgaya0o16PORQGA4FYCRr6Rdc7V80ci5tcRWUco6
6sxGm5HNsDOkI77ouv+vZzIjC3RjAL4MynLxF6ca+RPsitW4W7fqX7d7eTzg1+17ItClGCTC1uOd
1gIL7BDCLZu9bpNUXdV+29LhK0bktM1r+iUuzBbIlkqLhJ8uFKuJn6Zzk95lt8UeTOXGd+qA8rUc
xDT8l9kX556air5tkxUrixyv/JAsxSSdvBZQ30dm9mmp0F0McL2GUP221wt2J3J58HnHl/Gqn9k+
Sp5aiW/vAycDbZ2NXAiiG2dfinpo4AMT6Nk4KZn4ELH9XSc3W33N4Zo4VSVKwcu3DlFgStrq1FV2
6bO3YiAGBIhdRAwFssa4Y9jOamQqE+BvmE06tOUkXA3rebMa+vF84rEMhzOLHHwnEBBv0ALMKghE
cBd2K8OtTLwYtBLa1fsPllxM2dtqNa6xcz3GbFsQMGU/he0Kj7Vpfs6U54Z7dMoPBq/9Ydkpb/lF
ZQLDrwmsoc9hrQ8hWjhD4GBFSOu+KWsGZgUZjo4hDdT2P7mpgWxAjaiswDhhyyMmHg+x6/r9z3Be
poKrJ6QC8Wp6XEvEubLkaYIfiXfyRqRnNnoK57TlXwm+cgkydePnfu7mIm0budxH2VV8K1fQqLfn
ScgEqx6N68FjZID2WdIPvQ4FuKCKnl0kLZNYAejWdIuOJ/ZbwC9lgi2MpbwsbOMVvtJ4ObVh0ooF
iT0bfAJI/3lXauY2Ewrj0Q9q9RdiF6y8U3AVWxhE/rdIRe8nP7/Vx0H3n3u6cyku14UQlHl2nD7N
59nDjlE/ooaetSMvhTjCDqNaHe8eJbFqhg/3M9Rx34kWXUg37shuZ0QeSecwI7hU6bDxhgbctb06
/6Wgt1GnpocKBrQlULCMrJYFHmPoS2lf5EyWRj6osS+MZq1THeWBfCPgQ64WFfTBJ9oyWhG/wfQO
EPEVTRNlCk9m7LJUj88yzlysycWWDasELaxWXqrcVTQHqFBEsakLdaG2wVNSFqIU1cW+nBEg6wvb
l62B7ky6IFJSTHJfQXCTxvgLdjHfMB6e6aEPfSm3N162z5Ozof4tO0pNVAbqWVCcSfiexVauuAeR
ge4t8vQyGQjppkVWaBphglQsHMMUtd+wbC2y8J4eypGVCvRGBULK/oiMBH6T0VL7hOKwt9XkRKxA
pxXksytABGRXj6obwK6DHk2tmTtlnUZH9lGCn6jTkQpr6pwE9eNcoh27wj3vjN9zYh7ACu2yjUR0
1iyfdqCJrEtInHG/u89PQlkKS2rDMLydCc6vE2azGtn5kU7de/NHSwX43xMsKu/i6VP3rI0HmDm8
C26VnlGtlfrGrN7RebZdFCrU6NyYZ52VkUaTb1ZJ/WBC/bRToS8r7nNT8uIzAgN0kIR8Z0StK/u1
lEGX6/dS607pOvxeE6MMxmSDGKgMg0kdCQUI+4DaEI2QbFTOEwEcehbO8Jbi46uRkIzFNen4RV0C
JDwzUaoDHgRnbWISTQzaCSHqWxFuLdAA9LEi3kXiaocY50TnTjsl8D3F5Y4CwSOiyoiJkBzfBqiu
h8fhzdi+GGbutjoF37myFMC5e8hWMn7D5vdF//LX5BmhukL/olBecGBrVQrXU3vgA6dhvY5xJe3C
DZKBfxf2nHFVtm1x/jCmIhhnzSTBU7Z73kN4cuUWdaUnLEGlA9enmoLyViCXbaFGNvHZ4HcJ795R
DSoerxi2cksjeABARUz9JE1kE7L/V9az2JKXk5KoNVmT4p5VIePHz2E5uTq0qBYX8U3mdNtj9b6O
chmorTuD3wlovA1/9mraAGcgVbHbemnURrbZnZ1EyqgmD2kM1Ob7psmf1Lk4Uj6EdTigUks2Vjty
fK5jJVNY4ABp2mZQa6WMUoG/ItygBD7PcNdHqOyFNYSwwIMgbmdUaXsx66QPgD7LOvNGggQqGPDA
rK7dj6xBKVfg+Z6n5GLSL+FqJH7XJTyL705YURdt8fkzZb8xtj9suwVFdWHd32xsCYrqSb0bdUA2
MBWX0Rfv7KFpSEcq/2qWL/Be4pzSxOGV2FfltQL1+1y11h4uGbcgtWLohnfqNuvsmnrYnGxx9h0h
WwAXWnnIoDVge9sCfc4x7LYlZ+muh+2d7Za71NGIohrCjtHpiHWVunl1AUf1th7+gGUGBbFCYGXS
j8tUrJ5Q9eRaa/NcwolnL4wuUMY7iLe0Xd2gGIf76GiriIh+n/ER7iZapcREygMKRvTi6rlKjchA
ANISmnWMVuK8TAgP9kpyZqki7SF0FyGO32vGexdjOTqP3jBBgl2TnWu+MeBNxdar+dTI2R51FxSs
8sKMZXiJtigQSUN9M9V4WtE83mJUSMzzicE2IOFOR+FGCcGHC6of0bchsefNdbtldItP2nSq2WoO
O4B6do1uAAgybBM0WbdRNb81rQmBZCFP+MIWF+fo2+hoW3nWe/7e+UgnRCFozOGTKqxs/sg0NHCF
v3OvhHMW5vkbXB4158esTgnosk/irVBSROaUHE79a8UiGD4tYcW7Rf7iTPU8UEjwhn3gC1ucZxTV
0w8mH3Twh9JZTyMhaCq/eq++7GDTJrCN8Gp6qzU2KKd6XLcYq/pfBBIyZzeC0YXYK+Ly0h5KjbBJ
9APyW179qUmGFsTvtvx8p8HLVoNBHVFk5ImUVHclQIjgpcR5tfS8Q5Uh7e/d4JKPGrRBxzTVtVxA
KiRL0CZgjZvrhahxjz8SnxpjqU8QL+t7lyE59T8j+DJR/MONuWki7qNxCAlXFq2g00Qcqg3oyb5h
usK1wSckIOs/Q6RbQMIxBrNNy2IZ5croI1LrOkPp+9ffQ1P718jBBCNjB7m0+CiYkWKmr7LXgM5I
7oA9ET6gJW11MwJvact4ZavJePR541YIDdH9MLCmL7BPucyLKPgHkO56OkSWKsbMPtc6gcNY48hG
bRwUjSfIk7ppkjeCfu2YubRgA0jz47eC5zO1PpP2A+XRc3DLTwYl/O4+lW6tU3y8OkGz2JbDVr/U
VGzABO/MUPq4F/FgRoH6qcE2fYc7Ce9JLIWAOXNqiFjCN4unb9jwmi45HcNp7FYNd3pIfh9WBk/e
13Svqors4MExHnnqVlYRz2r0hnX0LR66TNvVD6Ml80avZJhLSLeMUzyp5yDp5fVOiNYdtK9d5KAx
ETK0iKClktoTnMI0PGlxhqbbDwhQCmklr32IhpE7s6NJJGop4YvNcSiM/nVuBa46g+UvmBAKcKkI
EWDs8RsC/3RjpiG9wRQTUc4iXXUaeI+AeZsK83DkIfvB0UL6coEeOkVudpzVteTcDQtkb4AVDkAc
uCMgNgOaNnYqgbV9/3M5nFJ1LRY+gwRcbb0M+2KXhoWxN7utBvSrGKMEM1KoATZZeJ4yv9wzNKJg
DkXGm8/xGpqXXMZCag+wv46l5SDxSA+Z0G2kcsoVXld/cnkadSMKO9/u2cKFisY/Y7uystU/fuTU
6hlDKZ6N7FysGAMTfP6mRb2ofrQ/sQIM90QPBSvDyTBrQq7popiJsBuciBZfXVdqZ/kpFA36PT75
YLRaIq0n7wqNtNWpM2U1+aGc2URBHD/YOkkaZot5w0FgpzyZavzAeEgamJ9j/2yN67Z2SRMXlVk7
rQixUBMbeUaBqyZh78IUTD3E1hwnf3WTgxo3em/WATn4hOqReTzLHmx9zSXy5V0p+AsmX5nvmIxj
bgYzN764MrIaMVOuvzwzgWM4UfQ6ulOgdpRqBsRqy5ZIwbThGsSB3zgENiYUaPWGu4GTx4Zl1fbt
VD+49pGCuaE6Rzftt7dq6Fehhg1vgaCsa/OsXmc7APXJrkVOXlFmEJNHQGHbCD6xpCBO7YHCtwzn
DFk0v23kyjmlmXObGgZ+NARjFd66iINIAkxAO2TfAoZavj/MC7J6+TAmxzHfG9NAmwPLPEUy67zS
DkpUtEAt5sveYYboIGXe+q2o/4qFCZowT5PPZAyiT7bfdaml/EfS3W5MaaACHZ29BLjZP4RRHkqp
HA+0KXU/9Ai01wTi3D29NyqxHFObhGo2gRFdZvMwwsRzj/QSfdcTJF2DhiQ6iyVjK4Vp35Ts3fR3
d0V1aSKiRgprPCqcJrDIbL+ft0Hv6SE+skTeMgcsukbYdClkJrdJ9HqiYgNEllrjDXwNLG89mNKO
l18f37JB/r52jvI+uy+xOKGRdOIdyLtxFS3bHy02XLwBShpI9Dl+/JPVpV2DdRqww/YTIzgJh7EF
K+SdqbHXMjW8bSqbRnUICF4bYZeCNBQoysnxqOz9AefsS48XxGhBB+qysFMs1mjwgrM2fFgjKEMG
dAyIL647Q/OB1YkjdT/4NLqqSI0dBvaD6jn2+qfhVVZtZWcLwYRKqgl8aq86v4ISesXTo66tENU2
mowDSyyVbUqj4EOZoWTU3czAlUqzvoy2YTPj81AQjYJe2eM3jdqC49aE0PJ8yfCEZHVHZVgturJ2
LYray9llgqhhjT7Xap0jkh2xkYOMj/iKvf33dLvRtFo2xufLeL4zxolEwV6t4X1ope7z62VwrvHj
ZM0H9clY++Ti74aZ5cWdafDVh6Y0Yqj9/GmsYwk6zud5N78u/4S4f//2eKEpgodaY8aXXkOjXo2Y
NtnZ2EVtRyOm/EOfD/2/7t7AvIeiUt7mQAS2K2tT1qPJr1r7OskVyjYAkSFebZ6q42STlPOU3Ifr
EQ3vpJveMHVKdnlThegiGbnKHZjdOBGUbDFsmczNC9wFZpuVV+4hTEn3jAsb/fA7UaFpgMIfb3hg
3LmrfreKMosIIx92Tf+8LrGY9Pxg3yXCRv/eMHL/ZKpyoPOIu8yqyqfyMdhmeiYDWc4PkNbrv2zT
MEkHJnFh9Tab90xZ7cS/GSqQRg0BoA8IeLvHMzCxJEJ110+aeGI4/l2SHh1+2gH2Z3jho2G6Wdbl
LHv59WwK323FbfAYwQFHkdvmdW4nDT1B5qIXFkamCczSfxv1JTNGpUXobtHXs1RF5ZA07vftjk9P
zH2Pa1MJli0pmnKM9owHbqqP87wj/4tl64/VhV9T3J7cOkR3/02BHmpg2EdrAYHfcBytv0rwli29
hjR0yr309td5cIvIcyA0dIoe1WggmBSpvfF8IHvRbMgJX0SVoJVNdIWsb37v7299D6CYU9RP6n2L
0gZH6KS1RzJGE4n9uhH/8mb3k67QPEaFLkSF5WdCTz6pzavQ/ocyvDLR6wKIqF2nvwLlM9MfVKPS
XMWrlun6TmspA7ORJPKB96swWj/xXjEzxUyzZkG5qV4e0hIugajFeSJvfilnmV0HRZDtsfTF7n6Q
ruDsCoa8eWENL5837lw8YVnX83Y9+MJVEwkF1bP+KWdG0jdbYhA+L6+UfJp0zvS8nGOfgxwobMOM
y2tLH9prWq2LGOHV6LP6X9WbOeNHTBFWQqx/Qnj8+uBqSB32qxLQnT8tWDEaXJwUJ9BNc2GOVj1e
b5Imrs+3gg7AlH1EJUEN0B9SB05kGUiQhvRlLKKSMNy6sVjAKUkxAuDAXmEle6tf5p0WVnhvOabe
u/J88v1Gs5CYq4BGAbr4TKuvPGukC2MZR5UMjiQco4JLG3N/P9wqO6x8zk8V6cMuKMSiG8//xlCl
y9B9XwoSyIam87m4SP9wRKScTr+eK5NWwYwIsu1FEmPebbUOx+0QIZooVza8F7nfhVWASJGZud7/
FWHu2zE78Z6NeOnmyn8pJtLiVFvyf0t5M7cHGsHPwtIdMxIVkDYXyf+iYLV5BiuicGDyCnQDCxEZ
PfDPFvqm++uXS0BDHkWSMlW/d+UOl6LdHc7bnfJ2st8zntK+cVWe/NCJ56mcUdx7/UfSONmS2hTo
8VCkhpeo0TD6X/EYVKbBZIikD8onZmT49vAqE62Pr55T4UWlfDQKXtRsMosTIuuBGPCzRrCWiCQP
7VWfR+eDuI21BiGbYaz1zU40bMc517dZLcmwvysozRfeieq5u3+/62+EE8OmsVMT/4aOECX2KQVU
1hGc0q1VBf6Uc9/GsZK5xwBuBki2p48UOEZRJIm1iojBsu8oK6yBKq/AJ82+CPpSFbCLq6m8qQx2
Dm69ugrJLSZ/L/5uVRc164Z/MlJdnOZGeqrITwgtO6l7Mo7SC2lyNsxaL0AaxNix6PsWRdt5/Z2P
mpV6uSCSM9V+cIJQSIzGqZrKTGOEFSmtlNzW7280v2EABLCAsCCKrsR4GjTMprRDMmvIpNjT8gYJ
bXGejjqw/0Q/DLqjbWfNkzv5P+HZ+OoSu7G9+5ajZoA+eMOpDpXhNaIqCRGHzqDLD1rALTjQ4u20
R2tuqZZMYM3EDL9/I8OfT3GeD6DQx4PGeORqpiqoGOLCypdun6h9/xt3U/n0u1x1dReXVH7arErv
+9rSqpp7J4CwJNT4bsYzzTd+VKSCB0xldHeymTVXiSIuLTktdSRNBejRBFJnZfPlFso8KHTv4uHc
YYuOy5ICaKY2IjCzKI0NlAJZ/ZV0iFcBcpqZHPDwCRsHiAhjF+VGgs8j0V0jBDCDGQAVjlTRIOkv
U57rnCKyvdILNw8+mbH7LIQH8K/9KfIklz1osADVibpmDpSMDyurFriyjuw/Xuyxzb6ktoRUl2Kj
hCB09xrZsRP8pYGQZTYDWLnvcVEuy4eoksh0C1H3Jk+b7RwfPLF04loPivzQxUlrltOo0M7U7nhq
Tqifu2siFFFRJJkif10Nfb2o1eK/hOWd35HsOWdbCdR5IPH2ttjRIJDc3O7HkND0FZS5uAUAo4Ld
K/7jdTBhoEcukdnJ77Nd8AAQpOXvcjosDEVUFKNCvMesxQcnMvG7oCJMsU8wAaFHjswhumqpkF4e
YCKJZfNK7XCB1bZssdxBvLgYNj2Hrbikw13wdBl/pdpmdmKmHC9FR+rWwLO93+VxoVGorHrQr1En
mIbhsS3Z4vxkbxMAR5qKYOeA7p0amIMIFH3CXfSpaPrXhrUNXqyywo3piqfjsZ2/oIwDLB/lig4o
W7pqz0HQcTH53GsYrRyRuIP6cK2G9p2ybECBTWr0URIfOzdTIhR2drKEmvL6pHAqfl6mdCEnnj33
0QFoP6IlQ/cwmCI6FdeUUQJ01pKK53VBQeo7uvvdECtbBCkQuECIR0/zgqq5ZIM19a0LtW4A9mBp
PZ6drEvIa/OQBuZTx5OcUlA8PhKNTW5Ah4sC3QKDmYYsDNmSRVZkgw1nPko8xjTx7TQeHFd1gZPe
JSQ5chNcMUbNFKCdhyNPGP5QTskTn2JwBIq0+ABrbW//0kzszBifgNaqBeO4HysHtE9bCIqMVunn
DR+TJXEd7u0Ow6NGWQfvWsOZ0r6EwQCmzNE2+EnYnpD97byosI1RP2ELqmHYsd7qumq7yWKyaxVu
rslHv0tsip9kc9jnX68bnVIaws65OkfBWBpWv9DbaGHXAiKjAc1NS79q/ZsCcX6pSFi5FTVeVkI0
8hsRJ3srJcXlK+nFcHSFCNevvM0Tc3wepn0QOPBH62524DlEDHo/sZXZ5Bd8E4kvgWpA//FAbJO/
P84JEi9uzuvloFQ7mgOkcOUqpaIimmYXPioFj38E4jTZOTYgzJY26kC94sz9JomkrAmcqdM09K9L
uDoAeSCWvcnzwk3BDZoc+yum2vhvJH8b71WPwS//0hGdx/NUU0Aq52sh+ZzVisq6K6ufbnHUeG4Y
yZN0hFqbmnPrJRVRYPWIGa9uhZmBARZQb707J5LzR76yKPqPfb7wvVSp2DqpnN44zBmHyU14isDV
DIH2YKeoee0W6x9CAturUIFOgN+kqla+2P3qiQCDBZ8IAFZbMy4zLmO517kxmRV+dsQZ140Tyv/H
BcSogD6PhMrfMp9Dyl2uJSwoS+zYIb/zU01vGobcj69sGb/HQVjcw1cJcO30jd0VH93mqy/h+oJ9
kKXG7dB8pDwIvNFaLcxECsZf4K5qKh6yRJ5ceYtjz/qKU6fQWM8twL5C7VhUOPhMw+Xj4bnOMll9
KqALU3aBxnuLzCnAPHN+hHua8fuqoQk0JReaDdgGqSemoOFJrc+YaxgeJZNzNrTXO7JH9mC7M5T1
1v8B+FMJQfJv+c4w0PVqhkBwlcGmtKu6tJLLjnsYLziOnL1A8GyKkx6war2yep9hEaIYvfi0rHY5
rhM4FVpXr+jd8UcOLYbpAYdzse7fhynmvz8iEU6TBsvN+wUoqC3Y3vSurTJSNpzLSavqksZnlsG9
cHrsZV8++XHuh/ytRhtKqwcSNs8kkPXUJbHO3JZJQrjFVy5mtjT6EX5GFt5orj+mLlUbPdroWscE
mL1k1qTGTXY0ooVbqcIIsIX+znM04zWwYpmYsx9oUSJcFK//188JBw31yu2SvF5X9JEX6tDzZpaC
ClhjPCAJJk9wcnLcvWHud49viS+rqsqhNrQvS65IFZJNBQy7LVlCH5MgbViCyb3DU9to0yQgpTdY
SS+6zeW5HHFJUvNM3WJ17KUevKBDMrUiOcgmPXrlGYsL5dnap5jVI7+2ywpbYLsG5kFyHKybavyy
VVW79FENnpjjiEIgoG3z4oZhN9msDShG19B0wwjw8dx+sWOAyyVUAEvFRrwBXAE6Ai7OwVTHhKYz
KsUH/98jnfq4bAMrqYxj1Bdr/CHHaK9og2rt4qnaamHCZaNdEBMrrQ8KGWiTV2eVDJG6wXEOUVDj
+dMM05/mNZG8TrwnpcFE2zHkMC6k+dm1QtMYUafZwej9l3/Fz2ulY9DsWFdJxuV03lwUyoEWxQgB
n0zi5PKwMP+Bwm/hripHj9HOGd0mVYTt+cQ2VGrpMx9FIUFy9fUJvS5+oSxownV+Pgm9CplxEo8p
+GRXfoVmJ3YymlqWya4jPx17eTHcbd7EaZLgftkWOsQMMZj/6LV2GCFOAJSwich6bkUlA0+wYzOp
dSI2KgaMVf0j5bn8QDHtur9J7rRNX2RR6SmFvuLN8uk+3DmwNX8UYXbaYY9VXCU1HVP2nIOA2dF4
vN4qf/Qm+QTg+HXWO6Te1LpqdtFGTKmO0BGqTAm9dCJjGzfmNWasPih0R9Jp0pJOt/RZYA6ylUpL
kngZLEdYXmlfH/YOOwJVWzD4szqQ3QjZu9ZXZIwAv2WE6fb3s1LBkOnp/JtJn13Ad/DzMJT7j/HT
TUFIL5/o46V/qgY2Li4DbDEK+XqFXaDaWg6waOx4egsuIEYCRKQ16mGe/yBpUdEA83bVm0LRwELf
QeDYr8S0Ev2gBInVgyH7gapRmL5IwJoIMWkEbtgfet+gTIBw5GpPgEkTVKhC9I9Qdz1r1+bQTC56
V8zKragqvRsnjFAIb337et92kG/u6hZkS3zIVEb/tn5BhRlue97dlsP453l6CHDWe23QNDA3nRlc
b3SgBpuAQHbt7zLkxwH1MINnUSTFvAoawaYwMBTV1AMRKaekcS9V1BsZ1d0n5F6SBiX1RSRRqSsU
UeMXB8WhB4DcKs7aPyvy/PVaAKlvrZEPuMhXBiz6wk+VKoDACI0VkIGefpALLlW/3DcZotH124wz
pPoeCtj7feiqKRF9UPc4It16XGTH4cmu3NYZDWme5qcqefLbqeNfJL1ZF+u0nBv+/jMH+bmk3xRu
r4NBEEc9CuSJV/QpzlCPTprM8+LNpTLtXDFh9YssHushd+1PlAr6Mi/llHjCU3vtvwjFvyhPUnib
Rhe0p227RbwCrc24gnCmLUBHn+2PWzEExY3xwO5sPgN5676TnHjxZTaPI01qnpy07m6ANKVpKN64
CbSIzmX7Skdg9xHHmOJnKNBBKkXkjdMI0pelq+WtLDAbN1oDFv6DTDM2hUM5yD/UnPybdBlwxos6
Jf0xB/yFDzBgCW02VRMWWcYixUdGYqmaegje6URig8ULZ3CMv9Q4eyKGQZMQSNw7PHJD5uWVGMy/
ffUwNCq7TGjPEGq4TvxcDtftTBUSWISCxfNNu1iA1xdezlD3R1HZbfDQImvt3KCvsLlrbZcm50tI
Kq9HU+FDWVk/ovrq+n7Bcewni/gM9L45MfzSyZnIoQmmbuhCMs+gl5YLvoLGpEoKEtqU7WfNGVpi
cAsvo4wQSuOZAyxKDbbwmwn5r9buq/Bd7yz3/o4WIK6cyxp7F6wAC+3DDhiJJ0BMyHWzd/NWWrMv
jxrF+xh6XBrzuY+88rmj5j/Wm9wiguNmm2gSdxU4ULQ2RWzUkmytsXWobJMi6ucWGo7Y/hbwj/0z
WLXyvapWzIggEwsE5r2lUG7xfP0wx8nJsjelOLw+lmD2IzPP60BGKLfDwXGwOkuWWNy6nwV4rdnL
mFpwFBUlLBVnvCHq1Fu2d92xYt7pz8JV8FFLBjdMcxjHIfi1GXS2yCR4JqTSSOh7324idPILstLO
cyypuOZ2Urcu52dt44uPPXLXkvxTXiP9DGkPmpDBzdORT3BiNogC+ry7iqIFJAu5wSGas0HcHXCa
0QuDRuuwnSyXLRM8U45uhaUeYXwe86ryDbzdpxjOuJliIUfrJOLtlfvj3Kl3z4IWWOCCiKCe2mng
W2tHeKbyge95C6wqYpdUb9p7h7YgGH4rLr6X376IYH8grl91XK5KkzyywAkcPzQWU5OoJc+uk7/j
TP8KhTZ/mGuVNKCRFK18OXQJSOI9Ke+wJHNThiiSwv0svlt+aGC8/11eS/V1QWGdXl4ap2k6wSTq
X2tTRM55EOLuUIFl4RqD042u783irR3BhrNakCjqkKfsYYvKaSFHSauvkjEycJuZCKkZOqQC+M/8
Bgftu3ZomyNW/0Tht4FM/mbnKQpV6unjScXKlZzbrxzugJTf/l6IJGVsaD++hw4Sw3xOqop6OTBz
RB8mMJuM7OQsYO5QQIQwKznCW2igz1cytpm9Rh308g8a0Wxu7BsZK5oST/E3eGm3UmcM/Wyyys3p
0WsUcvVix/yxjMxEbUQsHmIdFJ8bIdt3+N7NRg2mYxVHo/uNKnlP26tZ1xjbuZjjloxK88Nb78Wy
NcNuFC3M68+fm7C3XUXU94spNV+BNH8vGeikxsmiYQJe2pyOEsB8kYXc1ON1FPjx9iZRnIP/rNNf
pMd1Xnf6F22vXB+STPJCAnR82gTYS41oJXJbAYJxhCXr1yFOPhZlYOlRaO+EySAnnsaIHYMQLMyk
EjQvNIPz/MI/9Jj5YEHY3pup2m6PQSrxRcDic9qvAnFx3WRoYsH+FfAzQqHg+FcXsh1A5IvMV4RV
lIaEPE3lVuLasLMrQj50GycVa04msfDHvYLVJ999UF6BLCEAHoXUC0jiFE/qRxtA5FmE6slcAnHN
wHgPo38213RmyY71KBU+upjzoshgZUGqNt/v8blRbaWT7O7ARuybtqcmS8YsS/onzp7mCQJmedjm
cHUmzsuTUI/4zkxeqUgMyfA2b8jasXLMsug7KORKl+zhzPwDNFQbhrVE2sq2xYIJ05/iGxHyE/i/
t9P6/2xs8cvdkQ5cyUPdE0ppwFmxLSJsUyONmLsahxYOGHoqvHt1Z88oicL7utSqMeW66cZlLjhA
SLk5s8/ikRTtkT05Q6aVPoFblQ++liMl614UwIngDqT3PYqDJterItSNmZOw5JulFRAxlHf3RY/+
VdcbiHRIL9NwQdaIiaTC0VDkumwRASjqLX/Kp9aBtsA3+bTeCN0lxe66HnxPTkeooTZxEXApHcpI
uwflyzbmTzWGUUMdsUprQSwZIMaeqVEFMu3hYf1+YsQg7B+0UbJ1eHETGl89PNXbhqEExL+cTULt
D7IJ/4bO6d3PkHtUowG5NsGc1qygeVA57w138AeXKYChMvZEOEsCmp7zn2TJe9orTmBUi3esKkPb
wc2UagPqH43vZyfUemBWXtxi9ihrC8oIoaPs8fQVVmL2Cak7c4PCji5/Hca/5nTXm16dgPXCqDQB
rvNfwsI4Vut4lq7L0pVVodI/zHF/PH8MsYK68OpyG3CoCRRuC9vIeh/a1FMvJSomBxJ1APYweSe7
zztThoSHHZ9eMDXZYxb9b3rZcdppCweLcygB6pJdoMtx/TnvNIgeozXP4hvAkC1yXAgNcqlR3jhn
XV/pilI9W0eRBHV8/noR5DvyIHq+UqcFQ1Sj2dbT5OtkTJm7ISB6QwaQREau/O2ZCJlThEB3Pvuv
oJOkHo9GylPUw0BYHUCbs40m38pz6ejOblsycCMkPGjRjmejiPUafUWMOiYbFy+/pJhNkBPGBxEv
mrnqEZIDf0zXeerbnaP/QGxXiFcMFGhS0Rj3C4G/YDU9XHN9SXQ0FyybC5iZwIGHYScK1IZyCBEY
IN09yZS0s9c+uIHmRljJNiM2Oj84gU7/qYWjq4ITDR0DFrftRZ8E/dylsalcLGy+PbI0ypn1h/C5
sp+X/QSihNPEc1pElGhTJPUZENjz4KL0ww7Y3y/gDswYoj5IUt7Tr7qSgf7+h8zcJbO2+acrCzDD
qqeQITCfcKeovnZTYkbHyBJEW/WiFyUmG0k3gtSZ64niadgJOzzryzQPH5loDnR5wVbsVhj+jpNG
1+sigH+CNItg11A3GhPKBk0qPmSow6Gi2H14LldRXWjNKgeOTsdbnlVhcogMqvHTrU4lZwuDiduc
A3usoPCJihDoD/7Wo3JxhDECLTJ0PTot90kGIjq1z9M1hZp0FJijq+iI3Mlgwnqzalpik3BPBlAv
CgrOViHwNiytecyZfxTWE0yGC0RBDtofXc6se9NSxKJ0bt+0paqZK0bOkuNwTBr1yM1oqk2X+UD/
eFPNOIJmKUZLG6myYyKkwMq7SMiykPgy4+0N6a+S8yu4W3BZPaATpO4aPTRLHSMjKFRhlYieOH18
10/qCxsQ/Nz/rk62MzDHjuoN0/epQKILqKabgziy9J8EWiBYcbV6/W86w19MUc4wbfbzy1nFgTZ/
PBT0wJvBS7H0mY/e+m81PQakzAdD26wOzlerRJdw9PTYZJ431zSNdH53lHccDNjlAZJY8deYPKUG
COxlC38yjiDNf5wbZeCqIMOpFJGqhlDjRZ0lwoNOzB/mwFALbk8/Khaa3n20UgHYjpc7dDdA483n
WoeC2xZJu5wBEp6fi1a1CMzZw9JW+rLthZtbdFmvcBl9bDAJMm6CqG3mkVQ8eWtTAZB6QMElw/8M
OlTn2R6po9iVY/0jTo32tJbg4jDT0eK9+wO5mBmdDpF6odBR2g0d5/KVT4ZceLOX0hmCm55h9kob
kaGQ4Ei7+WxQf3sfQrd1xEI6UIHuhgE4oqbsdVrww/6gv1hEzX3uGTgU4Hq5Usv21+kVrHwR0t+1
9EbsqEGHe+LRhodd2JGGmw0mDyDm3nYBlkMaU9N8sMp5zQx+LSSsAZDmHIKk//gC0p1ItABTddvx
Qya781xhOwMk0tNndbFwANnTCmnpBNalf0vCrwE502gKkpmE4604s9n9josUsD7SCjTfkbQl0WdJ
qNxMKM7azip72JzkWrojiqoSA4TfhtmJ9CSLBZBoIa/rRfOSZoumvwwqME9ZIU6HS3LvnI+Cwi6+
6hy8v0w1BAUqiQ9x4UBMg7Ot4HLenCZwiYQTIAv7G2PbJgSzcjsK0GJMNqfwrgVe+pwguGIbFSCp
hd0UhnVqVzvtv/IdEXP+Ax6zIuo3zJsOcn12aViaVvPy5QXktbx7yxIz/f6GtvZhlNYWst8Xz6XC
v18pgcz+rvDAm2PUxg9Z2ael33noMTXn6cZZFln/2/eIFnQTYJ+OcMqv5KkBJWz7rVuQ2CyPIUEx
4eE8e7+njhaweEA5Bf3ZG7a6T7WZKodD2oEqu28UnTgmjRMEUr1a12u9cqg07HVljfEdxXKmUj/Z
1qX0TBMMXg/uBZYzVvXOo1NTlnSc37Xk3c90AEsixgaBuAGYJFV2GoP6XJ7xfryUAY9ct79Ak4zZ
hjnrnRfDRjT4haMRT1kwxUARPcPSlpKfpLUOMxGjqBPbKfCAP+nDN5Ka6WYI8GliGUSqYc+JxAoz
/h/dTbpo/gXdI/sszOTCEoihyJTLg7p4MMhiNh2Uyo4C8Sr9TarP1fQCP7poGb2lGwvNL+r3bDPm
TwUvlhz+gLZh93koYb17srigGJect/IAD8dTO0U27INPSFDcfvCd2Kto8b8yBBzQeYYCa7XaI4CY
SOo3LCI7NucQwCjRkAqVCosJpSac5b5iE8eWJctMt1JmB+Gs5XcnnuHDxm1E+AxY1RHwSh9GBUMh
ZDTS3iKxjnPyRB5+dxdoNc1kLT3ZGW9FHJ5XrKVsAAAHQs+K36QydXLRyybGGGJ1fBRcDe4eZqwG
VPL3t6zPzCB3rrnIMfaiB4ptfNQ/LC42BQm3hNveH2RXl8BVriZzkIKaiEL7bCW0gXh58bus3b5e
foGN3X+T3a5JVh6/I9Kgc9xqXKes2roFSXRsXweCSAfJxG6H1CKT9RxEyMWRKpTcX+IAFa3Vf2bN
QEGzRV/ladbQBsOsF+GwxBDHyS+myZgHvfHoEa9VMq8tBLtIpbTgszs36PSrBAOO5ZtPAskD5Ngw
JLgecmau/lMdjcA141/NzNnNGWgTw56YepMBcl7EcmjbS99v7aH2ThSxqWwQuuTf/6wTsZM1ReWY
/CaGULoEhcxNJiEhwhyFHqrPmDzKh6RBMPtkIizW6rRDcXK4l9wmBlCvhonXig/gIFJfL6jmN6tc
7O/SCtT8qCiQeWKmy0TIq8ApWtY4BfHGmXfiWmDZm8ytNtifUggwP5ykMIPvAcD3OGpKhNz3Q49b
7leB9/dnkqVJCJ0PsJGxZwc7VSN0KBxbzrifc0jpQnk0ON9NJh/X8kNC5xYU6dBH0j1agxSYML/W
wBs1TyAYXDnFFqeZldr7Zo3qjclD5paymvouFWGY15pQcvBY2Si1BNANYStbhIny6VTlkxFu2FHl
8hFwRuMPRz6dsiG32TyiTOcmQp5AzSIOvYlD5dzz1M54Kvqlhlj3mIbPWsIMzHOQQrJbZjhjFMnP
TvWK0r5w1CcgLthFOOVM8eNItytwngMP4eTCkNWhrDdkYb2nB1ECikVbJd9FeWRESOT3+anssuZ7
8Km0qPWifOtW99//THdh3BNTMnxQ+4SKoCsq3CgfXocKaSOQOq3o2o2dLEQZkHhqpmyXP/MFAgNw
LWfYNH/H3hSs/oE4MBC72X3NmP1SP9Of0KpXdNojXm5sdGPbJCzbftopFzZj/9ajH0KbaV8X4X+4
pWpYXBF3XvbKgJ32Cx8JsvgbPqJdRUCQ+CJQs3jnpHazxPfT0jlO71oRXEI1BO6NOiKK6G5BvVW8
/+mjtlmA8hPmwNCGciNb385cWxJRZLlYs2YnEzhyWCuote8tw2D+pVT3BDJdXlPeelnOE4FuE1tO
AFEjRcsDIvkBGSHYWQxcEGysEF83c8bJEifPFjNjgewQ05TxWKRKRY9wwhCpXeHFioTqdxWl2/aw
o99Xd6KSkQMuMyee7Re/NVk7XKZawiXvo/+krAD+jY6IogAtQ+7KDOx71rsGS/St7zUj8Tp8+HMw
CrCrUXP6w+wDo1hjLblvF42bwBzQeoGCLcPT2gmgHI2qSbC45YlDuTLPCSZh4qBU93UzwQj4zMdF
pcyn1sam2Nr4xqJpnZhHByAUmmT6CTrLcgKRoCAUdqUe9P+l6dRL6/I/Txcmm0dP3Y4x5TzzQKdw
Z3wEzi95Nw/SaE9XXw2Gp929+Lh0mEph7C8i2YsaK31i+F+lHYP6foe8UGqSkGzA0EaiYYuz5bUV
1XOIdsNN63YBaglEe37cv5JctNpprTfrtZvnySyQDviYEULw/RpjP1qHJ5/MO2fV4Nc2Q4JJhe3q
lBmUJpA2MlHDRRDnVyCuL1txbvLf4I3NxshuKpvXTunLBzKtPk7X9SFZQR4CBTRE+uhEc4koF6Ps
IfQPsAtj5hFOjsFYNA3Kwn9vj5U1c35XtUPuhVf9+cNupzpR8RHq6IaDmMYyt6QgdFNLK2tbv4P3
zfwXxOAYmNmnzcnNt68TK9Q+/4kxnQCH1VJzfqljsfAtNlBKMkSBDR0sifE5rjF7UNbWUxlVVnH4
e9mnh2PJOkVjHSb8zwifr0Crz6ulW8TqSUVfkyyqA1rKGILHhUNesh4bzoM5hEaAZ3lcBf5AIpKm
MR4Mna0kLr+uKEjFmNveRWkvvBtMdwKwLLXGaOGKh0B85OFz04N5MKQPmDXiqe3UjuFrU1PM4Xso
Y2BX6EdwrAYOaRd2AAx5Z28N/xqwjjXMhAoLz3OlBNLBeE5ZoOmX1p4t0vBSWqu3G2dgwbSi3JXS
hsGZsamzddaj/G/Zf4onpTnznAKIQYCSkndgNx7kat1OhUatDjNSWXBlZ5523yOJcUjJ4GNi286/
9ivre0fhtEBMELfGLj3phFRARJU7evzvqbnCtBAn3JGTmBTqMlHanyFbiL3vdISaSMqKRXmmbZIi
V9kGUELZBHMnGkLdJtOrFyYuMWba8z5+yyGckJISBfZlAoe3vEWFX+1FXdhZBeozOB6MudNvYa1x
Xm3p9T5qZSMSrhymgMEn7u/mfSACGVSSKjNXwMg2t9FP70ewYOEsppXkTnvikbO8dJgupAmlmdxO
3Oj5N5X+I2YMIxauDGZ9oZN6ZyuSlZl2CWjrrstTas6M7KO3KxOTm4hHwepkI0Aud90FyzvXdtE0
9xLnXcJw0M7aVppKzBIvH0qMlcPF39/2fxi013ttOFgJ3mahL9YdQGkEhWCY8ercF5lttrUwZOOQ
b8g2gj1zDN4UJhzw26wWLbcOhEsmFPhXxOsS8+7ErQ4euKUU0V82ZvAq+LjFgWZSBuLAGSZPK7a4
nsN4CLQFjF7kVH7tZ1arjhwQya4joD1Itz1i4wGPqH+S05Gv0p+ny3DBOTap5IvtvE9Mizac9JFn
/W2o6/RLHAiwXgU5Xcik7CQc6UJr/lAWs+xR1il2JXopOfVDEGJc9gBOdaACjam8vqEmIGxa0T9t
eGB6OlL853cEOsDA7HqJf7AHeHan1FSoHUkZ1fuDfFa4ZWaI8lCYJ1lDoNLF+2m//BHdcHC0aomQ
m3/CncSTHoBBRu0Z07dZgEzJtJ5fDvC4GnPQLkNZsuTjIUqyTohltWOV0iWZJLFyp87bQrK+w7du
sBsvyrujR29S/OFLkWGvof8EV2LbxR12rlQjTNrqz/Xfrs65Sx2LXOGkr2+pNRYxGEYCsUqDEDA3
2agQkv+qHEHorldGuME5GN5Mr1Rwb1H0Hz4+FMvX3FD0nBVtqGc5wQBeWmCzhqan4X3dpoiY87ZR
Tjs/oY9n9N7HNDHooUU+0Cp6VD29B4V6wu8nrMYRA8csQYHFjSHg5h8fXRQFIPnsC3iZfuN/RZEq
8xrycCbRIFIotIFdLqC7wlTRJMJ4VndE22kzI+wNn3XsrxmSMDmhf6ha1JOcQuY9G59+WspzbXL4
jpfuf72VoKr9WEewvj5rEYwq7CoIHmwhpQ09DnaODg0e2him9ye/bGB/vmFCu7obt3hh4l01R22L
KG1SYw+MeCkS3+mKIjwXtPpUWyaCSYDzhbTyeHSh7RWlK/Ul6QDh1E1h6Kd3ad53tnlOy9ipwhFa
sdTWA0+TbPmpIgZejFw2p1sEelbd1TKS5EPhY7S3tEAXReWWedewZjteDMilB0HRZ/7K63E2EB06
m5VC1eOr2q0QuRAUw8r2+wojkzn68ulyjI3rxuLG9TAiwncpTWH4LR3SrGWz7zKoykYMqsm2KKyw
AuqhgzJa/4Xux/qv4rNOSImyLAQBgh5vRUykAAIdS5GeO5ccS3vtK5VkHsHQfVfCzgVNN3NZF3ef
QFZFaTMGFjLWpz72I0393nr8AvYISRxFHJA9p4RSAspYydOtg4n64kIBsY8F0MQuVJwVNNhZBKL4
8+lE9p6QLDa8gqJa2k1e3k2WSefnWQY2P5yF2+T4RcF/4BdT8DvKVdhoTPnndtNAYBh4uD1hSImn
NqhlKXaSV30Rn4gM3pEonov8ZBvV3WbDidwrPyoWFlpqANigadPn5l3lI9eKKDVHmaJF26D+x+Gx
PUY18f+ecV4g4NH5oDtmYWPHBZJP3/3MlhteAB/+RDS1/R03Iq2QzKWDh+TavVTXL8wGYY6KpCWI
tlykvEl5JxPZIGNT55yB9xhZkOwB+9vrpTeFiF7gm8p8fIGdAIplYyMEOGqjlOK6IE4RjM9Ly46a
fch5eUhdwL7qd4lGGuwqQWJz8yONsIRK5mcLeatfmTqw8e0OTh7BUbWv+YsIN7CNdhJmMDB/MiG4
EOPuNitcYjaKFFJGsif8zq/r7YKrshY7jO26ExrtAl4DxD9CUzrK+ckPDiiEA75VKd7AzZKcl3DE
2+S+O3mL0xbV3MDVv1AXCt5f74c5mRtj831QqsAtqr8hgZsyQpTtrjz5M49qbr2h4xjsDAcf7B81
yS+RUfUUL40m6EFkUEAqmQFiFKrU6x4x8iEbGhfWDfsAF7lC8PMTKHyf9hMrtjNzYob61M4imqjo
vAsUJNCer4VzJ3c2fy1hGmS8sPnxXpmV4kiljMvahgHpkyLYMtnapuhMXj+9J1nL5t8F/1HaUcML
5U2jAtYnRjQTtCjO9o+TBv8qXLti5m966kc12rsDW9Dtr8drHqvHtRzeWViW6CAN7gmlJSl7moWi
JSDAU35Ibs+Bhzhx1D6c4QOCUibGDXbRT4R7CgxcW4fRzeYiNwgTQTfKt1wLCtTjiUg400CkBA4Q
lZVVrRPoQHHg15YuyCmvMrZvd1X2LBjlhNJ1z0WyGwanIcxAdqKKfj9MZdYLFlF0Qcznv0m3GjOs
Xry8nN6hc0ur46wwBzKABvcNsyTaMeb8EGWtWgqbbmGTksLogn1ltmIeJCmRPG86kP3TqONLujRo
R4avMLEkb1pT9qEvCFR2IRjRPVfDIZrt0LecN6Pctx1kseLXSZnQ4id6+UFjjkbmwpAeyIrbfvZt
30dXNKOTqKERY2NBuT06KED0NtwjB652DMxpHm6WR3M9U4cpS0BOoSSzFr51G32yF5QB/IXpCLgF
sV+TqLVYqz2X4jnV/OofiAuB6yMi3jso4yzds6jba49WGFofjkC7hNUKZcW8TMtVAufOIf1yYhbS
TM9LnjauxiaMun4g62ZYyOt6ncW10Z0Dtm2ReRo3pCHnjd4qAiid0qMIcya12Oz7GHOvDly9L5ZG
GwSoGM13NbeM+NfNmgiWZ2hSr58vUg+5qMnaU4Rw5Yyb3mehEoKtetIHuuPSw5qqGIBQCZAawNiv
o7QpP0yQTs/6m0tEkCYr6wUp+0rlIKwVWlg4ymHcdal19+miU3UWN1rzsq2rObpS1KyxNbUV9MlG
5BVHqr3SNhCoF7vzrj9lkP93IJl9hIGLW8+mUADyaNQe9UcB+FA48fWdKOgBBwl/sRSwRTbykp5t
MRO13ksQ7Lx2Wgd0XX7Dcb+xNo4jKUmjoHwk1VB5E5/xjHh8MWZBy7s7J33UKle+0pPxpX2aVC+w
tRiJaZbWR0wP+iiIqWz4HWZyVcLoHdxVq3/lI0WHufm0V+wmpVCMi3EORPpdsL8kvsJfI6U+c6p+
U4XZEeCJ4q0ZJqO8XyuidIruvbMJrw7vJnce/oP0UAYxQ0oomc46146t02ehHgUzwojsmzE/fs7B
E/cgGbbIbml6aS+jyS8jizNhdY2XhEICr/7q+c5+LGGEHVnBDwUrduT5RW78XyPstWB9U2kJGSI1
jeb+rSMCG5N30KA2EtRSazIM1w37aQZueoCqkoLrPPDRYXxDMzF3j/16mNT3o/RXr9bvVG07abSH
cGC4ZLjugn8fvHJa5Foq7M0PaX81qBy0xKLIlHdGpVX7/lxP7fKFF+ZIazQqnTna84kDJJjy5lhx
c1Pilc6YT3dGGvD9tXI5A6rP6mCD1yzIMopgFcWZCXOx0vboNvHgjprdIW/OmKCpKrcq+TBQlRxU
2k6H5aEY31anYWOymKkhuTJiFYsABoXr6pv9zCqUhy9aPjqkFZpPqASvgRuHBN3F1QbdyvggcFua
d38cxqzcV5v1MaJ32WklYs/l7LK+OPCfXnvkYD6qoSi6SmngvJeihdVvxTWJz2HcMDNOwHUQCPHu
uhnafuZESKELknC2wOrCIpAbiCC56juK3MZNNY3NCQNde0kYweE2ns2GxSFQ/XllyjEzn0jA/D+1
P96FaIjsoPhbNONE0J7nvZCfGq+q+WzlmQqXdJySFs+oW/cmV3GE5m1gnbXL0TQcxZ3OU/HjPXBM
X7HSKLecG9tvPPHCUxWVhKuoPc7d33cKE/Q2utbKqj+SIzYHU63h5WbeIu7a2gsm7P1i6wmNVFaX
ZOSgvBjgsyg4DMtnK/T9ZKHDodhYdyjq1UWFSF1En4hROpovov+we5ha0vw7fxMwValj8h/ENqgP
DBehgXCfybiYEcyd9z2GUOjUWyIGFQfNX7/VtInOkVFVp5ffNBs2JzXq2oo3YpU9cMbZH2/QoRJH
iw5L2/Pux6qGDysxLM41k8lT18F57SqOZMNRGc52DYome8Akn0R7M+8DkufBbn+6IThAiQnWBdP1
Ao77TC6MAyu1d28lU1LGNjc1blTvnMxUEyM0sNvDls3pEdiVqmRK1pZsyTALq7fsBZtTgLVF9HC4
zgG0xquMGEfmWT4CIKrJkZQzp4UUqLMbIsi1ytt+Lh/ouuXVpUjoUOx4TgeKMdOPmVNlYrtiDJ+q
W24OLxTg7+saX5Jlt7mgNGxikg7J67q8WttHn/FA3/bYQKN+QBOG7P49Xzxv01tOd/BDAu5WKK/A
bHWxRz44AbJuDF+qSNDxXy4hmfajLYfJwsP+3EaZFUREaxiIdaK8qPKo3mKhTymeqS3VO3jYFvBn
9ya8kIzgPUso2urNxISGtqCQ29SdAjv1I+Rr+62V+MLYh4bb+lxxKT8aRCl8FakVKl0ttzNSMVdr
IRoEkmt3CoJXp3Ls1+todEsHnUelySq+OD78ghncIEmc9ezZueHjdUuAQPSGCf8gXq0VQj4uRgOY
xsi2ye1DbX9s4d0dDrnT5L9hN3B8Vog4TiAr+XSsJ8uw0BMXUo4l0LkkeUerMYcmlxOjJqhxLARD
5jsVZaqveIgELE1N/n0x6XTuGWgTp/RQKJSWihpHAb7PurQ7gxVfDao321Bor+wr77e91DBV4pya
44UnBGfMat4erFnRe8XoIcLcyc2WY6XDI1vmMfl4L+ZHkJeTW7dxm4GguMpBkNBLu6/2D1MFkQr3
1/2S7ovtflSsnm9Bf7Z74nrIu5RtE57yhGocaZugNoqn8UZcibxOoOD09Sve59H7IJZzvnbG25aE
+psjYpyODccypt6nJEoe0Lt0aNGzRRJEck5Ir/VMRBBwasefx1q03PF1Xfh6+yZBe2fWMIRzkJx7
QyiTCJLVtmbtyZ0I6wic6rmO1fWxXk9Z7rcCwIFQ53govQdtfMKoYZpLRmv7vfdU8jiMp72T6ZY4
OV86yp6WzUSDZIyCLeIAR0fn3H8FZhshrEIbI8SooiOi5gI5sZ+6CzWj8g+wL1p7zbe6i4jDg4N1
jHHahoxuTraGP5FqQZRKAiIAuTYecxX/ez2hmr37E8ljd0OD6nCVIFSc8TXDyZ/vVzEAScXQABEI
Nx9kfWt/wUgXZytLiYYHm+23+FBlqHn8ucY2e6NpmRnY94fioTdBqHEy6QcLVYjX82Z1z5LTetgs
2CgrQgcLB74igILyv4EoN08aCcg4pncgn+rUKh3EajzGY5SwGv0QyPT3e0NNmzwJuCInNfIId8Mj
XiPTkPQfhJaIpx5CRtmou/yE0Bb4wtqERwcxN1aaS4SnfDJSs4WgRk6Jp5XsXDLi+7XUJPHRqEQf
WrNvTW8jJJrs1U1dIhBC2DRnl3pE3MjtzqvK6Ll5YYrBOPaQLKr1HbiWhMb3AxidbxQoh8HBAE/N
ZEJu3h+JpMTT8Ni/nqXU3eDieaG5CrB7bzU21R6DDoov3a0m3P/rbM840L8ePL78YaO19AqfwiFI
sOFVw0jYXKrrQrSMl8j/aS4t0a7o9g3ZMSJLWY/Nrykhksz6GPMGFYW4yl7K64HgXO+iJmYLXCPA
VptRwKC2kIOYK1BJi1NU85c1chnnwkP0b8rL+5nTPlcC21Eqb2mvRkuknOVlULNHjdkvWw7UCaHy
2RqB33kKKOoV9jliK2hpPAHPe9ZzC0sjpsZYMUXuQkuh5Obe3kF6JLDTWgqN8yMv3tyc13LAL+PL
vL4RE7Nqn3kmWP30iIs63T3Kg9qlxwhWq0TeQRwzemknBN9+6A4CAX0xv0TKBmBHZAL3bHvfYtUl
YMarqOyS1yQn+WVKmtB7DnbPGAS6P4l08lGgjn3+DoJP6+GfksLIIVrSHq+L8DlVSPFSKXIam4Qq
XzX8JIyeUDPg2lPucfu9zNYEAM5T95opOVfv+8CC8EVu1IHPswHghwL5wSjNuinsRALx1SDbrigd
21cIUpk9dxIbgxIeQ8vdR5U+o7gy/FhKI6dKoLlMu3q1G1Dwq/gY8vUx6Y1gTlJvkNNaXWyehMF+
GwJeSQ9dC8EEfKmWFvycHqGIRBx6LTrLhCAVuWWP/phXpSf6katsvaafajnqSSw6a0zV9PKoZM2E
jpx67+iwouwMoH0ZGd00uQHgn35cp/FJaL6UtQhan+v1qbILpGC6zTv5HW7yTyel0bZHFT+g44uS
CTI9+LGr3E+DiuSO5hIvXI/ZNSCrtZP7KHf7ELrUt6NWu+FDFQxDD3OeAKscD6F+inHSeqz2cQlJ
Oi7csj0Zh9oIxs24jDvhl0XwBaSzyu1UO4etHI7qIgA9UmLR+5iQIpIbVFKo5fz2TjSy2nCafw3i
NpE8wgp8avLzPf/tJDB5UsG3MoEpznJ7Ac/5Jpx142onI2M8CCoHmL7ZNKEB411x4xUxoiafc3iK
IVS0MiXC71yy0Zg5W8DpMutEBXqi3Fa4fdOMKJJasafRd/fgFPoeNdoBcnPA0ZIH3EsLbEjKGDeE
VJP+wp6MPssQQSAC4hrGTw0Oekq5CiQc2exuc1boPbdSuzNauvc4pI7ZW6r4CjVBwh7cvLqNmOzh
0WxZcv6jb+UOqLekc4Ae4j2ru+hFabSM2Oa7b0JP40Yog7gG09K6VYa/4sMR6Z1owcpYw14gHt9y
RpbniHVVwNULfdyOg1OZjFut1J06MuMSNZAojzz1OZTg3QDweNA+CruTsc2/fxC6zNYQepv7X+UH
aFDdoQMF45brc8HsYDTPFR1zeWASzKLobgH0eygacYG5u9Xu/fVC0zbaGd6vNN7n7lhWc3H77doe
+E504dMkFOWP3YOqhBx4pj6RKDiXGr0FjCa3EWKKDCnpwpmJcYz8JB1Ks5xwmycbraaIGBpYmeTM
UadvlkbjXAwlCu9aqOZdFFMLVrXOcXJTXJDI2SQBuAFYeD6vdmC2un0BaahTNqlGFeWe58BLRfIM
+yHS3tBOr/b9OFUComZDdFCeT7v6Se2/0OvWgk3XLdg2Uoy+o4fANyyvyecUBNByItf6RdCBhFzI
TjJh8w31oSCOmOgTuuWTYp22SaBm9+Q6ih8iGv8syqR3hvICOh31AhC+nbzZ56N909O3vXVBwLot
d9OxDDpiXPazt+jJLo57Cejj5BD2T31UCDP3slZhf6ZAhot9vYxrGQcqtuy/1dlv5EYIeq3vzbet
W1z+9CcgNUdFnhY5PhoLHpoTXYpXryCPqwfbgCAV6ht3soiS+pvc6gbFfVnymcXxfmUdneFCoDEN
J1cf/oVGxGPapvT5yjpMx3vrrer6HZIC34JZeolpmrCIBmMEMSw/4h9bXZlFHABK/zXoJwp/hWuF
pB8mVLlobDJbaA73DkJYVJKnS6JPHtemc3UZzmSTikWVjrq4cRY3Ghj6S+xhX1ZFee+ML30MUIwH
aNyZok1v8Q7ZPB59YzJkVzWnZVx3e2W3UQoY5VvfzZZmK6kgWvliiDdkr2nSJfz7o4nXr9+wDBAj
LBwTOHCHJrzwj2RGtU0KU92AD+e+MwFqipvBQHtKp5qP1QEBJ8IJl/eEjZc/XfuO/ZFhBk725DH6
7xX52tF95o0BaBNHdUqPlF3JslPIq73nt8JDOLlxFU6A8r0W5nj1Xbquee5X7oeuc5CTPuFtDMNc
0iXtmAkC8WVo9TS3YXuuO/R/w4Rn7g9aECexGOki/bduH9tinjr/WX5UHZVZ2rRzd3aTOFIIFRUv
g7sI+eUcALiGLedzbeGu/g/wfH1yh3nDvRA2tXXDsTeq2g8FIHDsOrd5A4eEcmA8qGHb6opwcqZV
sC3bq9xkVjkqxzdhwGsHZ2yLePa56JDJYvkL/EytjtdEEK4+bEjWDNNig62Ee19QoypvVF8kCu7m
5cEwUGtaEE1gZrLJkor+6jMcrzDqrE+2gSzRG2gkwlnWYiZINqWRIPnLuEUDSVeImNBqXBYpoH8H
Ww5plthbex8cy+2kRQ3c1i9DQghg2fRe1VhLLlarR1usHPgOafZWTqaokvDzA3hDwMdxXk93EEy/
0VAOinPuDagcxTvAd9hZ+hz5Llzcn3w6fkI3fiEqjm4qbWoM7Elx3aITrn6AlKyNw5gPaE0WUjmV
LxAk+RVfyRTCwipsTpcSsNyCAPv7FafwjHSwVn0AwHIhQX3ST5abkbP9jHI6ZSrAipb7bJ6AbPIM
m6xdxPeanwbWiNCJSeHKeT8VLV/T6ForcR8t8vgP16MXZVML1gAdKlXjygoFlp/oV2yE08Y+gNyN
umS1C6bmbkGvgsESGfZyHIPsX1aEpFcOFWiENU0t0v0YFYCwRjr2iourTwidn2IhlHUo1ZVrFpor
By1cKOU5G9F/J02sS4xVra9XGk5Da9PLs41nja6jv/v8fZmj8fztm/cNiE47689EX4jow5ZZzcop
1a9F8mRd9S9rOU5C2nBr6TRW5zBYI/br3+MDr8asE0Lw9pymIUN7sTqddUzQN8uyVnx2JnQGnSHi
JVltKdAybwKp/7mkLg4+gilQKFEcn6QJ0PeaNE7J6joSkc06ZMsNixXFA1QHUt744qjd1Ess5DjZ
rByRoxap1bfgpK6q3XP45Q29YJTL+WpBtzCWmeqChtKDg4/n1kwiGUuqzO4xS0o0nWzm6N2IdPma
yGlNzwz+9Jj3N081UynewTmW3ItOB0z44FeCAPXQJb+wlGZ3amL4KMWP/RH7cs1INZVWVVM/yAR2
4D9RTLwBomS92anjB0xrkwsCL9Wwco0PoqKUgs6NhixncqOMpSMpCKCsmPBdd6f4ysp1L2K2Inzm
kD50bVuZ6pfYeR5zT6pn8uSNWeo1DqQRyuIkbWNbpyh9XNzZKmlWU2133yklmzdm0uWw7EdxE8k1
3Shpa8EL0cYfdAMu3M9VxxBcy/o7levgJsajV/vE3Qdb3Z7LMGgW3Gn0fr4o0WPRqxKi0LJpC19F
U0fOl5C6GG3u1MpeTNZ/33W167zeW3041RWg4UTHrx78/N1nSNqTltm83/uNgQVlLdBJbt7M5NwM
X0EhGJT8fFnVboVRfZqnqSxD582hi1u1lG0Zg5tGegMSj+YUiOoT8U2I+Z5EqBuB3Ts8IEawP983
5st14lm6IDV+QsGypoHE7x8bMZc42fHocOyabws2mkWDRVBrn3M0AA8w29QUd0VfyERX9e4T3U6x
ae8yZAepTC4GrcTYI6iJlYom5qc255+qIpWi0Koh52lKnMAJhc2q5Se3Z3BeqHd5RXBcXDyqWJMM
b9daFIblSneTjhuabjFoqB2wAHTdD7H6huMXlPW9vVjwwdxFDAr4PdpT4CN1OpKVP40uptqNMdFw
u1iGTvaoP7lJqvqIzT4TTWVXYyMVy6x0sdpM6VFhTu7KmsiL/qkeLoCxlhdK2d9c+cebCazNkCxN
S1VoQbxlWLBKDQLnArYn3eTU9vyQxggYmrfnvQt/bEw3hYg4zBSbewepCTBc14kpxAd/b/6nnUGK
qNx47Jz4in7hpeWwDJApqMJUw7iKytqL+Cli5KbtQ3JIplr4K19RvQGxV8UzhGdyWUBEnu+dvZon
wHpoDWKWLavDOOkTN9ENLrOMUYOdLg3B51/5RL8Wud25LCrvQRbvuUvLBowh6q6fRyrDJMQXLQrh
VzfCxgivAnJ0j8cJt++1r0Vw/uF1zBiG/N+dWud9VRCB74+uUCNV1esxcc2SlmkaDzIW6Fv6EpcK
DnMlHq6VNJxoJQ0rwTMJYV+TrK8mQHA6b6lnk2JZ+RO46dhmhBZbSb9e7YBYsf1sLSzx3djQXERE
NPRgTT5746uXYXP9lN2l4OmPS3SCWF8Lp5vojhSemH88v5yJrleymtqxf1l/owN7o0kNXY22qVCv
UVAsOhIX2/sxIi7/Hw+n9u37yOiEkTXnfpbz5V9YPW49UGsOlWfwJ48/W61grYlm5nldR8L9/4q3
tf5vbFThSzf81HxYzxNjxIPkIYzQHXwJWWeKgJZiWf0i4PjkjQN3YUQuDfj7SoFrHG7OkrNgcRy7
mue9aau9/upE8gHCuD1/42t6Lo1eYU7NQAs/YHySObY/Iyze3RS/WAFODBULiQ0YKjDfu3LKQN5g
ugtfetkKwQKVXNUDMBWdSoIZlsaZzdtyBE/Es8uiz4EBP5rZ33lbChXIgwZG13lLu7WxwqYMd5iC
qCSvV/8XujHuyl6ALYw/QFJMh+J4fRYCgEF14OKX3PG/HVx8AS9FZPFL7Wd5b1nTNfo3EciKuEq0
92nraKZmYwCmHyn6ySctMnls+DWAXApcu7yO4tlj+VoX0bg2xpy7fi+9U/Ld5cwUEoiaY6FXYEDI
99BfFxd5DeZX4N9Yg/PFpQSWr0OQfoNVZj3Ly3N1FFhaG9utAs1AATYdjux39YdsAdjNgfx7t9gq
P5jgNOfOQi23YwFaEKhN+TDI+gatPHI/HjSBwk31iPVcCtIvrafXb/+CNrJ0AsExUyQ0vjKrccKv
bGAMV0R0u312HPhNPWchq770op0fjcGkPA8SZabyoIkYK0nt+lugDl7ncrLRTGmNdmqw2I9gLRfp
IV4/liyqkB5aQMD9DPalus1E5h/VxyMs0wEuqr4FKoK9HpJ0576QZ3YFAKYhpMoDfG7DCXBGt5dG
WdoAR2lcm3mxwGZO3NoSSbfaiXnH8L2TkqL81XVBu/PnViyw2qi4nrYsu+++Q0eLo3j8v2YTXvH+
4Vm60zgF5sL9YLyIDSK4rBMMISR2k3bnKiQX8l/SczPZ1837o81B8N/APouHcieTliENAXAYdMFH
IXuxier0L5gpKSJclLj3RRcBdglVNOMVixbhNhOKiGDsDwnaI91gN/Q6Z4WoVV9zdJRxgpj6tA7N
+xRg+tVaFXsgo0c5z1Rk/K7U6HP0Prt3XR6jmuqdiaqw0beuibXNNwbhSzHcAv/ay8NgbIoHFQoM
3/nP/WPID8b1TCYsqPgopIt0khdoTy1cTk8TFEaa4y+0XwgcSnXmVJOLBhhHgg9QgcAYYsoec0vJ
1z+N1pC/mMu8t1cKhKSpZLSGtMmRF+kUgn4Ux1slNi2eJMzvoHu9dsu+1TO0H1Tla5/y1QDm/B43
+NZuMvx+/QZKJB+cZH0Y6wuKfirIPV7gdt0SQbGnJE44bqnsBwsv8u4t8uwSzTw77aGI2SZVnHxN
NhpRoB6/VWOc6JwYJVdpyXugOqmRlUT4vrj4vywpnl3PjFB0kihN75Tsob2ZcFH63gDjKeotAIyo
hF1zmwT8LvWdKNKMGADRHftMV/IQjc6/dvO9MFKTpyKdxfnaSUiDoLUZwXHDOq0i5EBpfHxMF/Ht
EZ8lUqjeDoRSyWetm6GQJqqk7h5j9KYdtVbjiFxEn/P794mekNuM28Wwmkjk9er3JG2oHLwnDDYx
OoTVzBDvi1t74mKJd+zpMh8akw5ok0CzhqjsCwKVzERzdP04Vl/I0sbKYtJbTr31u0TTWeSDzo6O
mwOjlHXHiVu95uqNsoK1pudXnfJ8tuML4PJbyqjGmiLkHp/VwfHiyjRsdkmg3VYS1y6v+dkENL2x
9ntO5CcUvanJgwNtMr4pmSsntcahpoZJCr2nG8C/lXUKCc+IPL9jKW+ukejg3P4g2CKkGRaf21OZ
7YmB5KRzYfdy6kiac5i8g1NP2uY3LJ9wk8V/gp+oo8ETqCaKfnIXo9+/QtWi9Wcj2vkc/FWIz5zw
Z/sCDyetXBtg9arJlt6efNlTCuNITen+TBdOlEsCxvCuWZPM946oC/dkr+XiUzJhX8hpbfDOFp61
dqKY7k4VRIpoLryB1HvxOXzmAWuhfa3tkR5nJD4H8OrjB+T9oAY4XJbJlQsYS1wQTQGucCTLD3Gj
TsD28WlAB3TS7CfomKBLDH6dpKim67UuqOMyElCDOcE6gQIVBlT3a7k4DG6nx8P9TCvA4Li4Ancf
/ySPmrNeFgZQWGmGQFntuDxzP0Kt5WlCReTGosvq/8ylsru+lIQEFvqRYMPd2wJFJVXW7ma7ubbS
g8Ka9znE66K+FAYsCPhKxTgR4Y9cG4hFVDIH27pssS/uvMyT9qmj35fmHOa47GUXpANWZbD5PpDd
CcPOyqGeun7KywJ3u6vxOrF92DEm3YFpNVxvNgvKtsc4j0BwG43drRGOMsMDSuqU3fskEEnWw1XE
Smc89lX7y4qALvA6RzOiI33FxflQAqFtZgC0v7vcydN2ZYKe62XBfkbrZ6oF9Pb8TWyjyj0MnAr7
zUoma6dDdVPJVk/D9/jJxuHggBt93HM6ozdH/4UBvHHeXwK2TVXSMPT7zrI5XDl9vGNJo2QBxEff
U2RAh3G+rFJJVFj50iDl60FukiFwqaWjYYZcYPR0Pbjxy1o7Q4onyP6J0owQZi2w3b6vie54+XEO
gkC6pfnpgiMObTNbyx5bFfBkT/AHk2lrcnunHqubn5iykUi5fItjkUbK4GTaI+0zG1wPQI0KzYk+
PykizNqGVgjeDAL4aS/ChYSYVDwKedhIU6t0MU4y55ovLuiTLo4HYSMhlqtK3RBAPwHm28WKzyu8
K7hfiO9E7CztTfBqKVvam8o5I+bR4VyFp7x8/3k0h1uMU51JBtBjhVJuEtyEigbk+kzj38pSEevv
fXQV/eBNLbJuW7CY50b7jGroBV6uvkkqtDULm1g9S1yXl4azFbkJBfp1799oVSLo6T9FJpCg8/zI
8yvnAwG7HITMXWd+vNpWxKHuyDh9zLCeGLOscnHkEGl4HNpnKKut45ZRK3QfeIwRABiwLJxuUaLq
4m7I4rHMNEpGs+a0JCD0DwpTI029BzkiQgjBgt93Nd4Fab6i/g21ZD1nx5XnT6n36pWa9UV8N4Xe
GwkFCfdunaIyk1CwPvodFgaA4D1OoyIuXa1IZeJYj5ucVq++zi3sNyTzjYSHprLuoz0bg2OS1YVz
lYKMV4cW+RFAWBBFOq9uSF+4rUCp9Agv0V65egcsUzvAEt7mwpi2sfuNMmqIjAlN9kwb1f71FtVM
jcxd2RnauOmscU3/+DxwbLj2/acPDysYJm1ONKmMUZPYTUyI7CzH7xihlSEVXt3SJ+Kzwzanxrap
0WA4+KPOpVCGhxJ5t6TPvDU6+L+o1TceXtZQ7pIie9nZtDFmv+Yr/qSjyd4GF2C6N/S7i2acf75H
5+QxPqID1x2YeqcA3yCGzckirYct2vqYM3cuTkcd7vnj1TvoGJiHH+ovjc0MufDNRKfUngnNZ3PV
9Ht3VfWl//2i7/wBSijYMYtqTEIb2p4DelRYx0gCo2Q2roHF9Kx6qCpRRk3Q+e3zaRW3ugNqYRYO
1fR8pO1mI616yaoNLSHqzSeTZORODVMUwDVYxiwmelMLDz5sJoejIUN8Wn4esep7wanYIgOZBrpN
rt7pt0Aul3ywW0dlw5vAFmuL5LasV0lXvVINtl7dRHoLoMnhmOBsofGy3XGkyCNU0CmK4vW6Sf2D
VdX8/XiZjjV3FlGjpGRZ1klIK6T/qbBVpIm8B5rE+3ntZcdRvrak9Q5azqLhvKCBJHEkZZSD5qFU
BrFujE+Rg0QzVuywH1jGmDKXdf+XGNAm1PO4abih4o26i9/lkUP1mLwN+SQGH7O64PTnOXz9c4P/
3VI/1roiPhb86KpgFWFS0+/zgA8SX/mNKpc0dzvyxywAbG4/BS1b4oPgcr0uCoHQuwwALKvP63/W
rtjgeMImdNNzHRXoCv2lpGC6RBRjjxVOnhFSf8u3DVPR/IPQyvhZb/hJKIEt3IriPW2ewCEtr6ms
hBvSestwHptgck+yhV9565ElA0/EohPf7CkBdGF89ASNMwmz0ZmL7lt/HrWhWW4wCxJNZKje4sHy
6G5E8vwUMZKkOkoKCDlBuy7aMTJgAKtFTZZaJYplmsTo1j0pRuGL9+pyVUtcql/yVAZUZMUexvqB
JDazzC3fD17tFOFC18ij3XU3TUo5T/oqyhVXCjNGI6zRG1yyVG4nmkn77/Lc0Xj+DJ7WPTM5OV7s
7Tnbsa1P1tzU6ZJQX6l46SYAE47TwNNYw05dSSq6ThHoSaEok7MfXZMaGQXQEw1IjXoIwhBCfB9R
8xDx/21Pa4t0cTOYWoDIyW9hLHSf8oQ7RSky3A0yp4IP2vdB+Jpc7bD4Qq+QSCa/4m5wrxztY2sH
dSH1T4w/+PvReZIB+X1MvlgedM4UgR+gJS8l5jujAmZIgvf5eYXCzxN3zQ4EpOi7u3bZ6fftcN7O
WCI0TUZlbQP+5z3lQsiynFyVuNaJyjafIUG7LQ3IascndctUkuqZ5Yjpl2J6PMFGSd9bkclECrBB
mmewlaRhoqDAoHLAHrjV6O2+lHu/T5WLg+FC/IkF6XqgTh7uORaFMpCGikxYm8bz9FqqAAhv2Hba
ePmFHTIXS1EU2pzlCmfVqiLhVml8uozFXXYh2qWfV+KWuqV0Uz0db1Y58aWMqWnEk7up2rp6OOnT
vplNCd/5X5dEpmzRtLQikYB7LmSVBbhkqdiF/Qch6OxahjQjqsb4Y7UojIgg53D7vNpIUEky6K7K
tdBo0YYMtHM0tqrenQke3dKpPQVPuJhIfNCRnA0ZfW/+5okK1UXIP4NNuFbQsHSx6dEZrV6sF+b9
7FGlcDSEHQtsBHc+f21yQgckBxXPSb3gjMKWoLSWCMCfPn382mFrjx2aLIU7TW4Z4rUvVoykkvG2
7a5Jk+lpOmMM6doc2QI/4GjgRcm5M3p9qlg2BwPNd9iVMhvVCMuQMFXYjccug9Lwuuwaw5FEWFn7
jhV9pLIGBWvLqyaFGxSF1MTcJd3uvCDLeWxIjGeQt80X0vJNBlSvrLUAhcNJoIT04Bj/QdFJL2hP
D8ZkKgVaSmPea7nEPzTyGyWv2tgSgpqBBGXxUkrf26qC1a+Qt99grfZcZazW46Rt6h41K/6zvETJ
HHS6wYeLSTPdeFswkyf3DDiC0s83SKp5elPC01mGCFpJD6srnzkARTQfgwM2teUK6ShMPUBSb9cv
iNd6zEH1uIcowyVnTOKi4LBjsEx11fVXI9t7mAoqf7zlZLZ2k5mD6u9wkqJHdiS0Xtf5j1d+jHD2
Eqa1QzSmIak8GpYnZfetEyKdrv1Z6b+9I+VXibK0Olg1bafDcNghBGPlQtKlFdR85XoIHIrRIeDz
pGRkc0Z1H/J/+Rts8zMJgARwUsNLiu7FpjmiZ56GWzwEljqWkbnc05YydMtaBhSnTnSxBmbfBtoV
NGH9rS1AtnEfC5yGHsWHxIQSRxAjsqLH7W3QT4Mk/DsKKA09nX1zxJmIBJOd96I98mYIkHwXAbrr
kNqFEgnvJyj0TpWDOX9KlUC4VcIGIzPsabaBqBijxbUd7okmRIcRF83Y+x/FuiesiN0AbHr+rf8S
bNYn/JmyHVWqHVEjudc4J3eRMkr810xc4tkmhSfat+UZwJWB2SX6QKjy4Nxj0xrlbBp5l8hU3i4c
lnruUZ9DgVySmePV23ZaYp601Xhroz4IhWNAujhtRE3w9yhRmh+y2xlx15tjjHzTeOVpw+Zz0LlO
ifl6zVUaz3AwwHn287D9H4sW2XJdmZoMjCaqYKmlzp6aFFGyW9rtuELt8Bt8PshI2dS5gvRCpnzY
SSdxB4BMvN0lWhtMxp/YSBEnkFX8sthCb3dN/P05XKHyhKJucfW1pwofkDgYdIcN/FqPegcgFf/U
uDWF9z8iYFndzjqjwGInnPXEnvIBV7TxME9hseiSgf2qPDPNBpEzVmoe+AHFjtvUYfZmSOyx7SGN
WippTR9npP+0/zQ/bK9gJ9wMbWyC7kY1QihqsTj5OfHzAye8hHPpDKf8/okJ1vPgtQjfEqfdL09U
B4Mqip0DwvFKaDIBXG+jCnDbf3PagMKAiH5xlzfeirYXGYQSdH6rvKcIky0G7xkC22oZo3kMLaan
6Grchg/vHm5KwHKr52ULJ1GyhmkO5emR18aA9OiQZc/hXFXQxjnlC0Xtm//F21mEwpcQbkkaFWkl
Q1EdTdhLBV2mNXlKtJw2D5i+7YGXH/OvCeJ1yc6CfxfBEjIwDdDaE0334QLDdbVaJguW1Vfvyi3/
FNzyK+LYxbHsecUROnzfJ/OkxaKfqt1wZP35QFtnNE+NDjrr41hAV2baIw8wGRntTYDqPzmP7Q68
1Wu9BbbUFkbLovS/6s1JJ9En5LHISpKeX6JwiJnFTyKgth2L0/xWTZJk20PPUwIKDxZZEDk1G6zc
kp7YA8e4bybPW+1/e2o4fXhAhVb7592ck3TcD2sFBZd/whbyLHDp4ydDTqXjqJjon5PyKQ98B3Bi
o9RtVUjNF0f6YAHTUl5Bvx4+nQhbTBL5V2BylciheIe3mr/vAdlnh13OZbB6JVjx2/StWAFgLoW1
/0BeLJ/Gj/dA6Q7/o+1EicN5XjQLbhTE6KvSHvl4yITj1CGRTcf344YKD2/7vGmjfVIa4D73hlus
YByw3gTJ+54hh9Uveg7mytDbW4jcNumRbyQ6TQor15Lqg+vunK6iZ7NW9PpMI+hVgaW7gQmbKh6E
LJdo9ss9njB4IxAi+gBzTxgdTI3HpkmgeABorNOENYkfcYQvEbHJWFXECsS3qBVJ3gH2ripImHYP
my48csFEhdcK5w5pzua16NhI9yLOYprhvmWw/U9sPw6DEn+GW5UGfAd6yp6jfc3/+01TtWtGkOTp
ZomBm3VCNu/xkBNSlGbPwj5mcKsqdyelYPtJdOnXLSAQC2KD/VE6lYnhH4kbGKPvnTStM/tlbc8L
E5SwCjX3sum+EShLtgIOgNjlB383KmI1osiKAgsv4ke0vx9uCPjRmehSsFu04wZyRspt90iE8HVS
06VYVn3STWPtZLbpM8e4U733qxVFwgUPq2Ruk8dDh32YDG0zAho+qhRZmszS+MT0z56/gX0eMROs
fJOjGybi3bg67F2/iPibjNNQ4efcHF5WAoOe2YU5vt9ovPo2sQSd9QbqJxzqmu37tjtHxr6NBmoZ
OVMCVlYOerMYViNpc0AA795eZptjkl8ZcB0UABDOhRLYNpgXOwnu4YYznu4AIBR5GpxgoHayQvLx
dFje3n4AjxPX/gvFvPdKGaLlM/CIIe8QlLmIJ9m8vmT7ghaKyCXegzdOjvUMdALMAubqgpIupImE
GLGOZ3R/D9ZNK3D+BN4igZWh19eCUrdOeg/mzX9Zg4cK6EP058/8dnpYNpIQ0JKfj5yE2/Rzs93G
+dAOCD0ZE0M4sguHt7K4ZSrf6YnHilRDN/QpXeZRL+Y/n4FeoqCx8HBLHLJJaK/mDQG1rZ+g9svP
rqYEZC2AOtsXrD80B1KEcayqOo0F1kCePtO1tVxfmMUmqUm6FdeSDRo9fIlHWczwO13GjC7wOjAY
6PvKIEvRjzoNp1YeEdG1cfb7B/Z4HBBHfRlYakfv+7MIgqwMwMjTthBh8R6EnRYYyaIbEvRhqvi4
QF/f+4sHGXhz2kP42jTHlO8E/Awt7BH1BWgBpL6QtIhXgkKGnxNI5dSjgAenpb4Cd+w/cbksK+J9
217dsVg7xVJ/2Ko1bywAoeBjeo9OYSrZE7mZv8FmiFx9AK6gB5CoVFo13nyhvWHvFnWrMduIoTDC
l7kxtf2W7o9r2OGsXVCpE76MxE/NYLQAbOH7eZx80vWYdgHwMcqDA1osgVRSJ+ILpZ4Yh5gzLSQR
NVOgtteAQHlrOqUwaeTKRCsm8alZw4/nekPbygAObDzQkHj7dT+vqa1tSQUqLvrxyY8+KJu940Nb
h3GeRIRbenTKBY2lRS4loXpfec+gNHgb8U+WYSXTET8Ih1nUci8tvGFtJVfnrLK/7aZLg/Hq/NMR
Wtr2prscnQGXBEywHAe33AEfMAW7V+Hw1ed7WAyzOJwQJYmoPsjPoSrUV7aWm+/HGoFxgq3eon9A
RAwgneZm23eVaU95UezraKmmxo6yeW+QhgMHkFWUWOhi6hWy3Sp2p0sMEbjXNcgq20pSY6YHyHPI
KIOQYAZhvG/vT+LxYZGWnflJpA8e1FXqdVUsoXhVcNgLBMi2sldOfuTqRwGBqlmyPEwDtAcLDpbW
j+N4IyAZjv6wtB+dglE/KDEKuhSz4NDjbOhAcowDT034MNB1p1EJwhF2SLPWZBPKSVf9GQOe3Sj9
YA5zjboWdS6cpsuuotHkQvQUORlNwxkFJsLW2y5NsMidzPcug22ABfytKYd1hR5dEQAqemJ1Pn1q
6qKJS9gE3QrhBGI9UT818EOEjBSnf7st4YArp1cF4hk5miHtdaheTM+0/YrQyMorAPyPe06BO3DX
BitkSEyTjqMb12tYyrnY8CVBzCG0aUZbujb7yi0pDWjYnJV/Fc5Zx6FmzmTDPPwYByUo3qNMI5v4
bDYDTi+wxyZ6eRIup63ef0vRERaf2hOT+It65JWbudIqFksn019KtiZH39Za+BD5jerOdqeY+QzL
wdjxmjgik4NYY1WQgNPDmT+hUOXwxTLLn7C1Zm4CySNYNoyFJzM079hyRr5ZYVWUPDsS+ZbTeXkT
C63VbpFnEFJfBxuyo3FExMVD1uKTJ2VlQR64VSQx4RME2v8a4SCKe34qXl9VZWZf0k+QA+BMLSAH
iBSIjaDtHYh+By9WRtkhrTRHn3kdrMyqssiJj7Oz1bavhkSZjHhkbDng6usYEMVf0PXhGnRKifE9
pkKEibm2AYKQGLhd8KZcbFb7tphhP3LKkLPM1PeQWWmdMAiCy6J62lGg9+S5Ksv88ZyrpVEbSCLj
pOCZGx1Px+XhBKiYOIvwOJVUenvcMP7nn9vNGEBzZ9G9yRnfc62IF2ArvRP8qEWRUWVDU/lwFqV8
6uYDkHsG3OyrOSFxKBkfqRmGa5OigJq4lLKXmgXDCgzKIZcTXhrzvissAFkzgnz9ykxRe4dZ2lDO
NVGxFk90mxC6MEs9POTCllRKD4LwDuh8l5vJ9eDZDefFBp61zLxLP9tvoxdt01SpK9vHfjRCN5pD
v3VupeUcF9bdZXPoP8GIBLxqXSk0pNNvXc3EdB2J9zbgzr03MkN2VNJHQGsXRTOFNHdGNo6swaDU
FdrzlFWDwC26h7FHHN/b/PtUUkkqaQnCw0OVLNqmMB56JESisgoLMdsZ8j9IQRqZlRjoN83OMMrs
H9/uM/8iTsV9FNwU5Ve9iAVGQFTbs+1XGksx9/xbOtBW1G1tiGYUrXAdMqrYU0OXu5ZrTd9Y8s3d
I/tv3F2FHk5YXF4ObRAUHxCuhfkSQOJtTMMuGFavF7qFTl2w0tc1R++6A+X2X7qzieOLUoSb5opd
EgHkMTXM0ZqZ7+xcc1758idI7ITFUTN8p1wl6UXqJLP4oW+kczImKqFucxRRRnycNmp0TxPymEqB
re48MZ/zAIRQ/gwfKcF1lwHCpGg6lXwAr2YrdCocpAyFPYm82IF5ZG9/nnQCNkcLOr4vLOSEMl9i
3L8ETvL/G05bp8ZpvRD8/wjEZiCU/Qw/XD0pZNck5+YXlA2uR+F64kx4eg5CCO7R5SSQHjUQoWyb
cWV7B2D0ejPSxi+v9CYuTn2s8lTm2YV7ONp6ppaXEfzVdeFFCuociwWuphySCpGwKDHfxm4I3vRR
HlUwtbmiKV7JuhSSdPm+dvBScLFPDBO9RZ4l4vf2el8VakvnjhasZ2ODsfG+tDqNGe3Q1/f26XLH
hSdl4hYoUxehELYzJdPIJwPLODKiqCalMNIFs4RzuWd7hFRSxBVaTcfitK0K5GsX4iUm+8qUa9g2
7VuG6sWXxTZ1WIM64PlG6VRDbJQl0PLdd5VJ+THcAinQhSPqm+FEPLJ076YD73INzcgVBni/GUZy
9Gr74qeCSUwc8Ekx2nzmwIpU+jqm/4BTEGkCsAU4dx+ckVrxNxi9RFImPk7wxD6ieOp273qqAIBa
1fzp53SiplLS0TSS0EvykjMkwEm1pNOPEze2f08PPCG1mnzycJakszoyfaE73Rr5uazrI51vL0uV
duReT54okLYXhN+j7/fxOF/DJX39UG6t2McWBERGQ/UZf7yPXIkeziF7wKCxTyuhlsv3F68uHLi6
k1NLDklnSS4zPpTDGxP0V/ALHmjZ9lyRcMfm2FSKEpbwSXj/GvmGgKVVCXnlP15jgOUtxA8ECM0y
9a9SQbWDx6Oh7f3H8AdZBB6fcS2t+QR+YkkIEZL3WASbLdH5oa543LveY7K9VbWl/XNC63mCsGGy
dEGctTw2+UigGW9YZ2Rxe8PFMAAaYTqNpIm+bXgbyIhytJMbSTlquNhDvaI/0NHwhgcVO3IHyX/Z
MfB0XChZYVOJWNDrh1TR4KhMX3ke6+Zh15NwUYuWrMiY/UcqidlqNBvXfmkFxb/0f53zYSDnp+mu
jsboZu6mCmID5IyMsUIakam3vOp+cQpRHLql8u6Gor60h+sGtZ/GHXo7tFRl+v1oGbAvsrd3Daq5
krut03yKg5wINzL4eidUpgsomjc/hA5Uzj4BQMHnw7weA8XDfpd/vbp5wSRnC5wyk5Vq8Z/XZmiw
SBN5gbbsqsW2nEnTnVbqmzhfFtSum2djcNIm+peuS+TGdcN/5oMlpsI4zwu68kZvQnkRT0Af0C5x
1V0e7O81BSMnnEVEGxkJjCwpZ2Vb+L1eXxTLlT99XtY2FHz/VRN84Mv3lOaTiCZrD3vmTU+XloxK
4bq/gm4sqpSX++1cfF3FcNJ+z3x5A8Cpp1rHnyXuG7x9xx2/oqIruOtLZUR0q/s5B9GGA2ZV1ImF
PwDI6wTpbxVKNKopuaA/UYwChHl5B8IN/YU5Li7yhhkUCocN32H8WacYlpwheUPGIfLmCso4G0zk
IJcuOr28nW6jiBX/lr3DAOhSNO74BnhXEYCdtkXtdLo+AXMEra1GOqBbAYCgTgxFVBSWYdImvdud
k08jfwZ3zJguf4l9A8bi63KLSH9N4QNYxBs9NVl//KMMZ0JMoE+foQZu2ukx/U6ZknO30bbAqocU
doC87xXMv1nH1wbPggYks3jCEx+fTj5baqOStwNVtdIHrGcDjGorm8blJUaYGUJN5FYlcHckDn/d
bWEf5i3jmtvIuYAV+sVoTfEbibKHoiUsaP9lrDsj20s77BD00yZDi40YtGyEm9XUqk8BVkAwu7Fe
SkVPlEIJ1lGmjgZ0gPxk3U6xrWem4Xntwd47OBmqpV2QhTQ0PME8+Tqu9rBxqIBJVDWdi/A8oY9k
WL+QbaPiPIsI9Hb7bqX8bJsbtYK2q4qP/6uB5tdOpEqiDOymE2u13fUloeblnOnL8f2WjenaoOTq
TStHEg7AW6PlhT3MX+GDB7bOuYgHY9xIYLJ3l+YPCmrQ0N9PFS6cs6nx0AcquWJrEn8yikHFklMF
Ga7QnVTyxNie4UIfgsgKX+bmSoeNT2jr5cLgewj6Wxkkuo7xtpe8QpEqZzTD2s2aAcGTx4U61VGq
4CPs1PTuGjGstx004jSFbi/xXGRYLY7TDp8qINb92lkRqeDrPpENUKLUQ2lxce7TVcE8btPHI8dv
lwPZASWbvvpl2rphDInSrQYZdiGqHoVWQPlWpBpwwgp0muVOjQ8vpmS1OocISDxEJEuPhqzEYD9w
l8HtlQLiBMBtU0DoY5pBt3AHbRHxasVoDv8pVW4O49tKriZmWYMc/B6gYmeqFLHO73yXrk2RzRIA
OlplfGrnK2McVfCArvyxpzFZ886TRqKlC+EHC+pd0s7PBbkIAaKzPCDeAm8ibDGDB5om3PHRkKxf
VNyIacSsTUOl2HgmMYDBXZRmy1nbbaRZ3rQbc4FQu9Ay2zU0HgVcm04Pbjg67eEk1t35dM1YS4Wz
HXKKt2JNprtXtIe9uuwcBpk/+TMpPyNUC9zAboX/KVSQ0EcW2SNLddnK3j0YBLdP9jag25gklxe8
FCAA0zxp6Sna89vAprwLo4sHg7/hleEO+KpsxRI92trRAJm2HcZjaA3AYbixzV/+tpVroDEZ5MEl
nJ9VGlrC3MHcVvK2ABUFjSsBABCmqRGRNpzqOUF3LkL+1dkZelhCCOYZwAFFR4rMBODS1vakrptg
dBVqkAoIzBspsoxkOkRC1t/EOqixR/7KShYGrEKDHe365dZ//bgQVdUwVsrT7bXHkzqjengYMCPo
Vu3Sgp5TZGHqnla4mYMSParKkw74TdbYKrtmYqXtf1ZtzIc1tSdw83RQlocq3ilU29297LI1wNpp
N0gViRHYPeeBpnLvFlVFvhW4wqpPknIs9rK41qmOo70+JipikXkYe2bo7KcBVYlkCKDLgfpAb8kR
4qucQLk2NADzuexn07GJP23czz5U3ODYpHukMrJT/zMDsA/aeUmt+J9XqIYHSvNz4JJOoqoaMBRN
m7/Y+bLlS7pJLxcuMBoljNrNAEv2rtK6mskxVZla+n6qiADCcKxsezhSnNbN5UJitqp7NmiD6uVl
ngZXunBir5yWWeaIKN68iWrVd/zqc1XnzXOatgWC75yP9MjP53bxIc4AeUZhyBjNG+J0zFxhVYaK
uga1ESKTAG+A+FtgdB93ZM7mUvlnIA25oEehtkuUQxA6p40YLE7Ex9N7N0u2BddN6IjudfbC3rG4
eg876snTvIWK3lbqTKTQkkQpN0bOpZfMJB/39afGuAfbv/EVl3YYxKsvBrWIXym2uEO/De0gB/+j
badZLzBXnZAMXSxIauFyiTm+MlC9Qy5yaK9qVmJDYrVnxRdU+EGrYx9tPr45PbTEI//n8RCiUovw
FbQYM+E+ol2vWP0rViOqQWGvpBsd7Tt8qkYW4iVYKJl4KfNeZesBvWVGPAcpSmHC0IqtUHzGYcRl
9iGcO61HEnnZwSjtzaVO3eWnZw8rEwcw2hEghEUAV4W/0bHHxhtk6547LIFIerl/tkjer1Qx5GzX
TsWp3KjihaytMfaqA8QYi+XG2mEsCDYHI0/uM5ieAv8v4TuA6qKj0/Ux16E2qTNjVTAHZdNz9IBS
eNFddeqB6Ms+z6fh/QK5AdkswzU8mUS1/18t5Xd/7FOKO5ma9lcskWcvtDavXtAhquxhfHY5S1xL
Uzs4JepPrzTcnFGLIFOvWRxn2YLjtsHgqGfKwM5hpdm3hsVSACdi6lBHkuf28ZDR51gBy2YrWkqf
HigSJXZtS5gQVAdJwCE/R6xTmN5EcZ60evClA/Mxzpu/dCOOaNu6T8o0S7+sQoZ26ZtQenS2qnxR
0PZzhEOmw4lERmgiWLrLNXULlRR9ZDbjtVCSITIpGGdQYiszQtZxAninx1ya8k7DOTyXNKYEmsQW
NL2w92lEzdRptbPpfgPOxkjimYZ0nhDDXfivP4zm/RCHcU6MI9hwoBry/DFcuArgkxwat95Zqxb8
+iDHyN+NQIT3b0NpjuMh4yjq3W0uIT1/GnN9wzMp279UG63Wg9fYTn+IibEpy3mOlB8u2a9K1bXq
eMaS0zreV50yQ4YV8jq9fzNiTVdJtUMRJXhic67Jk5DaNcsTx+YMspBopxYA1l/03zrPbRZkeRhl
k5nXLYK2S1o/t5NN1BfEB8NlJ+NlAF59RBnYJKXMV0EO8MFVKPT4dcPX6WFJZRwZQwrUhMtv/dIG
4oaIg6STcwi7lwNE3+fZVaLs+ovtv8gPAh/wQ343nRt41u6RcxuRWv8bXDSUORBJEXpFX85n8IXB
PMFH1NPT2GG71loHtdZqJU+nH1sELj+/hG90ThAViZJPuOIFIkDREBAHsCmpntFwHAbCBjCbJqbu
UATCl4lwMeuxTb/Vif3UevKbxunPrsLKPBJsQolgJiJYt/twHKCHs/Skw3JtvuaaNdFYAJVYS5gM
Ly9QPnw19wMjIxXjsVYrS8JN4ty2IX1iyrY1qgXy/Hl3AuirZoQVFHSIWle1PHjaYuVHSVob0fB5
j8nrznQlJSj+oWaM5XBK3C/8fcpviC7K96tQT5+U9UDa/FDGl682NfuXkrkjjy3xsSlDOpfOqLr1
Yq9KAZuSbSUAA2IvRFBB4aEDYQziNQn9WWtUcumHMs8wBaOkL/FvT5bSltn9eU0md/epvCUw7wbn
2psxzZ1Dod+aCAiWQS/OFNj74iKLwF9uZ0VXwdNSFjAHiJUc02Yclmd0FnNa1Rfxi4vRbY/FkvXA
9/AveXItX2t/Yadw0xqN8ngb1XTasdcGQWAl+c/ThSqNn1KEYF8IlpxUwlSoz5oTiJM2bHkw4fXY
Cs0WF8pJFnmuesPbvFFsUBDo2JByeBCFTSSFtu2fZF110Q8QmSl43Z/N59NPm8iU009NffNsF8Sq
CsKW1m3yJ3AW1Xetkwh4eItvfGMMAQd/YKZZ6W9qTBWHTYunQhDHp7wBBuhHkHcEkZT+q+FdTpfC
aV600aQqfei53e20XfWJVSCAytH9dbEl50nJuKM1fkbXCWD8suUC0JuTpYgqxpX5Puo9y0BQ/OsM
Hzgmk0BLrgratmwqzJPiJf5KbqukJnmj/7s9kWgTzY9RL6ONUcvZzSk70AvprQEreZvO7Tl0Iv2X
0vboNGKE/SuZCQtrY7N+HAHP6J5fIf33s0U7ijy7lzLbTuJ/LfbxSITG1XX1v54h3XhzbEvU0m/r
Xyc/Lmb3YirX43GWS4rdfSon8Vc5LZNTmKO/MpzHvgvfbxoBB3KaBplmAI6TGuABlDE+3NTQ/O97
w6G/Tn0exuCiu8cmXAnVmeGodAR3o6epB9G/CW5fra0z65+Q+A25XrnFNNluvoha+gn5BKH8JmaV
NMNb6RZbas4GuOINZVjPguJAa1IH3Gwd7iyHdRW4LZqPzPX0nCYnJk4mPaKA9XJeLkLbl19i5BzF
gQ8pXeNz1rh4RLBz9pOwoyPraYhWU9DyGPXRJgQi7fZ5/ofLErfT04LsK+o7NqyzuFJaDypbPQVi
yiKJh4CQqE1+wIej7aujfckaUNNvBygul1N2i+7L/SrZyEEzVJNzWUDG6Vw7k4/I6kg0ag2b0R9Q
qel1wfFI0YQbO0w9A+FTXnyLe2Zvu+rkmn84x8CakVMFQVTwClzCe4UeFiB7lhcAqfA7hbisVc/E
QvQDTjYpesPII1TwTtpL6SU6KzyffpKkE0yKy/UuSIdBXAzcylZJb4fO18LCSerb1E9CdYxulrph
VQdTMVEirr2jszwp0gIbQ9OHw8cjoo9kYT1yYorPttxdx7hzfLDduzLqqlrsRc+lH2ZSUrzCOiv3
l2lJtsmZhocjouojM7DKMw+TxoSLnlBQqyOh76FyZ5HP/AS1od345eBJzl/1Sgl9waeCkQ5BHMsd
QyCrE6rvmIR0+wxJ3bfY2h1aFrQFqflWhrFb+fT4HfIRbu3f154V00OLYb61cRfSdJ8rwDG5kNqT
IIJynTc8R1pgTeFXU0bsV0ATpQXaPxUo6lY7QvZwnIBTzxUhC5kYbaUKOFdk9zgNCrwdoezs4icZ
RJGCA//mKO4pNT06o1JR46sS/olpASKkxnjDLgOxZ7bWsay1PiV0R2qRe4jUX5ISSgpwf5RJozIg
7J/q3Wrs0xmRwOV4FCmZTYMqIH2E3qRdDk6MrclnxD6loZ/m+zSVICHgWVeHe2fegVxZQQZdEGIX
uBoVbKDjj9AxQvK97MX1W2hzn7TwULMaWlg62iT0RwhOL/gLZMBqppZ/IuJQObELRBoaZ52Z+Pv4
O2b+2W+cnkwJdmvXm54Fg4jXugC1VEETXpPeCQt+ZBzO3rno94pF2CNy/YAg0E4XCntIAbYhCHZC
kaovf7KB6nHF4XYJJmdKM0NhFu2M4D6P7ceGNywjMT4HdFURsqTY728i7molf8Uey22rE+kKVvpn
9fy0741kMdwu7sl0AlSrtvCdtZVeWw+9tImR5H12IcFz55rmhfISz5TwFuvMbbAzvelHVzRUsONt
Y9eCKqyrQGGzHSBKArgHK6ZtgdfpofxyELXSKOwCfkuNdBlNQzfm8X9HJyhhGRM0NKV4QCjxofwc
1KtIJuiuWxK9ORy9rLbZ6KHC/mp+7mUCqkzeCvoWxvp7L5IxgyQlD3tCZMpKHMja8ksiHuly6uh9
iawTC8pQzsPs958MUN13BYMhL7kcNILpya43ArX+GzdXZwRKhPai/PB6E2HuW4MBsx9e1lW1ubZQ
U2wIo53rr9onJ6TYW/IpDkwoqSlY+iltGtXKy4awenQvAT8uTeecfEUyAInzohXIzjnooLzirNR5
hh5pqKPMSneJYIc7+b0xcLMtyK+hDvqW/mip5ciDjRT9HZSEo2HkQesw/9n7yhsj2G5+yxtybVkR
TG+6GHN6dr50dyV92DfOK0aplURxNxUhtICuJR0nIn2+mDvHIHasG3YK7V3c29CJVUJLtHZpFf4I
A/p9Y0BB4oSZhh6kqTqLJrVVKJXfS9jtBogHo1w4FxaSJBSTz+ri246O8Elcbc/+0vak8EpdSxPn
BEFt09FdKfyjVSqjmw6gedvZVAa3MEXrB3yJSFwKm1a3K3skK+wydtAW1Tg19wCi/Ou2YF9YjVIi
JXlTnAiwil7McD7ppbmuhvwmVksFbUMkH5chcys2hl9ZlD/wEQ69pYbcsMPIMSJEn4ouYySqOoXq
UfB+y9TbEqFv0sBLDDo24UwhMMkFrHwYnyCqBXO3A6UxnR55Z+Djais0N42lW6+pApB2M+mQzUgY
1e+aSCxvBZUeX/HifJuNKMRl48NZN/xfJ+ZnzPrxgwzA93ZcTmCNDXQDTTd/l4PQGVCAa+p8NNt4
a58YhDp99dL/iURLxpQV29NIA4mDMUQ4aydcWfqkzi8eujK0ZDO/kyLCVN7NEkMEM2e6TKsDw47b
FUSfzFNQyAjPzc6cxeS1hyyof4WaUkquERUwjBjDSAh2yed9yQR+nv8aAubkpAraxaz7RcewfMg0
R7/kEmfpubMryc195dXwzBMT9+ENG9TOv+nXdfxXmLll+MSR1bXmjzgb6r8Rb+HcNyePjwPNob4P
AtPv7yfjzmqAd9kbp14P+vL+yd4XLeJlMQXwWRGVruCwSZkmZVK/6B1k7xR4iWoQTxTmgAtn5t+8
+6fBSQ4xftd5s3/wNyhJlyEUIQZ/Q9cgKdz+nrYhHs1Ii+OeDD+8lxOkHCA9HplDCpGeB2AEbQbw
EPwZPZ7WKXpd8QLjlahQXrAUdWs8rN6EZNVAuh87vEOipfAh8ACYJzRi3xkMALwhhvWpJ1a1EoV7
s6GN2BuMJb3r/5CASHdmHYTKDUSICWcB5rExqW3N6q0hkiTM/1wgMa0B5JnecGFihSjSBnrRdYub
pJtUmvk2tBcrNjt2PQ+Hz+momf1ZSG+kPrylaDJYI2iMxjujL1/zYQcC79fYmW9xPWxI7kEiR7UO
Pubc9Vu8+0IEJAyo4N/pyrKnoIGKNm6pYzaF2k2WvKUGefdY0nM4JdsL+i208Q6f/45U2yEnh0DT
xQBQadfrO0oKLVy4EwL/bfDNNpXi8q0alK+i+2/c8kVeEJ+mWTArmolZngMG2reG+t13C1Lb3mnd
8C6pR0i4r3eH4ILjdxlHktk7VMbL+WcvCjLU9PNbGH4OARGHWfwoLkJOj2xhIBRAu/JgYtf6+prL
sEYtLhE+buGWCSG5tPaEPBLn+vPymlb6QOUVo/N3w7qUky8sUfw1gVyKnZXSdnKcsUvg4ThrnCOV
kQz9fYkW/rP5mWF9bHWezpznj4pR2GWrfBkCvaBAlosfNFWXVnZQ3mw/VrpWeQrarwkLlN3cT79N
Aji7HKC2JsBszekr7yDzf1ObIkCU8BVPJDlKXhPQDONH+stmotSZWYd9ekPkr2dzY/RXDBkHm/Xn
P8Etra3Y5uYAd3IwQe4igqWzuKRqknKLMgjIUxPfNzSFC+DdqfVgEPl+4PGibg/877GUXRsv4neP
B7/ReS3TKnxUcCPQMxvdc3Q2d4ZX7BULQLOmEGuQHy4JpkKmqnX7zy34p/XElLK9BeSM0DZBMcAL
63erM9J9cxBFg6GRICcQFdh21eFIb9jOoHOxnsmkU5RzRVhDkVmqsTY/gGz9+wlWBHIr3o2YNjLo
gpY1qKbj4WUp9cyvGBMKJSEph4pppvSZ5jDwKDDtoonqL7Eb4tIZS+l8JwrEw8UzfJhE19DL51cW
JO9hZ8j2s02LJ5yxFW3KvmYSxXyBq477ywXEMGQjn17tjoX0n/o+XlSWi3DWNMUXorM5G/NeJ3s3
gfmWkwLC5nAy2FP63lWXGxq4C0rV8bZkz5YIemyjsNbuWCqJwHF4RPzsgA2k6u4YVNh9BC+pXQ7C
MgnJQkJwVOWz7raYXSGqX9u4k7/Dy4aT+G1lEut+XYJSnPruf8KkrxFBtuT/x4RbFfVy2YrKQfW6
BaxAzTRDm5Vcntfj0E8fUiaCwi/dRniCtv2gA8b2JWoqZatkThdisEN3X9wqdNQQ/k7P5YI5Oih5
JHYhUUA+irpriBsmkEJx+84bimhPWSzzreITvD4dk4J7GZJZOxWMH0d21dslTfhWmbcOmC/WlCXg
Zjuy1LaX1DzervyrOsAwoX1a/7wstr+M+sM7WyALxATt/yEZ3Py/n4h6Pp3qVi6LUq4HcBhDxeZs
pZxvbDTeUS+5pCcLVD3OKv7jxXsdvFE0y2uBn/+zQkxnh0iBW75qJS4zpgtf+BleUAuhWTIu3SYx
rIo8hAfWlIRTPnJoqHFW8P24Ou0909V5E0PG/hUqDBQpM9KXcbWJs7TSPKsxYH2a1q5J/Vk3+kFZ
TzO/8mwsjMrmQzMwV2FxV3j3xsdSC+bLG2TUbxh+zROAqjSPyxD+bV3sJXxHaoEHpc/yu0XAA0Wm
nv6ZI+04u9/7NpBPUJxyvQBOX4SJ+SJkHoMJjvT7OhjSyPpEunDi953z1OwejlloHO66eUNM7Gz4
p2eXiYB8E5V16/x1vHfLN8l8rcY+4fLR/HhJsbHZGC0kyw44n2bw6grIVPIkVE4mmpniS5mQC8f9
DysFXi0EPpi5vm/2I+ByoqVPo0sk/8tc/59O/yv+ouXmG+i7NWC7ZFjyget9EFu/DYIPD+kBE51N
xVI7AG4abGrR1bIcpipk9MNBKABrKEipjJZQQvwOEXftRbHyM3om9lyD4+pauLUvBg6bQ5v9FXT5
0ExvayYuGmxahKbEv3U8UDAhRQ8nIdCN4Ns5dGUlK2aNG0mwk5U+A7M5ShIgS5WBsmph8ZklXWw4
EziarSpqgxSWE8myWiFQj7WSIU5yMBktVC8Uo9cXpZk/rREpO/OZez0xLxDHMrNzDMMM0gwRKfsz
9AKDXsGAyyLWyvmOUetoMj7Oi1andzloWvEJalIv7P5/kJOsjevXo0lV7Gd13cActNFiGgPWDS4c
fbyDWw3DguCL3HHk+P9/3fl5uSoZ6Eo1a0/7Kndso3Paj9fJrULBwb15n5eLGdWCYgCP35qMdIxo
xxnr16qHuhMaTPdDezwy3ytbUbQ8LWwfdI5Z4l5MZdXFrjZChNN/ezMYCS77eSsz8/SCOs5xTmWI
InaLXdo6Kv6mdh5wC2WomMrp9U3UADZgsZ4lddVmPbVwCr6HJmk4kMf1P3/bNKZnIJtKkK1NH9qs
C9B06Kni52VQAeV1eWV1aN0yeMOpP+s9appPI3sqOcuSdLINaR15drFugGEzzu+ZHcdu7BWddK7o
V6nMWpbr9G3R0fXjryw2ir6SFvsfQKfiK2fbxU4FcRLHEXXQ00jdnMHUOWtKupf5Z0OFW3R004sa
bimUtWCJv9ANEW8a9TtueFq2vGpjNboQfZzb7lCgoXwzrIl2GJ/UI4VkqlHORYf+5bDCE1b+2MM1
UMF5JhmbXq2ti3czTzgA2yeE2V2LKvm75s1g7XO1QTuGIoCRrGB/z4B6tkq9QlInL2+5BQoO8qYf
op780J1mtb1gIrO4RJQ/T3I8ztBKrd/KZNYLv1GU+CE6taZbPCC4mRbkvlTpzHI0Sia3QCWQbjB6
Zu+/6l56FICdXrlnlDBp8jQYuNlVni+3WXLWQVu9IaZY36+fBjJO26cKFJPPR6LbTVE5yyX6GehW
9EKccSvyIlcthAmuxQTaBRzsrPZ8wJq3Gi8vXGdPV1zAKYFtlX/VVRJgR9L/Htn66xD1TfNNa+Lj
mXGA+BILTYQY50Rt1b7V5JX3ePLVJxNqakACJrGbYtjo7LtpAY3uWBSZ4FhA7xZn5WmWU7/cMhaW
UHNX9rO7Q1j46vB7LTqH61ZqwGEmL5TccOGqOdqyPnDR6PaDOe7vVoHxPRSddmbfsgIr+NFD6jPS
3ABz/S9zDNAxaBxsyvCSlSWkuiAzkSTWRfXpGueH314VMkyKzcQGKE42IRW5Ldsm30fYbINfGEb8
rGKynxzC4mPwmcqlodqJWNCcmUOjLkHmE7FwiDOOVr/Pex8/4lO8rS+KcDUiO0IN8f14HWra04fR
hchuJsWqLGP0nLCs7Mq6UXyvoiSUpxalbxdE+kY2tRRKi+avdZQjqEzTCq+jdziY/Z7wUbmPOyJh
9LWY/lVJK5wLkVqAwhdbbwkSU0xDHOhz3fW0F4lGlITXGQ5jUNFnPjMYbGYIiOFqCBczQeOoUmbG
P5YgaTFxYOO5VvPuAmgVaEr0W99dD3gfXpRQXW2kMIY1nna6EXatxFZiLJF5680gj1tDPzIU+t7O
2jhVmHThEHjeujz6WKT5IIHEK+k7xDlETT/iXb8HrEgaUGoEPn8Xp0va4XyR7sOBZmxmTp8ls00R
XvnK3Apzbts4eGqZ81QG1G9jfI0w1NBetuk+zN/sINzNeUJrmqDas3w6YEWNQiNC/jAhzMRwljTm
3ZDBi8D9Ywokyhkx/+d+YfIGIRzYkoPc9sAnnUSlvGDIWvyD4VchsXX5rKpHW08r+zl1P4RzElKf
O0fL0DDDLLXoXeGBY35aRxpULRSd28TyNcxHmWsaRYw0XBM+NSI81dR/y4q9AbCIhXqGeT2kBEUo
pAWRgvJxDwZkTY4XNZlD7pF2NtboKX89Uyn9PrU6H1FNgcyq0l3G95Y1C+QcAYxVobmvYgwbFSrX
jo89wDrWrA8MFSdtTkBFGrrYj4P1vTKDf6MAYe0p3j1MOM7mMQpYSVsblbQ8lOOUqL9vqxbG1yIo
ENM5tg47VJWT/ZBx5ttW+XX1qKwTW8kcTSzWq6amrifI7x/ERxb5LbZGkTqX8UqEl9aO5lDhMIxD
kZk7XBnLOraoUH8+Y/CqGOz5uQF8GU4HqQhxLb4WP4v+SXBQZLBZD4923HLyySuQ//tt/GxGNng7
1xzjMv5VRdZite+Z0mP50ROL67j7epT1WhVaVgDryqPHT7J/VLQlnZSTAZCjDXg4Cwfzs58yPHzE
qNvv/Uh7ogeE/9sIJnHJ1tBeS3Gfdi+Izgj0yGi9cmrgtsZYfmXNZ3Q/w+hlClIFSoEoQOCRHNLE
Ejigqs+Rr+mbNm/P6wjLN2HVhYz7PmIIM3W2FEBAeGvbIZ8vEWItx9JHqsSSwe83tHc7izvalefE
t+U8s44y6INm17sYK4e1ZEju21zuqAUp/FwVI4RNr+t2n5Zwu73RT3GqLx8VgKzg58Q+QrG7Mirz
La+jWCA2XpnRjLGendkt1BKjuR5hIyfLMTqSi/7KanDFkNabx0Y3q6P0snoNxya38iNUjB0gFvZt
DBoaUcz1HAFAmS0ojOZYFlW/ffIO7u6dJsrgy2hGP3PqnYAJ9he8WzomYZXiHHfM3HHJB0U+Icq9
qXMCC5ckVFevHrUvKoeLHBweFAe5p+P+X2UiCn0bK8XvHKP1/7kw71mdS4AxSgR//O3wT/x/ib4r
HxvIUoGmduWUddYyOBOYX2D2Or51TNpbFQNbmBfFsRHQnPxj+aPIRxzbcsywQsAQnae5RJxM3b3I
70ikD40gOhBOkZf5zOy1jN3BT4F2NCI/+EMobPFgySUfetcxYqvAGnHvCRGYTryXyRwSrdh/cdZt
VsoDC8dPP1ILyjAn6eQZ/qmaoxBwTuqUh4b+7ZyNToiUMt9vviNa6iz7x6SaXUQcD7FuoBrR6ZP7
t95UQ1NdePnWKgH3jD18dVxLd16MsPpHJ//Y76jHR6CwUUvNZ9sTvZYaC35B785xR1w66L2h1sHK
otZjBJd4Py7dGjGxo0yMLR246DCFAKWE+8hGYc0/tBiEvznRI8G3QotfZYTUADmmE+I1owADGKsf
Izfy12rr7Ybqv/QXw/1uOiLhzdTmvvZfVuVDeT/VyTQgYP0M+3l0amRQMQdPfyUxOL75fBnWlrwN
RHtUF7KtnTKLyqX+7anQBQq4s3pZ663DAwHCjkWKE6eqSEAcT850WlHlA0TXu9HVqgEADRI+pFHV
pwGhDWV0sdA9829Irm09Q40SSCzFLpIcglMorBWSayZ3fg9hxvmnK6mIJ9KzU71vgBCiUlGEUgYn
zIefhwp67IctatMr53mrJs1C2iTu1NZIgvHZl8GdCpjDM4JPYzrKW5kc7PgPpKcgdeIAkcraqDZj
/bYcMbkRX4FWpSvmkyH3Oav1c8UKekApfXifXEWvXeVcvZd2R9yoxVpkVeQqtUzDPB7lnPpLpt3D
onVV3oOJ5OfLzLFizivEJoaTkmEpl4ht4ovTss8qTsVsPr7r/XbXe2Z7TlHpg7goHiz2gscWV7tJ
M2i+qeVCcOJzAl6MmUld0l8d6X7MOxOTzCDfNjFRTsX9YXzZ7yAZ2X1I+3s7mHyaQQuStgQQGG2G
nc3HlqSes+gvMfXWcnNLWDVTJ/TU7LwjJVuPx7HeIrIsYw4XRQd2U9Hl5ehip9HPkTxpqrzETznx
X3x9RDCn6d8SrGVlfn17HckpoNt+eqqnp5u1RFUQdksTYHqX7TBAqYruYdBzzUJoEv1mfSw7H+oc
x4aAZ9qwfq4Dmcdd2gBfnXNQ/HCsknbrE0uR1UlXgHfImKIm9gzV3fAs7iJq2IhAiVCh1u7BpXdC
/yKA6EMEvJroCkxBz7lVQ9bCmwXaQl9INQ1+kTlS1BNcaG/SEiNArlbS6IkYGyLur76wPWngRvtH
gjigJwOeTEnR5Zx462wuN9sZKIlSPiBw
`protect end_protected
