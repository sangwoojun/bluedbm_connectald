`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GfzB8LbLxggDM1KcEbl7vRrDiDva1Sg97WeOA5CkTU5Qw5tGcI+II+nqoBhu9mSnrTpEUnWRzFMI
6vObwg5U4w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZCu27aG9ipq9LPhY11MRetuaQ4uGCy8/ecc0OcrCHbViG5MJA4ugTmofaKcA+r2TTiCO8T76Ehz/
lSaoYpcpUaRkSW1mJUYEmwX0TW6h/LWfQptuEIFHiHhYQHyCvhZWRyRSHDCAFkeOQJnJOJ0BSyT1
X1/LGs5avnQqLY/XHCU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TS4w4W4Cuby03MYt/VDCY0iRrAyFPyxsK6fhvpJbmryQtwnltHOdvzz5/sITZTpVjyGtemU9KbR7
jK/zPPt+69Z91zLpNt6kXt90GPI+H3aTvLuHgGHejP1d8Cijbr25/LnKYpxy2QRqiDUQ85ls3pZn
5DjvrO5fFjYF2Ep31HHC1NG4N3exK4G/65nZfWuu//h2I4hxhFxGl39uQx7yEeHK6E1ybsKcLHvZ
yAp5zopThhqcoSFOSNd57G5VcACTwS26pI5C57ALmf1dssWtuHXWJqSpLA6l1GfqPIQYm52ZcBbL
1dqkWvprWFfZh6sSVofhdO/4rof2zJIIDD1zSA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L5f7GI1bYWVs4/pvLry6V0VdNH9EsOQWGKuB0CxSNzb9nNuk4asbgIDF8vbKn2X6tE5zdiq427f0
Gqi6upAuqRIFUhKKLMdXS/56J2gK6nUr43JZvHwHIfEAgC0EIMO2RRWuRO9U4eVQpVJHv/oWf87J
qjd/E40A2ZMBGyLaoOA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mdwdykzT2/il3gdk6FgMbU6vItbg3qa4j7am82d1vWAsQ9Ft49BASohcuC9U5bDu8nUkBdia2u9+
+s29Z8kcJJmcX7UTNTBNxReJJOfGFJcL81RS2CKW1Jv4PU5wdfO53i4k0Mj73ooucUu6Q+gw7+bw
MNfzqEGjlQ9nfQCfSIBkAGqmBjBTBfcNdziEFLTg/JjcolbiXit3iuSjYTCtDuLi4wxGtYWH6y4G
ZxHACSI8TcBOeBaMIUfo2Yhf+g/aqNaOTInGBanfAUjbKsViU9DOueIm8NeuCT5pBqb87G9kc5vQ
Idy7pQVoS15Zjc1NIAB0h6tHqT3yr/V4YYeWTA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47328)
`protect data_block
M7L2/MCGtAF0rSh7hEPUE2WC/fVAwUzHufHosvMTFic0Y2pSG8k+Bqz2siUZposigS7/FjEifYcp
g/H63DsjxMWIV92nFh8/Peh6R6KCJIhBZqw+zcfF/t6J3FlTGkK1oMzITOvgt/2MfenUvKs7F5zK
oeX2O7kZcFVVlOXRRxprh10/aZma8692fQI0XPz0NLOIZe55fJu/48S6ncEKb/bkToSVyFn9ULUv
E5CTf/pO5rWUW6Om57Tj0EgG0lWu7aoDxIdCTzsZps+79BqXKKErzWAd+rSHEgcQAMwugEiHjp1n
6Iv06yECPsZtuZRSx13vZYl5raFuWbIgYQ7dbRGCsbxEU5jhBIxaAIT3r6gkgfuqx9BbyTLNrZqE
LJ4rUZc6qjQ7lyRRh3W2ZKJmDKXKFQONn0HzOz09l50Zflj9d61UM9dH2ttINEEuDT6RIrcXdeQA
ZSuNxEN2Rprn06h7xC07ZjsiNb6rgU/acpYd7jGuC+rugy3ENmPJe/4tGWQwb7eS4sfL2JPXv3Js
umowUdEfBL+NzBwpYjmjIXwYi+BwdHnfRPaqYlTnlBenruJPkzRZNdvWfjDamOEo15HP+PNKdcdJ
X3Q/6jZYeEe80OlS889pEYyaV4v5E2vH2By0JkWgWmoAb4N0J5Uo8brPQOakyODL2cYYFuviK42m
nSlfjrcDrDX27ZSfBZO2uvGQcHCXs0lBxGXybUu3I1wPerlH4Y4muRR9W3koKEZQ4pILYMj7HC1O
PNhAxV7eY/W0muzvUBZ43SwtVKGojjI1lQu30s7SV35kLDaSjpJgn3CgrsvQK0IxJc4WIA+Idtfc
9k41EVtdS/RXcOmTzIxRCQ1o/GkCYpqI+1Dz+udHAfnvv1InkKyaJjEXw0ZPm+0DqFE9KtzFkElk
1OB983nXpeQ+SAURpZqVU7g+rZLM7BU1qc13J0/ADybSNTMXOirqUJ3Ptxg4NfCYWkQmTxWq4Dny
cqf72tyjI9upHHTYQiEqXEBCrSpZ7+I19nBdvzOmXPEBm484o8vL5DoAi/WSJ9nNN6QvB8O0r+Up
nxvpJjc6XiUh1NHJTHWS+lHkXaNzsNITzUc6Zmb58bxYOqa6hUYzuRq2Asgy4Bde9hECJvd7gWIN
ma4wE7KbKNS/+OTa9TmylWjz0PtF76marb0GCMzVu9l69aQST8JXTMrMVJwScByeA+R8zdPFj36O
UfMSXbaobfP2l/J6t++qRRbZFLcu79EOAKOz+dhGnfPnjz/0ERbABPfbOgHAfaqVP+ZYHprFyalg
xp18DtKkmImE+uNgCalENNj9WE1v/I8oHfpQDDCCzoidaVh7/+KRGDRwSONeTIcv2R6015rdvlwf
kCuOekbpnus2E6ut27K8egsqkSYgBUCWa6VYHAspy8NspI1RD1bIHPph7qdcOIlAD9ZUWyaAq85x
6WLmugWUnQtFvSnRgnRPsioPvZZPJWVYSkGAGkr0ro+Lr2fbT7+LC4JUQ+MPWiprPg4MT316a9MZ
rknm68p/eEj0+ST4U7dkGmS7P6YDYYLeBR97VpfnXmuMFV5C1tMO5AUcxPW+CCS7wJRP32AyQS4v
FtAFSh4+8Lsx7g89okLGExRVL+CDQ2auAJnspB2B4LNn85XRtDGYMsv9LJZUJ/G1AK5BvZ2d98K4
r9ir/yxZZmLsWTVnNb0BMUInuvHSG5fRLGM/byrVpxlHCe6yr/4ovxxcv2FWf9cKXklC6Kb6OsfR
EqCrnmjTMkHP4dOyir71ScrnojVQlboBnzjbCDNbv8jJUT/dSROFPKyc16UFQ0R+GRER3iUTPGAh
w0/vSAreupxIPKD2fGcoBh8jkqXxF46KgqQbikWIezdJSzfET+bheiA1z2vNVOdXzJ8V2OUJYt5y
zcpOlG3997h2e/kROVPtmO+Dqr5aBQSwEHmFq5owXmGF4k40ml9wrRuqDLarEzoBrNeHMFYXRQNJ
FZazeyWlNLGDU9kZLhVQOvMNZbXFCxbKumZwY5ZHx8Y8OrrUohFbJNlNGmJF4/+iEr3nTMa+sYim
GpIVHRjF35qGGHQWEM4vipa55Mtoi5ssidICPxH6wtW+S7+psBHsOM9blcvm0vW8rU4V/d7WJpUs
SvxjTU9v/VPAzFVOvp+gakO603M8nvp1Nx83Pg5JvbWSDgI6EqYzZsFF0ccy+UG9lrbQglA4kTEu
uA1zI+UirdXD5uD0rmbGXSxoEg5QKxdLjknajtGEn4AtBdXd5oTpiJNxZWiHrfbewXH7T1W0DZyA
7NvGvS8fBj9lL8cRu+hP2CRYVX3wf2sovu8nFukjIFOQpMPMl+kHF3ZE8sjip2z49jtdJvC2F5sp
RwMRepyPyuOGR6HcZVZnOwKVF1oxHeUg1v1i3c9YutG+b4KKNbw0F3eJitNl6erCHjn/Uw13L0uS
uGzToTMuEcDXg9j4daHyUZiCEBDaVFyPJdYMB+C5yoGa4VEIEDJ13aqYPEgm88aFA8FbyGK91+/r
2dajxXmtKHirJerd5ikVUBDNaqhYHIix87REzv5S91ichmjTWNoOMeH79fdyyyfRCQeERYM1Unj+
2btMxNLgSvBshQxuPnYjSjd9UE0YPKYriS3XFa2/2qw1hcAViHEFjnrg4P6bhrU6qm8qdpxQe1Nz
5O7+OsKazvWEP46b13STNfO9kKMdIN//Pu67IsoJRVuJSOsImF+Pvv/KPcHs4AxoCjTK0srijpjt
QHF1yrznTV78nWmu3scz//VI/1brbDWxrSR4OFmO0irjxasgariehzhyI7VTviLM8wHE+1C7QpwL
+qvOtxByNDS9KUFpdANrFlbqPWcW1ga22qEh/aDBoBeO/w3KZtTCmKVuBw+fvEWG40xwRnPO+nwO
vmbsKDEjDxi6VP952ugHexz6Ri5xKdHx7HF71Ti80d/kj3UcqhdLs5tORWLUVRHxR/4loqSRD9+5
Z5vY/QIVkJhSFEXsdzIMVMjK004D3w5N45679TtZn3UWMG0LBjM6UIHiaiIl+gXq+BRMMN0K1hqe
vwc1XwTyGD7+Qo6NgrFCbFzJm4T2cfTPwehORwNfO0BCTjMxdUiHhdaTqQnrfypLU0TtWEak0qzQ
iAPZzAkM13IDeD6ybz/jjbBfvHF0Tgvp+T7yHBX9FmXsmgLJ3maYDQmev2fGngSUhqiiQtcz3N+T
UlkINJTQggw6+eFdlpNV3O3fMRqt3X5tFre1Kl0mUT53RZ5SspHeXZxCXWfqE6jWADXp11qYfuwA
XE7EYdIzmLNcDt23BA9/FjQghLzxECncyb5P1AolIsdcIFn6dnFcibiES6QvwP16Jh+E8EyGbrqR
ftBeveTeHYZwZj7lOdZ8/gj7VXDAnCfYqIA76yjH0UQY1eA9XUC9LOdNqNUKvhz2Ic9tdf0JImVv
KIbggERb1KjKG+PIW5oV6psHyUY5W9HAIEQFpu5DedKQe2lnJHfuFvWYr6Ds38LQ9Aksse9cHiHi
6QTjPVTyQkqs/35d+6H14rcdd4C2uh3oBGVMp4srWwJlGQ2QWwEYClYerx5CmLCRTTOgIl2Ng5y+
+gUOGyI3ZWbr4LKrtuYID7Er97gUsOlTJV3Ft/fCTJJzhUqE8laaDf5coEkQNVQjZZb9RVFgbUlT
FPyhRqv7k1QJEjMvIHZFYymh1BE/c58eS54rhlXGMQzsyI0bIHRvdZPWQO+NPNqMLUtTzXu4q1Jb
pr7EqDUv4JKHcaWLf48CE8IDWB6SiTk8ka8oB+vNcY6r006+Z2H+LU1cYmDxVv+NScGF+DVAVKzm
wRlhQW2z8tkwNI+YIIjFm721FUGRNZ6Q8ZEXkLMrQlvGk4JDF/XXhwHuUMVAnxwh0Q0caxHa4JN8
UUg6KRqzzLe1RTcoC2y9EZkbOPPXGHV6V/gPWEbhYx+87OqD9NcLq6NHk07SEb0IV+BnzucoblLl
k1+Mhroi5RPyW6J6tCFPrEwFnnUzqF5NajdcaFBzoYVBhWTENxMmsmW5oLGL+QyV9hxO0ruFT8r8
z/zUdLnhBbrCdkPi97Aeoabr8ykOjj85Ko2izIGoSLE8pFwzEEj6+SweViCqOH4iUODRYSS3A+fC
9thwolb3S99sGT/AfzFOWZU+qVWIgIwgGEFaKouoGYCPotofvkLj3/fhX6XIaD+FueRcqgGS5V1d
Jboa73Ep/w0RRmcjmOjBMPLZ7IpePSwPw/8UIbBRkqegfXiXbcHW3Z7DeaiD0oQN6H0eDYjFtKtM
pFAveqHmoeeSzeKVPzldB1qJkNa2lXZfIZ3lK9Xka+8SMAkGDlkwXMt/Zj0AxaMmyzdhpXGDa2v5
XJqoyk+/H1Q6IxCHPRvR10C0x1vJGdGIWDmCPFsKz9+iZy0J+i0+noR2iTb4ZR4g9FpefGTxBZ7d
9elOSHTmSrOmazOwE2gKWsooD9kOQD4YEc+YMN503ibOSctMVrdFgS3f53tcDE0DxFTgi6mmVObZ
vuXLP1iYjJ1L8xl1Tc6KwSSFmCI/S30opn1tQqEHoa0CGQ2o7+swoDhUUEWnKBrumhGhFWsfq3eI
U2tItIe3KL3UMf15vJMcyXeba56K54V/G5nwmwYu8s9nyU8toia9PrZNMICyb8V1V8zqRBVbbGns
eyYj5iQ6i8atWIwCsrF8CfYqHl2ePhUbOv5MkO4rrech7oLJuXGcnUpHw5DPkoIZOncpUw0UKCce
+TwPmPTg5Udb/KRCpwWwkt9tLOSvsGMr/Z2TpmNPgVv69Ss4D4T1944nDlelWEBHMil7IP+Lyx3Z
2gOLCW0RCHoTQ2pIP3ZVVPGoTAl1wA5DMvGIpswjCOb9/80PpQ9uoJBVuMLSCTE9WfGyZ4vY1sVx
qxfN6UB99xJmAMcPZ/+xCXhU3LKTr4b6hqOKGsZUkvSa6qRKzKjMxGJpSuz6OsBChuij6S1p+GR/
oKoofVhXJUlzsDhrChKRNSvIl2w0mqWAGTwuqZNhN7IjwS0lJcm+r6vzaiyl5C0Wfe5cFdsrpj2H
iK0KoMEhAmJGp+muxSGpyVJhtydQfq2gkthCavJSY8jWUvHO0qszNLPWjJ4mYVofoFngNz8Pfz0p
OFermDrSPHmqmcbMZBdmwkCLjSn18eIe/6326sav3yr6BbNTXJQbYfeGnmdaTGaWWszM+MvTHHdK
bWlnvJEfafiqEWZG+N0C/JUZJoA2tLKOp+Ui9AZ/pxyf3TpQekpp6WjJ9ZHTaN+g245Fd+9+WV9c
fGod3H3C6Ps8/v8qo3xojDMr3tdYIqKXVTbF22RLgAFQJ5gvAnSLGao/4PbsUEl2vWgrClKRjUu1
ELbuj6rDyPOa4inQ1CuFFJ+CLf8dA6AKd2BZFrybaMhKa/VKT1xALoy6akILq5eYI11cgXdUkk6D
j1VAVdEeuvjmO5i1XOHKJNSJP/qfURQO+/3OxisHgPeuS1I0sJ9hX9gbpwX6zJWCShoptYk0FvkN
ms560GPLXpbpMjQ0/YvnnvB8MpIWP9hqBGpn0OpBtdlhm2UR2bf3sFS7lM5sopAd5Rox+ern5+pG
jEVSsoTK9bR/AL9Hg3RHyxqFAta2TULf1u6Fqp/6K2fLw3KEmr4uBIU5sZvwR0RKNrQpg6wczC+k
3Rw+8JKblL0pTULpceFqPzn8TA+LlZaZOZ+wz+VvKeCsyxRWjw/yMCWrwHy2wC5GKn6GJtl92pVy
rEoerZjJc3wrmfaCZjsni9ars27vGz+pVtaiR+HPZkL1MV6TSBgphnhJDM7meZ3hFUh7fQ/QimPc
XWDgmFBn/uDSaXlUQM171L4Zw9CSO1WeEVWcqiVJdhPnru41hbFcfW+/2oSaUskSQgZhAQA0wkUf
yCdgquIP1Pd5xN5BOQUxyJFEKNfdKbF2NWcq72lMG46/+4Y5OrtMdkmuwkm5XkNgolc1dQGQkSpq
pwKSHCtl+sAvCNMWRHoOOVFWqvsFNuCUpxfL5Bdxu/IR02MCGF8I07L1osXzQumgMpjEim8HLa1q
YWTU/ar8bQq0giva5cwH3fDHYzzVtfT3lIR2uy3nqTH1wMNhVcPlO1TfLDZqJF/4QJV5BFEFiMc0
OkJQK8XdVpGsncHbDZl/3QkWV1B5pUnc2ZiHGU3ZDkUL8DlglxxJBBzsfitOppzro8YG5AZpnTNz
6SWfOo3pNsURvrS0eAww2SPLxh66ASs/82NobZbZKBj2a+pUTGj8BSqgBdUpy+zyVr6cEYP7JGuE
P7UdXKUobtPauqZFZ9n8wvSJ/MjT/LqukBEl2qfIVEdD8gFPUd/LnVS8v9oItQB657fbpzxEBGHd
G5MO597zehhlzbojNMW1T3QMYU8nMI7CIQQvxX6sLli5Is4QinDJMncVcwPu5kbA8JmmEoJQAJIu
ke+BsIosaxag4c7OgxwAtFL1nNx9tjtNP0VT+yMcIAC3HBhIWc3bqnm74+yuxaDky7+pcfSPGI55
/CT2LUg+C848pVwREsJnBZKRe3ZGvR4syzJC9lMjABwgqpnOrCN461JJNM7dcsWohByjgXK2WDUP
Ns5lqgfCKVe0djuYL+encSErfylu2lQJxhppBbgXRXGuRxLwR3LcK/aHRle30s9vydDW+76Id5fT
5YemghDIxVhRVTfBGfOjT+tJhGOOGclIj7zQ8IYXA/SHeSTIkOD73n6ez+63yG0GDLA1lCqyDfO9
l0cjyR8wkaD/g2B2uWMbhZYmwGXoEmRmXeKBcJXp53Nj8/iBKpvUG5CEr0VrDB1K01O+pYm8Jrld
C415It/D7E/u0pZEsrrOXv8VvfPmgHO7TkJT/KkixGQK3gVL1CMGokv5mRGBioHeTKdr2EAnPj7F
3svrnr2f5dt5MZK5xEbDlpsId0yHy/Yur+J6rUUPqtmu/+3Nr+63yDJzPhmMug1Afft/cMFnTKRB
HJ9OdXF0yTclOZZ7B3NGgFXh+1mTYn4rvbqDa4L/11bhq/vFCQRtIhAisZFxi2FmwkeRAilJTuxA
SEKgz8/EoZ0l7scq1euxRUgaPDYr9rLbM6NUbl28ejcjYDEhnZk3htkF0nvVzVPspz0VOfeS0vQG
tDwqvIQdlQntg/5i4bjCdFzTNvBNPhFzFRuK7Ft4WBgJIC5uHapQbhhhj8i581fK7eMO/L7T85Ck
KG8x2qFNCV18RkdcZfbFKc6NZuHOWZwOGefLc+NXR4lpTu5EK2aVglkJBgbV6blQ2tWIy4GHts8a
sXVr6e/8wgzbaBPiWp6VS26rBzqpjExWrSeL8tccc3Fyz9eBw0OR9pt/vcwcC4mVx1waLFqZNXAo
RhOmqMYVdy5gLVZvbWWJd4Zv3Dd5SryLtoPPa1eGPiH1ZwG61/1Yi2fobpnvASqxyu5zDcYC3+8/
a/aoiMYAZx3OD1eh5cJZrvIyYtTkXavzaeq2m8ANBffGPnuSCN42FlQhdqyp3J8oD4t0ZRUI+Dy4
GOslMJXkoxjzkq8rNlvKkp6pRBpl3bYn3nR6uBCInKnhpbB0Y1OFkcMb//qwamUl32C/CY6jD/C5
jt7Bm7hXv/dk7Uara4pqjHQwDt0Ro3odgkiXVDPSIEL/jheLBcA5rwzUXHyNkVDTF1Ugzq9EsWKO
5rJuAWigNLcRhEiXCk+O9vHuxEnxAcnnwpz+COddK1hUZuhZmys3VIJum1+a63AyWAboKUp/F46X
k3DPloKz1/RywMeWu69FzCCKpuqQfVohqYurDzKW/k4IQhVIk0U1pXXaD3IhDzBoNAoRV3GXslz1
7mJjsupR26lLhiOz3dEHFd4ogjXvM0p+huuaE8xSBVU6M0S9dcE31AsQxlYtC938JuJJ8OmzSGrF
5WjqIlTTUbymbQCLKHs/OD54tAQsuzS+AVjIqQcl9tsUevycz5sS5tkBhqi+mMSTwSMdJhpzfmsB
whzcQB1ki6nfBPjOD2kwUXvJ8D/yR1fJ78fs8ZUslQW/s0sR0sUOKJWx0EIUchrWg5dy/9mLVNdR
QpOt33gIi0IjvMrop0W3uiyyDazkM0AQ0qkVmi6hESjCHCA7BW38JLptx848EVqyTUtA6lm+x36V
vzs5Cl57EU7eEQSibvxJY1+EarPVBjzGbf52cv1wA9NTWtCN4LJLFOAoa1SsIqbYpgtGC1UeKeJc
bDEjjA6cUjEeUdMTGSmvwW4ZQ+GaYFcc1+4HnK7N8GGS62UIwilexPnGcmvPMRtmLnxaX9LTDQEZ
tHSUaNlEHmacxhH3LCrTlKx7iPWnNvEswMHjdS+Ra1hY5VO0uBEjT85iYbx8foa9dwM0pLd6GBUx
30MbgFxVCOGWEf5PK6hawrr8NwRMx7jODNCoYRZGjP0RlwcAkfCZAUqGK9YyX5vk9lxMhDsTW6Cu
tw7lQnrkxRcun7GWQXT26D3+D0vNwdhOMIdMRz4mKL6WG6mvREnRWu53UNheM890FGtYaTaLypFI
jzSatTTOa2fMvZpuC5DTtk9A0JV/D/T3WlTp01TXOHZ+qc/n+2n43RWDhp3DK83Ve7C/rt/3CYge
6fhHc9H6hw13+f7mdvDL5hYtgpiJeeEEXVNSuZlXowogZ0wpkPrmBefW7hGA1WkV5kseSwSpPYgc
7DNii20V78eT2DOCh7zvsJlUwGVuGh7L0DllpzYxwb73OhT1W6hjQAmRopQ5ruUfX3KVhgL6MEkC
0C6iqTLpVQJwzoqCqhKVYc+m33cmqJZXPr2wY25dhgNvT8F+QLEzx892JTqIlJEKK8+odf2t9ueQ
xwF5CTXbdAaxWFuvjD4kcyapTAYeOmRD1wcCC3D5LGe8D1pb3ThnXdmcgprGWNijRb9KhftnsIwW
ul9/T9xke7SBuUd31QYhY6KpBtT8WMSEvyb3gI94PqanE00713Dh+6Dw08Ol6RZCvYev4RNWv38+
GlTzYGsHzc26/6Gp21rEBUVNBR1f0t/S2AWumGdIw8rA2gpn7H3LUhk+EK23VYa64woPQgfGTZxf
eeE0Fycf4Kzx2TLScoxnvvjiSpuJ3RcOXgAkYpNJu9cjXGM9iJDMKgelShAdRFZUuzONd8yZ3Zp+
zGQjLT/orrJJcbTEW99xM3F7obGkm5AZ/ae3EHOYqt9hZpWo0qf7FrLbvSA76te9pP88C2i/cJ8d
97Gfh3Su8KfWfg76KzsyogHEE2/cFtR07T8Keb6JLnTohCdoBGlA+Swr+5gHeFbTQDAWQYwNO5PL
jJIze1tC/wtNi3F6wRWIM1uXJn6lDClSRrVk+SQJdvtLgG5h1F2mfjgxB0ti/accOMX/2BNArCTM
4ZVG6UiO1p0FBigGs91/hwywzAogXbCvPlzSplKHt5DZpDAj9KvrFw5QSJzOXw2OdPeOh917fDRp
E4K7bF49g1ninPQviDIC8iuiy/MHKdQMFx6tKGtWVY9RUpQdDGnfOlF01rtrdYYHWdyxH6MW9f4D
6wH3zKxCfKmGKYLFXD475RpTp41WlBaTA+k90zRsTB4Zvxm8L5y4ioQNNPmrC7Z5+bYpWwGQygNN
uwtVts1DHUkUL3fYOcVURQTQsDb7ts3NOXHbxr3C/uPFumWc5yJSUBqct8Wt+uPvNc/fctDBF+U4
lbQP3o41rzTd+USNeqEpiAwQZXmJF2PT1BMhzEbam3xP/o/HtGKVtzd/msWpAYHWwFH1xDcUoJzw
t13uqkQiZPDFRI+V1bO1IqLhLlZQl/Oe0a7IUVJjatdkYbKZTT50mDavsSmmlfIghTqfJ3mDERH/
FWOqsQuVlaxArx+krlk27R5d3lHPoklcJ279bR2nP7O9JZ9nZ+0kI78mgmUCJ/n6WsZcNCdnOPVS
OrxjzRAOBJtixjGu1UEqkB2rn4GnBF4EwS7GD1RWtDKlk6u5OlB4ksJFZw1hFDDO8z72ac/ecH+x
k3LHa/NDQTvzLnINqdfoIdz3MtikFWosfDznoxwvvEFAdgV6K55mCDslBRnvUIyV08vnPgqk97/i
xsKX1dZavnAro/jzkVDC33ua0yZxFnGY1URZROB5CDle+Y2IS90Wu2Smi1AwOC9EB/mZFftuNuse
dQ45tTVzFOkcbDk7KauSc5ZsfKux6ENda0yyjlEod60XMKeuxNklicf8CRJH6C+YYD6B1NhPEMVR
5baeqy4+ETgGmxPlpzO4/IuH/ht0w5fdvIOyfd7o7a4/Usv1rXAvoV2NNNKyiiCfqsZ0cKRYtUqr
96a9uDjc1KxhrsjN91ILIB78/sCjMfVaPDYZIvQgQq9C/jekilIYdqq8opLI9E3PACvf55zHiAaD
g3PQ6D2lRcNAco/AkIb3PSWvvLoIyJIO+o8iU38h60wSLYlJH8Jt28kTSKEIDx+8r+TZ2PCpG3gK
ERbgq06z/WpxYgwTf9+Bxj4i22L7eS6aKMRfWyEPqiXo6SftPWtflcmFRXEGrO+tfwmm88qdBqtL
vV3q1QjsqqQzDM4xJ/Ft8wNsqkhkFYXAMboOxJsG57cOkBFywzbuVV1tsiAJXCk+DTqikJSAVWwt
1qqLloUqkFlFMFsZkTSdu2zGEMGK+7Pacdwo+hLunlTCVV/9r7L781DvrhHXUkdVLjmbuPxroD49
OiDfpyfk75tB2S4Ob3LR2kWudvLiCt24Y1P6azzpBB1+DXmsivJCr0tYq8wcAO3fc0gcfNAhGcCK
xJoyTA2pOZg/wZF7bp3UojLY6oFpZhEyiqcm7NDCyb7wcK4S2dFte4dGPJEAziqbw0L1bmXu+vC+
GGVEPDIYfxndqYNmNGwKgmfsAdzMvRdCMqhfowtKW4+Y5xeKBbHp84prO49BIVqhcds13wbE1Rwh
58pNx/jjdYi7b79Rexw9JdTOS1MuSjFbbM8+Hp/+3lKKsB+t+dJ5LMiRA+Cwk7qMGw/lM2dfcYcH
IrwdZY0vCggsHKaLTbNOv7GKwiygFFiWaVvoAwdVQiK5A/V01wYX+IR3R+ia62LEHZF2ZvLFZdKB
ZK/zH+ovMhRVDMPMdypQEQdDVXAeppjx5tWB0j/BrY5kU+7OMNrOcIuLeVoDUz50o3aveqxfzR71
rk7AWj1Kb4jJQHuKZBpao49C6oGn2aW7cEZs1DOXyKKzfSXOVK58g0vyiNoXpsq+aW89FFLE7sU8
+nhXdaenJ1AfTFxLD3fdjUBypNYvY0zWds5ZbOnZncHdLf1l6yeKrGDsQDsB3nEA10FD8ZfhYfWw
Y/bmrVJFn3ivy4gwNmiqNe0UHPdq8siXsJ7hdbxDsI8NnHZmzmCGR18+s4sblxphVSEDI5XWkS8u
NlL7JD9AdPagnCELl1TS5ZhkDPqtcd78tM31UPTmPd16VTrVyA2r2CONfKUN07ypQh0hO/1JHquV
StQSBNy7Iei1hlDk+onFT4aZ3ZPELAWZhiFkE4k3NtjQ7cH+MpD7DAziYjQPojnF26LIxohRr8a+
07pa3ECiYNGPE8gUwsBkDc8QeBLJIoGP1T3oB1Vh22zrYwkeD6SItjvBrrqcU114UUPYON2bmyWV
ZuP1xL8jOa/iQiLqc8cJ6LLCGgyxR6QxYb2FdfAn5web34y6Sl0HzKjGfur1lAI2Uc7dwMNpCWoe
KOOqiLJ8nz2kMrwWoh49PLkQ3H2qupdr4kzbNqFWcYQiCLDsbMz5Bzwpz8pymL9jgMlkgNj2GEnY
wJT1wTRhmmhrAt6HkfRTXakJXE8xyMUipmaXZCO8fEBlAx+xXFpOfnkkX4TPsvfMV8/zbkVmkJ1t
jdez71IWdot6aTVMJ/jzr/rxArj95r8qOmFGaWbqN9hU6m+TPtBci8pYtChl39WpbekeJGBKxlgk
ClpVGxyIxPPh52rRNygY5bhz8zC+cYEwhwOOToGVjLzM4zccg/KQANK0Masq2UrQOUyG5fONQCcw
qtA0vq7YXrxK9E6DlcEAo94zU4YibMJ5e+7LICRu5V1/vZB0FOo3VvRodCJgYKvK1YAZjWWeCAdl
2fhQrZA4yYz64XCH5n7I3rbDXUjJWyHaCJRhb6ORIpcjdtdsTE/mAxrL1oweszTNoVgbgtkq/6Le
QW3rowqrcGiIVVmiiU8JnQElwbYc4Gq90gEN1WtbiVH5JXjnsFocqpGZzOHI4h1+JvWB3HRTheDe
KbCCmq180zJQ2oAxynCJH5jpxJx8VW5eaR4JHrfRoPCtFJN77b4qUjzUvuxG3BY/5ouaGEaT47TE
ITx3OYuhb0y0kx/y4bfhUFKdJdwEa+WwCuLIZu4Xp5FH9N3unC8EU1eHq1EjRSuZ2pdZt6l8e/Jr
u+ARC3lcyCCRq+bbQnlloxcpKrVJJdRQEcozYYJfRrHxGuR4O38vTF/alx17K95K6gC9oc+alPNi
sBVnB17EePRnC1mD0iSVrnsPzxJJF5+HJV3RwUsETobxM8C4lIOmhm3kaHBzepQahFQHh3baRWu1
97b5XA9vdKWnot8y7Knmd6gQFLcKwwHXgbIMd2Lf7X8H7gJ6Q7zj02W8ZFN1+BZUrAUO0XhOeIb2
1r0dQiQArxGod+ejaJ4E4nLky5ePUmXazZ2tfch3GOdWBNVFzdCntWBlPoA2C3u7sjytuei9Dd1l
qb4rMy8rjJK83ukGTSlvL1M7F0fS141owIfIp+rEvYsjRtjwE1KKUNPAer1OATbqJHZfcNW1x/++
6ZIHj9XYF38yX9g7xgFhf4gJ73rFKNkmQfDC8DVXJQ0JH4dlrOcsOn+d3APl9T5AW+X4ACpjhvGC
o1cwts0h9hlv4R1WRUOCKbMogz32LFHyO68k/Rb+00bNndzxmWUMNvSzH75y8znT6fm1usTIJDfB
K2g1MC0nHPy8gOFH6G3Wf/+M+vxDPSfk97dvOsXC2942zsWskchIm7D+Xw/itDqOqtGXX7z5DiuJ
d8I4VgjRztGo+oh3IZm/4rV4mxuhWmBHXUJgmH2L3RsTRO7WICL5DeeZRY615DHV2iT5zvi0jQFJ
/gpI7hLKbDNsQRztpohkVhIXXY3FObv3n93bYAxqWE/vyQq9Ho8berVUOLNHGWEfXJTcfnQyccc4
UIBwEgQPBh9m5uAjB/Cdpt7JIkAG6fD2YiEin9Wq3l/f75kPaVmpdfxaVPIs+3eHOxoHRbl0PZED
99DCVgYRVspn39N9jBcU96S4JpmgoClIlRdKQgKEHEVlvsXRvRZCbsnL2VK5io1TYC/t9HIKGgIg
AYFrUQIoWHGZcgTpx4ZN8/LVFnzuPxquusZ3wOfKE94bI8tygAHMj8C/reqm5KYoZ0aI9tbzn+sf
jMqDNOBlc3YcNWQK/JbdZrETC+EmkYk1EgGG+Z5srtCnL0awtf6p86yfOWXAsoAbr8dFO4jL/D8D
HnbEW8PgI+MFduDh36Igj6xLb5nROjL1JXqyKmyirDsv+fWxYYA/bQq6JOZmLo47AhYxj62L/Nlm
/cMUxLjSGEtNNRt48zjN43rfumpXz6XyGjG/dGTx77JJ8jy6fZSGz+86BMwDEd1Sy2ZyJQYHJDlV
A4Ovr3xIXGd8vNhKu+uI1CcPEuAwmog1+QwILoXQmderBEd7SJl8fBw+gsywX/7bv3D34/sEUsBK
EtI7B7Z7rxN11LZKSqrJ1BkWGOXoyVXCUZ25GlkKrBqu068fgRaA7hpueW+kvdT4n0X5TvN2sW4/
BKXdbFo03KVRFMqFskIHzZLbxT5DQFSWc/kVN7mW9fASj6ksitNj6FsYQHq5Jhdd2MT+A1EnY0UQ
YrJFFdX83mAyNEzWeevMGNy114EJ1SqIyzjnqXpo0SoYR0ssOVRSgpQBlxZH1FmmPPLGz/0Dhrd0
e8u8mhdsWJvRE9jZA4fDyCL/KIQ5/DvCNdMuRIvcpfolbp9yeChTNBnXmVQTOT1Si59HRkihvaLW
TIgD+WcNJbKYa1uj7dZieIHZplliRUSAsc/s7QLDQbvv4LAskzw2Rip0bn8n7wCwKVpQt7LbZSZ+
z2GoT7UwzlrUuuKH6MecRhb0sx8/odHPHhNlsKxq1WMoqyHwS5rZPpSrxV3gVLmM3fR9NCvE6aeI
FLM5s+7fjevwkPb+pFZUP8fjC0IWawKVODtbDCVZ8xX15RPOb1ZS8aGOPQd/Lj7w17IrU1JdMWNV
gaSLW2XN+t0s1fCqrGMGFBLI2132zuwtKOdnvHAym52ZVBIasZBdVUhU+Y4PZfuCbvUeVsDsCzV7
MAy9hjoZps0juw3RXKzFJtLLv9UO8mv257wtHaMwDOSumjvg7HMbYgVWaoCBwriah/2zWekpH2Cb
TorfPUKpoD5n8jh5tmrHPnwIJbH6RQ4qQ9IDNzjaVbGTzTk63QHAQE1EbvcFFheSslVswAj8qN/4
c6W8XykvFWQbFQtZaxztfUemkXIdXu+z2L14W5++6INpOpDIclriYrQJNlhF5e7uonr7VxtCSvOy
HLPj0gi4hSOqcGUqaMbBVgEGpHX3nE2e/tMTj1h0/u5n8Xt+KNjqM0OgOqrSPyXtjHlYdKmybkLo
qRqdc3FrdIYUiz126Ry1OqW+nIQ3fC4SOO9FFpCHzyxhQr/3stvh8WMJKfj0LRC6I4A0o5fUuWCu
vRlx9XbD1NAC1Xuay0ZEgzNT8nztTJ26301zej2w7OgS702x8RaQHZPl9WJsEuaNuqVKOWCvEYN4
rDm8r0uNR8z4EBjNcWpQc74xW/+a9b7Orr7zIiq2Eafpfi1rpciJo6LyKsIdmFeqye9d3p+6BKA4
YSPV2yMc5Z5J+khE6uZElCe8wnEOP8zaksA8efD5bmmuHo+wV3alhYvytwXu8qFHfQCnkzwUbSfC
9qjiwrXPSWgMnZ7my4QCWQcYctix40hz/3TXQylrq4nuQra13qP/ussPwL7pXXOr5eelzW3GFgwZ
VwARWQuMt4x6CzOHtW9frmWTzPsab5UqmjiMwOYqGIXKDJN1HGV2aKkHGnn4yx7bDeBvXkXeHcVf
LNwVojXWZLUEH+A6P7bsI7Og5TMPdYzbi0AjXNYMp3a2fEIqW700DhkqS63E7/ukrMUQOvGH6air
9WfUnbsBmJSzMOootXs8uTdyB4EbrZaTf8+a3d63O1Na+w9XFJpwFqs40kvIQEx5iWURIocBpNCA
OBNa7yTbX6G04iLeJJzQRmts3d3a0oNoxg4StZuwDlWPc7LGV7eNzubduSo4UWXad9VHHJAqN5aE
iIpxrxZ8CgLElgMuyMJLPtpG3UeFLay6LE6hG9mjaVkIu1pkp6+zwXj7VApL+acLcoCFxkExU0Sa
IaDXzd4PIKZadIN/YNdatpkccebGDyyRmJ6QsrZviFZ4ZvO3SIzTjONRygEIoMsXWcVSV1dKhwFD
LweYcHcDh1a1BG20jGDLuMCcE3TNHpNdiZcftgFIuqHZFhdF3BbS61GDdrfLHuqF3MoPLqwhrD3m
cjfJ+yuH2uQ4m8L7MrBOlUWRv9TuWp/0bMENdFA7Sk9o35JM68dFY6IaTJk2PiecTR3GvSuB8XxF
4SoIwNdeigwkwd/vB6J6yOuKXTWhXLBdh5c1ZNhOEgn8kNMgBuvbEF347ulSAQlnw5JvoN5Tg6ko
JMOZYbREgtfS/TYXyIZQbC99wpOgdSeDGIAW7ng7msnnU44mJ2O31LWYaEYf+QNdNDOeTe08kCcM
UXl4wxL4V0a/qGjo9MGaGSONoHiMsweO9eGYsg442G9kAgApW0VjSiOIgEayqEPeq4ZDxCPd9+RX
D8mAAIkuZ/dm937JLoLmGT9v+LYBAmq84C55BmsJZrPR1xRDUIfLIVSQPrDXHlHfOJoYUZeeLhic
/keVtKFCWqbCqxGD0bKJfJYGGuY2KNKE9k1rFFK139asanLY1Sxdns4v9VyqJlXlghx4tZ3nqh1s
BaFFRq8I/UsUZp/d/ZzdWB+P3PcxkUbqiLAnkpreoUg2l4aO1quLHfiwC1Ov0SvlE6nK5wegsS/d
BV+Ec7iXiEyT5SST1OdGx3PPvzNb+Nu6CD3pk/ASxYRUqmTfyGX2vzgfVm0qz10hZq6QXWviOe0m
dF6AAfVXzPdiQ03WvGjY/ITFZOf/FHPQBFJUHXWe2fF476RapBg/yuzNwdVMJDM3Wb2TnyivybCM
+uQ/+v3p+C3+OVPwymQrR0BprumRQFQ6K992RhhAjZmDhrZkdZXYZURBAvx51rdjsSpY8S5PPnhH
G1xH7+C3BuQF3PxrHO7LX8Q3EkTI7mB1WbFXn84WWdqX1UJATAIyi4ak5OFXiVh4BNHSGn2hfjZH
uBFYpoa5Rqk9A4KoH9l6fe5C+DgfxxN5tDQarQhBZIJ9M7ydwmZmDnJQaCVUlSgoTvgy3eaBEPZB
G2UgOjmPA6UKgdG4auGq3tUKrPueBCRvMO/TPth+tXUmsEK5bKGEaRP4YRIMn3hSIs13IPbmGcjJ
ZpoH2Ka6CqhOnSmUdtTbew3MGc15dELduS01Wjun5MMzwXjvREU3HZeHCnd4ah8Don0OAqvmHTkr
JUIIozBh7NoSy/UkMBnULbKf3uAuNOEWsbqxdpDcI69tz4KfJ7EnaHPgARQqUzXQAtjgfGW1iBBE
v2HakbQSPt3Wypw5AU1hi6fNRpVDftcoFduknPqGTs6EyZimc0QcXjSh4dJ6n48Sc65lHV94OB6a
T9QkXHAjAxDcHAmR2t6OSrLQvz72ohNGXXL0qg97NUgAL5OMfYcWq5wVuYxH8GGUy5laOH5ptOlq
lGiUs8gu3d39fQ3dFFccRLSz/7+CO5WWP/1SCpnHk9zdAvawwy/yWlDQ+XICz7SygV1b79Ja5APr
JsfCY7mY6YrUmwf+49eBq2bM4a7/R1UcZQdTioUg9xUrKROJDrfHlsyh7AACG5ik2vh/ZfXxB4rg
kHSi1k+Yqpl87Zr2QzS+csjmm+2F7KIgVNWreTB7bcuUoE7ume6gqaub+HHOKtex7NYh/LlVPBoN
zUNAcx8J8r2HxPEl4YTWpJQvT2ad7P30L5tLveXTgUE8SB/T9BSKiKvIvivFN7N4toB0fxS5s53z
fcYfemFVV7qQbxLDPzM/BLz/NNwfKY2pa3w5gveMm4LubeI1lj+LuMe9Q7RtBnPbw+G5WAQwJ5fq
7nK7i/b+o+tWH3zzm9MjMTOejQ+FYwkEuUT56HLtnv/8cEwNfRVpLCr6NIvsyOAxqRRVVtLQ5puR
DASOZvlrXZg/WcXka4bSfahtSyI4xqknofFw6phWbbUwfCy4pHqbKi1xNzHeEEGA66GK5NUmiWZr
b8CInAHFUlNXhCJYe1Pbf6LG+hGpyFd7q7PXTGnCr/FG7pItU6mf7fTpePcmuzUx79lPt5wb4ss3
qgIlxluIUXRgfhtMLauQFV3yEzWrX757Kux/N6rCluLV9Uz3D5B6f5ScRxqIldE6/bsu7VPDCPWN
f35qfX9Ztp/Gm3ClHBMb6C3Y1Rtr7II6W/RjIQqy4kjVEJZQQqopzs6R9juMRUFDJVn1lLFn/XMu
y3h35zgfDOsoPe2w/d6v7e2GwdGXDdJOkjW1+Zq55ndGBKpuhewVHSAqDcO89fYcvyZ9D7fXdVca
C2sTA0wEwdGbBK9bxJa8aEp/LvrYsyiFO7tjw3rVX3vUkOKyPcoZJY09Wq5HH3xuop+DCznyNp6b
7tLK0t65yGqQTxI7BxPNNRCvMKBFi9tSXFjZ7JkXg0RTPDHd5g5IfTbEsWuwLC6sgPUskA/JGVap
00TbAW1InmKNg62LBpL1isxtJ86dFbpYDLhZTr3ZNdzdHTMqBH6fFYKlwlVPc0LfXeOXNDDoAtJn
8k/zr2y+xBw8Zs3b/3UL9iDs86Bo5Jbf/jf1tvsLXnX6FbtKIVBhiYEic4vo9xyybEb5YiqbPwmc
bLLytbUeYsfuZP480xs53g0Tz2diXskUKvkz/ImwMXL4+bA7GUZYbNgI1/KUFd3XO3eGCQuPZMKO
9vARQQ05iuT6mMz6LKi4D3S4UCwOws7N6p/qbaKgf37cTBLAKeuc9MujGwope1gBcztYI+qbRoHA
gOMbmyVwpFYGCz1w2U4QMHq/z54f8R3yxpLnhS6idV7RJkRqJAXhlmaOJkkhgvEY3egc1IB15k5X
XQxyvFjgP56J2Qd++8wLihKqcBssZRvy1d48yOdm2miXN5cC2LX1gGDJ7kMcWLRgjtgLjxa5BE1u
7xAEVQmTGGftH9Zb7DpdOHjdjL750etDaBVKMVGMyaKzDvB3bzhYh3HGyFA5ueApb0HnQS8ivjc/
BsqqqHkCNjKGhHiVOq29MWttI74u3OjSJIW83+mrQhVX+QCN8+0RvFKsKxVFb3tk1ZhXLLSGFza6
kkpFMy1fkNRGVgLNz85/9uX5IgF5loxFE7f0kBCSdCtxHZvXNwMgsJ8XDRx81InroZPDYTD7iyIt
nTwjh1o6eyUjZBtmfjuXYY/7+cmvVHyZhHw2Xla2ddm0L9lbR/AeEtetCx0fU8vA5tmFFU/4yWLQ
VkgeCeahBFGF9xgr+UwIHGbu7Bv7HYd22YJfQbgl8vpcdA9de539Zb8If6y0T4Xk6DKIWffbYLDl
7lxfomZoRF2LggupLC63ocMZ5C0MC/FQtwkvOj3cSmkgoprpejEGsvO4Ugue4BY1oqjsGMLjx4a+
r38pHnZO0rsTbHvCKMBPPesjvRvCW8oJyiFKLm8qIQh7bkuRCDvA7h/qrdqbta0vGHQ1Taz7y+16
QYnpKDpsm9LvBpokHaa9/gwqwlN6iOGjEAn69fKRynflygbJpcmo3iui7ZmzQHwvSQZpfD0a1ee1
UyFuf0LiTp6t8n0opogaVEV8G63jOpQZSDsy0axQLdQ+an5h/8o6dH5eHg8aZfynlsP2r1XjMHKj
LWI3dHuSs1wnDIW/KG69aywQHBIVUHf+Ez9nXBnSHeoRKcBBv8pu3Z2inK1o7O5B4z4GTwqTbuua
4F+yrGmczcZze2LgD2Qmrki4Si1VQ66bmUu4mhw0vGGl+FqPjiTlxtRbX3IY0MpXmaa69AFRWhAE
HHfRWrl/wNpng1j/uRJdBCib3VtGFnrabYJMlBL0U8aHPaTBYOiPHZ1rGj9J/OkukGrrFGyo8JDu
lWcBpl1hK1eElOx2Kef/f27q5WjlauDvcwdzqZ4yrHPEUdNKiDDHE+LgPxK/KAind23AO+Lc0Njg
spms+/0Vdq3vVL9663NCPwAYLFbCNXdXu+pSDXydqicgNKoMVyZDBcyaXttmiNh1l1t9xCJ93KvR
2J0cXqXzVymq9As/3HqnZ026nrJXkXo90m1VALBsC5qYu0FBQG3rkHwhQ3FA5Ht77TId/JAhg6km
+ryC50Cl4v4nNUBmjGVRb7KHtx2Yvp5j9Bpiz8/m/x9u0gq95x90bjfFm+PyW3/o/xy1miRMy6na
TxikVhavpTOj9+2wDNWJwrTPk7gyajnR1M+DII3PIrsFU/iW4EJd4z6TCUzIyROBTjE/B27kudPC
9HE7LS2D+jHMN3Oqlyg5CBUathhHFcOp178aaeI2G4Q6sHp/chDYcpuRzxK/p/oiiGt5bUS4Q3wT
A6gxyZU4Md7CxhmG33zZPL7pLi/hbshNhZT7zXsY02lb3bGwlaUOB1Z32brrgs8+r6kX+etxKvXK
LOt0UKQy+pq9oP3cOeLJd+gI0k9xVs6Rxs8Kt9T2TCKgTcl+golUWloWhhUBrxpzTkjrKJO8ni9A
btZ8vzAdSPVdYR306Ary8IeFtDtJXTMj7sdFr5C1DxBLpm4TZ06C6lrUA2ISB2RokbvClpel7U89
P017Zq6WPHxenDv44KPKDGCPTUvX7ZdwSWcBWPUHUsMrjiCs4G4UWQZe3KLfD6NgOfV4gHDbmz36
05PCpWL3brAV4G3Pj41uBDjeOnHyGEzVa/R/VBTInKjNJT6ZCnoBTzINJQ+AUDSxiSqcjQDVLr5T
+N6lAsKTa4+BJNlzHzo26XD06XJHWKc0taex0W43fSK4XsLQ6uhDDJM8hldAP4Fw8HrvygpTnVSy
vzD3uKFGPcOkkt7D5Qxx5vZ97prV68uC65PeEXovTzQ07A1Id0HZrH46yEjM8yVAixYWQgC8we3g
Q1dob6G8TxXS83/hI+N/d/1SwpYc162+7yGq4F9PTPdeqU8Ls/nkrostG5EVFDMhYHs6Kc8KO39C
RfgsFjRgMp5UJg7hQOUIQ+KRkJ3B2Cfabmdvc78uwUXJtLMPqqmNgien4XzTLBlMsK9Kcg2FmawF
tCUKamv8bgrHDRMQg8tkP6XGuEtyo8wnImcyOqwqNm1zfvhJzjQ3484Z6fS47mJZKy8Jm7NVKL7q
RYpjpu8PeKZFiu5PagNJF1BmUJh3A2p5cOXR2Ic8SIHQVMSiNe2wYQJQ2upSpQXKnKdcpUIscczh
uwF5DnsnR+jcRD0fILedaRBco05vNgB0BkMRJ+ZyfuaSrbEk3AiJ7VArPjjB8nEoa5o33GoiL2nP
6jVqW/swokbG4csaXSbqrNmZvQWWJsrmaYXWXkaW22pNXKv7Sqn1DJkYb5RNm6JfFoM3skX7cawR
FFv2dcRJw3k09jLoA7uKAZJIP2wQJ/NWW4bTCMZoKH0CisAJIcCAlFGdZRB7b57Cmx7mvlHHsqK7
V/kY4WCVmGwk8EjrGdzsW6zIa3MDCcpYrHoThquKobgDReLrYncaWBHTnOUb37nhrvEwgIoW0MeG
vzI9PIyT7JKLGSj/DUA+XicbwK1jdJLfg4V2bK12OpzIRTY7Xoyd3fzJ7isH44Xi0Cf7zI3WDKHn
4cS7GXd+soMrIrjLs4HRZVmYpZv9Cuw3f1iZXEiQ+Rcydd+ImwaN5mLWcnxjYMM8/HkeHZtrnZ7X
1ZqOuCMl6PkEqhWcHU9IrpgwxaUJbLI7QMTxLnuIKHl1nhQ8hB9sNIGrX+JAerObQKU3EqrcSjuy
6vj260DTbFLqhO2dWFGfc2gK2Njy5Sa4vZYeeZS4aCqsd8iclWKtapOgiBqczB6lLM2BwYhWFy1T
MtT8aZW/u6dsQKsCSLjbs0iCc305RZVbrIV4BqxQN7Zas54T7mEADDFsoV/mfibgXKFTNAjgx550
cbEtqQQM5XEQR2goXWAXHxOrHRJfYQmzJvN8UTR6WUa3S8N2HU2xDfUGTNQ+jZUPKOYKt2VYmnpW
+UUKS8Zes2H86eGQFDbV+eBOAJ480F0fzkw0CdNWot761yLNIvSxppQr1l62D8hH/y/BDwf8t66c
l7FeL2PJgED53yWkp+cDcdQukEMIeb/kw5EYn7yTz7dfdpbceI+pNL/DXRdZ66vQAy/vEAcrzVvt
lb3pUb6tp4FhSaKsElqCLWljsq3X5uPoK1AWkF6V7HM6jKZQXQbS6ALG0at3XUFAMnjSKWsYul61
zQawcHSWlGHdkE6aTBG1B4IVEivInHXuxQzl/tmadMXcyF/FRrw/pkEdgU1SqcZ/4ISluzcRW+r/
PSi+L8vV05phZTwQv/1MiyEXOIbehd6KSw9sdKXsq57uVxV2807KgVgEisijGIEGC4JZvEN3jhAi
7S9QGOjqbWTIT19yzxYdL4TeMy5O/uaM00ORBcDwT0GzbOLjhFvBRl2h4MiXEPNUtV2CtxffDa9y
VGX8u6rL/g2Co9oeXKQ6MRQCmA8BoLNVt7IFT0clrE1goPbhlOsXFYHeGv/eYK93seIpjPfz20YI
wxeeTgmTf2U+LqC1zvXZmGU+zkYYk79QX8MANSX2MO28IpgVNgqM+E6q76JT8FSMdVr3zArid/wX
UY7KcUGTRmKOYakJBYQBX89bw7x/pHFRiY3LU4X7YBowCH+KwrPxqZJiGIXumNSBMcd7HZttob48
jziYEcDh9+HXAC1iE/KI62pK0MI8DJZBB4+2AxmOPn+OGiAvIgJ3cUeebqYO7S0RTdQHbYT73NLy
3Ih4r5hMs41jYhz4bnbjv2LOEj87ARL0YM5d2KtzwGKM3IxDbfierw6L4B5xpL03gAb354DMREmL
kyFRTFK546eJMZS0stVTf/nmfu72ucJo1UGDo4Skh+ieZwcCyfpLBDO0LPft+l0dZ1QcYox5zXHi
sbobMChUHEJ6RudRvff/OfreicIdVVSQnc8E8sjJXHbYEmInWFWFVbkrCwGvlo5Bxj+NjijzBpHX
/E4zMs4NxvwN7zzfjl/5m3gakIfvgCzN91fzS6gPsiO53Ucxo9tzo0Kf4a6yJZmjUZAiU7YCB8GT
sHkBz5Mr4qwRk157hkTixUS2EP2FA8lp0nK9Tm0NPMsfapmepoLqCtfPI5yQLcpBHcOqqh+3tP+E
gNic4DY4UWzQ0wvROw8Hl5kVEQKkAWws5pxKbN3wmWfGpbgPEfaS7vl8Ckm5v2pQG+jD7HDZk6Dq
OJJK3cikerPuCK9Sci4wwmLa75QeKaMmTFhmenWKGVigfB0ecnaSuUSpmWTq3SKM4mwZ7I1O1wp4
tV6hI4J4SexU/ue23uDPccMY/9Q7BKjHhHHKssdb1QZa4pMmhlDgWvr3FnRROBACHuzc22cY0TIU
jve1VdPL13Gfx1+/5gUneXOqOzcfLmYVJscaP3m6LK9hTbdNiCT/gxr7fkoiMvJdnt6R8plxc/7P
Vni7f/Yrhwfs8w4JEpnx/83xiJjGfGpKB/YaoCQro9OmqzGDxu50m4fdCDiFG0Y4kxfi7fpukINx
3ffTvrPhqvA+NJlvMHm2b+SbyxUR8uJtou16GjwbCwxb6ypvd1VEotd6ZnIck6IGtKXs0bOASQXt
KBf0OAnZClt15tNAGPNGnwJ3j1brtoFF1t5lbkdxsd9FKSYPylD2qEt9bwoyQVAKKkOgCCHyScTj
+YOQousoO7GWlrIn8Du0n3ifPOQY+TW9tPwmsM4+Zm5vB8d3LERkaPNKH6ScQMD1ALTrJ909qm4Y
OMqp3B7VpVX+7S6xDFAld1uJ5sGaBcfmtB2MKelJxbxFr5JvOsqoHwuKF1U2cVDT8xvc8O3DOCF0
yR5ai3Y0kIgh8ld5VS5Zo9uKmVvgpLYJI8SxFPyyT3vixW+VWG0kh2T7krjdY2KiWotEK0EQCJBx
8D96y2LnkCAwENQD4GdvwrM2CSdLc2LCV77QtC5/I/UlEKenCmAg/jxh9gUBnznDoaD2tCrhaMb7
hW17NXoczCjchC35MZuX82cXOwZxIpOI6vMKDBXapeB108rBga/a8hd+JFK4yMmwINepdOiCEAtW
VkBLFSChI1KDD3XZfXx65BzbdUvZHa/kO2c227oHbJZ3tUSLkiODPIqhw2i6ipQAJDVKFyzmzRhQ
0Zj9/C9SFQhZ8afXxfdNCDXD7nSuW/CzrbxoGxsSApxjv79wjudsLzSd4cUi92y39NW9v3ckQ+GV
L8mu8KJXJfFKv+m76EksLbbefXoIxabaxj3xObgMBRIhIYvqMZnoP1F3MXi1e0t7F6GKTwHyVUzs
R5YpF2RJM47ydIRuBGSNVehJcC7IG0tSaG8YP+v3QsUSBbTrjiJ4nIrjJD5QvA+zgt9oFj8n0Ac7
/d7NSkDbJewQJOtxdaChaHLmTYCl459TTGEuvAi7AQ3/cg3/tz17L17MF+5/ZNJEApjesKXcWDTg
p+5g2errUE9qGXf/Llxsi+WQ5TA4f1KYqLIauvdV6nYwtGQavMcmK4EKL9f8RJ2fXip8oOsLvrD9
Bp9QQro0mj9iLjkP0sf+zMesJ9pPcnD93RA06V/zwg3QMjmqLRULRznJqqKmXCM0GUg6hYZNUMVr
bCMAT8dt3TNEkptqHLkD7tTrPum8JAs7/nyJh+uQWfsf9hly54N5gnG3FlaatgJudK0/TgJRr+4H
09YK7mkzrV/4TpeROvMcgbehk2WRR21EVWy8knZJxF0ECm25XeGfnOIRkqnkLoYYUnB3denlfiUT
tUHfUwguTrK+adQpJBY8D/qS7OyaHYu1vJe+bMARhTCGpP5ammMeuxmHYR7oZ+jGY6xTtr2gPWgb
i4wqzYgfhuhaHoleX30RgFoMp7RWLDSxw/TJgrlJ+RRJYVwg+ZCE2XeEXXM9Qw4PGvSnk6W9oE1s
52nTORkIHwPE5s3PUJiT9XkR4kxJ6A3Al0jWMNWj2QPO8OqJi9xwsvNtA2TdRvhPV5Vk6ZROAylQ
uBuVZ6QSI53WMYo6Y7UKM6/yIfHLtPtkU7jOPAMnoLrFzINld9x53gZPy8aT82W7Dq/uP+Ck/Fc2
IwHSsTkdxCdtgqzcTPh9cN7JtOCWRwOsDcy338FlT+TRqpRwuAIN7ai0qQ14bmQtiuEqwV+/CouS
UkrWOLan2rNnMPnNfwSwFGkgQaVaQEaI7iPo0oBxdnqjfUzBtL//bpRNr75tm06uPqgJ1tRn0/R5
i9qP7FmG5R2bIf9JKOE8op+gzeSq06q7hSF5RrnEYdElVM5ac2D+ZLMBUHsAxZ5hLJv8szeUDjym
uwsssv1iYK8y9EYq5XVLYom9ekwjFXTZCWdAiJwGt8Z3I6F5RBRoT6Yi14P34FXIHM93r3Ot0lRN
EnwpiLmxG40EfJcY6Qx+WuSX8s8ZMFGBOUuZM8RQO2zwt753TZtKaraWobNgZcAAfcuEECcqhMNg
MJOWC2qvgBgdGgqTMlwdL4kK1T/h84F2KpZv/427SyaSKk+jhmzHddskkjaVmtdYI8bjBXPge0wR
LevhtD9EKtM0Q+0mmJdifSN23bv3It+TObfyJydI8n+ww9qWonREDQaTBGvpu00zbiJkMmX8oqJ6
gMbhW1Dd1kcJGWLi99sAOiroz7Dg85yoqwSU7iPdIhu14/0wc8R0w7cPd8sWtZMsWRGSDDm6NIVk
PJIfwbmfQr85mx7pNjkklJ5uXjTUMtrsBXKCUnGn1M9EBZdWNrbmTug00VMipQNz9Juwf6Wl8Msj
6wpspBMVLMoOzPSvDT2KOgoOGSxRvjA8czP3S17AtZ5RoxjjwPwJYbD8FVNiy+DwnteOSth5vLxz
Nuxb7FngGSz9WLaKwCAK6wbQEovh379XhUzlwdq1AUhn7rxasJSQCKARSt10Vm6asG4NYp+GH380
cd7mL0nCMM6P1Gm7mxqqUInlU84Bxr/84VVSQHUxpza+4VaTD7dyTIofTJwSaVxmGRjinEEd8EDu
9tUEyVctyUnHjpKUbDZtyAlw2cVodfetwln66vc8azzwVSUdDyWPkjMJzQljSKTBX6Fkq7+jf3XV
3KKQ1j3drdfmpm7IWxYDlBDdaBrCH5T4n8XozhwDtCKnNiz5xzhLwYAJYv/rmFLFAhV9DNgvN7pV
RO0DJJDaZHgpRjUGK41Yhi7UvM3+7XYILoDxh977eEK/7h6iyt6IxS1y5kSChc+HG5wAkU0IZDKN
e80aUQkJf8MEdvIW4WnaBX3mhwntvm0W3gronm06f1SZF0MfiP1juw0SJtT4QdBeRKyyT/HBIz/Y
DaiIWzJI+CjdtgTNEJS1y5IVDatI0p8IL583oP8Fe1YaxYmfDvv9YvDtfVThL3dkoHdx2xhExtn/
il48XBnBL4/5wbHiz3QtzrybY55/7lKFoO9JkK7lyKTwpMMNzAkCDUGvLFulKh0/PeNXKx9pfdtE
9/9UAk89jERVrQbTfyLAF70vCDvytCgcB+jWfgzmlP892Rx6O5dSbqBAbuKrz3UG91U+jPw0uJ4B
Z4ZdiC15XIZPk5wHgIPy7AFzH82Qf4zh6xkt/KUZwvXdn680mcWQbM6GJmer7HBXTNOR+wKPBxmx
uXhED0/4H6fSB1QPdf1F1TvSKjTBmAamYoTXC1cUSq7VcV2GRAcvqgp9fsvU9JO5RjdbC/dd5mcG
hsvqo9mCjaQCFsiZrkkOCdD+FxGsy8fv/ufCilr7s2ylFouq4s6wJyL9RovQNdVtqs06WP2AkMmJ
kStag2lnUdx+OhFLnWnPq/n35yrM4pNctq0p/uQYbAy1lDAnWmLtS5cy5R2sdNIYxq2tTFO7BXNR
5rpj8Nkc6VanLqTvdwRmdCG83Ca+aMKEqEAGCHHsnir12l2hD0TzvMeWpm/RHFTEm2NgvNyJyfHp
FHQL3DUCmc4kWJAMoslLNX5dnO7mylWz2CP0lzcFmc9QLoP/35amqs6hz3DalHqIRM6h4H2vHAY+
PyoIVy3lMUQgbZHsF4KCmlYamFRlMxED7tmO4yjwSpb53EQ0TfTtbSVr9N480ygtSecVqyFGEtfE
ExEswC81iA6SWMyQ/6s0Eczf5cGVgTnTcQyGtE0mZ8J3BjW6WhVL6SZS70EnbQTtRM2GtgGjXrjy
hNkb65Qxxubl3Fkz8lVwvJbcLT20rxH6Kv/hlVtHSaIeg4sXBwYnfald2dfK7liQOz/er78b8XLV
tH9qIU7ADZaQA01ssZDHlm3mrYTdESSXI8qnGCtLkCHFxlob93iFUUktwr0l5qKekJS5J/DNP2pD
5xT1Wqfz/PG35I0j2HlcS/YikRb5xwPLnU59FBtOoa2kLqNis7dF/yPM14V4e8txcESPR/X5LExj
rpbBLwMrKYopB6rKR1u1y2inFa9LQrO8SSMsSkX3qJOAgqhljeFIpLYMnGo2g53gwUSqhKrIe5ab
bCkhlmglCJqKGQJ4nkBNrn/Fi3EiBqUDHTZ6vCVk+JHveHF9xuIb/RmUqSAnjo94fMXOrETA4mVi
AxLmeOVhfyk2e/wMS4zr/W7kWJD/7Rbiwl8ogKlNQMi9OShEacSy8+o0dP2yckGDn9s6+1lSXJ+K
89d3GqBosOnJRlSJ5IA/kHw6stO4jr7BCSxYr+B1G6jA4qL/nw3y8Cx19MaRW72nKFMbUDp8P6K7
Gdif+KVaTK/pYZi1PIOeSAIZkwcFLprL89GUmKdT7qyVWETozxAvUUwqri4eYWMaQddGp18OlIWr
WplcGaShIZ2F5XGM5bSbDDbyVTxBtAQ8MPhis7FfpsZU+UJGUmcEjTTa4YJT9lOMmXP1WK56E4wz
w2c7VOBA+8E83bu4lFVayK5L/Kige2lbqh2wbsrckIBtsegnSJSUkbala5KUrT8215qT9mqqRh52
LoMq9BL9QCWq4wIFCxwffs5wLbrQzqvHjlkexTy+ZHQ6A6oJu1zIOY1moURnC5AviT+RcevUrztc
p4Ts5+L4c9sarQGhE7Gy+/wfVNyQx4M2Bk3khWxnxtDsIUZqW256sfgO29KyF/k2Ifh8ihASvC0t
alLicSrmI93xKUBIskzOnz2CxkfJmpSQ6XVSmeaX0mB8SXmVdF/HdZs0DA5ULrYARzo/Hf6egaEY
5PvtjvzaqM6L5yWw1ElW6z+8RbOMIviF3faWcewC4dXGOnUuXkBQBI2o3xpK2fqUfuTStBnIB+Fk
3WFf0sKXOcyETwgDIG7nFTlxNg7VuMdrrjGVhL5NtxazbF/vwD40PLio+Y8wR/oiT04H6ixNIPQR
3TfU1ei72Ho9WjHqlyvKn1RIOSDeiJ1/ZMw2avZ3Vb2jXzEDfQAWL49Pa+MYVYPp7SuEKyC6SJ0l
H/VMy+prSdIbOMJDv9MgDvDU6DA2p7jOm54S3SISZV2S+BfLR35uBULCvTbvVBy3RgWG1HUpOmC+
rS3PhaMSVdmmgI42qCIcgGMDzkHw/2eYCiU4LJpOC3RBK2m7H+WbTSqghneRhtaH4jdEzOLU5NR0
VHVOcPNiode+b8oRSkqufXLUlUQmsjsxPi6+K27geoq/J3YD+SnNSlHa+QBio49lDh3boizhlQiI
MmbhfG8TG37UnQq8UxSv8txUkxK0ctq+JCSV3ofsM2czb+vpG831KqcBR+R4ROmmITpjtDLOzU97
ycPOAghQD5rClZo8Ey80WHXCAe/RT2YP02fWs93xXR6mo00yrbb2TncOXpsHGkDEOAxvBWiRTGot
/J+PB4dAZZ3GKjzd6MmaS+wsQQ5nhhSMh9e248v+J/FuMIQGodAS1XakDZN8tGdu9pPU1tIq+V3d
bwO3aGCKOFiFhvlVj7tvBQNW6J243cl5NMyaJkC4ZUyofutiO8UQ38ivZv795NMJAdAVRxS0ZG1Q
UcDfHBLih2lsnbk/REqR3fEiAiBMn90Xdfclu/LhO7DnJRJMWa0aTCa6HaQZy7r/pM+JIj4hh5iE
UJpkSQ2p85lLy0JVG52eIpqQ4e3scCIhjZef/MjDfrUN9uI38tUHIjqIpHDYIafdAE8K2qF4tZhq
Nd6njTXxwhlVAfwZYJfyDbnbVLoQaklMrgFzKXX0VIwMN7T2ldD68WE1QZR5U/oU2r8XGGg2vdXT
nzLdjItq9pIvsMOgREcxOUlIdL+MVJN3YUlZffehHHot1WTZ3qZtYg75KuY2nSblN0TkzPYxFOxw
qUpDY9WkGlZVbkQbJ26+mqFfvNVojm0354lQL6eP6HItuDfqyfv9IWbEMUbi8jouCIBAYs5ZySBi
Qt+r3b/4sK84zWIojKsBh8T6UwaQk1Nce6QrBrHZhJ4fNGc6sM4zVTD1Mb1HC2ca5gAh2EcUB+Jz
qksVC4yh3yk+Jl0Ciq7sHdV5CALNR+cZYSp+LRik7BCf/6bhY7ZEPkKjOJhEkF5t73+Lya7udh2g
tnieNmc8UFngh4Ala9fsYn+1E8aPfGckjJ/INJZvK3ykCVeUnsizx6iYXY4C1bki0ceiTjddnijD
4A+rZLk1n/6ATqI46/EweshwFmyt0jge26MU0EAkRiP40Vdb8BOAHUP2puwuMLEha+FAuiWDRVlS
afmJv0WtCHfRFLmHm7xTNu5uEUlU1XSG87MClLzQjKUoValnZUDafLNUX4lV0prXAAkRdaqq2mNy
PuiBgfI6X+RjcXUISgkpEiFqX9TEop98AsXYNmkwtPtpJEarRK9tLqaf4hyB8ECdIRWAXPyRoGw6
jUVfSxVxwZiKB7i4A0zKP94YABs7FITTOqVsjRsVeZjULThQl74yfMibBHyAJDapF8NCTNj4BHbE
bpQQjygOzbzr8y+D4eW2TtNzVX5h7wE25Kft8o0XUIS9QwsNgZkdrr0HGOTDBvkwTtLyAjJIcfyX
CFOXC9DSIkw6J+SZI2ADtwBjfRdZSKIaRy6wDd1ekpDzKkyJBL1lMAnnC1ObSZf2mxsoiGX2j2Qo
ChxuQZGRsFapO5QOc1b3hHDT5IM22QT84M0fbsKF4wZOCR2AiS+iXLtVeXyFMGBRGhu/KWBLW8mw
yXM09fi5u2kzub/ve42dMwUESHF1v8FmYg3gnv2ooPhDN27e9JtcSA38JOA1I+7Tj1WwfwLAzONv
Tfq29YDGZgJJIoYnouxxO2u0E2GG8cppEq+0Wd109JaK7jNGOHckHnxMDnxiIFKtAdKFnAQ0Yzw3
a/IbuwM+1ZWiDyNBMwiAjLvQxxia+yjZDFr1x+Xf5x5fJM/BGgnp/ITfSiXD4bwdIoBMTRZCkeN7
VZTvE21MHH4ZQD9iqWEvHXM2La29d9xESY0kSzt1WXwHVIXffS/7VeKAxZhlJCOtClZmMS2GG7uQ
pStYS9Gx7LhRKtYr9bnQsPiz5rAPNMJRMUYC1CfwFyAacmDLGUTAKf06q8EsDLbDUzk360oilUAV
T2kWo9aebW9zrKg/YCJ3zRuHoty6UPKMCsUFtpjZgeSzzrmVJ3/LuGeMElInr98pGpne2hk6iyoG
fOMYaKoYFQIlF/jm5JTY8eqNxg3QxpBmttjmu3WEyxj9folvWvXiETS6LY54A+bsKpmyDHznwe/2
xNLfhurYiLBazZtcuRBLc2tgy1TCskLrVLdepvMr1copDgAR1t/gu/PbEZDZ6zzMfDsuujlgBuBF
gN0e0EGayxkUQzrRo4udq9w3cl6DWwiRT+Z7TzfTWzp8WbJYwCCrnAqN24qPohVv8ClYhaEK2/tZ
SJQDIXxkxz947zaBdFh0L0VXZ1RujazWy10pe48ymE+8cZlNwljLTmwSRpd6TCipF7QaKKaQ2l6z
aUGh/q9r+fEIaHVdRzMtBxBu4/hIL243RtPHASJZIVxiXxUu3OSjEmTOJa6E9rOkfGxZgxERxZUS
NKGv3/JIbL+qj8MRIqtD3mfMv6jRQrjJ16t1HazYNTKon6GwvQ2w1Ueh6hLl/9EI/zkOribYuKL6
jcagJ8MF146Yg/B0v3GwttndLlRC/tybIwAnOpLlM+i9hRTgxvbTHyUgUwF5MRqIYc0T3D104XDh
GLaDx/aQm8fHAdEGYGvDiVqbGNvo0FcGn/pmNEydro+FPodnya3bsYnXcD34Eptl4r58WbbIynfF
Mex/T+agW8dbqJag/u/e6tBvYI1sQG17LCTzgm+Fvlm8507LAFlLBOT7WBBTvGOsjBA8TqgZ2nbE
Gos9jeU9vGaURtcRvQOS5WSzYwL7TkD723Qv/HePdWdI/g0FmboBDZ5p5NhkG01L04Wb5wag0KTU
3XHm5lfnWD7bVTEZbj38uipzapvXM3nxoJZy6EeKyZlnmaJxVsKJMgHxorkpav3WoXbKlfQ263fm
tVvTgoG6zolZdxkiecjgueRWcF72cA8uVkHNI2EaWpAAXAvvrCB4P9C5vec2BJYKii9rEap0Is2K
kKSnkBDwPFidbNtdoAnEplMop/0pLjwbCj8LGxPtZuUs/lhTX2vxcCQmBklw3Z05jG7MsCkZPnnv
S+3Jae5/SFBcVFhOa5BuxbQ/Bt6k6vXgK4Y+MetIkjIvj1p3du6RvwMY6KYgneqEvu+XsXZ7qOAN
EAtmkMRQBbAU+5qYGYwLYO33Mb4tMYpDwirS/J6tXxLNfW0x1C7Q/eec6zVPhBKsqRMtKwF8IPhk
smG8bPa7DqMeLpQnBJhji8BUCaNTamqRHPLeUEOYs8wEBeibGxKnKB3FHCe9bNh8cpZSeqMaViGb
5Lriete877EeH+fBJinpW6lYQqZ1lMj+HdyOjyBcblKYNUEC2+XPSLe6R9qBqAQ0FBEoNh7VliHM
KjnSCXIEJ+3dDKGGKLX369DH8DCRQiyUs2WUM7+iI/O0wxL3tlQ391pzCFIVxCXVHYGOQFlTnNoK
0rmCpFZ7aKm+ESZmcAd+G4uqypxdl8n2DCvqN7CtfBV7kL7UR7MG4Dt9hXp/MES8HdFFTxkLRswQ
YL9Y2KawP+0KkSZXlX3DfZnFmmeYuGBqgDIApazuRMdldye1uwVOEv498C6NBZpq4vDLqXnSYTjW
lNBHp+DiMy2y/FBFHAaocaBIU7V/d0AV/LVveztlZcQzTZ9sNyO2c/i44h848Z8dUEZ8o5Sdo544
OjMEpxL0zSSvYoaz7oo6kDFjH9AoHp+7lmdjEMinhrlaBm3FmxPxjHB23jYiSwZ5S7Pg3tEtK1y0
cY1HzyfszkC7435tXk1zOZs/jutf9bOTpztSfebKz+AepD+n/2b2c57WDloDo7muyCBoKTPRpHQe
/YMD5rCwX3zh2N+1NyZcVzSg94DcHn/SITHYpT8rbAetT3t5rO+u9RZ/v426S637tKwv9eM19w+y
HMAaTKXEHXhpuiJJSvdrETN7K6Of8TJBw29BlSWVqoDTVdeZ2/bSGDepI1WZE4F/Hs/wmKa9CvtZ
wOBFVA98dB+Ae+ZopCJzJe21gyLw6nzJji2mlmX5WyWqXFj01fYSL+ag2vAgzUGZ1IqA8RR9a/v8
fGC/ISlaeI26It0CJSpTm5zOuwCoS/+UCPQAgy/C6rYgqTjF87qiQvKLm6cLe11dF14tlKYxLYwp
WUgCz9s/sMYPwNahTwXqcQf6ssZeWC347FipnecdHP6uLJV9Lj2zdpALS6Wf1IM+qv6i2QOmQo3Q
KA1pLwRluGXIi4gzHK5Q3Bul00QKrF9TwmoHPm5iMq4TWq+yhyDuh7jc+r3TPZVlO0ywNB7DghdD
Z+bu6lpgCdUODYxCXattLSD4Rz9hbBwgb+qvZZM+zPnvOgcQkA2pwLV3bO+YXE75ETP/+Snvpeur
F6QCK0D9lqPVUm/rykO/+/S7NqNnuqxo7+VumSJi3DqX8Fwrm1ca9kQyzG76Dm12btQVRlmtiFuK
VlISULvMSRtl/L77KJ6nmvK0JCYgapuEfnyhkhVmtZq9j1/yvplLsRV3UAqz/TVQQvNo2iEGnu8h
rrcDzUIe+GU57DVjsh83B3fAoVoCD21pLPX8tC8rHQSl/tVfE/LARW8iM4RDP3DJcnicWkhR1B7P
QZjaRpHYMhqSExcwzVZEukNJzIf6eTYaH/yHTj426VEpalEsI+A1faeJeSZGgGOtkyIQgqcTfNw5
PnVXCZTxU+pVMIwfLjVSHgNbNo8lE6QLDWIby9+BjZtXZ0mlnFeJB6dqOxgk6YYL6381Dg7w9mLa
16Jgd9alcdF+h9OdCynfkyu7tFpIG/bTOzbyODpLjMD/C/WuYBfW+cnuf0FFYtvG6FKyeGupjQoL
RK4gNnitxU2fAhjYGAwG25j9S34U6j8gnAsg4NWLzfy8zQmSSnOdIrQo7uGAmDWUsVu/Jsf1j39w
8XjBevKIfSXsn2OyjT8QVlngewybDByRjpPYC1qDVFGi3j6l7mDyII4NGY2XruxSI8LKeF/sU/Qh
2Pbvg0DuTIRdSjeCOZg+6CaKk03kRFP4rIrVlCkiC/SkXNDawFGjMZofH5Q2GSPVgTUOIdjY5wsJ
J+kty0crPtJjSLsevLugWE70xVtjVx4c8MMswdr2RG07QGXZtaoBTy3rPNaXThQqvOSsnqvYLOE+
K7BX49mTefI488FVLZA6R0l+jsvVeNH7+uf0Fd8iklYAy3/NsICvNXChdoZD13zojBhJ9SN44s5l
Byx9i+ocZ2sEC17DIOeNtPaUYRWwmVG+TkGy+VLq+qFjNuKy/hmrh2kHavePN1ideZAo1DZu2YxT
HU0UxJEScodBpbyZtG0ufKroI+2bWT12O5SvmDbuxo5xAL6BwPwBtOJa1mbhUJ6+tQICUvpzguop
P9pOOz7+2GM0lW/05bOjdud4JvJy7hL0LBt1+rOdYZNRQIEGvaj9c1jn3SXqX8dbQV8fOJiN4Sui
B+iV1pmldwIyf3wZw1iCHmaB1Gq3oTdhjqgMvMDg14lgLYZ1leqwtAAlt2Rk0119yz05HT4DuTIs
3q1yVitRsnX7mw+ZHf33Kb4Ui8Pelu1WsG0iVVwtoNWpTIvKrWWf+QRV3u+QiVdgCPCVfvEPhwyl
c1RetaAjJU2wuAC2ZcqjGjTu377Cp+IS2yTGP9U15FzTtwn1i1gyjJ8pftmyOC3KDbZEMoMlyNRQ
kiNeoCChnvO5VPUp9/okuJaWcd/PBPzYwzGe7MKR51B97AbGY1KXU9vl15Ioh5Ww5mAfZ0lMbKSS
8AIEoeB6BYRCJxPG6NP4k7/U16poJ8eI/+gCF9nJ3s2U856jsCThPW0tF96oHlIJEhbzn4d6BHPt
SjrlxqWaXcS0PLB/7S5m9HKnFCbBKoemcrOphNecTnOZ6U7xHK+9mqKvf6T96q4nnIC9NaYnJEZk
bz35zRnYqWmsGu/Jquvnl+JOLKTv1QQfE/LxeZxwZibHkVeRrPNLoI4tVcYJrst8nAVh6WdnJN9R
NUvVYIWImtJ4ap0/oAZOeaoNYqxnr3I1PAJfwckJJNGdOMZPyIWDTlNiz7Qm6FlURJMcmQzEZBHW
5A7ZspQet5phYf4gxlTIQwhSh3hj4aDNJWPf+uch4lNl3//KtV1GP6Gv6qORw0mJn+lL/NkRzLh9
8xg8CaUV2c4DH4htam2sXJ0RARADG9QIzJ9L6F99ld2jVw+RddzLKALiGqrVD/AN6fPzgy9XwI7C
8ThSRN8U2PRICZWLgjCl5OQat0c2DzFo2IQBMJ+Yt5u4Om+RC5pVrR1bApFk4OvJPctnJzofuPDj
eU2z1ivnjKKfRzznLGauOVBN4bIX0+s10+TAwT7lGVaVoEnakUTmgRk15/hb4LT1Lg9wsP9TwBHk
ys4fepH9KkwjyakgES0H7jnnRBJss6hSD00y2sQkljNAj3TY6jqj2D3L+/4aamzGE3n/BgQjaSol
b5/Cmm0FOo/yHickQgtrl9qz0Afvp7EXXoXLcxVEkxac8DJfq8qQFIR6q83NscCq3qCW3FeWDwzc
c13J5N3+hELKX1SYR7cnFMGyd0xEbZIA+ddV0tGbhsYcjoVvQdWwzKLnVB03QzmI/Zvz82gIpJwv
IOcidjmVX+/cu2h1Ca+TbfHuAUuoTl6vnChp1VyXdcAwtD5hWDtFBIdnId6w0tChOoVDbSALbmyT
jwUeZfTGCiMu85SbWufROwpM6NSIcwF1x1JzksGjEzhSfaBUOESIDYARmocdEyAXaG+6/xIJdnnY
eaNL3cM06yIzUb4MiVlU6OSGacywvppzktgqiv08sa3jtoll0GOAUz0Zz8126MKZir8zuBS9KKFp
g0nhDKrQNZJgC2cWkRH6HCZDz7uVgJcGIiPFyy0uZOP3XXIgT3RzcC/FdRj4jzC/7B3YitTA+HI0
DbWkk97JcAlNA3t8hZ9j9CAmI2NPGW4wSJ3eT22sHsFrVYXz0Ysp6dae0HUMNKh5TlCpSaxHaJwp
qcXenhFEUdMOlj0SM6k4ln5X7Tx1WVqv7deRBXzYmfbxT5BhKgno4TGoZB2vwbpdBk2iyn+kN1hu
Cx40lzRW1mSeDq0pnAzeTFXKgzTlANAzgdxi57nLSYFgceHBL85Sb6QzQig9r2AjvEmTfbLKIVBh
DhuyOVOvfNSpCb6AY5zTh9hRrIvC2A2yMH9PXYMIm5KUW2FC7Uv2X+hVstCFWalGUsUxsEq+XDer
Q9073zfRLwfAYlL27AlQT+VaFCGuge1bOw2eOJYaDFGxr97ykju5iBLfnD40bRXOeTRZE2qUHfTy
gj4BruuItSb7Y8Dh2yfGpnw06V7LHGKxGIuTuEW5JIhCyaVOpZDQ13Q7MT3CU2Td1NEeXYI3y7Qk
A9vBoczxGOP6H2qpmresnLXEJzL6DqkmhZAloTYPDDcrSnYjNEt4fBcm7xScdoCYEs7Pl18V18md
P5Qo1YYSzaJLb7dUlPzZ86YlSWh9JhZVWiPTTdGD0ugQSGYI32TxBnwZpQta9vRXCJmmW7pNuTt7
OrAK3MzBhuTJrbvSeFc3K6fyYQ2+XSBW6aaP7lKJPihbqMd7js42ahjp9mbSsPkDdT+V7dF0i38u
jLWsgAYq+rsMcFXQwRck5Quou2x4an/t2xJynKSWIcstm7COD446isLpN1mrHU4Wc8cBX2Le+pvf
5Mg2IlLc80nvurtRPv3R4FVd6av4ckkBIdNLQ45N1AnlViWSidxnXolmDAfKLWQxPovT4GVtCUSL
7nJaIJZH0kwZKilhReARNvPj6ym1AXYqtBaO68bgO1FgTJpmtgSBfGgVqw5if7GLGw3HQln3k0+c
WM8cEITf3qxDEgDVVCc3e3xZbR1Fp11RUgH4ZIXGTzTZ58DdjVxUFD+DpiewG8Ceo028JkjC3uRK
T3ySb0zvbTDnFCktdrvfSTOJuF34tGlIFnHq5TgHan+g9bg5kzCgHA6ulgDvL1pFPU7j75oKtfkI
C0Nd6LWMEqPgPpUuMVus6Q68r5kMwBqp8LjD13FeBXLmIYZcjAafHdZl5HqRHirESwbRHbE7hzJQ
JiofG+MPNGnuZWPSCJaNixjHujhhs1Ap+VrgtTigsbPL0X4aYkOCL5Qp3EdrTd3ac+cQ1vRHj+CR
mci9bs5CC+1BgrrkcaBZo7mOWAWy0/jDwwF+gJ5GoS51bbpCprXdPKY77vTNmFms57EsseqA05r2
VaqxFVhebsYo7WM4dvvLtVVUCRtBt4djaymnt+WsMiYyQYBJEGwCIUJG7k/c4KTXTccdvLOjJ+WV
43wcg4dVNjgZw2js5w07gxrs30PzVIuD2hJU9wcWW4gA0nG3DH3dtMHg6YS/V6s89r7mvlD1tXoD
7xImfFKDFdWKuDuRUUXec072btbKUq0cgoDvcwYpJvgkmMayk7WO4p7Wu5ADvlxfU7DBiClnWpS8
ZQ0qL9b58FUvwpOdSoo5KIN+8Yf1c9A4PJM4CW7Q0Y3z4Z6vin3Axq9l1bjttbs4sBLdZM2SrbiK
D18h0g5vsZ4yBf96fxuOR697H6UEIxRjvpfGuMBU+UANo1O6s9NTG0PXMHoi049X35i/yVcVMzST
tjt8ASZe4R0uz9k9eQ6ksVDdOhZAmfVZ0a4t8y7MJLHNOh6hMrwyVOCg57HFizibVVz3VcI7RdWt
sDR+rMHtSd9ZPrmvOxsuSRewaGTd+i/QPS3mHJVVb8XEn/RClLOwu7iuqKd92dQ/RXCpg1m5K9MK
vycktVCt8nIVMTssvLga/PBPtO352/kLKfMsXy0aVrStmbUSF8fTetagMl1lJDo9FAMO/MUoWRzX
MTcxFIsHhWa+kxRCvzzTz7DabXkaSLuBtiTFhkj/VyU3U0+EYHx9usroX0xRUi+9SuTLsgI67IG7
UJqFECRoz8O1vn5Wa6+gxP8mauk9fLJFJjiZ2jBIdbRMWnnjtACsj3rNyOoXnB/XV+HYFSiO40kq
N2VrrcvmM700w2LKl0p6z6Hurq2kfuuJLjaopHYbY/KFb47G4z2gT1E9O8uRBFC3REAtKbfC1nL3
heOehvvUCV1t7xcronDhX7W1DVk8uaZ440hJmyyAa7i+z3BzvJGUMqlbz/sKhEeLhEKiT14psluM
Erot6ldBShVN0KpIVc70hLKxmC8d2C/IFj/MX6Ufis445Iw8PGS4Pd6pQE/WrLz6MiVKwHBNTGBT
EeXtZgEI7Aq4PZOUMC4dej2+29oIwCIVUyK7VXbAnZWKouabpPt89wdwWoltSdaEELI3NJzxFq0V
Mc7ip34VafSELmBnTHDJF8FhJU0nSYA3YmD9Cgfnwg7kdUegQWarNAcwCNevfqL9VadvYUTRqPhZ
CojaF9Zvby51LH1GhQ+3wUoedQbtCNci6YeUqjlt7inNPMmuz5iHQijr9APushR18CPqu75twXsT
ETUIx680orbRYgFHqrtB8cjhnZDDITyVoBhV5BSwHepv3Ff/O6utpzosFjOX1cvqCpILHxUZxIGn
2xfcZqXZM1Z75OHn/gunNJcZWXvP7pRAymKWo4Ir9Fah2PuqqHq6/mgcDyN4aitCiSVF+hCb7P7r
mNZBHnwWpHbLtSaFN6PE6+7+jAJPzfAidcbMvcaeV8B3b0T4gP5IecnlagfIb2Qg3m1lHiCBAtzE
4L4BQxc4kofJahd/Ciw7l7AMmuURY5pktf3vwwBnW0rT4M20ztxcaDjTEj0we3FWr5Z+XWaJlzdt
NPRmTRn3azk/67o0JSirvmQWj9zRs1E8cUfuDhkj1rEIZruFtu+KXElQUUk7UQAPHh3ks6fodWr6
j62tFzFcHAIqq7Epubhwa5EPzCfuR3Jhu+2qgAXBi4a3ZRq3D+7AKsGwWatF09+8X8/7qpIjiUlI
+S37eREDuyLTkZTJoA8DGMmbGEpSbyGN8HOxJ8m18UcyQkYjjWN6YFK9Zr5yJ4lOHGsjzpuiYwEM
tBMgnuAJgxQUPAXiyR5yVqiVkCp4eRYXCJprse2Y4hE0VJxePwy9vuakETksoRtqOdvSJV8MO5Gz
IReJQ5PTx2BIPeyVRkXGxBcP4ikPxA7/Fnhjq1Ds8Jv2UISuzrgXT+Md8YUyvahSPQQe2hXk24go
dF3pKYfHrmeMuny+llRz5sVJ5Cg9CtCnj/8PE7CJB3kGwwG57mvZEnLhaT2GwMrUq5VvxXfoP1ab
wCCMCkSYukeyXEMapJK+Xf5hi95LUCZxuu1R/3vjtLMRn7Bp0A2ljumRDBzanDqgc6EMKbQGK9tw
eNzEycfrIXc6E0DCt1G7zPZg0CTVMoHxYu6e5HqLQ5uz5YLUk7sVL4VTgoRJ1HkuaYwPDL0gwpu+
7TYpr7Px14usVxUHN6aWp+TF7he9nrRZGEoY1luf+96dq7YToHvQTXrEiPy5F/nNdz426oEw+gsg
hr78HjZjHny70wEHiquHfaNVyzqaCf9nZUVs+RC/5q4bxCzDjtf1/1kBrjcYinZiHJOhhUWm8GTy
c5FtbRT0OrK1vcNO0QDzt6vysu3JqZMu82w17mhlBLCwNRW+pjvrSGddLFPTf4sdTX4BafzRAWh7
i89qEqncigUMUB4y4XG4Q01GVHLYX+MuKWJicS9OQ/+ZlYvD8+9clJeRy74IgDRPvGDZ04qNnFh8
MDeIcMDhecPqgqZ0bzN5JJXIRoZ+mpWxauQwdc0TGuYh4f+3+TyBI+U9tD2fOGv/Ma35DWtpIHvs
vvzOr3tzx1wsu5lhZOkhedhfecN9B1bW5CEO3QJ/wMPKbJNXfjB3q27Ka6mcEgGOEQRx0V6Y1uU1
Rfw1hl6ymLEx32mlghp+kD1yAZJ9j5qq6vt03QanGuEFpn0mSwsk8CVBHvanqqr0vThIZCzFP/jM
tDjppBeEpRmLp2Otz74K86uRChps6EuPMLajibSh775R/rbsQeMx7Y/HkIAFj94EgQ2Ky25Q0DxN
YTjPtPgX8WWxXLRVxPkYJfbnFJMHcajQoYaj0ir/9HW4F98ig57gSyVKI3WRF2PXHAiz197NL9U1
c9in2ZXatGmhdNs1ZHvogTHlEm7hLVaWlahVrHN9bLzXw1OQjAZA8Ep1KGiryvpNZmUle+oonpCj
Vfai8a0BuaeA452qOYEral3FFeLilbsCc27l2ldDvYKp+MrWomLgGOccIlGOItShrOYUaYIhjMRQ
rv6TXrCDF/FsaYsV9kPAVG2icrpnLO0l0XmFvAGn91ZJsQuM25fktwsB1rcVp/mo/UibplpVWB0d
ivb4wpkCQ0hpLDU4YH5Zkd8pyRsIwr8Ufe2aDGDLwVWdEyA0vryDRrM2BfyDzRiTbhOPQPO7Kmx+
we46WFH9eReP2LoVsypSOWY0Rl0oOn+EJI70Zoj+zmV833/n2aTAT//vjEs4IRHILVRrIrMTd31r
g5V5AQaF77R/rR1I/HZ6Hf8xGCJgyFa4csUnNWLBU0wI338Ibmi7ftsakUqOjwHkiz1UsBXICWyQ
BGCD18+4htZYKDl6hqBQLIHtsqJn35CV/aQCASXyFFC7u/ACOyzfM3gv8YrqUvDUv9sa1n/8dYE4
Aci9EWr0Nr1Drm2jMyXT6Mxvc9loIrCSJwxa5zNDqIN81fvCRYYGhawOMqSwc3U6VyGFoB3OZMQ0
MYn7zdEoYCQBgoQPQJnMMAu1/b/Ma5LQvubaV/kcztD5/ZGRkGqkadRNqp+p5ZxvmGfSL+oPtrBB
IVFHtzdK1gqsdtj+jyHKXQaPPdDGXfwdsddmOTVkfcfeFaVgKEKJ0DURKFMWv7rqAz4YIj6o11D5
6VYK0OakuplCGH/6HhMBhFoAOYkd/hB7MQBHn0tg9s+dxfCKd5trqkpLXY34tCjpo8UMfsKw9INf
NrX5CbOElPIulS7TxYRLDPQatPju6KFJ5gKx9FA5j/6O0mhcp76EEaN7Yg5QSPvSqH0nZogGi4jY
INdJfBfhRTuwDVdsZdHtWefxDfaNBTrWwQgzTHYO7GfrmgNu+1ksPgFz8LXm2NskiwMvaihRtRGl
Zjhb8nGE2EyvK9HvCWBi5TykxMUa7h1RUYaTxKQQheDMHiL29/ll/9NNC2Ibo4slQvTHbZABvZP9
oAfcoY6a6xahlMoj2RXOcWbyGsHYbb2F+2SK9D18Z1v6l/yB4x7ie5iMFUcV9GO9dVU1hVEuFbgQ
1J8UAp4wMsNOOZbjOb4rborhqOf/3kh2rNt9PWDq0unY82xz2ItfXEL8WWL0Sb5ug6yQN7kS/jGb
vP1mxrBBKuyHfTJxXa0HBC0fy2H1HmffA1PtWXpFU+KW7md/cnvqaJgnpPhshlN4Q552haCQMDBL
laV1S9+oswU2ox/CgLUOidq+wea9Y+ddpEfRLQCyq/D1prSbimVXsrNg6EsEoBMGrJQyeQjth5Tv
WYneZYPv7jHGIXjtRLIbmT5Y1HaSCYsQxWHKkTG4UmkUoRF8JP7PqLkc7sNenMGuwps9Ul0AuZRE
4FWXUTbB0SYLTf8z2PLKy5bsoA8jz4QTv2ZSzGi+kOeQodE59lAuwZLv+Ax1r9+8zaXjFhmtoVNV
ygkNkV7+NXEIBh5V74ke9rNwlWdJm7968KmzO2WNxOflu3IvDQlUOwCR521Uup7j2v/Pa4J5dIHU
H3q3ZnO5zXZFfYvPXO7F2FZvnKxCrQV2IyHU7vOVIqu1982c/cHYVb+vNExsLN8sAZrLKwSJ8Xhh
pQAqL438gr5Ab1XkZGxdMakviaLw1bE0MaCZhYJVxgb6Arn7WTGi6yhqfP9lgR/qN5IgVInaxk8V
pkEEvKOvRlLPdqojrw97IyYQ0aLgP8Sl3HfaKgqd+ls0Dk1/KbmOqQauwcKKNQWKyQxjC73lnryK
fYszKBrTPUpXi2XnbrEk/BeyCogbhGVj0QR8YfPwGUJHOMeHn16WcgHm0XlLdOeh1h9PFs+Pt8Nj
qhzMzj/pGs0BJIGDFnKtN6MOetGv2hze+O1LYy0zUTJQB4h252XsnV+x8hlTL0YAlG0ZcwcdGOWr
TwE+hI1Ff1ZZJ2sMGsujgw9GcefbbIGTDy2FW/OPFhpiuOfXOkqOAOiNBSXhB3jnIpKJaR5Xs3rV
vYl/qG6juSdMLqiEAZMikBd+Escq5KzEuJbS4oj/7p2+QPUL7KGmy8laJtvINxv8PWO2nY24WHAc
bUkzOlWe9WcvsUGWjZ9HUizzCtCWiN5Ic5ehgd4ZKDyMf75Gq9uIRkKNkq4yiHD/nu4bL+IN6P9B
TCwMXkr38MEU6YAZV4mfDtqiJB9XWYtXqEYOu0JDacysMX3untPDTBk4gpPYwwK404MsyvqiQsir
M8H72ObeX+4HfoN/j7cFgC4sxspKXCQzMHOAcyyrEfOjVhcqiOFD6HPyUiXiA2/5RCwjU1bCxVBj
cuLu2y1q2DctW5Rz/NGd8EPU+Yf/kRiGkHwVzstcVOYkpeCTMuQiLADBl8V70NWSZCEo+tOJ8606
D/0W9Zvw2w6+6jSrKwCtWXVjYT6o6pDEcIb62w6iYDsCiAdbUS3InFwFS7+iz6gz/XHWLmeLtxJt
EIJUEkpM4TyP1veTdmNbvkVuwuLrOiATQvPssRz7FB1OZBydFGj5Tkz7UXzsdbSJIZrZCpk45dvY
jto3zo3wX9fzJvkWjxBjqQ4FfzDl6c5xInmvyQ8U10Xs1kxdObpyScidnPlEZufwuM5F9otaJPzP
ZpsBNfg/UKId70aj6YAfDI38lEu3iZxI+XX8rlK9BjJ4TVHk5mOFTDyBg7j41ny90V65WI6rRbnS
mx0Bo+KKPaRpYesIa4/IPhhfRtr+aRMzO82zEXn+EKnUrdjLJSabXW09nIDFVn7ApYyNHaYEwBlY
5l4svqXTMrw1cmdB/lQVXomF48z6DCK0JIU7ma295FECvlwCrSWhI/GfR2Mo1BcNrOj3eJMDr2fd
Qj/Z8i++NQLSwpuqnWD/yI4fszbOsyBQ3xAhU1d+JPLn5hpZaDx4OLNTf2hxtWVheAncFG5o2wne
cm91EBm+3ePCUTZDm6ii3iMcRgNIt8AJVi7yXDZWXwPxhfqZzZaqoC5I25PzKIpI5tjpqWqFcnzR
pCFAi3KpNtxYe8uvY1Yxo2ciP7R6D6GJs8A//27C2KZEVRhsAi+45EQ3fwbCgFBoAEqqafXdrCUr
s6YSxzL93T6Tmdrlkn7nF7PjRiUKZR3wXfeNTX34Eaa4Ix9BnR3l4j96QXk/4GtewLKEExOSSJZI
24PpXziHRaUiAX+HvXXwYO4XhLvmTeGJ4GtbiPk5XHA4irw9WJ5ObvTRqzC+Rd4KJJaZwEJ6wM5j
kbsnZCHIZY1RzJwEJzTdMTsho3/ewlSu0uutg8oZNUjHmy7/wrs0Z4T41VMmyI2GL93o7AzXmhCD
1QEU0iffCehcNAHUEgTuQfnSXjFPcy8cEID+Wz4CuZIttodS8ri9s7cuUstv3GCGxwPRLNgBbyJt
6coVVDoVmx+BQKADOVKULSoEvBbM5GdN0IKB3V1d5eoW8oxQdpjMTOwQHdDJ+reqD6HnZihxudE7
aKkTyhBDw4JbVM9UagXdFb45EP9U2BAFFdX90vLxPK0DjcXXEwR4xnqBCYllNaPrh/rBDihmmVMT
zqpkL4Og5kn0rDuO3W97wiEM9TRzVXoHc4ulEk6Yhs309KzSTIzgvKm/binSsx1xSJKsjOLf42FV
eVwBIlqng39iFaWgn42WtO2QaHI1lClSkmxI2z15peG71pGLicB2q3Knat8bqWAOVRQeX4XOAiPi
l3lOpmWsau1RIbmbIRBAQVrbM7XsexgUdu6g9BetRcEimjLkasGT0Q7HSacIC8sHx7nEoX2beqA3
ejCB3M1peckqXpvTioovOPJfh1zrffikyjDiHkBtlRS/QUA9/Ce8aGZ0SnlWlly43VYG39ny4kAu
RClCCV/r4XHmA9P5wZP/ZFOgd3hASrgbOvYqNrcAncf3vn3P+kLXRT6lKy19WaymFbnktEsmP0wq
G7TRlBQWlzCvEYorwS/ahsDXSWFkbKQYxm6bRWMokgRvZYssVn/jfSjyAJTT241J8ogD7w4nC36T
ugOxS7EFUFL8boTYpYazLsQM0QfXU80EzGi8ByobNwe2EyUnKwGisa2tPiPZaM/aCNvfgVSzIP00
yHFVhVQCadVBFQdqIhDJpz60aMuYpP3CS0oEWugin3//KeiBOHC6W6VAQjvQam28WXhCJPKaLC35
WUhGxxCLv7xxD/bRQ6Ce2vzLtSFztKYiTP3A4UAI/L5QTBsuda1YSrkMEJBGyITJ4kZmP/ETyyE8
XczQ1hyG7xGwuOOu8/w7JQjivlZOmfP/YndZT8LXQ0pGRHZPbcFUXrz8kaEA+CAApWh99qF97gpO
asK4afKWMfwu3twa1AqAGCPEFcf1lfXCgFT8tVuRQdzufHQRjroSaGCSUL6i5pe37lETocIrw7dL
Llenpd1fCAss/yF3lmu/9fw2ao608RfgptDzuJU9Z++e5VbUPLe7Hu3Ircnt1dRHe1kuC54l1WuS
jtABq9/1t0gRdbtGLew4YcZ0s/mr5WR95BBMIMsVX5BPlz25mb9S6i3YV49MtiVYWSjgLO4n09CC
mXcW2SzaeTyY8YjFUhlcEfZ5HZ3WepqKsbeUXmfVtQoTDJ6XmDR6idQeWAJu3JKxBbSijsW0WyLs
eXVyXbNmgaCdgrWRMdR0DNvFfNgXIg3Blb0qNDBPWUXxYuvSLcmOqhuDiR6svTlZU99E4Q0j8zeg
NgQ6LBpLfsOOMVJgHkqh+BdPhtxbCc6v9BYYs1pL0Qw7UwdcEHHLcwRanNRS0TA+8xu1eLDY/5ae
+28g3CyCRxSmID/pamjZBLy0nmg5kH6CxqNS2z1dgJ4sscV7W1Lcm04ozpnRO9PBiSb/F8/1HLBw
HTwgywVJB3g0dGt85NnBDza0j3k9qDGkXZIGxwk2v9DwecX5ZjMfTjU+ZuG8xaPGaggpO9gICyBQ
OI7s9Ldm7aaQ4qCn3Tuk6VL5ggBIamLbMcs6qLV/6Mx8PHyqpovavjRV7ad44bSlzDS7nnifc7v0
93tErxiSpnwOxlyLzOCEZM6Qp+IUEUmRsE9xMZA3PoP9/CqfmoF4q79H3QKlM9SKr1UmqZJ904TO
zDe6lDmToswk29IC2zFLcYVx90dmADR6ERcVyd4lSWWhcdh3FUibsn92Ej7WwbUrAjsCOJ7WvDHx
F7Ms2Jy7eHEavpoHYNQG/rDwOv6rHvq9t6/wa/7j8DhNGEICPmyH6yN7ubSPTiU89oxC//qBdoPV
N4StIVMFaaVgpqeUT2hyfdwHKKM0y+vNyzv8q2+RBBxblOT2RCxKyQkwilH/ImsTTdWPA5X7cxNJ
RmFZ3Jv3IrRlefevnW8Aj1puFrx6yTSFwCguzEb+uggwmg0aSbAs65JF6dtDenHC+2pAAGB32Sfz
mGCGCfP265TUYzRzEOe2rqVxXBbjA/gnZptVutzn+HUVjAjpmGokq1Oock8BWaT2LI74h972nfQM
ST+UTQLr8Vg900C5onsal7f3u6Sy/V+03ZFcgNp4UvJt7AUhwOLKtZqe9i8H16816FD9dQO3vKYy
xH312pzx8plN1jHfHDEOIku6gc41Wd6Ghj/gSlleDBiWV3GH3GpQC659cZkp9coPtWGNrwlU24Oe
1EfkaIr7hIWqOkLnrPgXMEgRQ8Xazt/oQl822pDtFgdizm6a5e29/SVNkkkUxrWuLMu6BKka7FWR
oW8jygc7pOheJg+eO2+MhSWiJzOyVwd98e2SVTGFp4rA5Qx7g5MjBGfiTq4w1EhP5aLS6uAfakGG
x0bQTXdRBIVWpUrXoAYCqFgriajBgyU2mFqZD0fE8lB9hgG09UZnLSpIAcm7BUDYvxBFyuAt1Njg
8drW2QGvukSfqniFLp/pZKa82fM9Ot4coOoh3HrKddU8R34XaJ9ybBlazQ8EnWmuikq0V/7DL7GI
NqNHGhqLHlGCwQ8lDO5qb8S+U+f7Id1xJTqRchN2vNfCxCt8DwCQ6sJXZgzv4bDLYEAJbW/f4+IW
Tfbi7gfpmLGChnQ8yE31VfLT1cUK70RryZ82ceu0zET9rq6PfxloyTFrRpU0UDa4rZ5xdNOvQZM3
QI35wrFkuugODlQTD6Psa8OmfoKB7nPMIFoJHoQpwctkly3I5m8cSVs/Gcr2k+XUPwBdIiPZ7R6E
zqA30mQ+/h08iEYfX4gmcsl0Dalj+HKf2qOpzfoG+3X4206kkK3+i2J3SB1gjycE4rIW0t1PE7dt
QVo+/8hq+1Mr+edjhne2iqywANRiXf+Bwb8UocK3iwnUsHHe7y6w0WAPTKp/Qavgy6t1qRkWPiGN
rfPc/CzYm2iOH19ljj/i6DC2uOyYpDzKeDClh3mSX0vIcxLPC+pHTCFBTvtfzDu8gsyzWExrc0Wm
ycWca83aXtgzo/O3LeWCMGu4KmuE0wTbvlJQMiJvOrli8DClH7EcQDTixu13eYyUtcAYe982BX1G
Ivs/PiuABYpZNtwS7Y7+0dEWDaf/i02DdjnVvkJCIfERQ1N5pklH7GEf0NlfIqJkaHFcqZRSXfyw
8o+rhVgTt8ssrNkIMOV9h3pnfxZnznvg03OjrRJgbAvAlM2IFljKgKAjtOYRUuuLChtF927mlQ8A
LY1KPD4goDQP6Kj/5CzfyvE4PehonBZ0rrnpIq+BCkyzItV4vcktdoXZ2LpyOO/OtHC4FxaLUvKV
1ueYklVvlCHTOjMIv9/0LzvzRFrcBnlaB8ZdPn7AwlDnnveO5xn3oR+u4pAc4rxPuKhEdVGfgEeT
scvUdf1B7+4KFwRHfFZwdvBPdxZCalWAosNCA6hKeOvv3sgxQ2XGmWO1R1s08oZNFaToLPyObYjO
kCwRo33bekiZ6AdU4++08MfGRFK7pmdxOOWUA+IXTo5H9PaJ7p2cQ8Vkhyq0AQp9zEscmAjmlbs1
wNjUrNhJueta7JiVw8S/y/SMa9dFJnZtXqcqKFuCVekY/WYl82QOnV81h86a732lRkQ9KI7x/+05
9xKVChQSz/98KdR+6CXlNmNatISZYe0cbNzDZvQ855qf/AmV0HYr0CAiwTM3ZibMAH24I/Di1hvS
l0EzbZdmLIe1GKKFC+ZoIUyMs+ZDubpWrr1HDDTkZKlNTOwWJ2rmC2u2cYpzOKNepNOR+uykSZyJ
lYl0XP3cx6FHh5CcnOHsJzSOAzvwX/pa9Q0kU/KrmKOSwkEqXKPTTfSmJMPYtI4ZKRXemKZfQYVC
WP5c8CgAwbMoL73rDkOfTJW75vYaYlehCDt7LVQiuHsT4HqYH9nZfkC5E0IECrApRKKJ8HZWmrsc
PkDdYfQw0MYHKoTnv72xI1UKMjxOfSLsHT2VhEf7H5Y3l6XVv4FB6YjJtpHyQPIBvovULSHlL2Bi
w7L83ViQBtWnN3y9IRV6BILC/hA0X5VYIlGZyDvow5Ota7t8O5GHqr/gf/Nkln7lUrei36eQPQqO
EVzqO9m05IUiFiLjsX6h3ffZ2I8xPJdr3MW4hS8BV8V8f90VWA7SNxLFt9DqRCKNK1cEf6U9KW7o
T24Z0XNUY2CSpkHUfEQKbAV051FU1/RUZcKAOVwieIXrTV8FqPJXDJRwjAG5SSri1hWqnuVbfj83
brZcIT+4woyz+Pn+AdYHMDpp/j8NR6LBUN1JWkKRO7ryROc5IHK5qmI3h3rA9dHWwQJCEHIhkxD6
awAuiElBXXFHASk8PFeNMtN/9En2KsP2QVp/g8WDlAJVu+YuY1Bl4hRuzpuClBaQer0BoPuCbCu5
pR0FPGU1w16L5qRb8w6YXPSunt+ThpOIPXGsNJ0tD+fd1NmGDmGDE/E7IxcMf6mN9/WmK6rys1K5
AW8AaaPnyzR6obGh0AGP43m26S6EwR/uVCUgMbE/2GEEybWNbF86aQi4eda6s2SwwvyEbqiOQL9D
bj0YiB4oLgqCPFxwyu6h76q3gqEd/pvs3RWUAdo+0DJeFEF6+nBvzWxkwWSAgDpiJuRen3InlhDZ
BOhax1v//2uaiSabU0l4N7r+9bQXk1Bw6sGt/3XVBYy+QpYrvT+TRXyJVzTQBUnDONcJLbkZKe+d
NZJCdgfF2Y3UnWrQBR3vOMt0vaDEWlLlIqM9B5CrtojrVIeoryOAXO0CvBVKXbOsduVBfTBJqdZA
QaZ3CZRcQ2sc7+C4pjhygCMQuvOQv1Ti1WSaa516qVeR/oFFCcDBmtn6w1zARdwsPMQVZjpTS6ko
aZZSBhEv5cwtRNimq33zhIsNsumlBVLFa64N92RstVVjDJtvWK6vG04tRyDgRcD49fi8c7cIXjou
ufEY/ICGTGs8DnMMq+49G5S4+hl0Su4g3rm+bjg3ZP1ScJwpILyi/rg3gTduBpgKPQOM8n8wW7BI
TubUZ+PjLQnAdnVqlVVq3AUNBW/T3IOu9Ipa8B2YfgjLqX1igHw1kg6Eu3SOC3bQlD74PHI9dK5I
IPCtBskhdQ47OloJjcvk+U6RnzNgfEMJvAnqe5Fdj065A0OnlBDRXU5FF9rFUFEPsuvxc8vS9q/l
Gw/U6bkqp/gprERfZzHkFNWLaX4ugvHMf69PSJc9cdhU/3teGCmXmY4YLhzL1yl7o82fHu3lRAdW
Zr1dtXRp+ps+XyAa+3KCPC0BOwSmOtxqA5XJaJddDIbR7Mgs93iooqCtL+JaYpkrkq7y15PpQUKB
Gh5d7Iqy5BhXnV2QoVALijEUKo5GV6t/IOhsNFTToujvSGFERi/muPVmlVljRIQ0EiazJ1OpMK/w
W4D1BIYvD4u29J1EekaHBZWtQDg22EjPCi+km3GOMqzkOpBHatJGYWeKS+ikfPUmq8BWn2CAHCHq
G98Jzq0NjM59lo3gqc/p0FQej9uB/7BZs81WHHDbwCgOwMsUjKRghJbtXd2X0zzwb82KT7th9Pv1
vwt0Uyb3eyRyxba3T46aMF/3I7dj9WQ8wOCkbXDIyT0lJLi1U5zvQu3uCDbyuk5keCBqegjGsZLR
6UHXLCSJ2+h5O1YtfHJj8+cujVT5VNNHVuVSsgPo5gIMv/zjdyPE3/4VnquZ9femFdUWpYUqxJme
v/X1sgPI4AKWdxDPciaWqMyxkMyyU1Mg3OrHqEMHiHL9Uck1AKXluvOoiO4HDDQqO087PhUrbyt6
o08BSxj1dPQhA+ZC1cfYiibHzKvUt1G/KoLEVr48yy+1Wd7Zr5H5loZozJlS6XqWUUG+0px26wxg
e6j6oFgrrI1QgC83iqho8vHPTSFqF8W7OqGziSDxxDdPL63pc/CcKiuL9jAxN+krYiLYr1bU57lC
LyQwPs3KpQkEKDMsC2VIbu+rWOKCkeyiH081wkRvloWDTIO0/vWn9XTZTxlPnZkq45UEMNVodj5x
//hZIAuvyAW4SFKEme/vhbwEfWA2fQh0/VEEg+SKecGUaWVx1C1BLDUWYE4dthD5C/+FmyLxI3JU
gOCfhG/8LYH63/VdCMjQTvqp0IsCK/pgmYpAjMladn3IdAgusdszsh5HUrHzIyFl0SnRl90gjLsd
+nsiEkCwQqVEO05MzM3B3oBqwJtfXRYWVSfmophV89qvX/brGprkE36C7E8eiZOs4EuMAP2NB2s4
ZL+XXTGeM3ivE1ky9a4DnMjSF5Bu1Y3BjoWCH3fmFyHTT/9KkrmGtjUfrkbYPDtOLmryzcfmSHSW
VauPa5TES759BGcPi+hK1mYZNH8vZEM/x7P4rUMOIEJkkBOcJpheed2WV22r1AyBOI+FrnNNkYLV
xsxnRE6bFtwbBFyCMVKDMEG7QyMMlY4lJjEkO1eQUaSwHHpi3rotAUey7LdiK+w15ThHTfb6iuoz
6uMkix7hJCSylbCPoKjPc0qbrMhAjn6LqsL6Aa15fOFBJ63ZjVlIxxky6p9Y70ytZNWcbHGWyffe
jnN/LCjdHWnn0MmY6EIsYIIZm/THa5LSyTpssIbtXOHQqJ5UusQ+Vq57C3nlcWOdDdXhO2KWPPE1
rnTgkRAuG/gpzsR7WzBeLtnfgQyqN9N403hoxHqY78mosPMVa8DnrGtsI9wBZwzTFNCUpLDX+lxv
X7NsU88izptc7H08WaghqqWEJu7PN0/oaZxh0qinj4FIXlbq7OrnBUTdKrwkM7Lk116DGDrl9TcW
8GwF9qGViGJMvfBFu8VQ5w3v+mAywb6zzRe09Q87X7BsLbHXhBc0rZXDQJUCwM9ZoVXIuELeT2Ju
nIaF53j91qXkIVrS8WzDZrLeJOgvD1xLBltUeOtJM4UV3jR0IJndYJvyCsiBFwYV5Lz99nM+Rj9u
s114naHLt0PbI3yolex706EEQb6U494MthDkkUCHjnxIkcVEvN4u6LoZGlt6nR1PKsEYoqGn7dLi
dytdsXNNSLDxnOchuAxnNS1/S5mo+li/LRdxisOuH9iRX8djPkdYdbHc5QMt4SHnWXO14+Q1waly
M1Z1m3HA9YI55JlLLM3vPTXt1xmKHJdJjgUHpAP0Z8wI9RCF9UbUvaufb0OjnZM3NQazmyI5NGjP
ZWcJOifMIKU0XrNIpdfMVzjJbX0W+wG2PO9n4lzawYoSpL3stM++3z6RBcd2EFILV4fxL1E4vf4V
hDvkeJlXO7iptBrpFJ7DmSTiZEbwhCb9CUP0lXW9HfU2acWlHaViKrk3FBwFXeTr7j8+ICfouAuW
HYi6JPunwh8DMeLXvxDV0firvil0dEL8Ln6Ul1W/5oEe3dZ0CXNMKHeuyllJ841wtRMLMs0Nfzz7
PLbdTNbHudAJJMG+Ea6xOF5TuGxk6FnNGgbYYTQtBqLsamZf/5NuGOPk8EPRR8vqoogD1cikj7a9
QomDlaOFa6EH8WoT/+GOHA9MHHWG5Qmc6nswGnRcTc1/0KOq2qDjSnrHsf4kyRn04tD2ay4Y7Jof
j1Di9KG/EtIVGSNu5mBMOsNXNOXcnTSs1HSb93GP9/6xNx2RWc7ckzaufh3DqjO6s0menK88xqv0
SQgZ4JnozAn69K0vlcmSjX8LN38fSp1rHxxFY810jqztDWRjUjZFK7RkYxbeZdgLBbFdhWH2Sk7T
IFdwgMvc1Wph81cLZ3O9R3sxLwXlGeCkaEYUxjt+YLTNhKWACx7Csxl76zS2jxOYaAAB/CCK+Qrk
MlOx5tkP9GhHa0cMDF9aOLmAFm01ksU8lWjvbxfrSeYPBo1lgblRxFChNvLPxbWx7NVPPpHUjudp
t6dPrXjwfpqGQtjD8hZ2aBjUdaiGwTkyvP0fS66puN9dA8sI3TTGeupObpjj+Ic5pPoH/SuWXz75
NGVkOm3AyAnRzxdQhzksy2FxFaFqyjuYC7dJsNmaakz5NbojSBoKDwQyLtGpxJg+EnjlY87DPDdB
BEx2NkcwNCfyW0h3FMHDM/VsqCJAXHbCvXWfjCzHFEm8zBA4UWqVaBy1a00TbjTwY9F8u6qnUGtZ
2B7izOoCxXf8s3e3IiNKTSjL3157//t6S51rFvjIqTdN2jny+r1gCt/PRgeEoMkUBk6cbZHb2tvI
OlJBW/CJArnrI8+BNzB/OgAruNYeJz0JsMqfwaesTWVODclICRT4cJSIBpzjYcDSTd2gy7wdzMNo
gb9Cij8n5PehRp/YvwL5aCiWcRDmDDnFEejKYgFrkvXfyxeHhgQ5pbkgTNn4d4Wedz1+PZ7hndVe
1avzlAlmuxIRfiuhUUbIVWgKh5HEgkTx+PALMusHZk4QkuM1TJCXTwCCXr92lWbgNHcvzZJ5+WXc
yCHBY1h2rtlPpjiSj9ut2MaYIao69BUKk4trkpBXubXRSJ1DD5HN+3xHy7X+dJsmH5hD63xL5l6q
ZLyny5C2x0v3U0UTajThXq9fGG8qPJDKO5VQxBcCu2MCPwE5az3jHqaihQj3xBdRluGDZB+0ndck
cAAGhkszXyjwLF54NMm9OStWwBdsFrut0c8iL11CNFj7HspivG/igx+0jUpIAwMZsyTMHPwwMxVw
GJPtBWUQlkHtisJOG7MGXdUIJ6zpKLWbYpCsUyMol/LK5uSll5dpRvLfgcS0Kk1YQqFOp+FIwNwS
IWnrH1KMze/ZS1S3TscoNuw9B7dDXMKLM3U/hif+9lEynFHqb9WNKfhowXA+6l2+wtfh1KzrRLPM
VnmqpxAU6EQBX63VnoY3uHb9AQxIjVNmtNCu9aw9Ji6DV7kLjiXAFmlk839Dc5lE0USunt8VWVRE
0j4c/teo6atUfKNU/jE/XgqJLOxdnqYXBWh9+bqxr7Z1KVRUCOSYrkqhScKNJXeCKeT0n9eAkpz4
FQlPsdkjQ72cA0YtfpNVwqC9wxy/tH7jqngtTJPn/IZSNoMqwnOP7dAsqLYt3vT1Lnelcv4MOcsa
bGZwognGAmAqlK3l/wSYSmfi6PgnH9lEZ8ANM67RynedSS187FnbGseS0oafXK2kk6f9QuTDt4l1
X5BSW6Zy5KGF4VQHB1w8L+GTBbHCi4w6xdp5rl46BjNN9kin6Z35o3ea7fEtO6gZZaJb2F252vb7
MoWxRHGl5o350vYcGRnjuCuQiW8KGO7VptMopKZ0++GOsqV9f7pzLSToj6hA2d942KBw76wIBeMs
VI09xTpvhcxX99TtYrE0SzN+uF+W+U3YJohFEI6h1KK4APIhETc3NpDHKdQpjE0Oq96I3cUyr1uF
/l5plDT0rmP2Rxi9CclTqBUdEw8PA3D/zWUKHxXNi7zon7Lb1HaM3AUkUOgXd9UzeqLic+acWB8B
cpNiOT+52CSN+XznwsrfeAi5WlR9BObDDo9xHMj3a8J068SnzfKeQNoN5wpoSuGsXU9sPgimCpK7
kUK4PnG3E84axkOUj7kkYkCNAW4GyQdWj+gDQW5hlxcAh3+K25TzgQ3t8s0b6K6B118icEtc24Tm
eYSniBdGzZ4V10293NqqOb66FL0b7eyq+GJSnD0qqz7qkkJuL7B8bVncqZVa6+UWjBdG33eSy5G9
0PFulmhvncgp4xPiK4VgRpUgOihTCEm2KJv4O0dhsBfA71POGqqbOQRCRyI4K2uVBibYcNIWQ+dK
iRX1CfhKwpldQ1I0GkWa/CKS/IIbE6gI3lWYqDn1FswPBmspYmXqTL1WxyVT8kGH2aRWob1LxUhw
PqwW6KAPckIhFpPgn2QTwt2AnZIMQACwFBagyYjdNvN2tos5sh7rx3fWiIWQLIrwFvLSAAJf3IqJ
nhGPhqrd4Hef8vSNYQNuW5QwhvjsFgj/RtXlXwTRobEiT7JdUgl/JsliomBeqK9qf/8PM4rVH1hV
iKTLK6pNPP8e4u8qLUHpiCdnw7mbhruSMsBScuv8kC8iMl0W1MREzEg4Llf02mJbTRd4jyNscApi
Q39GkskdbMFwTcoOheC37d5ulxiO+GvJeg3s+ZJtmJUunJ2879YsaTzX5s4MhL7HvtPkqrITEs3L
KeyxkjIJlf/MXdm+18NjQ+HdBapu4/4pzMNEiHCRJzBV+f56+sbzUHoozYq0Zfq9A0UavPcpD9mU
0s4WIUVrfFjjgR7ZkHsqL2OHu8bRFxjepUMnkZNtLEOzhZleE5y8jKLpFjLghUdBbrm3BwTiIIOa
2g4ZQq6bzPRwWLunLMsjYjB8H+u/YXuC5DTkBH5KDiVMk5hmKFM/ZbPncKCooit3b8ZMFeJxYWz+
RU4n/GwwdvcO2g8ylcUuA16qg7C9gpY09IBCzc+ocR5OFfCW0hqb53SKRBe1ML1YeacCvkQEEg/W
8z9GRypyKo8k4SsMEtDywl9rjYjihR7UE14Qio7yvmZb3YQSXrNy9gZBEHw770EoYtfUnHP5JOjp
AHBAVMzawBBVB6/ZlzF55SgZtP1KCDLmkH/sekxnmSc4ecMjL7dpVCnZqIyQRf2+uIUWGmHFokpb
o3HBuw3yjPOR43RFEeJKrdPosPxBK2ZmX5dhBKa86msTB+2WTuhjfzhbO1+EXWVhXYuWc5gFSe4r
p7yvSNqVDEQSa/TWTDWfTVZPB58Nciwll432+K8a2Vc6osRFNbII9lGIUn9g36OkkDk88j2orJcI
j+OWVDzqnBYx+wdi+gajtc8aZpQR8PaB05io0ZhDemG/JLAr02CFN3a+RqGGUEJqcdTNx4AFLqqV
g9/VtC/lUg4t5kyTKrbL+kO1GXnm9sFJPn3NZjPRcGnU7pa8RtGustf7qVGcetqNPtQBuVDlPZ+r
Wlz/eGAcAnYW7D3/msLkMor9hCVpOe4rB17ZjasJQ9ZxYZOhJkoOFohbuHjvLZ8V4Wmj5539FEJZ
PMdpzBB2Dx4m51dfD5oIq3v8IbbG2vzLnC0AoX6GlSMu8xQxDKza0SATMZqe2vBXulnA9vWaER4C
47YsH0FW3U8ZdIJZF1wJVdIdAmsWmdZ/ycAZlBoBIr9qCpdtB9vyXUYZamoRdI7gz2yGy7SsXeRY
2YEZZXeyrx0Zm5LVp5AIM8gZyEIOZ5+twbq3P0kBZj5X/dAtH1CLK8TozH5U1fZVM9c6YyaiwCqK
hETNERp4kmDsAthUMTWLGd7ozv3l0QzpPCQXe9YOw6/nigX4KcTMEjv70QTjOaUmMC0x5zlHN2Cr
0wpTrGqz5I8+J2wJtfngtJ+EG7JBZcyehne0j0snqfrfHeYuZ2Z7lCgNbHUa0clFBx93JiaPTnSK
hcga1to+ChkmMM90pe1dXvYJxnwtldzd2tI/d3uMwDJvzUOnLfTbKKluLTULtPxvJORoqcdo3rFi
kARTSPMFGKS0jmeE9aSJu99k80GTCSAF2hcE2Tyl6om6vxArdm1XdkCRbctciz2oQ1texFgEwOy0
v8qju/Myk8WIieyx/wp/A5mThEX0HD9J+EvryUjZ++2o73M+s7HpkBYZkS0F431ymWaOn7rrzwqN
YGavXoyJU41qOHNj/lTIAcwSHareUjjPZWxUq1+xFRkBA7EKor5DGDwaVHGisd3D8Gd0NevTRBaI
qTIbjWadR4E3nZf4WkEi9GPTfXz6MB9/KVnN2ZUp1hb7UNkI43LK+GEh/cHx57XMxu44lsdjyr+D
e7VdxrcV/+yag1DgSEU965bbIOVEWbbuLIfXhRA5MSNX0xrmwG1t/naYw18SiYhWAgoKxvulzsiP
KMjAahShzGRo6fv0SMKwfy0F1pSR4J6iYjlwuXUp7rZhbfqJV64FBlYlxPt0vEzQG2udHxYiKdQK
GUlJnPadGsmZ7xP+7WOF45+sqyZ8XWvrIPrizi1QgDlC5XhvBhM5Z2kkBEQ1sudUiUMf2+jl3zIx
VRPzXF569yrXgOnrc0v3rDEBaPvRgu0xlJYod/72KbNaa8R4gZDuAu/UargVXs1iQR024RwO9dLu
dCUCD8FjwafOV6ilYZQde09X9pvvBSuIxjla37B7+Pa6jf5hMeBPJEg0aOaLuLE+TFoI0ToVUOas
gXOuO7e81nVBnNlKur+dEeSehaVPRw0/ur4yp40uvj6txIqtD47GYfDI0TCLAZ32BqY6S7zvuQPg
LP49fUuRrop9zefu/jJtdQnkpX89imSVkC6t09g/hsXKIYTPvXUoEtUT7aC09wKufBJGHbDIiEvP
bVb/DQdFi6JUjAnGYy7N1CY7gqexZ6NEnRHay8nSX8phNasO9BbJwJNR2OoHgd+TjgBHC+LT7T66
Cq6+N5MVgkLGGIo0W0rpBedUIVEHBttzjwwJXuoW4X7hNsua/jBjhNKICdgB2htyY3XEteccgSH7
xHUosGZFTCYMKx5sq4TNtzATd9R8hmqk18Phlhue/eFty25vp/OuvuYfq9DLjgEI8AJi8FPUoMW4
PQUY5708BijToTy1AeJ76007v3m7J4yE5S1f2iPJ1yIWZinPOspkfB+//ClOCkSlzH0RBSc7GtRE
x8rYqtaIgHLqSYTGxuW95r2/5TGlWXhNI6lTon5twP7J7UkL73An1hhEebu9pqwF9+uKjn1cuNaj
LaQDNy7YYieOQyIKuJ2BaLXKhv/iEJ7V+IEUfqbria/b4wsaGskYiH3TgTe82ErSl1RcnhQWrj9O
JDZXTSa5YTHYpPwKMn7KwiN3dqnJTVtegWRKFbU3fRX91dGsCMPBivR/5PsGldCN9JFKLBoeDDCF
q2SNYpheGKSB4LEjPJInF3jq6mOTJpgv31eFo6BiNI6OP2by9H9GS1a95HWRuoKu9ErJb2z7FcFE
6gPcIEOxSPS0hfcsMuOQ1PHClS8orC9SfUjlICSk3y2SUGj3Ksf9eiPLMZUV3PChxR4KSQ+kCon9
MvgSRulFFL7+cajamSXylbYuczxdKgmfKDffMKLPNtqQEp5zThuq/9oKXZ+WaxrThEwz94H9F49h
5cWCOpExXIB4LdVlgJyHJMLGwacB7F+TplkWIUEU3TQb+8KUTfwgBybnDykrTk4PGV8R5OnaJCZo
4spPbCbFDVNvtaGnINcLBmYOyaYBJHwRcmNOoEn/T9f1g6diB1764w42ZJdNAuXEIt1yQwovT515
F/4scbtwPpK+Tu7Kc9fvFdp1CJ+aG1TEnoUcJASqrTK9Me5Rru+wkPl9TCUwceAo4FocYTyTsQKs
aQvorTJxMvLMtgjsAL8LwCzic+7Kiwd+LLfWSSbWL+TkHb+DxdUTdWIAD8Kk5Xk3D/3BTXr1Szt/
/lZE2miRJ6UoEKsWalXCsXpHKN0wClPyAtUPMNy+YYPBCp/nkiLx05uVEsBOR30r5o7+umRznWJ/
QZPumXcJf6UcWrooMegAQJp1WZRdlThHcQLTFglfWAUjYPds7+8AGFT6CwNEdmviGjhhY9dkjQri
bgtt5TREfn9R5jYktGzPm4jRcQ5cWPJKqlZr9Zgi+WgXgIcyTVo1G5mtHqzfeH1h3MAexnUrlbDz
0FXRZSMo9Pg/P0t/VyRRyYnKMLg8hN7Uvcqfybaj5nORV0jzp4PbL1suAp5T8rQXBTV8mlod/OKf
OFAeA9EWV9abtbUgOlvz8wB/hipXHKbW+R09H9oPsmHZ56/Nlp/zcKHCNOGDhZUUNWMC/2GPZyqv
PrUhKGcXwd9rZb2Rdmw4UllUc0s8WHRb19pt1hUpJ/hdsGVpO5cHcUC/uPshwCaJh4dfz2sXCApz
9mrI3Zusoaqq1mh8nA3rLI4QKZCLW0linFN9cLekGzZTYbCI+DWTaJ5gapkNuvb2ySJ4xjel14RV
TyviANNh46ggejHBysMhOu302GBzWFGAmcDr01qZx9diWDOhw0wKKGlS1WM1n4IiBGdQaq46Yf+H
c2vf9OV0tGV3uk+Eg+PKHZ8gaB1b+foqCe9TLWEK35s2ZSLO86rgW97Q6VsK1Wviu97z8Lc8IvLK
fCi9rZsjEIj+37ywYA3ViGgaHBcN9WsBMyq860Bc6XtMnDKkDSGn4o+moCU3PMOLKSPle89NTX2A
EmWB3dVL7cbGE6840ilZnFWg8dzN9TepXYCmxO5D9MhFJnjO8z2cAULKc7ElrRyHCBNWEZKF7yMN
kS8mkbLgCsQblaBxddBt9kkOca2/SMuOggrDjFWIOtHBYD+2UntNQyS905XRi/9pAU60DGLebjHX
vewc2caC3uAdozGtY6KzBRZvyNpdGMj4WdPldvAs7s8pYS+RQmAQYG2ocz0bUMkBgibfirGu42Xe
MMLcMi01POneUWfIDanI/cyvVXYeJ5kYCPbhGbTJPvJVuEMZREFReIjke+kVnPA1WJSmchjnA1oN
T/aUv17rqojdIG1f0h53m5SwGpYXom07AHOS3V1NmrOY2WcC+WSRODXMXidv/Sc73IbAwCayB9XA
pgyx++YJJQg5z0KoSVonfbC1Cw8IQL4RLOiy9mxcfv6Q/1z+2gO61mIoekIO407hxD5FhKI1WZee
SDxKlXw/jZbSpE/dHVivFpAc0JPp80+2wqO6Ecf1iloCMPMLJepKS4QD0rR1eZZ5WnAxyGd+oZ/s
3Enphg9VCwAwP2MI8GCed3uqbu5KJb6h2Am7hK8UHRQyU/cE70fQhjp/LSWk8X60zvQIRAL4L9Gq
+5uWQ66ve6i4rsgNMQH6zL44Y3dGpDVD+jD0ilF8TzvZ3PrtorqoJXvZTNgCT5oUlzX6xJ68+inY
jng70fB+dB/MMQb+xr5LoEeV+dcdfkLhoniyVuD8YzLNlS6GzFNbYSU5ieWWbobmCxwBMxJG0rCM
nyy8GnC8PPaLKcc2KkX5/f6g7WFBuMP/aVsoY0YZEkx6Y7AZEWzM/2/T6eNkZMyCqOiD0iaNo6JW
YONfezibO4gd6Rt3iElr7shWRlvVuNTTMFLmA7rvE+6/FWyIWLHYFYwxjPuFQjpEf8SOTw2ug9aK
JR1ko3dqQKrq5wfGm9pFxJjA7Ht/xBCl/JvjRd8IaScwnJVdLhRZJNBu4t3iFOcXKqgj5h46TpQ3
Ogamn3JjEzQMXaHV2wh+zcrGernk225s5jOticvx7KQShc3GLLxeClZRkTAE2O3p1Zfn1XbQVnW3
5XkWZjv+F3mf3sxIvEJwOMGQh2HanurC3ohmVkkBxW2VeDH41GNALDiuzEN96wR4deKHUnhCnpAW
eYILUKsTuUyrzdOmSpUtHA4obM0rGeURiqCieUYHx5vxspmDTshHSeMNvWge09W1KeInCha7NCeN
4aKNBDxii2eVZarkpfMOEDU+JxDDTKC/m6Nfa+rbebrJwcdGVUPgy7rGCKWij7E6Thj02iP10dda
rNbP4icYbq0XrThOJwFm2BIYvRVQqkEAcLGSDHqSogiNxnQVgccFbK7Z6L0nrdhn5KK5MiyPkZMd
cFkUDpvq35mUjpDERJfJe1FB/WgsBwFmDlWThXDzWoS49v8G9ZaahE9/g/Qtynlan1Y5sPbJ7vSf
wZZziQDTNBYfK3VrRGOg+RTGPqRMx6Rq77xKFgFEBWb+XZ0YOryE96qjrW5isfPzM3NBAr3vEdyu
rj/JPbOdajJ4Bka8mROy7SPwJzxvm3AQmKaSRHS4UrPmfvtsvbIbUsPgzgukSZUAL1+8qAozAFTc
G/MyVqIe4fpyMnz9xIIrGfksa22S/jBwk62T42suYrG/rp2Gu0udbveY/76e31xwokqysM0HrPRV
keBhKihXoGj/edx/ONR3NzkFSWYNR+r9glmdpv1BaN3De2CPkx4wDc25+X0n673wDXo9UCSdqvcD
9vaLUdvvZCbODQr1AWIgH09ytIfl4klUpWaD2G5qwSDtlVyQAKukbyGjEJSo0kQTNmhfeFKgqb8B
sHI0bU/e3cjeyRTFRtQ0X7Tz5jMkci7EJp4ZH4Dsb/oZJRTd0tYv5wI8xk/ic3W/h8ohF3vdzP45
/syzFHyt4wz64wiqP748Kyk2qCqfGqOtMLqiRvXAVIb5RBfoS10V4IUyYSPsEV7pLWxnFW/6tIVF
81Kz8l7ATubX29MTnMD2xRVb4xRKB2RygyB7bEJv7SELvSmszfMpIlkNF1sHZ+hvRGyuM7d2y8cV
bS6oW9Th/dk+h4BsIYJA4uYIovEwORvlETV25lQKhDdHx3wA7Gzu+Fanb1ti3f16jYhl9OQqQgAP
JabrvIflpBEm1i3LOoRZ+crcfOh6vtr6ia1uqrznnyRL03Yvp2LxxPRqtEH1mkWYKKEQycZuoX1v
w+Qs7Kvw63c8aoW9uDk3nxvPl+fNcw5pBoZGLTLF9uE3RO3ZjOWjHZxupYX42hPKy588L2Ae3t4u
Icexmts4mdwtLK/neYEm1LuisJh0R2JwIac/QKpIMLxUQOoLOOEdVwZ153WMqff5riBLu6wkOuZP
18FL32HPhcan0mfs+L8mX1CbmxVO8XgPbhfP3ra3rTnftG+v9J8+WI9A22fGF0tMBo8YHGfnzlhr
DqWKRMpr2hucBtePeFdpLh8GGgkTJ2OB9ZOwI/VBnCKN38jZXJLFiCk3I9q8vuuNdepMf862+Kqn
os4wbHtjF9fv+49RN7ukT5wEd40nq25N3B5wGob1muqVIYdtuXRkQjyp8NE59ezHQzuZ8TJqV7Gp
aiDQCwfRPoLLT8pjXM4TqeNXKRxT1agaTOTsQQ8Qn2z/Rw4XlR8Rq7PGtIXqKTqHrVglBLw0hn8Z
yX6+Tw0SGyl2SDp1ezKjwZWgFavi7Hk+eb6+5rDFAia4s4Iacj3eqdHv1T3BHK1RB9IpygOhuFhS
Dx3xWMHnSYP8jaBilUAAQa8NyLdaFjgCY/REhOP+yWk3hsvkdniqw4Sg6nPMmFWV8L/yxp0Nea7c
uDHD7h++uYfezpb8H9eeYfcuPOTAtLneUF+J9oeqiw+LBnOQLBULRYDlNkSLkh5p+EEYv/WdezwG
dBuOeicEuIbtFwJD6p+CMAd55FHohI3nD5z/sRmb1HtmZioSUVQybA91nvbD7Ij0SKFYAFPL0yJ4
yNDqccqSFj6ddWxP6t2mB7xUx6EX473X22yImidVoCJcpmV0tauaJCDPr77NdVYPXbCmkCCSVp98
Pq3E/3gtCiWPcAYDSJ/regaMSqyvjPZzn3JQkYYkEkOXROMcx5uyb5LQOJojW2Iv8oZaDo0MXPtO
8J19KVdUBgM7JXNuEfsPYt4c4JtXFt6qpzutPSs9Q0BNcungRNkFUsKgG4sN5ZjDCen40ZScsPed
3T8OFr/uWBqkyKD3AQ7a4o9NoZbOeAvPzaIQZRvtNTlW/uZbN9EG2J92NID8e9KAA4rJexlSjCaf
p01u+mFuS7kHJOHKh9kS8hxk2LLSKSdQmEvb0TNeDtn0os0cKIztC93ulDpYDjmMuGbmEdaEXjkQ
cWDSMXhR7jn9VtXbj5VY5a1jPEIrvLogRARWeznJ3BnCN9CmvLYUI0M49bNdb3p6lQYAZ03d+4PK
Di25adEUDyLeI6DTO8VnT4+Kj8EoiaJiN8KqvRfJ31nmCKb1aATO1E80P//dURc792kmcMqQfB8n
GNSQQSJqjjVHclh1tuETw1+zwonhUoMdb0ZWbYPVGoUO7TyuOYg45vVAaCJwGadiguPJniO8j1Np
voPxLvKMrSbwE3S+fR+RHe5jhaUfNRNKJc4mJUYE2sL11cRFbDO+BSBN6eCIl/dt3d+GS6WYTUXi
svy3QoX1Og2BN+GpblrFS7DCYsaUyANcW1OPayTVoOJ+JdoSyTYQUt6zVDuhnEgEa5snTpf5DBt+
ZM9Twftxctvug8IdsrJKZDe0CW/lgXFLrHXbQRDbpfYDlPvi/NEnvkY5XW2ODr7NHxxiZT4/mvs8
3fW1hqv2MJslQo1DuzsPLJjf5+RxG0DadfF6c82monS6gu7/nI50gZaBkJJcXOjRjXNOaWMaGq5u
hQsMgUkc3UxwncJVrPCM6rqKUvqOa+1Mh0Q0L1h0guDTbzkzixKJZjWY5A6ZgBFKocH7Su4fabcw
xvceP644J6cwlQVsJC8e44Xv5sowhyw7oabResOJdFtJIyEx3m40M2buAl5mQAzJ6BQIKSL+f/pj
X+xiTawOxPJxcQxAn2zsc7h+0i5Pbnd0VKo22fyqWukHYOhdP4DYEmmvd4MJgxkSkNXpzE0FyWZD
776D52hsmnBiufaOodsY3+CrFb4lYeHsaZCRzWOUGJgsHTBJdWFt7rxy1BucbCE0aB9ElDQNAbEu
vK1LpKCqAJSZ7XXw4QVsvSGvTmNU1OS8UjftEzVLaOYNhWWQg5UgPjdfm3xsI19xtby71QyxbIDv
wj1/8je6fzyXuTWfRKsXdwuG9K3mdRTkAyuhpVFFR07f2DxNU988sITgUG8YJzikMTAGzwsSaJkc
i+StW49YONEVeI2GCKs04zOBR5Hnvx8ekwGhpbvKGoObxt9B9N8hHnUdouLDRmZ2ZQdvKbWvek6A
hNccI0Vg73Au+JOmK64QpRJYn+EoIl1huCKm2js8eu5NbtzjCwA8yc+6K5N0GxZRW8voSEeUhXYS
dDrHa0pTWQkFX8d+TfvDfUWowETzoBsKwhFYrzyhvrSUGIezC5bnGB8oMsIMJLFoILDWlIShIb+8
3P1V/AuhvJ2j2DgPAhsrfWxH1GGPLd8eUm6wbNVPgzYDPgz/OsCQAwdtSoLVxxkFKRBhsWUYxlqC
W78wLlFbGLFsJdS7pO0N8oMK3GYjPCc3nBMFoIllXx3yPTsy9gidMEKBt91TtGRoWcxbFZ+MDWzB
cXGYkv2ZOX/YjThlyYZsyDjBBXbka5Mn4E+6ETgU2PvdtZ5saE7vnH1pDzJEeOAeFskXbZ3iNCsu
OBhW5fbkQoagAeAn77show0xQpZX2d7H9meV1qwcnECU4e9VctuFHs7xmhwSzCJGmzpmR+DRupDk
LbONU6z7Dp5KnLeU8nHSB2ca1lfFYxi474SMBvlzbr5eGS3kiroLxHyyVKpUNDiqI/qZiLVd0tnW
DmlZ8hiOPMDzjpWoqwKkD/2QAnSXwXBz5QJ4C5USe/OQ1y1J2e3CdAxnl+VWUZoWwp/rxelbbMeg
3WL/j4Udaz4ckBunzlnWBVCwGmoIXl67IoevHsUqVMGwxD8CDOz9fjKnJSvn4sSCFqbSfMl7c/dt
3+tWNs1/R/Shkm5eqxLfYLifqghghLzAwVI6AVdykTdIr0f7JsB/j1lXakzEPAuFwIAVw+3jhIrR
Qd9JNDD5nrTkKPyRi6LEgtilqDgPPpCGLi04xqlc0eEpogiJljV4gj8yRB/5gjgUmISJLDwm0877
X8Go/IYDr7p5qapGApjoZ3nkX/RthfVNpzBQd3nqKawlKQNIhtF3LKO0BOSezcNq5lVGW//fdIDe
t6z5OsxQHE28yNOxneRDaA7ki3dsTGj9EeQNZu6yWhUqhxS9P57Gb4G5zogdQyjcAI0/dpBqckKn
NEtVH7JFksLKRp2Jv54ZuVIQb7T3VZrujDwvNzWI67Zc/rADYEgZ4TO2Zva4Y61U5x65HgaKJtgZ
WhAxx+wbKW9JcXm35VEuW4sknYB0QiuHemxW3KWNVpjFjuE4RYDoROQVEAVPvE7KmGkpguorgrqT
MCUe4hy8AP2BDeTLs5NPDrSIzOKHuuZxHwV8Iuh0dScrubGqP42BreJV21Bl4sOL8GM+kpz4OmiS
BFP/dPPIIqPyW6m2Pn0fGgSeEM06N7qV/uwjdR/SpnEqlp3vF/48VgZQnPLoiDg+Jb+fe0MO0eYh
oDdgYe1NeVshfvhnle0QivgZSHfFDSMCP/oU6wV2Dt3f7Es6fiUP9jgfPRfoTws85lsNe8FktwFd
NBNYvNggQ2NWgYHYvjcSyn784czakyZFO4dTrbb5LmKZSxk4cPV+yOrLE3LLC4RFFs1PIq41C6U4
YsqDpFYHIADbAJQeA5OEIBObjraaYAwmE2I3gpQxDILz6h2q4Q/SzO75mggq7vGzVQUxgsjaqyP7
9azdcengf2kV368vQBIFITZhIZ0LlXxoiq0w5vZ1wIFu9OtUS537a8rBnhp7r605x9qo4a9nrck9
jpbufFmKiCczIN8pYBIKPzZOD0plPAaIiPaHNow+9LYkNaAfQgPFsp5I8iEbzhcWQzDjrL5LmisI
pKfDgqx4IyzvUGos0TngLzaA0398kHKVBk/Qwnd+wr4TaeXZm4bbJsPSnbHoETK3K5UEH9hwNnuL
CZf2jqe4q6ndoUIB0DOhtCtt0730rieTWCYQmlUkdD9O7N/XxTrsK+1yN1WQG3hSdCjTe8JCu6w8
VVipk8yk0zlwTIGMnaYbm7zyzW69B6KVYhiBxM6/LO0u6yOmf41stHyv4UWNV3/dA9oKwyY67sJv
zFK6y0lM70Y4FLdteATsnc/Y87Iyz4HMiYMkwY5tiaSkIt6adfT9vUYy3Fn3XG8ZvZeaizEmXVP8
NahKhyLTATcniAiQWZfQWJUSwBvt3uG6FgXxHFt1OrfG9odfyIhbUUQ597hcM9R3qYu6PofA24GD
TutfA/ugpdqHCo0q+Xq+hg8GhyK8Pbnzm9qbdJfmOIHe+1y/BaT1H5vgQiPUtdGvLMzLiOmiB9/i
MFINPqhy17KpyFjcX7d5+rkpe5OOTwn6AyifiYsuyAaf7p1RlRsL0OZ2HYXeNpWfoQy0zMrzopBn
C2XydHHiKF9r984tk68K1O3bbWPVxQREsFsTByBjsgN5TKrnYAOtIQFaV0aeHyPLrkOecsgcp5Wp
kamT9GVbeuTR74OWv3YNdTiBUh+14AjvOlCToJjyqwLBi1tnhIYMkTmPvw3IluhUr1UDT3cRovEg
EvKLrA8MBnaRBcp/OdWjLGfvY12snxezIFKMEcWXWi9On8WFeMT9e8zFlD+UiJ2ec8TP5d4MMfqL
en9x68o/mSBaOVps+UG+GNGUgrVnjr3VeHivSOH3XLdgTGx3LB7pyLzRsf5s71o5xPIPalgaHfvV
aNxOiED1EeT5u1BuhvhJXxp8JNQpvWLVuKI2ju5m+Z+nz2Fgr3w8NhnFMJrP1Z6ZIVT0oj53YonE
JSLNsHp4P9Q7wOqZWDoiFY4eGU4W68HO2hjuu/FdjjkYhJhkTMYL78/Ml03oKKxGFzhVdtqElrc2
fIX4XreRjjWAnsGhsQxdBbvwsTrKm0aiZkiSGjchwBNAnP5nHf/2BK48v0twN9yYb9DFW6oW922l
OMKIkFrU64iz4w8fMUKZ4yLRpmiDZ70HaT+JYVXEgO9q2//ntSJfwnTfuATEIM33aVeWvVMLonxW
JSWr45jr3j846dNB/Nj5ewPRdiKbEo1fpg6WaZSvJMduXEufg0QaMEqzZ0cafV5LYyerABmORfpp
jV28fVMdWwMmdAmMt3IochtHCBcAKGc6Y+8GMN5R/ucJLgsxSlOo6S40K4zl43nIe5y9yoEXHuA1
giCDiN9nCOAA/K7QIhH6NG9M
`protect end_protected
