`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
f45ENrOvV5QABsdJC3zTHUbe9o1jN7VwZGbBctIFXgONXmFKoluKjnssZYQ3ujDTVackCAOgpz6i
0lKkL+4PIQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Tg7itq1EkObSd3bxV14rdSogAVobg1roGdDYpHr0dJu519nSPuaPTZmDNHNhLzIWUacRXyoY5YgE
bfeWad3oTy2+2ffItz/cP9VYuYL2iNxZlHMJdXkT1ftVjxZR8I/c7aiepFcH2Pq/qD2ZTBXioXF+
mqcHwCrMf7GqWyCUS4o=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IJpuKy/fQ7NaAnKyhMHHMYAj6W1zGYlXauDwQLCkXyrMEsrlb0nK2/7wuaTRaZBC9Vv69PBbVcoM
xMCsW7EhTTXJStnvLI52rwXlAMrpvJUa2lv5EhaONDuPNVX2WzpxrIRSFkSB9ntUsiPalivkT4i8
k3Td8EoWndb7qGiY+IYkYJYPg2aIVfBYu6HJko2P7Eqeqx92Yd3XnKlQrXfXjuSb5jabI2mC+0Ew
r8JNK9vO4FMMRKQz8ENjPRNgF04UE6lyu4T4zA2OqEqCboQTwr4DhdSdALq0bv2yy1cH8cNy83jq
7diNwiJ9bF9LZHpfQikgcEGKxitaG/R9W0fU0Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o8NAFuMo0CWTW8F4wVU9Eeh72FYvPu+VrG3dW0B4FgdvYFoASRdE4JkEeE9wkWC4ua71nSBd6SKk
6/N2e+VA3UKMYrTHd05cBNCuuUtjn+uKNQWOBFDg/4/pvxNc1Y8WYmaG2GCHhR884MqN/r8Otnc7
7lJVn72iDXbDwhGFCTo=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S41yIGvZe02y1u84WGjj/bxV9CXZJULUC5F9HvB10r1Ize7WDCIzNlTazEV+NE+/TTTq3raSNMrz
VaEWilhsLe2NP6POpYRyqacnMDwAek/WxLtvlB0hYoSDHIWFDNuKZhbqXrZYxtzZuzGzEDFYn0k9
TVriK2DW8F6logXT9KFMAwJXd1pvdERqswRr/Bz3fV1sfhE77sGxX6c2RpVWRk7VieZf/5hYDlTb
IuUjohB3UU8/t3x9xm4/OqZ5aJ4z3vd5/w/Ospp66D/xu8jtnbIWXc7r9gmpZy/u0ZINmGxUrqzL
+9emK942IZVlVoTOystxGHHv7sZARc0slIcL4A==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60368)
`protect data_block
D0qMayPWRl711dknXv/XEW/stvVI90j/8bBHAOdMC7Yc2Z7B4GwakO/TLuGwL+9Uvx0CLostsCf8
mhB3DHGF/lY9LL15eE1rs6OibmYRoznwP2dz3eXbrioOMDHEyxc9PhAyLRWdlydShc64qo375RuD
dEdRd7wCRIpAQNRGAgfUIF9Tkg5O0z9HAYP8V4WsEebEPHCYElXaMnhGoV5x8wwUfBhWG+1q4fm0
ddBJOUhdm+I+hDvd6pllNc+/4c5Sh7KFgZoTKDPEHYapNmeFufZMNZ4amm5k7cwN6Yyd2thgL+Um
Y+Xw3H6uOV+HX+Gc0V1s6MUdA83cv2ywlWrPbidXbiOX57PRssb9F3LctN2Zk9Tujz7UZaviKKgl
KeJ/E4wfQldJHugEwhLJWWlLAS9BZdUDWH+JtrB9+ze/bcSQhqcwhntnboJz0t7rxbnYFtUZD5+/
HNVDHlNUtv1hqmqKukK9FHJsCRzrG21gbjCiiJCPj8lDk1UPwLHP7MzVQ6CaQlb3OidoWrBnKwx1
CFZRiwk17YLTBUzeiO3nudwUW7JYEXKLwhga1vXvQ6ZARXFcxksGb35GqinV0ghEEIXbdRChxUYl
XVYYOz1vmUW+t7IzEtKxUyaXadnbvuhT0OT3r7nG8g3UWHV4AfNjpNtapmawrHFyXGXJREmhKTlp
czWt1E1RlgH2s5152b3imhPG/iWza2Wj76RxqEPOk/+DTjScmO8bzbAO5AfyZM5k3c3+r7Ove7QW
I7mccrM2WBhdvvWMgyr1YoYY4XBqMvmro14lmdyrBMsOVfLHyIClgEoZ7ePSpYzKCR9bEDn01uO+
fJJz4IZCSay0XsdAh572gFhVyYHLACOWLlVCJY35QsjAOT8yBk7R5m9KJ1KBuk/RwuLfz/HXIF1p
OMqRH67XWejZMwQyVbR4UMBqV1DBpEaVENG6ya5dWliQo4do1Q6HzqsPqHyXXDAe91EcH71jHqpY
APMMQnymaTRaPm3h8XqedDXKa5Xf5t3QFxhLGpGmMLyzhh8+8pBygEQITDafaUQ3v4cpoJ/USZEv
kQvkWiB33mwwh/53J6hCp7/ldZMhBs7v6XPpjfJT9Rih8vqRlZZFdJj337C8Tk4IKGCNHILSZ6HY
xYG3o1IgQCSW2xhE75g+7dpVFhdfxq/ll82xdb8/GnztZIULix8I8pqHww22gR8Dk6nVj8nm3Pnn
gARLC1biA1GDfZTXc15eEPaKnWLsOiHHgkxvSczui9eQnNm+e5WQB2jZkELbQvHxyisAlpccLy8v
zTZGMa4ZxkHs2T0c63KQnF5rPGx0BhE2bhKd0Vbb4BqUZecgt0lNnjmYzFv6nawchKKTFBucsREI
BPTyqisdzPOCXxe6LT5f2MiItcg7CMsT8COirpBgzfAA2RHm0YIUx/AzANsUWz06QiOmJF7IiRcg
wcKCCi3ecD3G1h51I9TVwI0YZMobGNT5LflWHHsg5QC4ywDbhuwZ9jxViW7BihAToVwWUAFCy0qk
WM88jpsashJTwcgWJtv1h3F9JWuuGi2q6c28gSW+BUzG7ldni01qJtJQJQZ8I3MtZeiUKYBvPRrH
KjmS557WMoK48parF5istlJr9+DA5oowErzCF5jPpNi5t9j89tvAoVgVxf4LZzckFOgXEnOAwZIZ
LeZNcXbCDDyMa9rQ+GGlkLdqsDwzzk2wE4GlrovssIz7GAlVNWAoeYQQRyyZRc0wPv7IgomgCMpG
RIxH84hFFX5eu4rz8TZ5rKvQQClZ1RxQx9SekuCxlrMJo1TkKwUxoaKoXvMuS9beayMyUf/5KjDB
rGQe5ObHoHl4gGab9ZQRmsId8I9svDjlsfDhXfvUlFGfHSXDqN6p8E4GCUfXNmH8TcNbR9DROdVB
ZxIsoXbV12cvzvsOw7d1okRtqJ/9la+vAn2FSR8RoyChAcARj/bF3VHvk1rg5B1qbVfhFK+JvR0E
BM3sN1gVUb1oTq7jI4WyQ1n6E6eeaA6sKAR24P45daXDw5eb/hHRZWtqR8isXjWcNY7m0r83oQ+u
W3nVJ2319lx4R7w1Ej1SjMsAdgyvPPN5RzfYeSJ9Jyg86HZZOcKdVdZ5HwfZEywRIZlmunyj6cgn
EQ6KQFfSEb0IktXMbY7Z5HOPTKRYUSVVvNB6m2D0LA1p8jrpuHD7ajoJIIE5t9WzcEW6zBW0ldwg
c1ptKpQGUaqx4c1CE4VRXFn86u4fLaA4NGGoh7e8G6SqulHQnlU2lFCqoPwvRbsuo7WugCe+WCWm
v/mTOrd296SINWYEsy0HO0lZIVC7zTw5XAsTP2Vfiri4+WbLQuhT/x0PkOWb25BQ/Yab90XkfBq/
CS+kwYdplp5Ve8nkQ19EHmAKueC5rjFfGWua4K9n51BRleXeyr8x5IQ8zL4L2jq6d+h+8FA+/V9b
YLK0GDdGw/U5X9bk7mHdcUoOy20oiq9kitWsHugRK3ID+pFQ8uUBwns053CqcPyToTuPEjeAOJU+
PFXrIbuoxg9aoq2j+NI85ZC65hQEZL49koorbHgF8ytD48zT5r/+AZ+lNU2nsv7qRHyCwCoJkWoU
PL6oOTi3KnUKK9PWl2jhqpwavbpUo/gpIb/TerrfWC14aLXrZWG0YnWgPg1Qyu+qULQcV1AUuIBa
CQPSwD/MTXMlcGrJ51suFMgnvysBxylIhjPZ5HGV2LU5jGnIZVkcKUM5RXRk+7Y3ievm1uIVlA80
Mz9wktTcqRV885TtM4lyksxOh8g0oZAvUSAzGjaNgAM6aL8E/bfrWdon/VmjKQaif8fZYoRl5hrc
QLel/F+bIgJw081YEQjuiwQCVJkuc11Nl0XOQq2AAtWbJIl9XZ72erRjyz39j8wk46TASqUHwOp6
30ZG0PSKbZkakoU4t9aKB0YPcejeXqYyAr0kJUZUwqiyH27DOO8UmgKPYaORwJs1lw+o8UuPkB4Z
a36Zg8l3G7B0EaPTIM8WoC7fBXQaxNMG6axp2gIg+v+FVw4JuQcMK0OA6rgHNjudoph8thzJfxHQ
8Tg4B1PD2/04Qfug2BuP7BXcl+Ax9TIHCmbpdfr2F3eLkVbNMwM/uD7CrJ0WNog3B+5ulA1iuMWU
KCmxhzz9Ounj5cIiMmJ3Bg9juwn4QgqmqVH5X2MFtdpnyMd4LEfkg9oEg2rLvtlamZf/1kweW3Gn
6SG266MH9+RP6EspJVSEr0N2PpEK1+wQQk5qggp9kgxwvHINk7RPoWROo8QC29KdTYnnGXGhPWkn
rSOH1mZ+iVeC9uHTuaOearF4BcuEYMzy2vv8HmpTVqg4iRT1Q3JdxnoFYKWuOTthgB5B7cccelS9
cytBt6Ygo9zDuXGgHIzaee/y3b1iFeEFJNboHFieNpoTpeDSfFEABVpSP9x/kiQdRPs1mSQiwNsF
eZplQBbxpTmbj5DOy6h1eluEK6zl1TKt7Fy+Oys3OSYhNQ+eJ60+7Oy4fk0usOFOroaLLhqG7g97
QOSy9zllG94TKGIWSKgNC4UYiB2rTOyuMnIUowScVRXGlUm2DbAP26kiDaVJCbRtvSDw0+udqyaM
3zx25Vu/dYEhMG+Ou9P76xjFJ4nK6auw2wpdBAgaKPiX28QILO/ADsb2Em2yXJdJpw1uU/tkdwTj
7H1S59StKV4QE8JZ/lpP+NEvAFhvO1xBqmkcqZl58W72gxNA8GMv5Ybp3W1x9Pz6TliaJUB36EEj
MloeWz8ibesqUtufzXMtvcbftpCOLmFLLCuZAo6m4ByuFQG3TTrQn8zqc950KI7UBJZu9hld+pLa
TmEOyBDUN0JKenVmIulHea27DWfFLvgKjRwPcRtroWfnwIxaUlI3UMONfVufxo1LDmH+Xnuesj/1
DxbVta5cwNr2z3UYFu4kNgiXF3lcgXWWP2hp4yN95iD0RgGeR5iapCV+V9fcP5Q9oBpK2W0tyYKb
lwk4n4+tWyTuQnPykf+nwTAG0Fez56ivez4J+7AzGAoWnCmcWHF/MJJjH6oLN26fpVgWQXRdrATI
4y2diOCbXVnlhJHpIU7FBKvSaFy0ih0v+vHQTX919Sox0Mzreh9VULsF5JdpnUjG85jx/DECm1pw
pJ5pZ2YyLASnEDrveHRaQLWtWIisF/nIRjN887eMEFXToW+fsHSfUWxY7PvvDxeKREGJvh20/zv2
VOFkEl8Ps/IXjJp374wSClr6RLSk4RNsMUZ6t7VAcqrHNgPAbUYgmNdnLlVPeuidiI5Lfwmm3uq5
ohg4AE8ar8jpTAYW0O9Lrc9blodfn5lRXJkGe7f8Gm03wkDPSBj05AH1NXvnnKqV/eEv1vpW+NP1
o/IoEWS+qtVhC2kLTBpP+6A5drYURMlE89ePe8SQAWJ/9uRZSW87bOftpRdo/1wpOGZjXZdaDupu
W84UA/ekR9Dh5vEJX1L5vm5jk50AGWaWFlNCEAc8nrxqg5sGduDR0BdL+mK7xpmcY0kbdilVvE+v
wxjoBbBXqdxM10IYWUUO3kh0jIUV4vgqY0Qonn1WQJH0IwcItKnfrdVycKCecPDf8YTn2VOxnp/H
W0yJ44hMhT6zFdinzSPfIdgasl98hme67vruwxyGV4oiE7HpZUbPlD+JsRsvhf+YFp++L5iV7IW6
b6ZnmZOBO73tK8yUcITa98AkXosjoxeXMCSHpx7kqnPYC2RgKX3EKsA9SudQzZf/RRUdPZkHZbUr
WCEPGsrI6cO1eqDmVph+Ms8D+tPlXZZYajBcOlyB8S7vXGuAxv1ApWzptqdd7LdAg81dW8lputou
cHMnIWvo2fZpjgRzFMpfLvcKcvbHVp5Qz4o7hXFM4bgE03Z7qPRpOpBrfGHLrm7WV8/jGNFEkRAT
B4eoG1Zry7J6O6JkmVH7vXTElk4wM+NW3x20+LMD8srG1ASd7niHQu1zR9DPbCJZKFAteTUBVHy+
zCwDjkv8W5EOdzAHsakKZ8tNOxExK4AhpsnrZTs/A0UeBgJJ+EBCHUsa8wiUt6CUams0+qACscmJ
onlttr2RN0jsxZ0XL0MBxb4Ku2/IGJWkQ+h95D3RmG0JCKcoqLMHFzsuRRGmJRcX6k1tdt1OmGyD
05Ik38kXhJHXluDPUdEZthfxmqo1aMLn+QvQ1ibMySqYjMWtsjG2QtKWYHfo1xsjzp+TqQhgOj/3
tSgjPCXOYThqkdsKsICTscgBZ75x0LtPVddFvFrSx7bWbkLFb93rTBD/DGvv5BxsDBrf8zdyoo2s
j/vcC3rY0e56scKwrQFhHgru1G5YuwSGxGA3fKlRPCp+DGBKjm0Fevzuo5lxfQNHw7tmXbaiMgK4
ciZK9/eU4LX/UFm05CpNRtTwkgVKMu/lIX9HhqZGiGhNs4Bwo//StXq0u/1KAGVp930GIYkh+MC6
sGjILs50ooX3wLIWccUKCso2f7uoKuoBGF8nPgEte+GPmayIkZbWPOZ7TOH87e9vNEs1Mslo8lVU
ojDk+FWte5uu7UPY8+DZNhMOr+F9AyMixrMlbN8CILerPUqOZm+25vZ7xg+lOaAKLRx00tzggcsp
574SHKKRFRYAjYXkNJ/yHvnDW1fwviHfugYWMd9jaqZXtCROAnT37f93aTKNeiAM7rBgyN0XcPOT
aST9bLXvWuo2P1OVdIUsRUvFRFbpYKClI4Q6z8xGSywHRyAnJD3UNdd9RMXaGqvHAQjs7JgE+WD5
CduJwUJV9kDjpzi59zecsPmbmCoLOY2ihrGyzWD6wFz0ofzuZd+Ts5O6rwZVojVdLl9SZKnQRl5N
kF8gS5Hx/ljZJ8b5XjJ50X25F7q6Yvpk7fHQasM+CJbWlLgm13gURtHvk5qE6XpeZ+gZH2QHr3sF
FKSd5qXpYnOTN9QeNoKW/3r0O06Pfpnj/4C/6AkZnCo4oCzzCS8ungr9kHXUSHrzspVXK7tO8oHY
hzX65BPYLU3J/HGpCkDo9nuNRuPIHxMpqrQVf0M4EJMjDJrbBJrPbLaJkYN+R/oQ3lTUtPmca9WY
4vqFva/lRp/N5/jtcxfguEZcAzmbPmtYyXpXu3dsp+vS1PuYyV/28jq8SgUYREuHjblIaJfl8bK7
wn2ZZSS++cfnZc+MxA/BQ1D71HDWdCrgM5hZAC28+4vdsUE6W/Asd6sMMMVFOf8hTMjFs47dVKcF
hHdBym9vs2CX8wSgfaOoFGMXthwRx7S/fZvBJf5iHxEIsF1UQ4azkkFWoQWj7wQzbLEvJd8ZgXwv
bJXdFLDIiyWcl9y29ME4w4Fy73G+M68oUcIRlSWm5tsQpK0fUmPeaGEtoytAL/GiAJTTTQ42xEEK
uDdBJXrNkD3vne+KfpUrK2775issatUrQibuVjAVDLMMsrsnNkwE5ou9qPnuCBOSbc/3frZrf3e2
kMY09131yFb+MZWvNlEyLr25GBN36NSFEK4w1bqC8RZ/LmKa7AhNt6OcZi8S20eEGEkrq9bWjpNQ
qG2nFky+EtB89g2GnuVNn3uUOAcn8/r0TZTO3xcdQKBwgSHjkD7/zP0t9xqGvvTholkT1CnEOrp9
5QdHi9DFESB3gifHwh65Zp2uE63Fce7sOAogpGBtEh1aZd89uXgDgTPnE4BObU04x1gz1TF/aVH2
sBngObXcG4VDrCZxM2bRazY7Mc0NTR011F4uX3VLhcazq5E3mSlmbXKvbfrm8KUhb3e8nZVzwwJD
cVW3q+U1U1aWD9CPU+kwlZepxyiB9R1wNzVNDkt1O6CP8o0awfVCpTfdDHMYj6rfuF/I3t4aB2Tg
OtWfNrM0y8KE+7uljWO+37nouSwTlHcOcA37disnHdOquaQJVwijDgNpLTY3WcPxA+39RWN1F4Vi
yxzaW4FybVKDNnVuSl6lXKPrcwcbtj7whB5dC+zPRWE1X8YhTWgVHYRspnpgxyrul5T2yJeAc5Uw
WrT9d1xiwn1TEFlqwcALZnYMm5nixSzOCZSoZDE4ZiLVJo11ovah5O2U1+OqCVRHlR5M6n2N1snl
4GVjIPOY23SoRG+u64m/0BI2jL5n2msFMu0dZIsfyHP8uHcCFuc5WOd7ZRWdOpujz5Ob7UwuZAZt
+LaYMu6XFUEAhTinwGS4QqRgqJETfQ0zVzz1s8CYeb2zig7t9pV2rjwLCts7FMUF0zfcRpyWOS/J
jwYSwSH+QXcBCKALTxMRZJAqLjO11+kuuqhpPHAHl/vQLnYH2zn23deI1gdw+8yRJFBh7UIh3R8g
Mg+9tcM/2csoFfGG+o9db8aDWDTasXtKUsFUL5/Dv4s3RTTW9zVTJHlAJanFwlyeArsawabbRGlB
keAUvEkZM0kCCVMjuErDyb29FvTSMZi+kCvF9J7pHbRjF1NCfUkaB+F0M3wp8WXubynta/tO8UZd
+zKg3oqn/FIM2Le0HP8tV2QmGj1eTZIkstqewKWXTircRXNcm1KUtv4QdgkX/xMiRKvv/zoWquPh
E/BAXbyFYbzfppxVA0WcXf1v0m3GP4oP1AtFcJDpABHoNzwDIaVIyekKfXAb6JfxnSw/vwjbjsTl
UWN+cKpIUKI4Mrig52IcLYI7BrFDL0RubaoIeL37tCpw4ix4dQY9cxGudebLf9YURgtuP+ckJ2gk
RQ7nxaX4D7uYJUqnK0ti//KwtFvA0K7uedR5E840df/vAYkM68sJSU2sxbfamVR1BON4K3EmRzaF
vdF+LdS8eLvZuM1I9MQ0QqPHwquQjerEWNxJOcuh1D5zkSX9vDWNWkW7Koo2Q1zxW5IYLLAUvVLN
mHm/SK7s2yB8TCiVF01iWkt/D45q4D9S+1kYcrbMyoTs2f735IVbdEw+k3DbYHSFMkwteb3lXV2X
5LTfuvsN+84U6S3PV0HFBkgBMBiHCh4ZGdW+NuTxDDu5+H33c8/PoC+Lar03mnivnA5nlTCRnVE9
201mXXV+NOPFNJV5VGD/+VEEVqfXLnXakpqOLqvWI/tXXi3qXRIGusB8OE0HEbdf+7HrCOB8+gcl
OIbS0sD1JdtBSL4M8rMwaaXZcZ8lPrQr3kC+fLCRlkEc5J6Z0RB34+YjTGONkYhclkQVdomVnfJ8
fKNRxMettp2XvZiT0nhjSWvrAupCnbwlbcAugJ6OrcrCaOHxln36qEp1WWyVQLwPrjhZ8qWAsrpL
MO965n6w0w+CB9eIL8ezK4shEHxuIV0F3OOlfTT2ukNOOXd7fTh4idfQAnr1Ca1wAYkUprZ5qivk
oP5SfTUc4DKNa9PZadEThWL7P2I+bKssMDCPM1RFkGIb2G55M3QMryfBzJQ9ThIfaVSZnsyoScLr
1bPjHSNP1dzeUiAzANI4zdiBWilODvdh1uleqhPeCgIrTxJM04QN5UIVe5eOGsg0RkQ3VKZk57M8
FutOKEVOj6GRtTNTAhAgYs2YQ743/BkQjUgMNlT6OctXYT5jVEPz6EhkGe++7pitkZZYMqNOk8Hm
/m7ykmqLSn+UCB4LDlIRcP+Y0rRha0xVePAgf1j0/4zq6ijAi8Jq7LZfpB+ZGQNr5gVGtoVJq8l0
F8e6GILU91AewS1DFtgDfMLWXEG56yJnegZgcX3egfAIpgzJTuGk6wtpJahR7T359MXjHcDoHpug
kgVSBuWAV2Jq1Oy1pdTBZRRZUWmbigWs2B+Ag4klNNnNvwZq/8nhuoHpgZ7s/riVdZl+AR/2PE/u
5uZ+0LhYUV+McmTscLCnc0IJa/RwEhobzGaXE5pnkCDfsV+5oQKz0Ie+tpyJ1U2r131pm+esYzZz
KyVMrNLR5QeEbxQh/MQ1xMYcbxJCv60NnUQDU7mE1PJHJ340Xz+VPWmPo4Eqy4dgbxf3pcBdKRXT
Hf6DVpIKHQgOOZBHGM6Vv/BP2w6xfCMnrK8lYcPHjsWYsfs7DNWOBu+0g0hTq8XMFCcBaTMXpqz2
XA1359LjE6bysIpQWvCf9YM0K6AuwyA01TNmB5l8hlvRJXY/05xG8rDuAWcuVI/XJTeo9fq28/+0
ZfMTmQ95LOwZy6wCieXQ7bxslR9TJnd3cWrDAlDYWDMSk7FXTn06IyjLEuvsa1jDKdnly7VT+yaL
DVctUEZGNr2QSylKthp9/QjoS7RA9/ioF2r3t7HmO/1p3+HSe2uFfyrNK8sXkRCXtFczWW2aQoAe
7s8wwbP0RmqsF1CI1Io8dvjeF86dsiTt1/qY5KmbgYCvsWRu4bKf630poyu0FKokbRnf23UV6ZCC
gWdSNNkWK3RU/j1bGdk8SynBcEur/P96ai0fXRRVjF39DSsQ3Ud2mv//eIEdO6vaPZfov0d5tz5t
JavJ0cvWBSC582Hn4XJsNR7hJ7m9qvvq8+77o8D6graoYRwh+lNFmKtFst7iLUSUgeB6R+J+shwI
1KujVnPr5hT2S7IMx4pqPkVqrJPYccYoW71A6B16KaLbKyvLbk8X6YN8VaFvBfLi4xb8Ko1IqHZd
H5AN9GWZhYztotwiX+67dEuGdQXgY3FuOsNnuSckL/CKOLinCJXf7qpwyNOXIy4rdrH+m0+J91pF
XVkVdk/XGHvEhohqqPxRx6twodbPOaqE682SYQkSHAXAuuZ76VVuhSDhHfsPgvNJcTOipok0qWhq
FqJgXXHF0Asr6EXAwVPo6O66FPvawYtJbDf9EVUQ9O3Lz5qZF4l623407HNdJaIxbN7s09koLIrC
zPPG4FFLUdR4mD/U/VY81m5BTJSCEQUPDaWQFOaIe/dOnc4RzgDBhTGVBSEKYjF11NCi4AX0KTsv
biPHakXBUcKKM0kkc+rCbr903pCknNKXA9fHhDVkHragewf7v+/rRIa5Huj77zKXoj+AaEci60xj
ICAH6tTa7pcoQuXWTwK1Nes0ZQ2NCrEZjR0rD/m/uUMyn9kM5On0AKEzu1dSWRL8P9dnEz3aGtPi
8BAskrXKDDf4Oj+0eDfCvfLFXRyza5mgjloYdyBYJ7WNpfkZYJ+FebMaSMzR+EhsvP9Z+bkFeiVN
lAO4D/w2rQJaHba6xD+3rMmCyVh70inpc3W2QsYHyFm5u1sKX8Pxpvwjs4InjMSH6C9YeaZ/J5pY
7rt9tH3v13CtGvrxTjJyztmYot1+LxmvuVM5ujWnaE6Hs/j3A0hlmRnKxB+xosxiEP2lEFpPt8c+
HlY6zA7OCGCkAYTSSE/SaKKA0LtMx+RxrQeglbFJkhM4Sr3k2NRDMvc0kleJKmwNhsZqeFaHNxu+
+9xNplyJyuYo4bxYaQ8SKsLMmrvYB2T4IJV1qINDR17CdTGMLkjrEhWOknBrF8TWaZKYG+ioFWII
IpoCg45REmk/65WHjuLmofACP32tt4uUXoS+KRp9qFbX+em2rl9/sIGZxrEkBjS8t35idnJ2kqqu
S8dUdmNLxHirYJu9IHq6ygehiWaBbWrkygt9migGetpPLPtaPl5VwL9XBDuUfl2hoPaG1PKPviPS
XS6P6f9TbF0coBOE0PYiX9xFShrCpvB+TuMGZ4l093GCZ+wVh2X1ps8ZU196Y1iTcsXWKfkEtfv8
AVe4wA5/jYUpjVUb3glZ+kFnxk+pf4vOfBhfhGi5mqwI5dazE3eCQktVHFH9SsXMap1PKQC3eccU
y/j6Fk2574TrZoMkGawJWQSO9U5gouPOUkOgiZlMGDEIYwQX86Gd8dZuulzQ0eR1oxHVzJJDz49j
AmHpGUOwLxQ5pLcIDLyDjOs32j32NR42VRsXYLxMpF3Yl4Ds2tBeGNJQj7/r/UO4BVYb/W0i+TJl
6u07AOVhqfXuzb7Y0fs1qz3uq6FTbq5hZT32qur6FA1kDhTm6VqikeDElC7nVvtq9XdxhD4c1xJu
i5mX3R9foUqhdpXnEcuZfePYAf2X5r6rMTtgpDsV6CjbGUgD7JTJwNFPpy9LIKL3IM281znmFck9
OFe2WMY8heHMyK/jInXbmzhu+nofOzYsrVPhE5zGHFLfe9a6Qov2/3KNRgUJY/sN8QZO0X7rMgow
TIj93u+1ffzwxAyPehA8JiM67lRsZVo5JLWj45UM/HpSUYyKa61t0LJXH7tMBevZxSXA1xwU2LKG
2eJdrJp6wfDhhSpQ/Sll+R/2mMRiIdwAzeQ5Qor08TfVhLyZ6wtpKK5WH4qZ59zk992Z4tEe5A3m
0RGw6Pf4mT49hFR5HnAAoLpcOfcunCSEpjBAZRDEkPflyOpybsmjclTFmZl0jI0l2/NtXLSTLXni
gxODUGBYt5buBxHzFtOtlvWJg2px4Jy6Vd9UupsHiz3QMeVszgIF9yAcHybapEZdzWQ0wxe49fZd
tCOZIbYNlYYkGJEcdu6z+Ff5AsINpi3k76tXsfnNPZcZxGDN6hkv/PZSYZHDaPUpNmHnNRdZIe64
POdwVFCafr8xgKbNlyOLn4olWCdYwVPA1J60qWnJInwF89me+TdvlQSvK5Pdyx2KOe3psNF2wzeD
HYDsh7G0sOH67QdAEztqCNmqJBpq308jbWtgUfT7/quoSK6aMrV0EgZ3IREiRIORY/ikvn0ssFCp
O2iPuXXTDL7CnpRKbIRQmAXpAOIAQUJYq4Gfwq/7KdRbVRYqMpx4Z9xyYOprm9Q3v0dg/DKqfiGj
ELcGPWhHtRlYKTbP0LGe+TIeXk6FqSIgoWcODz57Tyv9Co27N1BLkV9cLqHXxbNEQkGqjD1IJMQz
GNwhvLftKhz1xj7R5GVf91NAica0V1wnPuFppzgplF/zsVrfslspe10wcWGCQ7CUi5nNjSu4oAKf
8k0Xnq1/WBxseNE1kiftH9ybohobdxqad6QLMID/KGDgpSHhuviinSpsoc4EFPcjv37TN3sRP5Je
sQTR1HX9DhvapEyrA4a0Zog6ZG23OnNkVHpN6Xl1V12HaNwf453AeDoWIr7LXSmciW6pMc5ucjWI
Y7GQlsHK6rvhlGRq2ifO8RWpRrhkkWqlZbDOfOm9CRQt8aaFjSjW8/CgjjKcuYTipO1NiW+sSt1G
r1/ZRaNPTgyw1rjxMDU+E3E2rORu/si9msIS2bvKF8ABqVfb91TxCgjMEi8QUh6j3yVk76GsBirA
eniNy2DcBnq6AeuacTllV6BCB5MKBd5UXPqIb/mo+v/jYqJPl6ES3oDR0G4gCXo+NbHWeKPUbbNu
F7d/f2THUrsuEGXyVAShkADhKrnBUA3ZkWYykzgzOUYbP9VzCbWPvuqQKJNKR8mPsdm27KI725yQ
S0SjmXbYI6a4NtWZtto5VWTb18107AEdbA0AX+OTHQ0jkpPJHdYnqSHWTSoUICcswWllt0aIAb4e
qjcOCZOqgN8kwjOsVI2osy9DksTb43MC9b+4WS3Jors7EwjS/5BNceRFRxBKceV6usHTBqJ0WOzV
vKZIeXvzKNt3ZoRYkPbNmLMMsOBR8y/Mor4a1U5g4nZk35BKwy/z9MyXTrLJsmhaku0Ujnb35ITI
kLDO1GL5U3KPupmuwp8WFOPfgTZvkLtrhpBn/QPgGiP0KvjfLQmI5ikNX0xxII7oX3FI6jNxQJM8
RVAxB3la9ngHN9lZFlOr//hhdJO1aovNDBPkHVY309LRoHOixzPhl/f78bYrBZyaMhwoHDFDSJhZ
l6A84KufL3blQsKxoyVDHw5+iBMixlfMMQ7PKoXBtG37useW4CGCJUQVhO1QwwbCXrbXouAYKvMu
HDxnm99cStYipySHt4vv3mic+YONXFsHFO4ockqgnaYVTF4IcvUx+6HCSB5UPmXCbq22kdMfU0Ny
xG1lew5VFZqoFXqomUCBjM7oY91l7ZHJIq+kIbYw9sWu2mt17bMuPrxCtnghekrMpl7+xaDr95/Q
crBg9/PfhR4ncFOUNVivqy+7qCX8HzPUu3rkpCRx3gsu1LXPALpyUPh/SaAA9SDNBAHTR/CKeEwR
KAsSATFycgkSCvdg1ex1aRVZ8JM9jXupQlkh0cuHrt/tDWcoW8v593cQ6NYCbjdQBJapuw3UJwAx
Ykfj6UFyd6KO94ujHSH+HueLzKl7yvAg5ap5qw2CIlKM/IHjOVioZCGv8GW94CqMSvPaCnNuv0gL
87MsqIoL+lZmolX3RDwYvNd1Xb7xRn0K7PfUUj5gLL5vOfp2YU19B3qChfFFX9sQ1T2ZdN586RwX
+3nk7OAVOBJ9ZURxs/60TeW9PVdtJ5z6nEb9vtMEbOn0CB6BayeEUWcMZr3kB+ITec00nQxMkVRI
tLHw25o4+AoxLfMVmQG9RolmXr8U0Wlk2Xh5YVnqoP5r56+hl7DLx+JwC55/RfLi6U6zBt00ljLi
Sqk/9b4bkqf3qnbtyvC97k6nZdm0mi3OGQz1G8WoYFcUlS3zFH9IRvMomZ0KkRJpJ9e7prqRdRtM
Dlnl2rtw3UV5VE0M3UGOVPbEnScG1+Aq4LRpNruPFXBeviCZbA6DprDxsWSDjt19NEWyUIO9hSVL
GBoSwRNNZ21r7fPA0Yz3xKeG/29fdKNjXo1/nDqtX1cEnpY5eC0clroa0M20PbO/4XHjRhSDHeL8
Jeadvs0ttVSf3U5mxo1FsuHKe/09UAyBmfCVWNeAL0WbKJ/MiVTUduyQaCeAq/yuIs2q+uRdJpe6
8FwET55xaF5uYL69eGN3SmrSOZNcnn1MMC2z+98SfBvA6xcxYZq4253vhy7dIUgyX/EkmJ1ZoD6M
OaL0i40ei8cP+k/LMcZclspbK8XiVUbZMHuFLxE0QvLK6OfmuQFVii+kNSgVTt0PGcpdEnnGsl3Q
Ep0U4MwC3j4snG9PZVPuyeta9J2OmmYcQOEswgMD5WYT6XWS5D+g1VFyRG5o3adpN6vzE1wONpAh
kJcTWvOWtVWuOmrYgpEDOto/05U0AQUfddyuk2DOsGOGuMjnpuz8kyjXwQdZK+38A1rL3WnY8I+h
pzzEOICXNVjYBQDiSdYX5yn+DaZWD+4+vbD3I57GOm3jpM7CL0viKGGflD/wtV9kcaHVpUcbh3iA
q5D1QcAygO3QVk5Kz1Q+sAGf+bxwt+F/75L3PjGJxGklXV8goIqSRhX8KhBW5XqDehrlwob/ycP6
qoRZ5GXlTLLnw9WPCk3Foo6aeY/iEe9KRRNw0XUcu+bQCH7azbwtXBV3CHgezxobRw52Oaa+UfAK
Y9XwcBFn8V3zizxnY5lt5rLpUZzvUMFzea7cELceZptEOaQFo/avFCaLZ//U2zqNfKY0+H0NWXr3
3kUAbqGxdFwTf0JSRJTbAwGuyHfniSFoMlgpW0RoVUpxFtqWNBhjQ1aCd2iSIGDG29XZc9gG3lJ/
Ju1uO1bFHmwVFGFL568H6HAdl50Lmc275sxEjSzlRadkzrxBRXly9DffXx9NJpRanXKOAaP81Ngl
hlnCHNR+XRumyyj/YLKrxAy9VHSr9xVV8YtLAqrKrNPiLA7I7U2FURPn4UKgbautz31v/UMKDzHQ
36Q2HUVMDTpgBQFZfoduZKo+/71IXVFxMjdY0d9qSjWsxFPReQDSoKCOpjsshxzjCRDyHzC71spc
tymW/mpfq48qNiiDjz4pIacXNzu/g9Mq6o710CDlvvEki0ZYj1B7tGw+Z/uwBwXe5PxNKjyzs+uw
leE0mX9BVY7UQGsig9XiCDboxies50Q7BfwZoyVHwRVYsfJJJR7BjroymjAFNHd/LnW6qoBrDg3T
A4RGJBw85MFr7KSc4afIAVraEglBz0icxauVpUzeEctpN++iP5Sqia1oz6cdJocOA11Z7tjZ3T8v
WnzVazr1TMzyVjD+Z+gCGahOEitR5kZE1HohqhjrJZ6KwZMCmLPgTA3ryprDYOB2VrpynS7FVAh0
cxY9m4uWbchS0UcFNYJ4wy2ECWr69P6cnGVpVQvDkIK35RjYlSwdqW0ezm6x/aTpZRbAUlEt5gaL
aWLLlaf+sCY+pyGRpSk+CnZT1usR9qGeWGgcbqZAAMW2ATzSyIeOJ7NhhRFA24dVKGSasI9HDuYg
617Fsg6aZx0MffTSH09DCI0xemGja+2meizuCDuTzFu7zdGADNMpXOb0i3AUBbNR2uRyOjpIJPq8
5CHl4uXUrUMleJIDkZcKgpd1UII/CNVaXgycCbHFICEYPbkgBN7zKGM6qe4WWWz/Zp/6RkaXwIAV
sXA6S0O9sao2A10/GdqIORiErCyX1l//nSuRFcgTmqZhxV9SM6TRNFP0D5VleEMB0EQtmQDM239i
PE5U/DtKafYEIZOSnwerLnyCJm86GsAG+wLQDHz67vVS72w1+vNE1thHMDJvUUaL+S9KJRcZhBjJ
wFJT4ZBQUJoXyofcmHYSpxlDbXW/2kocQ2LcjuREPCko9BqE6KPEnzFIiDFzejblogS3KMdO/qxS
Ma1Nq6yA22MR9dJKme7myT2FVcIOPhtyUYlZAa/9puEhgSSYpicerhdmxrLMPDOs/Xvf4QFzm3XF
PDxmR4zY3BxxKObpxyq2FTM8Iyu8pEfyQu/dNBnpZWoJYsv+DICBdtE6f4JxhzpL60/ZjyZ/01uN
PR7qg/jOfd4DjIhAj77nKNzHE7qq8OI5U2G73GqVBpx759rLXcx95YuXeQX0NlwM5TdlFYjTxVha
wpqQoTPL0tAZvgv9W3SllwsGS/BZfp+MYOjb1G/LHeXeR8sVpiOfxv7tEMPmj9ve/meaI5eqroSb
ro+ECa62OSgpsSRHSNY4W+ZBz28gNIOt6vfgibKjHPqHUDc86Z4Yt6ccNgwuuB/JiwQXXIBSZedS
5m+QOYxdExD6uoEvP/h9K52d8cp+f5k4wxIZ4OmRVqi14BP7fzI3yFmk5TtvknLrgbQvIeEU7LSf
QVh003CyJ42jckxxQIHMu8OXvFOZz0hJLPBrv7dR3wmmhwQB1Qbtxvuuv7Ad8WSeUfPswZx6PwmC
7I8pJQaxxVp0QZGyzvknividEVyJxE5/7tW+DMmuY7dw+ckA96zRR9wDW226JyLifjhJVGhLrB6E
HosfjoKVWTpBY5zLKFIZcahW4w+EPXyd0aPfqcc3Rc43NWNSUUjS3oyZzIuIbnQGbIcHw06xeHkx
9nWSq7a4Hkd3ksCiwsKia0Z6qxzF4sXMKOqLtp6HdE1N7VZSawTi5XfWrNMmni6vhHjO62gQBp53
LhAOVkE+pdcWmZchTUxpB0vT1f7/KxZH0i+X+CJZSK/LIEW/P4LTYOlPbDzAdLLItIHs7vqQCEOC
NrGLfraiyHy2Q8sxtaVM9WJ3qUUVxvCcTD3EVzKPlCWeXoe/+Ol6cPLrQ57yUy7Wg/Tuq1OsIML5
wp1CeXMr/u6lp6daL0cSm7Xm8o5GiJ7upFD33KcrV7x1MLMnE9S8PgdVyhK/6C7BO8bMbgeVR+Hg
OwPvKCJGOBtB9Mflhq/ouez31MjjxZ7dKDCrEYSMyxz1rTGywX9VB8SXTtWnMjF/hOYhCwsoAoUJ
tfjbw6R+Rirsqba2sgNNMQxtxB+bWKyplTN0Fmrq6qhkbs+iLAbwSgsgrwAtRvRZtvQ5axOHqAtW
sNff2dEJD/0CaO5I0dDN1/Cv7dWwdpkPBhBd2r7Kb9FjZ/AwdM2+NLXnN920qG5eB1HQBc1UrfqR
wkb1vKF094oQnMCq5ollvrPcjS/ZMg9F0ta5gDo3s6W+fYZZiVTdHuvthRcj7BfZhK3HeuyhheBq
o2gFfQT+2DdGu045JPgaDW9RaU1GhH5NK7A6uDPwgPO5zSmbApVabA7av2NirvnWl/oQmUUeIj1U
DLY1rvFnC7OEtiRXuL5amRUqyxMohFOmZWyvu0ETmlI2vTQ/B3OQob9qjRduzMD7HXV6toqITHcW
Cn623PZdhq48QeOVRVOk2NUKO7oAa3VgJK1LJRuZoegi8+xbL9P2bmXqk7sfpCWoFLv9KYYriAbb
74II4KUelitmNFtUMsH5LBq6WE0kM+ejwX+IzxjUWUdAa5W4D7K0LcK4s6v9iwqB409EZXOqRxgR
khEy4Pbhrlt/LpzjfIx4ozLLRjAyjhQ7E4+LbmTJmiQd0XuCCxTZyrSCQioXmn0PWpNNb+V7ACv5
hwP+oDywornfZSyV8lc0mHNtGNPWNit4pRwAHTTB5drl7eaRovsS2USkYClCfPGScvOMqYpqiFs4
XE4N0wIWwDFC77AHNTk06AqOHtOfzMwCDvDCrd6I4xMdmjvSeVHibD5dHdgDZwOMOdverzb7uX9k
BmcwaXSyzktSHztNnxQVcyzIXrcOVfCVX63dLVxkRHtKs3hZZtVXf1AmMoSMR8oXWXrfaNObDa5x
D91koWZ0BtAc4za4ZCWhR0akH/jx4HhtRv1raBdJ1anUrPdquN9xdaSmzqpTX5GCJzksre18t5fy
PifiCHOQZzjlulgoQQhKpaTinB46zydbhG4rP6FmBwwddE/rmXjxEYgJ+hhIs8Jf+dcL9CZZfAA4
Hve8GZHWmyKDISgm1vsFMH5TLA3V4bcqmU9H6CS/xEBHWzsgCp+AcPfwdYLcNfsmwrnG9YVRy8Yb
l1tAigtooJkDTJlgEQRRwE9V7NTYOJXCfB4gilqhwfnHqqFqe+3ONP2KH5k6tDFE1M5qO5s1gZga
cAsr43jnNJGtvKZr506ghFoBscL95Ijp9p0nP4k2YYJ0ldsEwW3LikM+RU8j8ePnGt82k1M1jHvf
MRZpqcrfhN3yrjhjWcC6R6jSQ5DI/AlDmmLuzyLXdBDnpA+8u51LUg8lUEW8GzE2jWzkY6gAORLC
Gsr8EcybHnkqgFWnu+5abpbm7oGVod/jYdkI2P6r77B53CmG2s9iAMlExEaodbtZecG1BIlNk5Bl
gML26FxX18N1+irBcyY28+jrs0ZaH2g1O9KET38izIb8yG+8XXf1TppM6ozAPXxAHMHfkPeYyXaj
7vfAEqB9V33X+GFByEVtw4ooh0gvUKR8EM6Va4cjIXDN6Yy5PV5R6Hmxe5Zvx7FB3pmSCoy8SkIT
L4TzfbnB9GyrwXgNEYeblFSOq0PeTjq9L6vtxZiybWKRAbBK4+vk3SPCPwLfWWRwhITua/6f89ji
CkKdyd2GwpUml99+bYBrtZiW7EI+shpom+SkbaZRgKRTQQ1H50igHac5HN3wKyrJUIEX3pxkpNjI
3SYIa1FahAYrvbgJRv81u5fQ5ch3w798Xs8csD2+mVarjMQi4DwGrcuUQozoU/dbUiUBfD/ClPgw
T25zNLWt73RFkyd2MvNMqKfoOytM1mENNJ9d2GWjfUrXpNSa2N71BoDgzl4hLv8bjEUqJDtd+j8T
Sm6fy2gNzXrDXy/w95KBTTY/3/nWsGwLJ0DcmgHL3O/+prolGOlVEM8cU0wJsKjlZ7FX6P5OqRqX
jIwfqzYvun+5X+ugjqQqY/tHWFqdjodNruJ5iLVwt80i5C+IfGRfLVWcpObjDJom8Wk4KGKARs2b
CdWSW4vBzgXa0o2dUlUk0YlGIRO30tl+Gm/tEmg8QUdYfe52H1vQ4XN/y3MQAOI0BqeSJxU2Rd4x
g6rQgIuRMa1Pw9w6Z129FtSG+wPoa4s8FdG4cNp0IyNdpH3uppef3VMTX4h4vSKI2URnmRGcNKWm
EelKvqDeWDQ5o07Dv49wDxLegfwnORSYCLoHVL+KSJ2FEk1hnXiS4XksHrltGsVoRHpPRUFq4vBl
EqP3RirHIOvGtDhc+TCjK46o5Af+HzHKB5mfwIGEtuWI32ew5zsXIdIZPgUBI+4sJo24jc1Yiycz
mw9R2+fa2FDNJMiE3Hf1rs4hYuw67r840UYpgywF9z3+QFQOTIE2JAVvTEi0444z+0XrQ1njm+Yb
6bvXnmsZzhQK9A6khPImzNd1ElTN9rcPU3wr40KO9UTncDAUEy7mIJAcB1MJ9cEiz0H7liN1Ff2k
GBww9kKcum1uPaqa7r6A/mtmPMa9lgG5kUvbkwpDVemZ8iCNBGCXKxatdx1SgzKyz05dkJbBYR50
yTd73epVDyAi5xXshDRB2wM9URgPx2pPTdMmoO2HVFqd2YPTxW37JXbSS8Nxtn3q+udWq7344JGQ
rc2xwSgQAKaKBQ62k4qtfRwlxlz1252jvlOgMxp9cRGoDbRcd/1IeyEpQZlSjTkWL9hIJibaYYmG
XvCii6hZJcPwQgTV1yKrSko7UWJBlFtHhlDt5Wh2LQe3IDySKdl9TLWZp6vA++GakHYh8RYTlu5e
aGsLRnz07nQiP7N3sAj6yzUtn+MZBctcmc5rIQr2i23m5EJPyyAVn2q4ZkiVPOl5cOJd5uZ9Rwz6
ZXYamkiK5Ymcjdy2iTX6kruCpdd/I+AgfFqTe+ETGHIa3BLXCKlUfTXY6rzQgM5ng5bvoXo/er/o
PZWq4oowV+AUTUPRlX+7vbwSzkHVZ2frUny+GMZ8w0Hdspcacowl3esGQBfX2jC1duZOPsLlUss+
FdsVHV0pnN9avQN4RvvfNr48UmT1fGe3ECpyGXwcppr1hXZjPLTS9MZZcuysmi/AGiBmH0qia7fE
SRvBHDOZWBrCOm0pqF33zQiqkarnhYm74QNnXrBj5YBXj6gmy0z2zvv8tjDm1v6cYAvyVpLUnvMY
9+bsYuD/AlAb07mrtnEVdsQgVKdHVOpGWJNOjLGF6TRuKg4o2qTVuCdvFOIJKV/IIDn2XDvvARQQ
zcYtBqaKIhLQtPLq730IDWASFtyn1GSrfjGQFkbbHBtyQYkOLQrmbNVEDEtciLAfS4RkYEaPybEz
pL3cDXcFUkq265/uekBouNuhkUf/07L+Drefvt+DywufBAG5/YM0Jfo1Zh2BJmI8a+rS3Qy1xLP6
a68NdVDXuhglw1twDAFNEzLz4z61hT1iuD3BhmSOtKXMbdDZcA+RcLnvtXXRsMZpRb3I4D0Ax/1P
sj0OVGYznx/WTLOFfYeBIKUE9qUz65KGftp9RGHDPG1bh3OTOnCEQmSmu+2qaFex+O0WQsvV1rf/
cV5T+dNfBbuG7g5dOCYKd2n0UAo8AnbnjfYpgkn2RMEE6+GTcbWmEoQYXDMNSQVbH0FESjBRwY6X
KrcdtwC7hcp/r9XAToYP5r8Y82WWrBFP91/w1sqEhYxcyV5lZu0HDNXlkFVj/0W5FmErb0OvALNF
3F4UQbiSTLlZzAeNiRvvXUNnEGXLGQ8OHPZAiHWx+R/QFbVqiMUu9CfQjYQJW+qyMS7A1MyTIY9C
db/mcuWoG0r4MM90qVE2dwjk1IiTZBavFykTHm3zB21Znp/ue50CVNu5AugLFzm+VJSsrJ39uw3S
vfZducqHY5b0Dhep3EXSsc19YP+zbsOCXvy9rrvLUsKyrSIMPQmDqmZiyl5i3rbQ04BiVcrHsHX4
5k1DeRYTmna5c96gG7I25tcGzhEexN2M49u9/gD85UHR35clsF9bhwdeJWvWpTWakHn/tRS1n75q
5G+0R4QyD0mpsWsCi/OXuJO03zcvmUBp28sIV4jM+if2AMfH6xpMjHFIhsNX/C4MoHa/K8mkgWo9
ce3lUJyUyjLVEvRd/0KTqSWXXQv6N91WtCDVSzt2zFmT4tFlfb0jTLYhPGO/BnJPe8JphTJ3yMEB
L4W/ljM+yEv9Cl/ZCvg4oAzk37WIEZ0zcbeT1ZhJ04milxWlGBCiXhULYM38Z769IXG25UXkn7Jy
Rg4K2OE/awsmdKFKPXO+Efy27gYG6wg/qXM/qpUMaOAsGxjv/b0sqp+GQcOYZC+N+WvTZiIB/PEe
YIZEB7lHPbRzbVcY+WLBtTYfX/368+R1te/iOj+kyks3IiH73GTqew7suMHv0TyAbyNqBM/Duk1/
lheP2EWLxn8k1/XFP3otPSATqP7MV0eDK4jwXtDY8LKbxYcZLovaF4CHr8YA3uCDGX4Oz89lnPaM
8ZmSIg5N5UfBuIVNXOWf3x67DYMHmt05Id/ylazPM7ADW/RMlMrAMnwdA4AmeFsXDVDf1IOqT2CA
7LOUy/uc9p3IYOvBSaC271mK9KXjOqcAWZRjXFagAxsoakVheQPlP4IIoWUfwbB4Xq9gA/etFMUl
3O+tQPZ1fPlL+BlKf+hrb00Fqr06YXyejPc64ED1og2F7d1h1tVaSgh5Wo2Ujzfx7UKVPZXlprer
nHdTVeVm2NWBvVZ0H3OSchnRe7k+3HlPxTIzCDTYC0tEsqqpXjx8Iv429887hgeCsd/YDNwGYk5v
hResCpc/8JtH6V1zQ9QrOSVlWOfMIHjhFBjG0lmXtgpyYgTF1N7GFBHeZZQwsOizAz7/jjuQb8hV
32umm3C0f3VHfTiB2mduG9r44Kih1PaRCGEloOkSfFTOBAuq1rE1ASLAlzdxErrp0zpgcv2w2f7C
MrtkAv/pFw3tYizERBHALqfytkNrxZUmZ//Wdbc725iji7ryud/nQvIEwFxf+Lg7s5JwcU5v0lwu
58ZFm22xM0wfTVSLlKiI2qBKw7gacNbxhV7sukP7nIfOgD9X9f76S0HZqyATu+nk8rWEZHGQdFeW
nasUvLhlBWGRSv0e7PO48N12hrVZHturl4zW5u9+Cg+5/PkzXmVtT6dwZnjl79zhHESaoDgevtUk
GP9PK71Xly6GBbXtflZpyHbCHx+m7/n1NGv6dIYd7NT5dlCnUryRi9T6kzcin71SjBdo9Xyrm23A
CIxi7iz5EcY3yUykgY0fYCUatr2/Skp9jpb3Ly82D8RIvvtmPbp/+9TAQSuwLrBc9G5nz0iUzHDq
+Z7hkrD8ep+8tYf2X38fFuf3S3tvWvM1HFkvKPYmbNvhF/4Ax/4mykSE+59cg8WasycZo7MBW0V9
Wnw+Vjzl6PY13xkV94FBjhp8qpd6k574EbUsofbJSlXmyijTbsjSCVuRoLOjADQdLWTAHl9dMRfo
Lqr3GxRY29PbFrx+NK0C0tfJMqpgRgMKktPTG5sxCmDn7mg+WPA0lTO06wjWx34VMAsqBq5TJUpK
gKISXbhTZxLUuVceBUC/oL22svoP34rqigdF3fNIl2iPbQj5/yDD8ScSkAKNMsz03+TqMUGZeFCS
UFbBt7jhdFR3NcBKvQ5FvXioxMcJ7+N/S40Q/Bvi4sKZQkcmZlx0aYlgMiklf5hiAM8FeBWVFU5z
uVTZoB1/XEFzlH8mlO7vTGx83db+Gsf2BfbWUA5pKNFyIPjlGBEGlGleuFChA+CRCxGsKE/mz/bs
2ZWO6jOzGyvfoTC1+Ht16MR1GHDSTlkqQP8ucpIer1lbJkfl2q2H1LqxKHqD0js/pXo9gidoOhyo
Mg/aJVBqRFU7DcXCPNNJNtX4mghuj+3jbMjU1lRO+wFP3JVqz75l95jvFTRR0RRcbvXzKAPSdiBl
/vbHXcpwaiG+TNhBPPWI0cPaMVEr0LxJ7W6QrMY4bZ4ZejB7KG7wE8vimD9I8fcQ34wMGu+Fmumw
PXKNUpkDbEYEXPyPUIjf2LvG/ZCFMAurBPRsBy1CDfibuj90xnJvGKCV2VgpGOgtR0bAYL0jjSmH
6AyBPflYigk3sjzG3tLdbcbJ5MLK91ZLyDokQr4CV9CcYiOcPENaz/LRb4KjBxPkfzBz19Fb9ZDV
8Qqu6nYKFabrHxnDg26xMSFc/OShXk8wM+wvJkYmqEROb2eOYP5WqFWgx0BW5kODuuNV/gvlRS6B
lEkUtOYP9CZRUgYcbO/iLvTDxbTtM5CBkkuzYydOGueh2k9vnXbvm86dOPRoYoAjU6MvMuUTQfE6
Cd3MCWwpEdpiWRVfvJPET1XqlNFwgkBNxHPYaPu0RPsuWghAYxNr5ydRbGJBQQ6qnkR7MMt+/VNL
lrf2od7wEAjLlwfFisW+OICgByULugmFsB5AD1ogJ2pzkXHI69D75eOJ1/coLWY/r75UAjUu5zRC
Mu8P7mZ/mQRq3SGl+nBiH2Cb3qzwUIs5mA1P5JIt8M987rSf6ueG7+ZZcxKws4zFuhWXx2t7bBNt
sm+5W8tDEua8BDvSznDAp80Q9j52H2LgXUx61QDSDduCE3orjepKPTHHOTC8pM712QNcrPCNzlv3
rPIehSCZz57IV+RG7ySp6GQ7xNi0KQqISNeBIEbRPil84I+aK6kkJTOsiyvFvpU9aNFN9J3IpmPT
UPkEi0DpJlzBenH6zrr057vW8csA4vl+Yt3DNkup9A5PjgWylVOyKxyY6nOGlvsh3TxUKwDs2ejA
1qKOhNilVphxyLHOVesFLvDYfDcEgaoTfKY1JvN1z77YA1rudi+PabMU4xmqbyvOvrqs4UN5nFZ/
U6VTMU+e8WtEF6lpBje6IVwz4HTPkx2O41764SpxIdYFNRcRgf6uXlof9rBJ5ggNXIayyNq2MRhi
zv7mvLIHbB3wueUND2pTfs9sKxx+oy58/Mbvtndl4ofj4tlG3hhgIWTzIrF5Jt/TYDNayp/NF5QH
mHUGloKDKYlS5ljMZWnqHSfJHb0fgDvG7dpNOkxh8tPJD3PHS0yxiEBFT0tI9i7DSAkP8+jS7VOc
KMr6NzpYlEghvcYrcCfkPrmQMi8n2c3uHGu4Ag0PR09xhG4WTfKtWZVsuhbfzi5tJwpXOa5dJnu4
9OTfAL89Q65MWIsHxtKiKZ2zES9xXMUt6EUeXsxCpPI5S+7yIyeOYVbTvvyKofCHWDFjrGYA3T2N
fANLXf4v+Tw7Ed+/csbHJnWIf+WHVYSqWOup+ze0bUi9F5aJ32WJBn2CiR1rBgYWxbosxVMtNn59
wtecLanVQA3zyprwnjZR9tMJL82f3kGOskWkHkdgQdVicokEaerbVcMJ3mmJQmf5UR+If09Wqj0g
5ceyT43SFJ7UUnw91MytkAexP+i8zob4DNibp/ghNwa4c8uWVgZpPHQmKybLv9QE28yITOA5jWiB
tW80tJ4JWwncUb0sgLFgJCeRads9+8KC1uo3odyaCAYy90gTk22q7Tqk7x+xQIHqV+ms5I9XvSQn
g5zFLAUva2Qi+yInxntrkbDT3bBMHmiyqOX7rODyW1fDGLGNaujdXEKP7QzOym6ib5C+SfJ8OcHU
7+XUEDa4o6wE690/CSFzXfpefGMGEq/bdWjQdgDlYZAylKGBcBIXqnqvmEFAmwdKygnbB4+yfPMi
kK1Ml6EL5qczWB5SLNcHEihzn8XoOmPKKA32vRnN/JCDQeQFhI4983G7xEs6/7/vf8viPaacAOMq
xuCglHaiKBIxW37IaALxSSEvc+34/527LWUWu+q7LYh0Pz4r47BlfQoKVzEzRddCpQAoBU3E85bg
XsbJZYxNsXv93nn4dDxE7fJp/sqC5iYkOzdZk3gkc1KAIenTIQK82RUFwTJX1B+8aAUZ0Wm10biD
ttlTyR5SL5+a4WyYP+pJd/QMV0yWys75w1PPmlhpNdZum+lwHfHyIpssfLcLCRwYlKD8Jc5qTNTJ
SM8NLRG160HYraYbQJND9iXeACBqKrBfCeEV8Q+7JU37TtZ8kcOuMFzodip3xUVbAQl6rJt4ileu
2n02uzKe7UDnbYcjWCYO5ZwhU7DL+upu/qusBhxgX42ZnX8ozfzSVNkiyrC0KUg/mqyQS3gSAvHX
bDv+wd0K1M0e3ktlnijI28tBxv7tQRyPlFOOHSXfCQ2PnVPHtnRRgyPmh1iBKmHnMxLfk/zBAWiO
0NZDlcRRepL7NmLXI+M58WbptLbWNwn1ylp1CFXUtRA7i56icfCZO0tlTw6bIN3viP5G3CXdwVAs
FQOP4bSZsUNpXjRjqGWtp1KPg2kfykqmRFTIcr9tRGQGU6GXKUerxr0jbD7UgSDA8PLONUMEU/Fi
MiLE4OZYk0Gb/txAlCDgBNXJM6uEDAT5YOHjXrxOMlN0IFUkC0xJNbuHmtmgFWY/1V+HKAAwGBTP
Qdc1HhoFloqH1z5mr8ydvAMunUKbXkNe/dpqGYDK1NICtaj0DgNN1l37BM7mhEKNXu5CwFgA9p5Z
Dr3fbMCDRmSUMhBil/BLm+jYptS6KKXpMhohp0y3cdyz4HhUMWte1Zh6ZGCopSppl265JpNsP+iA
BZ9aR2R39gVTbWsyQ/LiquT/F+1hwSLlRziU8R/CbromvfCXy7JU3SOu4AKndeWnTGPTwfePtNW0
TiWyenTsx+GaBUxJXqagxbTBcEDeXwuQEoBbRdhGPRRvEfx4BSsZL1+ZvuLNhm+wNeU8ovUdenvC
awZ/nAiqfJhMHjnHQh2k/dC7pYTaybeMxfR+YHJSpeqSOGBfjiBuKUCQyWzKkxivmsX2LXVDy7un
11MaZNlY1AQ38vbs0h0CkWCyN6YEcYD5N3WEPKuvgbM3GuVhtJg1FFSGKGcMRMDG6Yuzeej1D243
QNoNgkdBijfuC3cllssKMvq1EZ1CVm4psvykShXgaVylL5U0kMidlyScOC6BPK9/CCpx/A/O93bS
r60s+/llZLm2rAmWWwxPpZ/AcBFD+cZgx5TEmi1+9sU7yLZIO+osO/KiNbZQr21PanGc59+98QSU
IgXkIv4qEi1U9+2mY4UY2O5aR6oNL5LSaeok8QoXJIOYguXSascYFuZHBhHHSwH0tsqMgUgmeY8G
opgysJJgyB/ehoQUY+5OxlgmBo/hTdfBL4kAFEzm9+TeTFUW6r0pdkHWObFhZ9C2mlxvixm82+7W
2wGrd9HWUT+uz3XjYszvo8kq84Hj6o+8MTdtzGyeLcaQT3TAtQiehiwoi71219Hv677r1A93PE0O
dNabbJwkdDd37yqLvYaUA0+KADDQAopALQv48wOtiZNwKPJ9XVyx4qAUa2z43mmX6LHoL5/VcWGe
FIOZsNuOdxPYxf/45YH5Dl83PnNzXZDAl1ph1caD1bDMIYHdKCY9ESGyNXd7mwGI/nWHbrlIyafq
+9VScebXgFXcdkK/aY2KVD+iX/W/zxu8VVdsZZWW1xliOAAwlexjt8Y6s5DKLBs5q+OrvxWvCGNJ
ydG6olgG8Ta7wbbKJLBl0sRkuVrIqC7tDHli/p5wGImBUmdzxNpvuCns4e+ZgX0dwDPII6bvJTgZ
U48aPvebWV66S2JSAlXliDb8M11wbKHMIAk8u89BPtYe311jAUcSfSYh/EiOS4b1ajEnSqMdAZIS
hoyeGzt70vliKb6d9U83oGtboH/MOvT1vOtwmDoi8nIpRStbXfXixVHQyutsMPJ2kwFXTVY7Ani1
N3ShIojvjHVJvufVz5ioQUMphWZ0FQtcdE5ArDX6mKUQjM7XfJPlZotcw6HS+i7sxiq7DI2W69CX
2l8pEvuxteVccpVQB0/UFnSJABf0zFCFxer5SqE39w7ASEB4tdlil4FsHkBVIyAbnodGcspDCIGN
EVuXUE+R3I3+hI4WsmRFI3pfc+xK/Nl8IBt67i6iprBnhBKcNga5jLtcUCiNSiYjbzpCEnW+Q96u
wbp+DRUet4W6W8gwiqFJ2mNuUqSgQVwrtSJ7wPXv1kGLQQ5fNV5Ye3bXFZCo05j7L5WnhNA5DfVX
rsV59uDP9Ao00b9+DytlvVXja/oSW0Tc/iOlh1AW6+sB3PyqR2EtmcRaL+8eFlOgElEu6hRZ9RlB
wYhB1rRSWNokWmNaynbcXRgsEP7fauVyFMbpsrvl9mbn7etIei3MmnOQFsms7K74alogMT4S5Be5
hZGCDIslP7rbQXESmdNnYMCYd/8pujwuPXzLqNgJlX7cJhMuuR1+zxZ1IBhtELjsCWz1XDt8zPnM
ru7R3wUZ9jVR/7fK9VwWhBz5mbHJ86jQgZQXFg+doVHrt4RHMySVMMHxAOYvPJzDiLE0FnZMTi9q
rfXFUA/Y1s0NARdFWVLc/VWzPmCKe7YYGzXORouzrdg8lLt/kjLdCy8eXEsVwij4EWsNaDF5Oja8
WlGBMXlqKz+c79HDbPvCNIZxx30n0eVWNQey4oALkCO2cgrWt6TebdNOFRxMJMQmmP9ifna4mjBd
sXs/2TZrmK5j/Z3RNZ+xLZjFrrUjNEZ7tKV5Y6gjnaou5kWHeN8hGWckzxXOzuF0nlCmi5ZdjGbx
yBaOpwqCr/HjTlY2N+XeI3kfc4qsXljb3wcEqSxB57EjvLDVxYKALvmMjwsmMx5Nu1mVnDHzQEpD
UTaJ1hXl0zrFYJ3Yl7IKHnqeluRm6K6H287kBUFYQ3m7SIxaCUNkAFIhM/a8I3axciYsakbNZE8W
7cS4y+d8Cbrj+lvyMfXnzWP6e97B1+5qH+j+7DCXh0DXObcYytFWIlWeQUrMls6eC27TJ/xOv86F
J8qJa8SCQDcwQD4SLt5hU8dPjetg9u8iO9twKiMjAqQXbf2H2v6/AebfLXwDnvgP7I5KIOnp/Dkd
4CrpFWLHflhN7rZE3SAbYqh8ofR+jJk00L9Onxj7jVv7BJtegpvpk8wOnMEV/uPBB2v/malrdSkF
hy09z1HuUK3B2nvJ+GeHqTN76Avg8QE6zxgBqxdFBhw17ef+OZIk4dRP8T9qs7E8zgLAOffK1Bk0
HR+RY7T+8oRLbL7R2BzkifiCHtGnq4Y9rKgvKH6cObNdZPhSmN52gphj0BbRNnSykHYwjPWrN+yK
7ncxuif0Om9G12m019xf8vsl8E9VT4HXb+ljKEwAf2dZ0u9ox/Sp5bE45sWSMjn0iUFBBuRQiKwm
GkTxmhmKed4lnLMHYwL8D/KSpy/UYRcaFn2v92wqRVCkNYA3FAWJRRUUf8rprLBM16hAQo8XvIlb
/WBaHGVsPrlN7XoJ8fl/CJkq1yRBPJV6XB/veI3KdaJXaK3vwnjyXBI4vamIAW43BW++Ocy1UZJX
LkshUW8W7mRO0s+Zxv8ObGRfuSK8hrOKnRehW9MoUUIe9O2y3w9KF1D11tIukLAi0SnKEa+t4OhJ
j5K5Dcocf0rgNaIBabvxZJ0eKSliy+VupCcLoeQsRqE4gjrYklzphvAdxSoBRJpwzU6Wr2cwbT9P
laIlWHdnDtDJTRRQ8TEm5vbOPm4uP9yhbWR925dPvo4t7aU52vogjOH4Wqc4+SIhKXw3xnmINJQu
6j4QAiIfPkAEixQZTSms3mpn1C/uIJskbmpL8fz1UOj1KEWgmGbvgHEdcMF7OPTzLeEXIPcrdKTf
bBx4xAK+EbRMYP72K/ch0s1R1kqH3fDV/nw+KhpOzIz+hItdSqHBe5lrGw2WqEDkTmOic3Nm2eaQ
XJpUPqKg4CDqvFUv20iIe75tUCJXcRAXJA0i7Nar2TFxVvBGga1x6G3olqQsouxUwaMuYpzrR5Nf
c16nbmFvp4SOD4Qxd5+CXTlgsIuQHsQBs2vIq8lvOp+mzjBUbODEq/XHX8dfnZN4GZw9FnW/Bu2k
e9OfY8Fa9HrlsDGa+z36O2l5ZeaZUKm3AYKzNPA7UyHX4dMmv6T7n9fTNfsGeU4U4n/K6PBsupLV
iobx8xuAc99RB9yPWXj4PvcOe5UGAnuKH9g8BXcSex09Dsjp6ut9+qTwExir4wrPwrDteAV/sz7+
UEj4LPTSplJHuusoyKJPVKRnxtp3a3iwfTFq+92kmGboBpVjEbYg7FNaj4xy2nDHXsQ4RgSuskEP
a0TRhDe3cJE3Pxh1bU7C9igcpfEdrBjFasX6tAmYGiOmxlne6Z4jxD5KIoEtucJnfoeDKyFsSiyZ
e0sg0Y9eYVA962wUdqJWjPhxi2isqVNRS/HiKPtTw3YgPzumi8/0ooYKXj6BlwTs+doRP9lGzaHg
fC77F7sdwQRDy3JKf1GcosRQEPVQZVwDYdksqYjh64mA4y8YBCnI21poxjkAqIT9FgPMMJpzOpR6
Gal3w6ZiNNMrQ/Fe5Jx1HkiPuU/G9YPRle8Z0NBL/KhlIkYPeJoWRrQo9c/mG7Kq6d035Ytf72Vd
iS1REDvmQksryidJKWmrJ7dnkan/UmwQloJpK0O0TTAacg1zJkeoIu+QSnhn6yK+3BTM5kfxUkZE
mFxnWGqS8k4v1WUttkd0gDJ7q+3EISGyIrwRigD2nHjEYwu0SKMqQDBYOOiCDdf31TcMTGlAAUdX
cWKmT6tri+iXe7IietXRrUs8HO8zHDWqqruc8fsrLEWSc7acIzkTVP83UPZbUrU0AUi164LOlDjf
2TPq9IKOKv53anmLudf2Fb6n9p7TfYcKi9Cd84Gck5KBRWnQFSnD4hoRTcW7E+dOMGlJERl8TG8v
TfJCOUEwtKjzlPjCewZpX7aMMOvzPbOZ+82ygUQ3s0/xkvupCTIxDMYYyh6lw1Bh5O4KpsX6U43f
vI7ULLhOj5b8yCvLNualPtlZKXtFxOk1FqESPqNEOF5R3dxWUaPgWqXeAKcB7gDiOGHG9TENN6N2
RLtzanYVqRu3wC2N6tdCqLJdoa3uQIUtCVFZcwVzennbDl14EbWPqlMTzdN7fkG5CG/GGDPeW8PC
jbyJqTjeyKRfvAmclkfS7OAGLe1ww0iTjtmlt0sVjI4JYg5ET+Nvo3vQ18oAA2/8fHEYL/bmrgCm
78Kc1gWFo1Fw90mEcXCg7e9uFZLyeeJ53kyD6cclg1/NO10HJi8vkShczdshB40IaFfVbvV/bQCb
8YY5D+pnEbZGn4/DBB01oKsO+oyBKYdqJ1FnX94DebVeiDuAzQqpfjUfFTvF02izMOlDS3FesfAZ
IKYfabii1INxy6W+Zrxx0YCeAyBBRqL5ufj6X+jrVbyTY9uuDp9YVM7cS0TybSUmVMyqtLcnK1xV
4FSHE8bQlwDALg1hEZQwfm3RvenvIkGluJuZ/5aiO23rbOcrNgt6mP/KLSoDBuY4+bvCkQjsIjX/
UQADK7oC6BrAL+q1OKYZ5Qot29c4PGYmCnwIZn3M0HaHSyQoStFR8JA1inGU/E8XOpGj0DjsJQRk
iW7e41i0PiUMYsMtCEslXvRJ5laK0wfP7E5KF2y304xnzpFsl5j/h9vs7/3TwygrKCZ9ej7TtZTo
r/88HQT0V/c3S07L5gHz82koPWkocEdTDX2KcP0HHmUNWtQC7EJwznAzUPh2kiNVtXemW7H6qFKK
D1fkbMYF6U6B413J3CKyjTlGb3nkyKJOYpwL5PzFK9F8W9jPQKNe0mRLfJA6g86WW4Av9wqVSEqY
gSULzQw6I6fu3uqI99ClRm0Kp0Wd2hBkX8IVUkNNvoLlu3WvjK8tqmSttNVzIYHSCFiMbz0wSx7K
dMM4YJylRDWNWZXwRo8u/+lOcNSabsg781lVqy2lnG61FSvGsm/u45OI1fq5fWt+wuTrztOp1K+3
1eFbPN5+KYkHkCEYtIVLjPDgxl5lGpQVbWJCyXLuhFlGd19Rj4COKIiYEsOmhP2RAzD0vsw53Op1
VgXT8vVUnxQ+yPl/qiTPxWRJH2940huj0exbPjmvogBHWozvxSdBwPvOKgq3VfeS5b27gTwnZjVy
XouedR7xwoLZZiEKmb4uYeHfLdJF6Y+SCwutctmMu0QZ/Gj+0zz2zK+p3d4bQQRhPwRo2IlPKNNs
6UFyVkvTOiv3fzHd0t7dZSZn09KBqlVtNW+ep7iVjuFa6tD15tN3YWNAaqTSnKzYwKtzTDBZMneY
mKu+p+UIRh59k/wHOCuAh/6CBZFwJKQpb0uXl8YhyegC4UEjaVlwk4Jx8pefXHdoN5gV4gVRnXgR
mEs1TBD/gSLHhsgiIislmSSjdgg3xB4F4pIt8Lv83GW1ZRSpzLFAV7St6L9XpPgWcx4cIuWoAY/l
Qox8e17RhrBjDYC3JhFS+PRFc1FFQaGx6arkJHYQnDp6e/LHs93Q9mmydAQMoHGgq4xWRPYTzFyI
arYqrN0dX4NOxfQCTqY84neR/pzvc8SGDIB2xQrX7JqGZMgE4RI+YeJqmSViWMBCFFIWJAfvkhRB
0sv6iXwyEv+EJ+IRI8jRQtPea2vYj0349qH1etMUszPnlPZ/d5ZOYNNSPl38lhztzhkeoCygzlPe
nCx+LwKrwUcQ8RV8KgoWYB3FDV83pigiwZoDPtLYwZ/23W5isj+vuRoazyIHkKNJfhRYbPbCYbVk
DF82yMp9cDNXN4J58J0aDrX1d7agtzrohLCEi+j/cUvyyvI3Q6kGkX263gH8eiTL3JN7uOSyxJjV
EpbS2tTP+ikT2n/CJqsaTG5h8xWmW6mhDy8F8nVtbTeoIokM1T/K3t3P3CC3uNyV4bALiRCD/j4z
G7NJpk28MpP4736CFrxRNBxvyKGoy/xU981HOPMVdZrhSqs5qzZRFuBYOigWmDJ5SaTQKjAd5qZ6
jtvzWXWYJvacu+LxOd5SgdFCDz65hdi+T4kZu0BGsZz3ET30czveB9O68LFovBkBYPwXNxKbkh2C
JnjVn2Cgm+OSNjMDkj/MydjoGZHel97N2Uo+eQ7Xo5HB2f5HpylqzyGI4koi0gTgdwFpo1u6m1dV
hOd4v1UXqxf0Tqbu5ASbqk65KFx9R0gOpzqwCrqestuS+O+vxEH9kLS1kqgka+42YRMev2hrEHD0
pW7J8VBSPEK668ZngsfymQ/8NjDkkvZ8F4ZayF+S4j+Q6lu3Mo7oCZByvCjx48OdFQczmfZelYTr
JLjy8TfJfVCHWkmi1GCcDPcIi80ngerfyAVNmmDqF7plqMnuBTYMyWeTVAwfTOx3eI0AykgUA57l
fWGMIlTp1qzEPUjj2gz3bAIX22LTy9nNkfFi9MpL3lb3x3T5s6eJMOYiUB+Va3++uac9y1ZV20gV
esunfikgx18aXp/EbrvYjVn2jm08z5eDxlvad6g5xX22Y4S0wSbbhQfMhxz47ZNoMnZLLvuir6FP
9X8aBPEN+oTQ/R0+55fpFkZHP0Ry/kKFnS2DPa8UFAI+bzjDFsW0bcffFhKxIU7SUrwJ4qyCrYDl
GAxA5H5kNpH13figWFiwpdjtOX8sO+f5/OOR8DvaB+jvmTJcCv3An1hozW39HzzaS/D5vVZpbxKs
DuUSCLjus8gfTJga3zUwV/Zri/4YJOKYplH+/yCLFFasXUDKlj925liBi2Hm7cstINbCFmzKCGlW
sQzdit/w/t15WVZN+dlFqoPd9L5dXzGrNhMLkuFIhAcrmKOHcYGLwiu5yicVsUfVX0TASqA3LXLW
GPRyY2SS5UDul3J5IrUc4erEPkfEpxmP4CDqKF/JMftHcwHgAcyH9sZNeVVlcAWsU6TsVUkwoNN4
HR+T5iRBCFoRb1HmwPVNZKCliyp/o8c/aipxwLHAfUPBuD7drbCFc9kVS2oyi1F5/QLPGS4I6vg4
bvRTU1YXkozCMkhemPPxulVpmbTDOk5pguVXd/9/8yjl+KX03uDOtlqz67NzbaZ2d3V+pqx+x5Ke
675iNQHd+D/GSrhZhhxtAwmt77YRKPu7ZiAgXu36VZDYELBanuBGca7DJrQ+Nm1MtV0EErg8cMmm
/XSn6NyCNy8V1SeN6+gjoVWv4p4sHrWofhZ76563OkvY0NnT5frZUzVYHtpzMic1pfhkBwuqHuz6
bBYLvSIDXsUXvpnMAFN4NfYU7pzOaUIoxPl2fEmy0fUmZlGX1lLku9ruOw8/QVZLxozwkPXCPL45
Cd4xSynV4cVCHFzwqbjMFq5RTasPgKMxgiG1yp2TEvEb+5nWV8f6mrjRxiZoQLtC2qIxw8JIqHPX
z1+RD1Fhnb5lt4TwV6GTbt01Oka0GDe/eILkWTo5QGOd0YNuV1Ec6FICFpKnA2uoJMJvwPioqZMP
kSasg6B5WSNg1wns3otJehLF0K6GEgu6LKaYQS4DWicwKJ7B/97uYmdKIef1Tcm9zFXblHQzYqWf
Zwt0he2SfmvEDH+oXs31xMWshAEC2ewiroumCxVKSCUtxlEtd5fcowYAgmInn3WQ2VEg82JGZG1z
D2zAFDKWMe/Rln7e1qeKt5PSwFRyx63NonnR4SXQKIN3C+X2O0zKvLrylZsfPfdUt9E0kqmrgO2+
STkePPzt+qoQwnx56M4Lv81mlgzRCeUIbwZs/kQU4R4i6D2PpmIIlAWH3WWdJ5QAr6qzli/1t37t
WyDU8+XVxBkmPS3VZM6R/YW5rqQuDg14gJSSD/5VnWv74kYULzBznDFbDZSDUimcQG5qI2iOOtks
Z8tr9AYq3eM76cvx+vdQeO+KSKzVo/joU5xu76YV/w/+iBUr57JsJ6F03w7Aylbk5rQ4Du+2Q+GJ
NZWRZ/YSK4+x4IeaQdiIisvrAU+gb/vomA9pHU2vwoSjCrODFH7+knMir24QpH6UTPaMgIpsrPQF
mXgMX/sHpG98wACuHNHu/MFNf2Ai7vWeD1g1UNmbqgvMkNDuxTYgxrHTh0iHC9gnWDCtdaSLYw3X
9y9LiXlZruTI3DU8q0jTIue0PbpHQVjodVjXQ9KzERdpHMgawIqDL9sR9Z8JkafGQdKPayxsjmn8
/cQRAe6BbFh1e4BA3KhQseY08Js7ptWcEICErcX1v5fPKGOaAtpmcQWS6GFF3XYNDBP643W3w3mE
dHw8v3zKc299lo+AvSe2i+g1BtVtdg/hy1qrAM0OEJ9wasc4B3JqcelUCOVbpwnNHGl/3Xk9DM6L
u1LXPBQdTXEaJojb/6y1iQ/I6NWWMhPVGWgHmF0IgapW469mpFxi8nAMHLRaqTu23At96HANwAGG
MQ3jj78k2mwoczWJRjf07IhLcr96CnLLyG54s2/h4qjL7OJr7ZAu00ndqxnhxF2qyUGSq6/u6IC1
O2CbRKQZYh2FhRWfcdK6JUJd3D1EWPqQwJNp54bm/PWk857uR1NM86igehQujhDPsvqgmP6KpU5h
1b48qSQe690CtpRw1SV+Gh/smOO//KTS8Ky3imvnLs0nJDQIlcIwZzwhfT5HeUcMtB0kOIZsLv5z
d1h6u/0YIzgLVcZydoF0oDVuu0+rv4PUPsFWmhpaPLjHoSoI6eUXdTjGPdHuCwpHdmMC6xJHMLl6
v3mwbyBqZ3PXB3/sLl3a9w1Unie5ijmWElR0jORMfoNoRakJMEPgP0sQ0KVDF6KlswY80wG9BuMc
oeQ82R/YXwQfQTQ6WqIDG4VK+s6Vihj4qqfxNO8fbrnZ/MJWs9QWmFxkxOTPQOAnwPSWd2Xh4VCH
LOJf6H6lTaHP6GeYQkruQdRohv7uHu8qrO8tOZrJBJDcGVZbahD2gR80/WuZozLvLirWwD4gyno8
CyjXgo1FVIMcKWZnXNxZ2NCHsSbu2REre7gY+LdWv24csWpS1siFhjxiZsYyZ6xAJunwNXaWquFq
Q8o2oEUkcRa0c559HLT1vpb+7i+cwoP44uiApF1YDAterMr8WRiW3le4i/vqz+MBXiuwtqRJkh5A
qqi6WOgvoJJ6U2h0zFYsfJcnIIgKLu8IckK/WVqKrcFkkq0ovd5TdfvC2YC9Iwuot6cX/6+2e3ep
HruuzwQSwYbr1uHflBnT3Fbme7Elz9qlqEnbzj92Cz+8fgpWhhSZYOcWLSPWzKfNP53/pNg0L7d8
gI+okJNR7FTIgUBfs+VTSzcyISA0NxLwqOXWjmcnshyVW5eMOeKqjnr9iME2bOdsmnNTsdSsqBs2
ThJnZeCC58VUS6cu/lWuJAQ5ykeW6OvWunbpAQBbTOlvLJXZEgT95sN0sKxURw7bh1037rIjwghy
sSUA45J8ytj9JuCW9HhFsAAYSIiARW5wA0YkWuQvF8z6xQnBFg4K69jky8iaFFRsOTNZtIsPunWR
HwmFmEbEo9SkAV4HTGT5WQ9nXlPhYwgSDFGfr85g9HVJ96q5a/4U6mBLn7yUE6YRZiYemk490OfU
3N6B4joTlFOKwKLeFdr9YxEf/ByAwA8gP73TKE5hJq4TEp4AlCwSWmgzmVwcdOv/l+HlXPgMfipa
4FNhOWevxLtsT/ZZ3yLC8T9K3yvZAb6f0h5N6Vx/lfoe5XeUB5R4uTQnm9vHolDSsk/r+4Cn06oa
e+pajB7MgbDtBdQanCwMzyi59MIZpxEd8RMDwJh39orslqlALFHtr996kreM5paQGOtrxlp2O1yG
K8mcfJOzbMNjHb/8spMaSdc5LxOIzkfAv9mNvwJgytEJLxz+V39ZySUWLv92/44W4dA0rq0LcgyM
U+zH/XaIdICp2UKkQIHo7iCBakuuqyHtkY9Xuh6LR8K4mZluHZi75drZEB9+7jm3gAKF0xnH8pRi
6gt33PGlO8u8UVg+0tD3sT16rHHlFVmBK5bBzkzR4PtUh6mOtOAj6qNfoQ8L88V8CaaSlIdXGddW
Owdf5RVm11HvHkzj//kaeQU9pUM0k6VoiUmn4h/blkiSvWXrBkPrgkyW/lwKze7wu8G08wrxF8t/
1cFXD91Xdw1595+T5qCwvR6pa9WaVQcSrxtD58F3YI++KFjh4n1xsdVqp1D2qXmtZ86cuXESp9jJ
8qUzE2BfQ52l0CekSz2jXDFB/1aDE1tj/IzEoSykEC56R+unClfu/+AZvUqre0pfPm4lKeH29uEw
wlkI2i3HVOwyBU3fHn0wXCeeJ69GYsKRkSOGdkEBBc2iAu3gShRP3Z8iBua72VxN69SZjpn5iNfV
ZP5KT0V22HnjTwVl+wnI8ZGwTyXfEDJGCMg1+7StNS0W9m4cubu5jISKjtSrmDu1POEEplA+cq7p
o6BPYf0Ts/w6RO3lgH0bHBJC3x7WLXQXs9ATtyug2HE7nYf/fNi2DHjdhFu3ykgDjby/3L1HyZx/
1znFbFFz4y0385eupnTuwYDRLkAz435C2cpNwbqa52rZZqVH+pY4r5MZKTqikt6ozywLKou3xBMx
uELX2WxXAr/VaRpqwf+HAFmL3hAhCHvcz2dqNeffPiTZZ5lijX0NWhFUK/uN6S+AX9kRsXS+asm/
dnEqhI6cHNXeQ7qeSnjsNDZXFLREFTSDhNCXLLiUJmg+TQ4XhSGadbtJlRjOngvo3IDWjLyddlt5
YH395xwPlYrHpUkZ0ZNwZw1IV+79esudjw2IudO2+1M5xeapeX7oLP9NfJgQuI2jZokWbbfn4vga
knRV50ecn10TJRd4UWLQJFdHvGSjagsAZZe46dkHZeZ5zWvTVAB8bQNN0eb96oaf4Uy7NxDEYc6b
VIfs8ssTu09MSMImapdGZD0XPWxJ3wNSivhS2LFIkX8fXjP0ElQaZuuLPbBKWF0PzN6SB/A2AQbE
svmM/CsoPGGQ2SGOhTZmN3pCrBAyoFl5yY9yLGF62Gq2KYih0oUb8dTzraKomdFIxvSgb85HhVOc
YoLNnEkvoEidgJkY8/DvCwIFI1if+iI+nITCS4nYwGFtef+K5YwEf65EDTeIY1jP30XidFbRsqPk
CPC1mfck/j3XCdUmGurhzAjdPfCrztXzCikrUH9UE1/W16vTKBSqgqy/hIga3ICVn1bpKbj2dVsX
ZC/J8q7wAeos/BJEzkKxbZ8bb3+mbDG67mStWRRC0wBlcZGCmYyeeDuekFHqzpB/bOSkP9A+sDvK
HmQs7Apuj2prhL3kSi4v9Y+iOPy+t42ogfcaMsIdC97r76/IXRVp5cNqr4ngGzOZAW0VoeENSfY2
qikHP36J2LjI40zW4Y1D99cGoFnWcZMo6c2mc87iwm8zzqBcTl82zV6+0+mm9KC19nsuXp5Nhw/v
cKpprQoX0LFHiN8CCrOLxc+XbQaFlp6Q84l65ublZmfHmKspzmGXMue5Gbn0PgH8fwbpdsWiBedX
xU/rRe2kUgMOTaAbaqaeEU5g92QjQBqSDjIvWugA/I9ng7AlYrY1UNJijL0rii7RtWKvaUZZCdFb
GK3wu5oCfkoWYG6ZnGhZClZrTE176AuhUcLlITTgACmCuNvPulii6Acn/VxqYvj+EXHeBzHsiser
BIrXyWMMAEwCRjm7K7u5Eraw/3m0wdPxnxTQZjbLay4fRnlURBVd9jGn9ptqDbFSPdb/C7HHACsO
vhBm2erPy8LPLKb5gi5PiznsrTzD1KBXy86AZ2XpZYdYySirkAlxPQjie1yhCpiDjfc+BjD2ozp4
ZbYMCF95Hi49qDIgHmB6MHp9ShnWlbThwe2d3FUZliufFfGfyzRiSLVCgS3dZdA9xqATNZYYFO7+
OCl2hJIBgZB5OVzpPw61h0u1csyLdtq+95XG3k89RG7MlAJptK3iRlgILsZ6VrQoOjUvCKULN/Pc
yGYd1DCXvEld17wBA4RTCySIlNzJlkoSYDKKxhzidVpCDQ/jwuq4Fq7ebwroX/E1MT8wiauAgp6c
nXvEns3b8lk0e/0+t3g0vvn14Q9Mc/rj9OzPYP3Y0+GDWcD82kLIvvMSYRRd+5W1kt2mdYsPHsKJ
HBMC0ceM083sCNBA/rdRi5wIvKTjhgU08U8wekNwuNZhJG0lIR83jpkvqAzjoJ7hzjvEzaRJRP9D
MUmQ4MObqL8DyyV2BciQOog/qWBAUOTmkTdeLTq3aHZAitg7lX6DJqUJahi0cbGPhByfd6HMdJp1
QNFNFWWIkjmL4MQRI+VCXfKixS6CMtaEFHbMnQGQhNnBanpqikmbGxpXMLwon9BOuT/OGE4ergrP
hmIAQnj9iUHqjqmo7gIPj2H3MWNbXhaDQR1z59HT7hmfc7yFClKFfl3Dt6R2a6QmF8mIaaceDatr
3WZQBH3vzqVsTTjNiLI7n7v0Y1QnOAcOddH0vui89XKaiVbU5hFBxYYR4De/5/CwyaZvDkqXXK+f
oZitzJKnoc6Iu4mKmWMJ1FHGI+3iZdQI637ks4ubeM8/MSFxp+m5oofkrHU34mxO3t85gBfXUzy4
w1e+uF936P+TUQoM5A4KJ5jroSKfTIVHwPgDcJbd2n+3uR+RjeM7y6Px+697FGI9dpyN76I8HpRk
QYZEWEEgsDKJrYExq9AZuMU76fQqtGnziYmhYuUG1Bsr7o/TYmoiOT4lOpTC98MyCRuYTRIKH3fS
clKnlW2QWpvOUbi/nQGMrJWaIoOBIeMySkDItXU6idViUZRiguHfzn8oNv1IwIBKkmJWGd5kD2zi
3LEmgzAQT/9ctvz9q+oBLf/0cT5rXSyaQUr6i99tmQkj+JIVC+dGtW9Ba+UPLEORcdJ+YdcIFH1z
8IhV+AysI6LmEmzhl2ekkjFlDIFRYs2da8L1wQ7Kb6JHuM9zjLyIxYFuHW30vy4Ggf4XH7KqOkBt
1x3l/fSPSinP1h0Uprdx1ucZCwn6uUJmlOply8yRNx0mTJYibvZDIhQFqgmXDSgq1YQ68RLXpbZd
q2FgYaPFwXRiqcpYUhisM7Wd9MCqnkx4dNuSpZau1TsQKRmtw3m6X0xRo95ebsg6gK0zCYfpNX5n
Zqs1f00aqKqfFteCsPv/4t2WsvS6BnV+ttXE+B6FU9zrM96v6oam+Gr/wNu28afUpO71rEGsS7ZB
w89xVyaODZ7GFpmmkVbC9JTfW55aBP7wP84KnkgXjvgeQoia80BmxUPOPtC/doLxDXo1sWccZPb0
HsNjXYBPQxfTAGNpF97V4IvGzKZKXYm7vzqGs4YF478FBChOSGj6y0rxUsdkUDy7egKa/ZN394Og
gqejhuCBEZldmb6wI8G3cjETXhaBILvvL4wXxxh175Hv/565j/WbvGP4d6FVXl3fHDdP+fQ07931
4aTI9QQDmykgoEgTvweaY/iPgwRL487UqsJqecIStcxm/r4sWze3Ctqb/N85jJd2WrvucFMefVEN
SaM++Fck+fyYjYH3wnCsfeUATqQgP83cPdH2zYDdqQ8/xo9qZLoBumdxQTCzYXQmZD756gG1LlDE
wZSTedAHagG2rqgs0in5TYgWRobfgzaEdGKHieQ4bdYlgyBKrrQDReMSE83sgWYhK7CzakvqURba
4mA8xPhUAmMDV4qs71KXlefZWSNavnU6gODkiWWMBOQqY65KQvVwBGa1AXwmUwCYHZI2o0ZC9daU
xZMngFL8K78FKBeIvFSFkyDQ6TK+BXrH/odWxNZIHHR2sBFKYY8XarT3HsGtrVFzAuL08L7G7nHJ
khpaCer+NgHKPWaiemIhkzkyRqLEyWgS70+0FvXzEkwy4Brtr1FfxkVUlAvAF+USZCwFulKV0jw9
/8NralsPrdUuqRdYGR/p2fH4tJcYgStG8ZvwN2wXVwjtLygqCqSNdNNhoAAhuRNA4fhEOcc28D8b
FiIKaDpC2lxInrXQ4+6pJNxdU0dAudJReG/PbSB1jewO2iSa2f8iW86lW1TfQ4DbcBaVZrwPF3mS
EUsfP2liqpMouu+rs2T+v5a2+hz2LakfcoKT6/c/71Y3QiMAMFzPmjZsmH7SuS8SEdD3wTWXW0bl
QFZLPpbbVW4Pzu5dgKZ+ox/A2uDeajGEd0emNGf0E/6pUXMVc4wFL91VW1no6MBZjTzxP9ejmdst
mAS5PbBZw2Oakc14mOIrJXb4chke7xXvV9lPzIC58LXKU8J7P+xGGWVbYdlwGXhRFR5UUXKt2ijf
GqhVFbm3wHA7JLMcLHsU3Jh4jEn7EDG9Cfxp14U7XmBZKkkjGjxvRHtJH0lHHDitA70U3lmpfhyd
Wo7KiXWtx15gU11Weo+cMXIbWmq5nbT0OOhIwtQTw+QrqxLGT4Xqoow1ViPLX8f5zloYeB78uk8Y
HIjh1HtenaEURWOlGd9eEzUIVrRShG5EZFJvjcKtGzWFgyBqSeZTn8X6XokWMkpqEH/nQj122FPH
O3UUzI9JXHA6ifiPeWM3/Xl1K/FnsMF9r5Jd5ntin7N7rl/vWhd6xZn1eRtVlNqFvwzEdnt7WJsw
hlradzPz++jyWz7AFBhStHo6cRxrLBVwC3qB0jkerD9DpzaZaTqRDVAOL3Gv+KKmGEF6H9dTNmi0
fV8/nij4CMB/HsAb8pyUpnFqU31uc90nlRtfJDpIqrNItSKeeZjZ1ip40K4S36/spQgzidkgPr7v
jcaNnly2lZVEDrLX+ce3bxCg3a36usUCZC+aY4X9IjXqNvboFsb4qczDAaL2+LxqnzaMuTPuBRib
AzCBeD8JKX7+Zkv6yvxIXfS/VZQu4PIXZJbIQ02gWIh59L9bWSxWKOz0gjVTjReIRTghjQMulZif
ZnuqXITjeCXCx1gtKLxuRILPal93NYKABdQbZv0eBuef6rdIxv4cvemjp3aGRuOqFnRo34ng3bTr
zQh0Jps1JcSmLtt/mEVFt4Q8yzaTzGPqA5AwHwuas7VVI+y8p/tuCy+QHQPDpIPElDvV4DOKBnK5
l7o9M323L3OPyswuMT+BLvsDlPpR0RuN3BmZ6BIuD7qxe/tNrEE39UytiZ8trfMtm4G6YAweNPPa
critqMR0ycRc/AsDdUk+leWjQMJZw8WJGC3WOauC3vIPJzn27rvH1MHI/3NOzO8FRssyW+x4PBbZ
jm2+///92yQyJo3vGW5jtY/NNevCsuUVZkG0HnPlYfuwNtZISGNkIWqpjvbhdFx3hNeGoPvh7E2o
JTwZ70/Mva4Qnd4APMdBBTY7hYFfzVokXRf4vvRMV2n87e4LlblHYWBRRHtIgQr87QAjbKNosQc9
rkQNBd9oWb7HEHXnNQSFLWFOySBJdE0hp+tj6Nzz96y1OvpxAtH08zXtP/WU77izIRmL6sVphiBF
HrejlfpQlLmZEoXC8e/LFy5BaEfD9IcOnHogvTnRgHZKE2NabVUY5XBObQHIvETVEDCaePpe7RER
OyhEgZfF0veR+9YYmAFrgGdEnvNZfo0ojvWhvYCYv3h9lpJIwf0gGIZmv5mDwuIzL2z/6d3l/lPc
KAK2tqu/1n9dyga/Avqj2i0WOiaUrN5/y+CwD9w26BW4O/b0q0zJCMS6iGFUnzbnLi5IB5ELQArg
lw+1Ep7yxHDHfFIF+3oOEZQicGi0y7aIXIlF7BE7lKlbgBdXFlt8z+5xkTLyP+fYe2p7zp/wTP//
ugrRDKoSldkKG/6ZsjFWHKeWh0rSUb2em7M8JBPVaNN82Au14sNWwVZ0Tvd0u9sDtu12FxcOTTY8
2P91bZLzX0+18eNswz3aGodiSHUHDHGXrRVj6DidfawG6sDd1ikB+1AynB6YJHlrJzeQdSkIf/d2
eBp1AIxxadHsTKOcebHevr9VNSBKfpXgHoenSkhvN6LKrOqLbxn34tI1XncnjhziSAWGT+2act4j
NJYf3KzRQEX06YxleLS9zYtTfhKEdR1CW802+IqxDwUVs2dUt6M8f6jHt6HHZd21eVtujp8T2FZ2
Aas+fn3ThoS2SlCxiqxNqiSDcCq1vQuCfPDwrdmWtMNAWeAyUcwB52U9sULuQ66YUkUAlyU+cpgf
zM618rki4Eo7AVIR1WadjJETa8Qudr7M5OxxllGZREscnMk6CsATveHiGK1iZmrpEUGagt6hi5nB
yAf9ohNgataD7Koz1VXgUdE9rzt1IcDhJfSU6vKfdAJCfjtffRk8npc+Ye7H/KDzktcQtj4MBgZ0
gQ1YWH2kncTRFdDfiUaY32pC4HqbuzhMh2diNpeSFlnZJ1HxZLgs+DVTtChSD9Td82AFwHccer2Y
7kItYGkek8Ymfz25/fqxhoGoe9dplurMcRi2Bk1v8PrgcblGghllNL437QAuWW5ItcbrNF9fWxNa
fGrNrxyrLEcsU1QTgE8CpL3cUFHpIqCC76zRl8TL4uCJtduNcOSdTApn5SVJuDibddx2CnvjcWsH
oSzNmDC2Hie6WkzNrSMuOkVsbte6dNa/Y2IJmvMh8/71cDUt/CyJPqyixvROSI1VrHOBfLgSZSao
tl/T5MaANFTm7K4urIyrt64Vkb1+NaBLer7ehCOydm7XTDSC+sJrVzQyVC+PE8dZdOAHLr1P7N5B
qSTeWfpufHEvJdtH3Uz1oASUIo9UEM0XQ9dW96jyf0DQ9O2TkeaTNU1oBgCdheaiOtkGfqCvPbLV
NYnomFJJAtQfqAQDRkOeILKxduQ4wQxBspCCbI8uohHwc3HSNrhfyp63lArOy+hGYDuYV4JtT7pv
+yPmMa8YH7iWdX5dyknKLPymjniPCMvb6Mbt6AbKX4KVNr1BaAAcbrQjGeHfim8UBaEz8N8SHeRG
hyIToCRpnsSePeZayJBPQwB8cgnsiK4Ps+4B7Gsdm7q3v/oYftG2/byWHAu4HMGNxx9dlRYIYHFD
Djn9HXOHXcbP1PAgeFYLY6Cs3jwJTBOB1i9lZP7MgcQEwORFWyofY4Gj4t90R0xjRz1ysurlttTG
zc76Oi5C3e76D6sdXSDtWMd13E6WLmTfmOZaT0mO9B9N4yBfqy18hEOULYval8GvzEmRoAS4rl0I
7fO5ni/WNB/UzGzTMsdA4BBuCe/tQHpQDXACA0GQwJD5fvXqjMSte1Ry5yvf1Dgo6kpChvARbuQA
9cNBGPnK0J+PefjcR7jA4h7CbJzbQ4q7N40vq+gVjPNVl+/WpAo6utMv0zwQQp5EDNmoQrxZtAqQ
pN2BtgHcbcZZCZ2wGwTvnYZtceqHa3XrLYWNSsL01ik7cXyvFJEYMF0n7qqvW/HkUeKC5jcyzg66
UPdeCSse+eL5H19pNMU8eWueMtpOsgiGwcbe0S68iWZ84G7q2Rr57B6eAMmDNbMrsdHXogC8J9j1
pQXIN0s4oAY5AQtuNRtrWSIBDGS/zot2mInBCFbX2A9K8bAlnadoLmCJYnJ8xR/fc+HG0ncJiUg1
CjsRx29FTP5V59NPvn3oJRp5wJv392fL6Vc24wlDFKHV3Y+2Os5KDwlfRjAW/o7G6YgJQdng/ox7
Go9C9H1i5i1OhPeI7hzDEs693QSWJHrbBnStd7T0OLCQLvs8KjfcpNjhPI6Z+QcQic1PIMEnOF9q
Wew4m54dq1H1rR7eh2NLgzsA0HOF50l3GBrFuSiegQWk47r8HZQNgqNoBteHSfGkngdfmAbxU1VG
5bKEZknYK5GrXgJKVqFn3FruTmR2mDcwiK7ibKVa78gFh18yLHVsosiqcq6DvyvdGe6we/obxusl
FKgrC34D7kMu/uD/YfafHhYLH6+S1UFiPFvFqnzuszUDlSBB2TbhKPtbFvNLXkndlpD7spcsg6Gm
K4hj9s+EiDQ8QHaUnz1vsigjg4y6jQAAOvY75gk3DvQTD4Ps5ESQ8blRRE0tLvOzLkChkSi7ttqI
+2Jq75XPlL9aXnyXk9eSNO/utsA5IJWn49j9VPpnS8I8tCz8UuHWCuTcC/k3ogWHlOiDqhJ1rcgP
TN+XrO8iJHZhfguem2SDuGwK3sG+oV4aCdaM5NWhS+p/z3Ci/smvRqr0wZqnZyHNP2fmvm2Kex+P
Z3pQj/vJtbZiiyJqZ14bgZE3BL9ogysMjPmqnaJLEUvmLoadDVx/pPtZlCW6wAG6STMduRNWR4Bp
F4hUP0cAq+C/+liWoeW7YWeH+r81eWpUumwJie6W2JiZWies5OFwV3sTgoYbzsj9lwIVXCVdt3I2
SLSq5DabhTFY6hAITTOv9lu0KVMq3S0d3P209u1AYjFo5YiDTYjxxvb05ZEEL0XGyKpkUR3oU7H+
aeeDM8XHdxroIQAgOM9fEI67aNq0MDp4KJmuCNFkGcOl4rNpvLOcFkj+ynKpxJns1mNd5zMk2LW5
txdT33JqW7+Hn5921dyLoLkAEYwa/EDqd3pzUWq6elvVpzivsi/dU2cmo5p7X0UuOGY2HSjESEyG
+gjQgN/uESgwBx2WSe5wpVFuNHda6z+PMl+PKGW7Dc0joZkn8FD9BgDG02KWjz2LeSH8K8JeHqWz
bhA0qf68MC2pqPzVBIHr4MBAh6iUo5DEhyoWrj7GYZ4wK1PAJRlll8g4V69uwmLZuBSdUv3ZDrDb
GcWAvOZj1wGvPMUUxrVScwhC/uOIjVVvwkb3KT7T+ki+TvdQIJHSIdABNE2qxnFH3vxJWnqx1eYX
n77+y3VzfMVwIt1Wtr3TLbvfz/t50p6JfvAGKX1LBwWRFkN2FfnH2N2HHTg/xIiDBIVlL0fgdyUd
ysLy2LuIdrJGPwy0kH8Tonm0f9EG01HYUX225pCrIGn9HFFyxjqkAmT8kgQhyOoDjhJDBFgfKFhy
heCSCu++iMedxhwfLT1qPviMNiKJaQATwjs+7uwUMWspOZT/FUPQ1jJxVMZq71PkyE5GVU0E/D12
vbmmG6gmybNoMZsiYYquqQLxxDda6KPPVBTRvhBoBebCOBuwolYiv2+sEjmGgB1nivBzWBvq87FP
C19ZjftVX4Tdzrnak6VdVTNAcLSFF4GLtcY2cfE7htDJsw947by1B6hq9FoQtlMmPHK0xV62zbqX
iPIRHdsrWV5xmJvt9neioMkycx0jyUL/JdkgdITfzb/WjpZ+O+15PUocPvfN9uWQlM1gXQcb1tcZ
/eG/QcBh7RRbQ/oFGAd3ntbmkIl6QTNbrE30fbYXO7urtygDfDFDOgf2WyI0ao3FOT/ICgkAq/9A
clS2W1mJKaLRRTnHR7CLlQwWpKTdks/aUZWVGUcUe201y31hMSEP+S3bgwWHuZIC+Kf07SZCisfR
qOSF4ev1/p4cvfE4B7VMZke6vQUz/9h9kVnZ1Lxy+EVgb3UBZz8w7QqMEuRTyP7LTs90JW/ETIF8
6Rio6u2fNz3ySL2zarznqoX4AHDX8Wk7XZatcm4ZmxOfvY+uDrFbylkBnBMa85z46C5DB7EBb1Aa
EcfALEusiDxXzRgU/TZfrPvaeLpV4RIQ4p8q1+cMRPicay4aC100crXuNN76u8edKK71npl9+zyy
5tJ8cKIlTAct3pQX8cLSaDJnscUFNqttEPO1s7EUvSft3LHxF5JHgZwkxXokymB6K3faGuFk3XHc
XY2bkAUBS3EgydW44Xp9k+ilgGbn09VFgfDTkDJDlkL1qfDEQRHmfm68mdBz8d038mGFUwDVu9Mp
nctfisrho2FeuRvU7UvAfBFF/1qUDkVHfOseAPO+C6Kv177Pp2siPIr3+He66TlDmKKXM8dj6K5t
d6DjujtM1yjMAdB0lbJOEWA/m9oQuCXJs+dR3oT0LQ+6BdwZTTaONw6YX4MXzB9ClonFpixtfLJr
DpyMrwLI1yBoORdhpM6MT1ZBffA9Awa6NPRAOub8NtS8d0ePDJwr863qThTzkXEgCyazBEUZk30Y
aiq+r3V4J9yxdcBUkvbrZCNXYd2JhyZJEG6c97is/YCsfpCMR7vUHU+UQWerL9VSbAE3Y2vhYda4
ujcuF1l/FThD1QlOku7mX9n+OqOBONmem48rygpgWOjbCD1vmgwdwD5AJysjf6H+0PqqvUTG5OeY
/lh3bgdsCz6Buu5B+lOA6+vVMI7x/oM2Pgeo6D0tDL47oLiwiCuPPM7SC2pSM11eSWr0+ODQ3ila
sK5TIpF/059fKcWSpORbTuiarCEeqbu1Y35OgRaINaexGJkp+2xDKgLCpZ0DySYwqsZMOP/qCpIQ
sKICVBz4JyPkT47Fu523IoehKwy3zgXj5uGgLi935sK4GSQtCHBSPXWnpUR0sA29/J938rYQMLQm
7BEFJcHfIcmskVc7Ao/CteSOZkFwIR7YkqPsP9qmibLmBipH3bHrRTBrzcbcLF+MROvRSWzW+oYb
tais7DTYt1lfxBKiFDpwVQwnCsA33jyvfjhJBNrn7mYF+fEAou3k5CzV1lsxAxF8R/SAc8okN4D+
m6fDfdJ48yKviKJibqM6kNoQd5S4aUcXM4zsxRblHU0/7pacOBxO/lQv30tJloGeXMre5/ByhOuk
LUlHdrE37PxRvw1fmZQ39WSHWYRqtCb6d3V8wk7dqouyF2wbmONHhgGeEtQjax+X6HuP5g1Iim/e
7oJ+nXTkzhB5VZ0h1Blib3Afz/tZeyA7xPsEaedNiCLcBowj2DfwrTlVxnPelU1H531I3iHVRkpg
Vj3WaQt/vclrVXK4T+Js6p+XXG1eS8CEnqqcO2q9sMpjeT8R0Bt11K6nlfffcWJ6vp08Uk9rEWKA
5y7ivfH4Qvq8F/DFMYsp9qu6mpRZos+yRymg9mPyPrkMx3/RArXN29ruJ/6kfBp1hg0etFGZyEB1
iuoIUiMqj9mNK9FrlJxMZBuDmcTKcdi9ZC3xkyz9uTP3NaVKDAJZgHYbIYszfaFY15jRVYRSdzuk
p5mr7CJ7FUDCjsoTdmhC7NkQFmzH+Pvk20931EtEW+1wA+fmbtlFjsiOUwXWKgziZEalO6PUgwUA
aTiXO+OY31/angSx1DeW3BGk2p9cmIf77Gmcf1ENl154Cr90fHeKxwqu8gGkbC/F3ZgudBW7Cqpe
GeNVWnpYbpUbjxIxMblbMjesLZHzERIVnqcW36jYEOT+71i4jL2KUsDZSRtBYddJtjRhXYo6Ig8s
jggTd+DFAP+Qcr2uwesQH3lSc0gcPrUEzU+2Wbr3hzGxROTv0hnYROrHUf4AtqGXoLk4ydYdbpUj
wPzCTwD0dvkXsswEksQLlBNOLSuhy81jZiQYqho9lwGJDNjdfTU7zTg5Hgq7VdnVP8w0L2e5hTZ3
TGm7mLpRJO0BjIiqVMAyF/RI1Lkdcb1yx83uvGpGDHeGfhc8sgDRMdXXQ72hXCpq6drYDd/iBaZz
YbFNfMwb/CB8K882Alu8IKJAAJxIluqWdWXr1/RQ8C74nIVFk+5wpL7SmNJi19MEwr4bgEVyu+kz
MjTJtWAJJqgp558izjNyN5aDMhnAYnUz8EdQeBveb+H4VUbtgF8Qqx/PF208eJrSX4yntpFNGr5S
xIEHCJDi/Din+ynfIVRItph7e2GaRTerd+qlURKBLhpD5tjcAQEyLvjbTTLF0Nsi7O24iDiVtNfc
N4V4Mi+dWPq/89rPyCibppTnt17oRZ/3AWxFDt3+K/NxODAy73yRzQqjpRGMmpniVElgbULfO3dB
PojKPOVokfyMaF1R+0K3ZZbdIdOAxKFMG7Dh/MvjJvQhw/+uHmYZlbrALpf0/8Prf9jbTgTu9kQ/
6G2j8bsr91vKAn6P62v8Uq7Li1M/h0Pyi7dtUlEs3YqaCLWHhcuPSicoA8zArhQK2RyJOle+zdTL
KrYCu8jIuQQKHFwP7YBl/5mngCUfdMOq4L+u1cTyFbJacEsEA1BjmrsPF2WMV5TNyImQ5Xutqn9R
ZvGsTyv+vSDIQ51BbE6DPG4tKCpxLDYvumgjiqQp9XuEVGEqTU+8Or2EULDDsv3laUXwYn8FiKUe
vHIkm/3CNCugOP9qHbvG1jTmeW+lBjMbgrjzO8qSF4THh9ICrCzaH+mjNopDs+dSREiG6uvYi9SF
R28BHO0DeNnvp9JQWiUXFl4Y3nZir5gjoRsw4IWNOXnp0kmBIdXuSFsWyN0jAf9sclLZWGjtWUzq
pjVWH+54hcbg8SJf26JERhTsk5ClF6t5LT9tTIMwR+yrQPYXn6c8TUWuguhUAdh/b2oZXdh9qHDN
Bcwcw4Fnl+uqpuD7KSrTTLlQZt7vQ7+Ex95cLD3dZ1gV/AFkIgB4JvUScNrH4lLoDIxXEOTQ+C+O
hvy7uyInH17dQXBCAXhWpBbW95YiMeWf1E8cCbfXL0A91GMzUvze2l2saOXqmKugqwVDwNOG1tTM
tTMp+hJLDRLSYTegbB8zGcv5CG/yfDi8+kpyCKncxR6SO0z38JvaxPzKdQDSWW2kDUauOlRVQz3R
0gh+aMN0Itzphes3JUy5Lm+Ca9vA9FIXTWQaSKqRClbN6+teg/MoZDnvvTNK3YFwkUoNggrSWrq+
WWF9CW7Xhny8Hbee5AaeHcaCEq7MBDL0wP5htLFCPPfq9oqZh0RuYiHEnI9Hr5dFzQd9U2WIkrsA
qvS1IQqkGVST9LJ5pwLaqYdZrU+RevN36nKOo7epGA9VYmn8KSd+DCqtum57fqCMZICNI+PgeeBI
aKGzCSXAiPceo7sVNlzgSRAxJfeXnbRCKlV+CElGfVX/hossZ8JYZs/qeAx2ZmzqZMR6pZ9j7HZH
QZ8PFLU0FPZnq2NyjDqcOpDWpwHpCZK5xma6cJjOygQPp9kH7cK3a2kr89lb46bhofmscbE85uAS
tzBQOUWAK7wCVq3RjvCKfFksIqeQ1AoPQeZulByOHFEZEaUSQjh1CAhCg1n/q0/Svrif/Gtwy1Eu
cYsy7T9FBYmH9WfLZg2wmdVge/ucZCd0Xpxm7bK5ZSE+mV+IrCYm90fLR/AHbKSquRjo7PlA5xcM
ANi/glmZfwrFid/juorTVuxQqG2sYqPdyIibPDOLZ9Ngz0IIPh0yxtLkUqg5clSS8F9sehoraJpw
ZfqkWg/nPbaRdEP60zAWIpX3bAnOsBAVbzyfDyhiZPVm8AeyFzvHhCZOQLjLR0TMi+j36O2sdExK
kgmHoNyMRaCApZGP+yWmm4q6ZekLe/AxugEz11RxrWKbOITL3cqEndnEcR2jH4c9NUHrKjdXDnGK
H0d3DIMwgZTfSqd/l0a3a0P5bYgPnwfAhhv1ZAwKDiJMuVAHZcbLfKc6HGjmB+G34v2X9y6ZSuAd
L0JG117deBOJNoVWh9SWC6VGo97x7UKuzWjDa9edt0DlCukIhzt7C2clKfAEhb98CEZVjHtVDkfz
4Og0/T5CD57Lrs772HivyA5UZkSygyvD0lBDz4gUAVSYoS3MvoIC0Hc1csMiooeJBA/4gqZkFkY2
yacAE8Rng/aI/uYONXe90byyGKRqOEATFvk6jyuzJvjz6wGkAhLVrV+iltgxSjhptp1rgBgE7V3u
kjfNnaRMl55WWLiOY0SkH1tsrj6zrMciX+vr5h9AAjlKTe3kLQ8u85v6L2r1DZvESKQUZCaDs/L7
rvOXEeQUzFQM9bGv2D0BPQTbsIh3jaK8RLdVDKwxrJl0YQUoQtbgD3L0/4OsSCA1e6I9C8gaUaLR
6Y+7tpGOMSelYJnFOCWr2yKS48O9jF2tb8TQJGfSs4MSaF4iU77I9JFeQNc035/Er6nLQdhM06jk
3Bxf89/ZvmfSafIO+drVidudu17t/wuF0gan1ELDX2Xb9y+5hTQld6b8S5lZqFnD5vZajBV0Hdms
/6+pRJKBjabcru1KGR9CvwjiJvj3JC1QJ1Z/YrGtJCo5Ge/VKnuf5KjLQZplpR6Uf4CcA/zSnuZi
hRuySSJFyIF2XTeayo+xC8jST/eoDfhofow06j9MeQyDMw2YWm9QWKjY6bg2sC3Enlt17r2jz9rq
gAkNdG+3nDGfuYWiMPTAuNX63Y+2JT0KGZkjq/m8kdVJyyKOZ1AGLkaVu2hwRRSfJDgn2bsK6AKT
N/Rl0CR/baUcex+ax2LqHa2IJWyUcM2jZD9qBuLQ5eA9TKHZHEsa+Z846VVuzctx23j8ozlrNbbu
Lc1/HJ9oJY9ZK/XrcXekDH97LLoaPmokTnTMWgAqSpmVxtkh6VW+LSYrlPai1cL7Kxxq0RffWiXV
ChpXANkQ1z50goJq0d0hyCzpJ8RM8k2wtHPMI9HlYxK5eLUrHHsBr8G4exf4cEJhOf+JKxCl3Ev9
DeDGxB9f/js9VVZp/saf72r8npJwoNLMoSI/L4u68L0YOBlRwivgFVeQEON1ebvHKsLzxmGmLZLC
sHtxfUnUjTwu/MXq1FiEQc6LY7VDJ2gnaEiM/jpdQGtqBmIGq1iwmLQhCBZYKH12FPfqUCWmGkTa
MIqSM46RQKw1gJbNvZdeCjPUK2sJJqAusPSFopn4wAvXLOCZ2D82hwB+tsg5Y9H5MfjZkBqhX3vE
H7kz7Hx0ANE5QiWnx0aRPbYIP/jYa79/94sHRhzRztJwLoCac66UZ3La0Bd3Sh9kwNRrJD9l00gN
79QFwUk/vQXw4PmKdbNKFy3gBYsI1iDJdimsGl34mjlYJWEJ+4QdwmsRus9fuIUwEwqxckUf4MMm
42dcTP6tCYzMxADMiAP41An1o19c30IAoH7O5FIUvqRbKvyAti4VNyJpcmMqHGs3CIIQdp2dX9E2
J0Jjz+ODY/AxxSunyqcKfV/H82X5KS3rt7HMUhOObeyisv2ebOmU3AyaMzSuUPb+SyXGtKe9blMG
Pd8EGjoZMFBQhPuFfGRwEJb3rIuroIK/bXqPkSxG7BpQNy8q7hKQtpEhTlYnK2ckW0uAdVMHKGdD
LaPS+plSI+Sm4kNOUgWW8C0Dp81U9N9g9nbiiChnsh8bauZrH/AL83b0frDgNJzvp5D+wrQRgL6s
bHwS3u2xJP/sWuxUcH/MkAVSloNRJWZUVyWb7FJY2ZCdEfZhLXvMOqbtjNIVFWQ7pSxeOZPvo33K
LCnlSG7nKxPMCP4ib7bKxzTnb2IVlxi5zBu/h6JDN7RiS1DOp34niH0rV72bQPw902kOI8GB2szT
eTn9NfJBS3j/ceK9uqa1wHrSh5AymZJzPKU9AGw5G6vM8b6f67eGWC1n+14EXQlB3xXHNWorJXjP
0PSVwYZzmQFNw8BYwz2tJEwx+dljA9zgst7LsX6vCzM7zcMjzS3iXK7MrDyS7V+ZLL3eQu6T5ak1
FMyxbs2AItqXHxUlBDcONd7EdDTDF8v5D6U56ygWSzdjyMktB3kt2RhVr1dJ9YhwBFMUseo7ObPM
D7AEVRLP7XKEHC4MtbUoGm3fZPOojhAITT6hQX/rsDGH0rIT1rXZw0DmdFRzidfkqplTq2WWF/M1
00s/jxstI0zt7P6hQz50y2oPn2Ke0Y6bUV8FI86WltaPiD/14AKBkwY6QqxDTJVmHF+rErYGDNGg
wO9/yN598zD0Qw/UL6kzlQ2+HW+eW8Ii1l1EY65CoXltlPZy0BZq3IOq0Hqq0xiZnfDDiXVAyWyA
x1OaSzeytOVOghsm6ur1+aykLqXYzyREDvYxYkrHViBneaX8BO5+pt29QRL8gdnw1SmNLGw980lH
ZPXat7NbPr52XeDXtB9s4pHLXOhdSdkSJCu5eVxQW20mt8Ioo8cAtRsxP7SgkLXVPwkHe0qmm42o
JR8jJaSoKt8Sy65byAIx8Z8oVJcjrmHoPwRS9gO3LNRnNTWaRBuPP+63hY1CSgYaXjH+NOIoVRqe
pLVz2yas4o2GD2w+4En4nTcdSSDdF+G5VEuahDIObQewGBjJzm5A0MjQJJfoSe3p6Cq1hrQU3Y5+
qkd8nqYJmnBLftoK2XYvsfX4Q2C516subAlHqRMMIyL+z/d12T3eQbdrRa+GAhJGYIeyD29yDPRI
8IdD50DURoZxw975k/wYL3n2l6LVwWmNESvpXW+7smNLS8+nijynYK/ABF9nfnVqEDvHjB89dg2F
KW3v/kIcwBKkuHyvO0SVM3/GZk0Hjw7eNxIxGye1sGGZQ1gT3X/WShB8xgzQyG3OhNWMRtnFNWtn
siUJaVw6kkMOUycXs4pBTMRwszUFfdMD/scQzI2/W7mjaVLLa5iAFrRArYDU4zQw6eYdSzkC1rIO
Wih88vnlBhPJt+sSWzG/iH5vbiULkhlf4CersTxHp33EjNLi7gapJP+yb6qUyUtcVtZwUOTLbxeZ
IKP2nqa39ThfzKqEkywCgrMg5XKWPhFrfcZv4qIfi44ZeThq8XFqIrKBkCKsbzrVUXdJ2pQjVFzt
mAtuMMR7HmXqzEkROmfXZysDmlmldbCyXiJuXD3x9fnmE/k8SG6x+n2SNlOHf4pcZJvJznE4oaWQ
lp0RQSsyV/AF6Gm7vpkif/42W0b+sfW0qAzaj+x9pNunckP4YEdIFAsXDiFErFiYIK6zVfaRdoAi
d7/GM8GOHlzDUHTQ+WZfQPeNJptNBndu2yW1yt3Aby9TOhPpHyuPe4yTdlH1vmx8ZpOchuSAurV6
ujXDgOw6xmsujUSnwZbmnlQalrK+bUyTCZLpO0FxNnidSPec7xVNYUdFxGmulx8gj23J1HAF5GE9
GFm7+5NmzvHAQK9vw3EVL8+NybGYfXTXFXV4FMCIw5CcpX7DD6vttxv6RnG6ap+tUd/Tp6IAIz7D
NmlePgTfwbPNGg6I/9fRWFviMYzIg6jD32WSwfinxWOCyJqQDb5bUEQvdST0y6NkM8FUZWrL1j3c
4pZZhMVHi9LKK3bfrrhsM8ApZSLf+I/3dmNJcO7IcnlNjMl5Ztjqy0kirZSobhOowpDIvt0sgUT+
GX+SR4Te1F944tBRpt1gy8NxItOZxCy1GuNmx9qhIQv8f+7X8DZgexCJ5GdjyRKUUOk3I4/lUogG
c1qBcqqICCYcikNx/mrDdj66g16daduE8hlit39DRcR1MiXiDoCRhzDtY74xBRN5llfwB8oWtkSC
YyfIHagVD38yRn2l/1rz1LMxtjadaqQlBifNDP6ppg10iDNkE2R6wS/+PaGiRjUStD+750xwIHTR
H+8g3IWdIKJFBjU0NMEpwsq9/H0P9AbxRglYNPLn0Rwgx3NDbVjtJpweGISReCa2G9mXw2mz7VPr
0rsQdwLpjoODxFp8PefHN3P2x1KfPLDtXhIcjX2z7aOl0Sr94nnEzldd0u7SkOc/FRAWQj6CaCvC
WbMJ0oggy94uyXoJvb0XTAR3lu/uqZxg+aKralhPW4HSOKNLy3Kk8854jwgs35eMKAhh2Vdq/OwR
ZPgg/mcM7SCvibPZyoQWXys49AQOSEcevMmiGyyKm5SztqZB3/eRrsDiDOO/CccUfEw5NFfSSJ83
g+zTXYkPAb+U7QfeHqS8AewxJAKopT1x5CXNhZ4+8enSezoJPdpy9i+t24Rz7z9vVBHDU7VbPCCq
GuoH26j/f5NDo4fvg9LNbFI3XkYfkg1hzEO69QLEOLAz6paNHGS/rpK3x4LnxChhuqPo0F0T4kHm
f/1X2k1BMbgtrCE/eTd9QhemRKm+B5zOMkapfYi3TXmWLHsRQtvFQQqQMSPkbCZUXAdiyvaHAtYa
ahDYsfZohlAQ/KLa42V6y46dZkZ/v1tNhqLXkd5LU+y2i/sdiq2F4eKu6aYV0hfc67buV3U+TrcR
rKwOlsSc2qoQsh0AVwD7MbHbQe7VfM+wEbNplXNkWGFwBtrnlfcVl8ip1AeMZ4FbJ5UUrPQFoTSR
UHkkUnCMLgViQ5I5SXCSf0+uvXSJUAi5E34btHtkzdp6uAtjbdpu4/IUsF8hkKLbhpMLQcdXGu1h
6bgcJI/tITRrJSB3A4P4R26KoHHfOKBLyWeRJH9+KDVh7vKNNiT28t86KBHlHXn9rJCx2EHaJ67X
vJOLBQbRtT3yqG3OEf7ecQACojFE3enCafjm8/IAXL0pG3FQcBFBZr9XFvrtpeyFI2nqRuqux5kN
BDIqPaJ+CJ+Mca3LHsBLgUalqRXQ9XZK9ilpcD6MelhbDCqgInNznuYUYAqdXGyy1So0EY8ywZ41
NNhbDajIFMIvyBOre7apD18Djx7Zzf47ibiBtN5T3l4mkk/HwQSWVPKfuDPCFgCZszPJhmEgozHt
8TSG9PuZb26JI3XTXjzTcV0bFitYvEmDuuE+JwldIMKkRTmeuqavwCNFTpvztnxW6arPtZI6+kS6
WTU9grkp5hA81HdYK7op8MDUalJh4sidOu3LSu67f6+HLBZPjNqazu9JCEMqow1ewuywB9z72AbH
MCGfAijVJgh3uhdF4W5N7uoda0NNS9UIdom2r7vbr2kF4bYhM2p+O47Y4yunBcQuqwmHWB4yvRD+
Wb/za1357InU8sNPmPCwdB8yEBG2wDZ5RV44DOSrQ6cnkkG/cMmouk2iXQeVOUDIKMZOBHd7/aX5
LMz6gni0YJdjLUFjbQqXOHaLGI+lRloNB6pRH1hdqNApZoLPtSPh6CCfks9bSK363vPT4tO/e2+h
r/K0VuwGn5GGX04fH4+8mKiTBF+uyGFEgvgrlKBU+OKWQ/MLB09/mRUS6hcYixI4z0WjrThjia9R
Oo942ZI/71vxDi3ZmZHrAPUN2PLOvxOR/ufeLtIby7rHdrFISpiehdkZ10XliGd4ulQ7inItTkAy
OO6PNODKLriVhyLBJm7HVM/JNQvBoJV4p6sBedJ4bWqgCnyI6GJP1k1A/Nj0sUkX5++bb5ndID0b
ZHfpos6e5ot7WGBxfeBYwUQ97TAxhtfVievVgr4XKNBu921lyrFt6XMptGZO44zSD8QqenBE0SFV
W5e2CF8RW3f0ZgtWsfeJMGLfYetWRyAPJNy11RHnX+rrsBrf7cPC4rKobuhWl+W5MDW4sjaoR6Ip
/C5Osad+cMRKiC24VtlVd7vCP2el8a1fZlOoqqntglfBfuUXM1GGTHYgK0QdNYcg428/Vzfa6Mq3
/UQiTUUuc4qo4IqK28QaFU22QwJq6Uft4iIidr2dJTHxDkzWhK2sI18Ee2RWvsqDf/AxRWPVSGJ5
I3i3DGmwLDJIlZU39XRuRMwiGyoAyG26gmWS3zdASJDK0MDKFsU+LR3yX4M4H3ixY60e7H9bhDaH
lDEwYfua9y2GFJwsYf3OarH4BbX2P1FOw27qoJChgZU8mjbW+CRvSbwsIgxNf3+0o6aYBp3pRu68
fCOsgmGi4D8tcaLcl8y/8I7skkKD2NtYcETd+EXSXKflbSIb2TB9+P891Frx+xySsX7UchLjrgOk
MAkRL4v04OYgL4Nrul3F+FBgrtomC1Wbpiwqt6lcyWZq4N7OVA60DCYKLmpc0dHTYSNkxDZFXluh
0FAG78qvLc5GuTBTpcbo1RAgI4dyDjQL1SWsHcfItxrEzwlm2dEgjzBiqWXUTCJKc0HwFLQXaNXY
9fqxEqszQYdp5cQiJEmxMgl/mDQVJVVYAE8UhVZNU3SzPccZX6QQqcww8a8b18Mo+ou5e5UsaDU1
MpLOCEtearGNxu5T3eHWMFq3o3ac8AbIozItw/VYai0WkcGjjfVpVYkY4EDw8TNCrT6rPR9/WJV+
j8t/rdRU8Iz6sbbum/MWZiTAuawLN5VNBQjJBcKnkE347OG3WVYYNJzYc+XrpnBCR6rhE4pob2qP
V3v8aI3IMUyKWN2nfGUXHTHNZKcZ5X9ztVspR3qxHIrFZJ4Mo8AfC6vqPfm4v44K0qH3Rwocbg67
NUso4f4eA60d+d1S6e9tBtiCcCManUAnbdX8BEqz0Fkz+eeCxV7No2XltkX04ASF+BpqpZcx8oFf
gRHLKQcURuipm5iy9LTxUh7tyn346v5W66hE8KWVrI2U2OPC3Q8KtZBz5+uY9ecKVHdvkeFWMoIs
0C54rc9wXn1d/wz1CUxoXOiGekM1nLZX9jTeOzMjueMwUSKonxaCogDPW8Yoyz8fn2TZkcoPgkLx
6vRZ4yq7v/5FQmGb4N3g201TBIv+mYEudxfSaz2f9jdlzcehCWs3ZAkqZZV34Jy4fCLKHyWyypj7
4jpXJ9tvRIQB3fmhtTRQQocNSEJPatxJ4Q45M8u1wSjMqcekxR+R1ewU0/Mv374U02+F2zL0obCW
9LLUdYTLO1MAVDaAGPp7SOxZ/XnufIlSHQHdlcOqd3TdVbhFh7bACyUhqo6+ghKD/7euRZp1wxla
iY6KQSOJlUMzfBCLkJJ9Mh9rUCuaqHnHMYIm7L/bJzxUKW6L0bNIV9H89RK6eEW4tFfAZLMCOQ8o
Se3rNei94vgk0KUl/9qziM6PEsWpNonDA/+vj4P/Q1EplkqHoEY/7KEUBa8JidE4PY1zrFWxjPCt
KAx2wUydnQ7Qe0nsB26Pj340sEoIGKSC4zdopsYMbUg4Ztc7U+DlCVACCAXQC7KCNLj0q5JeUtTp
c2hbFyAI+ZDcHpy6gpdQXsAjh8cJaUXTYaO/w/qopQ64iMtUuMfWwONHtMkfCTMrHXDq618p237U
vZMnAbthcf8Lj+yCU4IBRq+C8isa+5tP+cmlnFrj4cWZnoLiCdK/x3vRm2ldJT3gDelKXQ7fU+PQ
2t9wv+/4IYL96ZQgNjjtUz5VW+vJhxMsd3gsK1EE1YZBHHGm/gick47/SMapP5j9yzoAHqW83roJ
5x//L48WBMkf3lTsXDUDG2bsu70BroRmcwsK0PxyYUlpyEIoL2J/EKQjkhuHdhIrgBFUUwgjhnMK
watTdOe07Gpn1aktU+BvHpJdbgmLfqYyJPpSaKNvDSCm+9OmdWTR5sVHaal4Q8FWAiIvfgG56fKK
cGhiEYWa9DHVuyTln8+0O2dJSXGhMbeH3Ubri19272gsrNl9w8oKoeVGDkWGdmDDw6LWtvtGeWVE
tDZRt+nJRfl4rQaisVjyr1B3VmCkMORssKrl4OU2Qx8JbrLxHXPumsSuSTRSsadIjVwQGqoBsjQu
kNdruFRfnwenAZ4QZOXxPK3W266kKXYnQHXB+gqcNHO/hHc1iJmt4Tu1775Eiwfxsf7ld9EetQFx
o3OgvU0UzMbnsY4qzxKwlE9svEI5sBcTawNd/xb4CBpwODfAfYMe9JT5GR296Cmrds5bxUEr0SLb
51m7Erv21jJ9HzK3Ui1F2YCuSNbpD2KsHLDhCsRvnYxsJ5aGwuF+Bskkf4mphEzbxqcboCoeQJBS
TSzGWYkpVRAkDJi/orG5xeS6Q9ZJuKM/HHncVVbGVxSth1q/tgMWAJaXv8HqML3SoH8zxutwUJaG
zewIEm5vXSMsgxbx6quGz4jLS83MgzjiSbiZCKceLZ5RniRsqKfESAz19sDvpQE+MLcRG091PP2U
bOJTBLuXcqcji/Rqgs3bDtGbucT89j3HCf8TVCFoXBxw90T9H0VsXSQy499QaYFVdpBI4cHUhH6K
zLoKXx2fbtJj7z0QyB0H+33tXzXHOe3drA+WGAqaHtyhRX92JW2R0BKqJL5yqXsC3D0oFksGcmP9
CTyIFov9G5kiNgpiItAkdFh9Pq+TESJiYPGHR+YDR5zhFAItB1/72HW8aVgyWWfxuF6bR+JL8LXH
afxHoCGQv0VJ2yNbX65L9Dxx4X/cWMKNvqHOy5xRFTEj/GjgBHiyxpZdlWXQuFnk0rdpGszGOYE8
wRJRUXu7l8CQtNfLRBMZyzAiVi8Rm7hH8z4VsOYVMK55mxMUA+Da2CgIVHk/zjQ109Ev6TLpuIdF
lwf7HuIOVb5lJB3iV3AqqRKpb0vNrDNA/2LwPuRzssZwlcrKXGm59MDUEDV2ui8zRAOAV85imunE
mB4FXpbM5GBGqVP7hsS786dMtJmIXlceOvR1bNJCH5uayJJCUYeFl2K7q6WY91NlYSdNV0KcQlxL
IwzZorxC5334V0irUJKtECTNQHhGCeuDv0Ib/+C3z0FZFIJ8Wgx5tjH/tXrAB4s85Xocl6WiZ5Nt
CzO0rNLh47csKl/ZlX064m3wbLWqunrGOHK5TH4ZbludTd0vITxR8rV2Fby0fLmqCPAHV0HMkiHz
W61UDr0lN3xwlk8ltnaWu0z0vEH9y/+QJhSt5x5xexrLnf/4cJlDCBZ2HNlXSjB6rSuhJ3H+aTcn
GUKmrh3Pw/dK7LP7mnDztcDmQZPVARXLxJuJXSHNVozo1GpkM45NZEX1+6doWeDHSNgUoP3LMmnk
u1Amp38lRtPFJ2EEsz1MjWH8iz0Xo+KAv/CobcFMIuJUizO4yk1+W51hF9RDzVvzAOysneKDnye1
6IwgsHH80zNevI5h2L2Pwlf6+Qx0DNfDDLESEJhT6p3zHPfJoY3wU0I7T+BxFKI3opBcLLcqWtuu
Q79uqVds7Cz9KobcSf9h8YaSXVghjv/SoCRgDsmUD304Adw4cfM5UcoOIdDT/wFsv/9XhumbsUIB
HfNT/ydeBiigeFJIgk99HCaWai6eVacqj6L4mBuklHwKFhuMNWkts3/O7ENYptpgADod51ENammj
6cEn5WSvOv3CqFYl0g/C3xB9QtxVnOXMCbyUdrGuWv6C1wAaVMZX7tt71XqVBfwf/CimyxShR3g0
TZHqcw5qos8AtK1D6EZ8bsCpzt8OXwO2r1aEKTHbQTaiKWhQBAc9E+lUi5NGrvSsvjBgenE27HfG
WlMxMPV/LgPONbJhZSovJD5A3j1VKdMTpNZdp1wt7GpTcBxzV+KRORBOtvMxfox1HiZpm4KndTwf
RkNCyaBMSOMhvsAY5XaybgHbyfpODBpxRADQZCjkvV4zQekHHk/ldkIRJSL6WdPU1E+WStEAlUov
XGE+OxrN8FkBgsvRHe+g95rXm03BFKvExVsDQmTFlzTY1uE+14QN6ArC/teyX3fDYG0R9WWOwIwN
PUfvaSYgtLMqf9DVoJfggeN2ppmWfGf30qaSo0jyO0v/zNFBw7p5LBdVj7RYQtiztGwZPPswW89v
vPbLYNayv8Ai7hrPyiI2a74OAU8rt0hutDbpxalMrTvVHxaEr423yBXjhSSKcnidW4LRc0BAh7dt
v2tOPTI2uAkeiEX0/fPg/bHUhOtlS7YUu6MN+WiqWkMluszFCIvWt98nH25/YxFmHac/gdi2WfFv
SbWlATIGNgkT9xShF/0zluAv2UoYEAAG9qcDGea0dF7mKH3QviwzXsoMXlQxUDWtKtzHlKUrzf+6
bStpIwJm8fpqdjeKLkJWE3jYtylksa5OkkJSvoQZ7kFe6d0AFDvD6972exhlgFOiKCjHWPuOUaQu
KTK5l/ydv2EFvKjPcVapBUTQoNk+gMMpIeKk+9TkZDCdCycnAZTgXQ+dS1QfVELDHErlmk2WKUph
5LI7LNuu1dXLF48PhYpaEAj2k6VIpm7IH2lXeaLEMEICpOGiPSgu9ZLWa0wdbrmhK3q+hQXqwbJg
S+ADjmT36ZqAtuVYdvykJS20AshfOZD93WsZtFAygPi8lJmczoWFZkWRWsVheEypi045GXgoDCYU
oUgUipcp6XWMtCULZguX7QYOme9z8ahkc8dPh5pJYUapdWlF5ZqY07jKAoj5qWJV8c+w0Iu5Fqpc
Y0u7hCXNH5Lmb9bv5hFAD5JRWCKdbUjLrnRvKn7z/BpHvitUwSwQt3QImAyzHV9Xi5sGznHT03gw
53+HaH44kSLlndXp+vu+gNeHUjeY78NyX0uInnot748wmrtb6cdjaVNUmKFT0TuoflQko2HTMx98
8Xq9+Fx22/5n/jvM+piMCD9Dv3spx/F33LiWlY2EjW2NcJkiIlLaevGGRWl9HQfjdvvsQZG3FZ7n
JxAHn4ZwIn321Vr6cpJV1UBTbf7GfNee7fpkqr22VDQVEqVjnaEKdNWTG1KvhZsuYJ1Dgi3oITT7
cXwjKp5Ygbs8NB34kB/DNN4j8LJn8JFEMgI5XXX8wOOO8YEPszXcS9yqofoxZgoR/78HjQpUKwkE
jm0Xy/TvC/KEOeOsmYIpKhjRzOEmUo8No+qDweOWkQNieOa8NLlm3SfHiiW3ViYak5Ba5s/Njy+U
PvAAmDIoZJhokYCi3pk4KgoXSzRddLWSEH+PBIE0T6tTbas/zU2AZyTI6XmUZQyZxcCV0bW4u6s0
eqHjvtYhZ4lFAKKosmZsHh2DnUsfaNVeBAIPBZDwRmF0PjYOitJm3Lff1sPRPSlzuGKK6VfWN4WA
Iev6JT4KEfTlcpbsLxrc0kZHw6IDRl9WCBEz2mBoJ0N80VqJ9QfYe1y6ljaQKsGyQg6JiTjGGrBV
eOeWmoM2mg69Xh9333hLYDsceHejeii7XPI5PkvldOE4c4ro8BS89SJ3gvwFv3spngrNZMnPo3O4
k157HqMjGYdOAt38zQ7EKCn/Y9E9Mjxo5SigkbQ1vQVcuHW+EtGbN3moUuzryBX6FDOk5vGNRpRv
72Xf1QSS6191J5G5NruJYGRAgb59v39LxFI+8iW8mg6MP4T8fcfCVTCFiAo7yD2FSn4W+xUmWz/W
f28YB5Si8BgL/NcVyswPaC7E0Y6aUQS+FRyfHnY2BIuYJQoV0C1V0Y2OOhzH+F46GOLVkFms4/X7
T7LcnxALqJiL9HCbmolRsfY7TSgklc1dES4rUh2VRwMAjDv9WScAqsZ1OUCMh3lDMrZehjwhwM1t
jufrwWqywcARWpNyVXK2qU5L8CVmHKCpLGVit7QgS/qhpyvUPxY4OgIDyW1nbTj52AkQje2GZTxj
gTO8ABd96f8v1vloiK8dVTUZPd9CnkqiLILux9OcD5PU5073Nx2ZVyFSHAP7VNjLm/pd4DVl2dvS
o704tvjKaOc+x2ZlylgTBSnMvDerwhc5g4AXZy19Fh2BIb5w5aALalp5HW8oDf77TU3ufu0Mv1cb
H3+MtYoht5HWpZyPYaPWfF9wZvqCQVstrTUKHiU3U3fifN8S1ZWm1TlLspHrFbHX33SH3HuA3OqW
fiugKwfyQoIo8BI9p/WFfKytkwVYB4MKE5HFt+y7l5Yfg4Cwa+dkiCM5gsjaVHeUwh7sPjsIDZ0f
m/HHKfeg6rRqL6D/NbmNJJJdv0i3XYY3xUWQixcagJIKvHm7LgK+y8PwATQO+7eyaYSBtqje4hVK
3hlJvxGLsf397xWL4O/CKqy+bQ3EJ2EqmEYzcyEegQRSe/GpWZQ+7Cja3xX2fjp6CjdK1kROFaad
vrWvtpGSjkO8XtzxJUufNyhxgKcCyypZbCXEBSfhxsDKceIZuKWkbDVtUBide3CaJCjR9ZteVGcD
BUvVKVvgm1OA/4PY4DGG6rf/Fsj6tnBx1EtLr8U4x5exLeGrDqohkBVZrk+tjlvpEx8l3RPtUNGB
G1KMFrAvwcYcPsaGuvexOu4TzVaajUGNZAPf5kYU7vQjssDaazJ8bTQ3EKDxnb2mYrAN8EDOtZLy
TeQgESdzo8V4Ttnu2UeBh1ZZRSrcep0+w2LkTt210D6SPHguofCXg1G4xmw4wmMk50zuNORB25EQ
IQEBzoa47ZYAlELl4XLQ9z7BZnxxMsPiAbNbXrL7W14TFzZhXSc6GdPzGSzccX3BAWcOFZLW0XHV
xFa4Dv1yxXgxf9skpkmB/Gcrb8sBEcEWwlOcgp1lQY04qnI8fihKW89cae2TlFSOZV/7Avn04Z26
kNT+NdU/zU0QmAsKxcJo//0AsrsVpdPEGSZZ5oNKkxW2jDSAugDcWvRbct+gxmXGVd68DMFrJgKt
y185TQJXCFeQX52lmWT7WTgvLy25LoXzMybEsCBcSliqpU65ExKkm2dl1AKbZh14LWGESPBK0gea
x/hy62IEeMakjkin8KA0//URqcNBe4ViK/jul9Gsv2Zhn/3V7BX8EuiIdAVSUTXDKePzaonaFLOr
RRMOL3txqFtWo3QwhPQh2qb3Z40rTFG/f1K4Y6+JODIXmZfl26/U1tUuSGgDOz9r2eAInUjoTk3p
7cKR+z15b7wzVx331Jc+mccRzlt6hszNwOc7HcQn7u5OKLQ/rkrC9zKesVy0C1Cc6BI94qZ4dnSE
ZDLFqo5fjsHjraUeAadtdFn9PvtjfWU4kecKliKjwmMz7M4rXvrpgNZxs2Vye3EeNh2tGapyN4vJ
Skc86bBxJUDG+POxlU/ioftzuCDdy65lHPP/jv3Wqt3ipSU5vXhzdjLk4JjRpsUIWXpGG6qWPTiY
G8/Ea4yrqCIkvbuJgeP5gb+Xus0K8pN82xAg2XIDI2IppBvDE4zRf0UGrNz+6BCpMAjSh44R0fIE
pp586r9/cWgwm7LtDRqUv+w/mP9ktDdiJBd5vM6QyPAJ9o/QOXA+X8xX/ihaM0/8+mL9gwUS+B9y
aJaFyRI9EBNYMHgaCSefS/ptRq5Iln4yQ2bAq8mZbl91DyoAD87NhIqBX9uuFiRzUDy7R76wxbfW
o2+LcCyTO2T2CWU+ib0Btxz7w1XgcCED5ViMYlpH298FwHa9+LJEajbqiC44w4SauJDyr/zY+QY+
vcLyEJ+08h7KFHzpnG54m2GQ1R+94aH+1p3YZeFUKlZMBkw8FBPY2l0ucqacuvFCkCmiG3ljt4t/
rVwiuwNxvnzWQJyyaF3ORCUm9rfU6d8eli7Dl+Ri6zJoDQ5rIIoA2dmcBnmhW+wz+sCu27u6R7nv
4ryZIKWlsN36g0turyRu38f1XrLFCbjLG+n8ajZ9S+Otio6Ax3rxEBBzXQG0X2Np7m9g6cGMXnir
pbBFT6IgyRyqvd5+hu+e5+kBqezVx4O5rrVqVAoDvln0mOiIbwumLVCbEAloKuD/nQi3OlRS3p9Q
0QNyWFlm8VTdkPYEOycCWp39DRq3Mn8WaWZuIXETvdtrvIQ6cAZjv/A9qIDo1RGaoz11xw0wxtRQ
Ip9TalrBv17CgkOTpVb2xZVn3QZhEsomgxJr0XTacErGDzbCiHe+rAcF8bX0/dhRK0GZr2Zv3AoV
OWJfhIGRYovTgG66wrZohO51M+54R3jysc51qFmWxuvJvJ94UiSKombgzVbFNmtET/g6T/3GgG9H
95Hozc2cFoGgFI6J/3fPfqW/iyT3ibsxIFP1n87Ec4HFuly2QbNT2XsNTRNAF8B4mUc1KQs9qF+y
Z1mWj/yv8gEzuCI0E1AjO4LfY0xvMUsRPj1wBIzYRaKNqQ7mhlGWD2ca8DqvgrcxKZaDngGvFw93
dPy+q/vrxafp2WugcSFpGNR2jiQEyN6Vig+M9LnAvcq+Di4LkS5NO3pDrARY8pdjW8Q6QLx5em7H
oaFL9XHOwPIxl4Lei5kIr8HQPGkOECFwcUJ1O254/pBn9HFcMmMKwbNiHQppyP9RuIVni7e60GCW
zpopFEMUMTG5GXdRax6UYIKXKo/YYnmPmK0YwNW6FiLWSN2wQ/UF2YlNxgNV0mnMcdElanrqOL2W
LPjy37/qvsCvwDvSC6JCAauUAwAWMRpN3nrsH6xQl7eHudOKp8cTCoh5YtB++LsFgwa26EPwt21O
IwRo/en191Jam7yM8FOxy7VDTWSxO7yDSSoXRF3fIa/ifl6I+ak6y0t2jB6YrSLOUJ0OO4DNmng3
gZxT1HM/pcTtqRRxqZ6tng/s/4ce/yqAdnCB6JPGoOyx2Gukwg0gtEne9G9v2sDjDhVIGiUd5jDM
72Ztq+ChyM0+JzeoabAlYA83ZoJwV2dXGBC2soCnZ8g7eu9MdAhUNsF552udUV8AyJkP98LwJRqp
UqBjILAPKeErfxPIEOeZTfXVfoi86hZVhopqBffQh1Lx+d5N0rN2F3vbe8/8wW7YAiDk/3CEzhYt
iKdkcHDVDbRb7SxBN1PbOYCuC5/v5ZIVlQZMirk9qvSnw3BUsD0x+rLonfNBsH2XSEKRRn22pjm4
1xQ7hdwNBZjHS0SYVgmeQxEiX80PYkxGsczBsXVH8/uhON03gKXLjEya2JKcWoqxLiBAqfOmeww4
JBuMmIF6ZNAteJlqQnWsqnksLlVx5Q4UhX896tBRAmpuSUr6NZKie/GjXMkwzMEGnRVypdNKZ4yp
VBcJ4mcIDV4R3w1rrEt49J1Ubn1Lw9nXSVch8lUrgT4VX2UKPgtMZdlPOs1icgvxNepKOxNwbFvt
Go01GT1J32d3RztkDI7bboDFqFiu57uPBGgIwAwJ1NV9v1QU0gyI4me2QrFQNw4hIK4dC81eKtKu
rKYGc3nCEIWlDlu5ofpFa9LutOvcimkQwiHz1KaCvoHCGRPi9a4lwGvZsKXiV4tyBpu2CgUMw1R1
wuKTWLaCZ/xyZeVphbp/7PL8jgUvWLbErcyv0iiAwCbZseE2e9YuXHpfnZeug+AEDVa6Ps7wndfE
94B5MJjIgitaPfD090dSw5YbK7bt8pR9ScXCJLK7ZLfE1RZjIymK/a0MzXxKKVteyZI/mMvHfTUD
S9oTh6Iv5TjvKfS1HOwNzXy6BLwx74AAyMzcZ0Y6LGE/Wveav4SUQaGbTGnGMwmHuFtvdxpUU2nQ
mzgp2XSt8Vvyv65j20T3pUKpxg7LOilJzrRuJOPMawWEwpN165KuCnXB/1RPbuUApE/K6N1JGcJm
Cflmw0A7/+xi2aNp7UAQg22W/rA1QDm3T/jjbiCZHfAr9jKkwSSOOPBPbEWnMbVrZhwHmtblWBxp
yxabs+EaQVYLe+vl7JPXlUqutoDOZCIS1sY/SiixfvF/EAbyWABPJBM0cINFP+dUqNJsdJv/1Xss
DA9bCUJXjRPgFuqr6z76jyrq45OQ9FZIAlv2+Ljzi2IYine7kkRed9c+VARPVJJoeC+XlIOjSXm5
w8OunDZObv3XcQ2NWInBZSOX1KmUoxMw5CeMo2LnLEWr8jevrHu6YARkPVTDnwGyrT9G8zZwEYm3
E8yPL6ygEV9N16qi0pfjSa03GViSKk3MRe3DD6KlzLSHPkJaKs4oAGztZuiqyppoGOBQR0qAPFLX
NdRK8fBqm/xuS6YTV1aR2qiCQENLbVS+/jemThqa5wT4vWbUB85lWasAJuJnGuHFVuuiBHKtBDSl
JSK5bDX8HIk4brQ9wURAD37XMnSrcoFxQGVbaIGU9OHNBHioyIhBVH48K8HcHbrafBvigaDTwrkQ
uOMtamkoj+6w6hXa5+WGfZoMnfggvyO846Gc50/51V26+xbr8fWgh8IWDwLSLmrBhIeZ2ncsG/Wd
V5ZeZWJD6Pjcdz8o9xij90B7yLk9gOGRqaG7NQh+1ptsxRqOFiRJFg4EN4JJF4/W+fJJEQsRMr6X
CWQHQfnJhDc0kjX6qcGkGxg+ub/q5J5aUqq7IDxEeNGDMqM17Xa+DfmNi0672AyVPBysFlJgAPCs
LeudysbqLXNgmhsZs/Tvb5LIVNtU857E7ew4CMd1McCQm0a8e87IpMz5o4SzvFNDfm3efGqrZ/Su
1PALS7i1aXgv3nrBU14uomEKvYmoP9CaHKWel1pPKYWSm0Bi5By0etjg0Zw5fkeICYkz88Dloioi
kqUILE1O6IjIcRweOtSc3uWOJmDHs6WNKCLUg2RWjDs57HEjDTy8gMBQyHrFJYS5JzNB1qIpEeID
OS6TsAsYiqr5jlHjFSp2r/6qWRJ4++d4sbW2iYfTKqHnAwS5XgHaKaHJOQyBeVF+ssZEkzxhoBEc
qBUJg4cj6hOHj3RJaPNjbBqc7zqEx6iZ3yT+QDZKj4WXqbB8TonUAd3iksZ4GI+Ns0pLZAbV3FOI
SwA06a0FJnTKqyTtif0tDz8dGdDJa/O8NZDyZr3vu7aBTR/MfNfHnIGQU/GkItVLfJFjdsmlNa7H
dZSDRrZEdy2Ib9k/QSBB0Yzaf9N8hzuU7IDQS5P3oj2aU9kqCTmepgZOg7x68Lvvb2hteV3LBr7X
bIiNlHxuD3REa4U8/6W6t6dOVdfrBHao0y428enX1Ij5ksFYumzemZbvhQcj34cImaeifXkoPOIb
GiZawqEm5usPWDB8Ml7/qMgHAwU/fb0FJTjQPdGCAee/ZlEmIq8BxMjn6arJPUeeZ0Fg9mZwjGr7
mbHz2sRUvX+fA60RQJKXSucIvzIn4I6MLoE+/Zq1LoRaUd05xP31yWlyBhIxQxngzDmJAO72nbHy
bEiJ4KEXyniXIMN7gajukYefxRSFeV2OzY4rxSr2AhBDrwwiUKdpG8+ZTYbdDLOnonxv+ab6Htq/
qK8WhauLcwOCBGBaORF01erdGfA5xeFLBSxoY8G1cOGR+fh4A2jVSg4yKyeKmenwUXVgHP9Qh3id
aelxCQuFZsyVtfeyDtq+bGN77gM6CX6CVbevv43ZQ9ka6XMTEqrE2q3ma7HHry3wVcMqY8WRqSn7
ctxLQH8wl+HXzys3vWsMA/NrUxaES1VoO/T1Km42zLO9qkOU+IYk9ajNGrp+FRaEfiebp+CwSOzB
14u+OsG328VwkJMbsZp8yeyEyJ/lQYcYgZNP4dQ9EuNCS9YxVaMLf+YXYvSPo0ZVojIfBlV+XeaG
68OqrGKTnjf/j5b+sF1Yj8lRXcgdSRJXJzby83YJzNdFouTNgXjoM8tpSFkJ6v18QtKcZcdmW/SB
5uFa3qbpEirsA6t1rzQUNBV4H0wsTl7KzFuLoARX+m1p97Dr7H2YD2Y8FuzgdF62Tj401T+NkB5f
8zdfCHMjedHHLi0ll7bKPaeRqTzj6n3SfYzbiuxTyF1rraCprdyQ7I/BZTT4iGf5FRS80JEuxBfx
m7rlKLuoT2LtryElLssYbcwfScIZOPzU0seF0E0ggAKru3FJmoeDNouwSx6Z2bCqbRKNSuMtHYDF
kUPRVkI/jSNy5UjsmCG0Svv3UXeq4AoGcDezKSAzeHVuBtwXCLhdqqv2NesbwjVQp0ujOjDnlZ7O
EeEw0lMxID9gMVgODxc+QEvRXJnryxmArIbNL2z0RvYpfbsV+ZZeJ/sj47au6OxpIOJChzYZNdGq
4v5Rd6TAMvGTZ34ZTEpztnUza2xaObldngHFElTGDINr4uJtFs2iqKoGF7mns0Y2PNniChiyhxqJ
meJ5Vi2lFXmOJpRGpXalP73A4OVBpbWsLNsw8mL6Yt0HLg7oGaH7uYdFvtz+YLs+WRaG6bNPMXFN
y9QNSqUDBWtg+irAeVYHrAhSjkaEHGmrZEkgpmcliKaXJ6CK1aRT76K+g/QQOS9041zBNO1CDocN
cGYIx8bAG97WdFTwdo6BEbHu/8vHDZvqsu6YDqOwZqcMTOwmChYRIU05TsrMxJZ02ORY1os4mJQ2
O23JBkkfvtAt9PgflweO24KSFbVA+FGiKIRXPX+yPlMEw15FZe3iKdwgLGs5vlC7T0QVxXfutgDU
OWvaBK4T31hS3NfhyG8D2fH6j2NGqOa9oxPrKFej/wVfH5WJkYKNCoM4y32X4V35Ys4N2PoMMKSn
j1oBw9L0eltTiVmlHwWRHoHhoyAJS4qbwzHM1F0XXNvxNn04R05jpgAzOgXwJ3pmacPfRaIVUNse
0Zmjm9R94oR/IjFs4pkzTFdouglHugYrKQT1EZkVDsCZAY7k6QS2POi5gjaTlHzZk1VYpGldLeZv
Rt7y5S+ylONtYk+FNkVO14+fWMxVu1Qdj7tlMVIj0xMqHXpEA3dUWhBdRcGvFDxwGqsdI/8AES0y
RlHlI6MBWmTBurdi8opMjzJwJbL0mxB6iwv1xtuh1L0aWYak6GvJGY0jR8PakC0nMXacYH2eeOvE
KfahZpp+/oe+lAq3i04csyNRnLP5gZa0QqCTuREvueM1kDVNRl2fsSpJP1vCzVg4FSjCe8hjtgtE
dFNd+B+hoHtaPqF3B4ppLbrf433QyStWcirPKNeV+SWZ7cZBrp5N2iIgdBpWdVhXuXkCLx6GpsMQ
6j/9fHz73tTolHJj+CDOKKfZRVUHqKdidwfepX/+2jDXOrPwL48+Eu7jSIgbO2ujRwi11lqR/E2l
8TDi+mZhcPdRMt9n17Pn3AgMRTjPEMl6RvcRfLL5fTOITnDJkXnu1ysTVCJEw+M2O2MXcZfQkn5+
47EyTiaoUjZC1ldiwTu3d2bpQBpan1Ro5PP6wVAN4oEQRfuRkrAk6jdAbiibK6GhiYioMNqgkkij
f31cgl6MiMewyma3daUU3oRXE8AlaeBPxSWoyvEY99JLGgHiFfxQhiMVgm4dRIChbpnlLrTxad65
cjtAK2XYJaZ/ATVR825QUr034PDvJTJgaT36LXPZs3dfYuiDJxlTdHt10X17T+XRZ1v6xLVCC2Kb
GZ3LaTGM+ChIV8peBBtrv7zvOJgi/2gCmKHXV4x1AOnHaBjpO28od6LAuSx3NOrdX2PF5+5tNTBB
qXNrgqB22jbET5X8BpX65RtjFOvWcoNWLbLM7eVenCV14EJNPVhG9daUf6HVW1/xhsMU+8hzKx2h
+z397vRB7NFVP4xIZ8IdyFL12o79TRQLY+bRI3eTLRYLyOxvlR1oYzuzzl20pqQQx0ayccqs1nOf
Fne5WjDg/PKSXMWLexmoFD9brN3dCAm9oaK1+XJ5WxRTc7zmXtzXtvOdGayC1ioZ+Qmgb0CKSU2I
GWPhsYB9HIyekgjgRUz/lVRa5iA4voNwdQgaUGrE7F30vrmqI0xd9XAcqAG1DOt3qJ3ySQNU5ojf
FZuGmZjQbGqmnfJx2yE/+vMlzrvwK1CD6ubSun6Ahv4o6Q6b4a2kzU0e+lzESNTuj27rLBiBQceP
x1AIyVH2zAylRRMi9Kcq+wX7Gc4XhuMz1WbOVhpmOadRCWXpjccQcfmtcZlmt3QgpUlvSvMfex26
EAVI4DOvDsqkJJJAykEJGnuXRO3nCLOnuuc0tIxj0sEflhS61Uvhc6K3zZyPPQQJQba0zl7KMIID
yDY9dcqPrvR6TUAaZDagXsukTqB6IFwrByoAYHjD8A8va8/RnSuLtLKsddO3qISjFRfmzW8jkA8C
UA1ImCxmL+xRAtoPgmikf/rk6zZoG0J+iyYdsDYA5lQbbzRAoK+qcACoFEoqu4g/+la3KlmBfGDd
glJw49zRvZ/ZPYYpyzhN/ogBy2DpIXblDw+jWUaqVi7ppINGsOYO6STAG693V8b1bD6FIbLTQO0Y
yr1BUKH1RsqusLXaHtQXWSPUDcnb4QtCMp6rAePzLeo/T05x5Php5zJEsxETi0Twh9Kfh9OTaOL0
vkt0O84DvWQQbc4YD1Sy+QfTJL/iYYLg9z7Fdy98KtRagIdkctncAxa7tRvZ3TuFd919eJQXkh6l
PEZ8VQ/8xHhuZNevEBW1ZHAbdHlFauEREC0RRo/LkBu2w7/8KccesrgVYSB4kk4oYOT8lAM0zMYu
POAibgPvmfFx0jQOaqybQkNdrQj+/zmzjvuGSni9qCZuHlspmpV3ozBoffgfy3Lx01dJHBn6z5v5
l+gADoobBcjnAj9de4Nvd0Y2S2xUmc1BBeCEoLOYD/tcfM9q8u1cTxo/dWVS/CXy42xRJF7tT7Wt
RX2Ul89QoHhYfvo7mmP0D+g8WBeFmTly9CrEfvyrMYgEaGvxF2GRLKBzLAosAkY1Vw4a+5ELm9il
j1OUhb+ErTSvRC0ijYtBYT7osKLwGZPvd68sUTHUW0UvmLO65QrOJtwHEFZSCA3M+sK7iSh79Fy/
bHeP+NQaD1uv6enXEcHC1jmJmqqlSaQ0tGRLQOYlGydBb96PS14Sr9MHIhcS9+rz6PRjljaPlBaO
nsPhUTcEiURbhROwWJKCw1BWJm6hTVEDnLuoCoyKxhKIQ1aQ8rS5SW3vr5uOlHarsjHWVxs8tuGB
oVXtUegppKgKOC5vzYGg6Ir0wcOlUt0lkmtxGbGsPjzGnaQs+Aq9GDcTwBP8H6A+aERzTnBgUKtr
hpjJb6ugw9fk1Qjh9DeUeUvzqZo7u6f5pat+3AxAPjV+IrXI4fdjavblYyGo/ha9kOF/igXzx4iv
JBXrvKJhPBP+jmONFUhMZDQY8IVtCSm9U678VyaTkNyisWJBhl8jSlmH0vq0AHbtSB7BxaDZ5p7H
KAK9JLuUoGKPbTcU2zQtZtic+kPb8UAs/8kUFWLMqzdSsBEiB3pdP+FmQMUQXNlav/estW7n1B4W
mtkpZCJFaP2ZWtLdFaetgEmtM76BceJla2fuw4Rg1siDE6GsAZWYEXsYnpuoPSzzH36+shd6I+X7
ENh1kio6MUrg/+7PAYgenfwnSg4dOV5oTQFLZ2YBaoh1SGro1f0xLjWwdqjU0CkT/kMiaoaqS9BS
smmO8QP53hYEL9S5v7pl0wl3T4CwXPp/v118Gjk+LWYlOS1CwjKLjAb1WDlDkkxDRSm77bGrGzsI
8MFVwYbBB4nwarfQGHUpwbUSdNToHHL0l7a2/SRwGi4m07S12hT3QJtNPu9rPGSYxEdq4mwoWegJ
cAN+QP3khyjo8NVG3aFEX+YoDBugQrNLrFKOtImG+ZnWnHALE4mL5yEXLE7waso310ze3yxF64gV
kQfLhB6AZedXQkkR9nOJYgil3Jf7yasXCRV7+ddidu3GM/iCrlLp+zPBKulUEvZxpl8VSqw62itO
8j3Z2EAmtrQzcVBMMJsgRcgtu0FfiPClsnEP4tsDnfSQsA61G3FhMgWfxxLCsJR10XBV6gidGQ33
87Y0s4VEsvgpEljUYGfsZQb3mhc5yvcdIxafneMB1TA3P4WnFdgDIJWh4qhKJNmfaPwkcLSZ/nJN
Xzf+c7bwOiiwlcVUjg3/IApzGFmgEl3G43DH3LiqeScG/A+OLJ2Pidm4uDy4Xj06Zklaqaoe/UuG
qwvq15oqrbspVBwx56pGx6Gbz+OvMDIM0FYlCTFi9C1kVEQI3L5HBLeQcqL1h3Wl23/MRVpLH6Td
292y3xnWKyjiDGN+X2EUBZtrDB79GvL7MIe7QQIFTtJ+g8k02Vy+a/6LxMQ//3kW6ADaqXtmnyOC
pcNS4wwENlb0lDyDHMT+E5Q+wImc18nwWhHjHp87ytJ+RR+1DmimFHAbonQqxRulBFgbPOEshAUr
zF+f/M1BBf92JRJtTK2feMjzF5VZ2m8KziU9GdPX+p+Q+RieVNt4gg233Gl8Q7B2ksmg7LEHZjQZ
ZOLDgX5r+R5tITYzFuqJjYVKBVRWjVaSErnV+chlIv0xDsi7vr7KfSnox6tD/NtMPFIcX8JetNnB
e/0c1JgZDUVxk+rUZ9b8pe8wOYzRlyrUo8HbmM7eLlXUUVGK3wnxcnMzXQk63qfPpkTDIl+T8ZV8
kb7k6hLvQNcs4cNNNCnClZ67JU8AQyQ9yvdjbf53zrflRxvSNIHunA3ScTtw7s9TutXYnf4Rov31
HOPcVOO6islemDEib5x0lciOzUBLQlXWWPL6hn5fjQ0BkpP/VgPkQ8oyQi+OqXbHQH2TVSznmADW
XmEqTD+n1jCPlc5XMq+ZzLwdbVWMnhGUsGDVVcQnuss9vG/26fTl12Lc59YC2ljeRYfTdHzPGFDW
3Naw9jpt2NfVxzMmoudkhrfJxL6LUqi6t5Ms2PQrJIT6IM/bHZlCdcFSJpFvc/70JbU6WWTR4bM3
c4P90B7DGiwkHoQQPoEu4Pk7jf7syIf7uC5QxlpHvU0ngQSU3kITJEP9u1NldbDkTVYUXOHDyRnS
Zab03qwjZ0uHgw4OG9DgefE6v2dEAv3WcOTseTrKKt5Hg3yw3aVklmQ839sWPtwijTTTq0L+mWaZ
XAtqW5cVIkV4ru7i8PxQkLdTIfLgTVk9gdvcW/7QtIVbS9nijc3w50XZHnjldNxCUgLTKOgewLtb
8Poxi18IuHYguVczuKzaNoOXHSe8Vw5pCFXNlwi9NvAmVv3Pq1VWNiLcGyp1eWNybiTOAmyaXncF
DMUTtGXmaK9kMcWUJF5SzpuyJL6OhJpys8tyX5TA3msolDwBf314SCtd5eE4vF40cPPSedGLPh4N
7XwHUBHNqxXVj+lzJj0ViRZInw5bfvSXkgZmfdW/yQw5IQd4xjctuPp8glNsXjqEOOVP15iBIRWu
8w2z2S59MkIcZFR/I3AwF96Ou8zd/NeYCK3RBeZQgWG7Fv2JPXTxq1hQyId8Yixteso0qaM8PJsC
c538j7vLOZnO+aXIeCB18tIFjyql7B1siw25F96ru4yg9SjsCCtjIfWfZRqxifE16hJeKUMYUp60
Ve7rgoyhIVztwRB4qYZu7GnAHMRIT+zn1H7QZP6fAr0LRIzVGkeBE5yGalplVBm7TVqPaCUyIYq/
FNog2bZEkGWT5LqKg2U4/NhPwtlRD7Urzc/j+0UXaqSJhnFMpFekdLWDHGOdvSN44kxZRSigURoj
3okR+a8FttHR6NpiyfipHRHozpxKoXoYs1RJQRGpWTPi0SjipT9X0T+WTAwm3dNZ33htQ+8w7aEh
NL1LcBhpHf48HdOOUG7CR0Pmk8CPxkqHBdwWYNkqwgm8aEh41zpZ+dA32uQ581tmNr6Uh6GFoAym
SDaTHUUpm+1M7hhZOFC+RoyF04KnHev046QKfnRwylNzwhpj2bP6oIlCPLiqiMyAAL4dmwEUfOWZ
Fq0CcbgkPHbO30k/RQMDt4Q/TET899JMhRofSDokRdABoZR+shetwmNIrx8Ga0vEg7sv9iFLLbuq
sxzOHTP0DvOhnCV7H7L8Gx5rAbiAHDdGrDjpYTILuhhIfJhNzV3wzGqhpp99VGQM8AOQahU6G7n8
1sVRhdC1WLamYx76WmckxPmsod1voqRiCGpxqoOkjibRd4CbilWikita52qfRBc0dh66M7R+Cplk
iFHcmoFUoiLAByJL1jb6kbVO+ILpW/7NXt+YfH+GjJ4EZR6TKvFZgE2/MkxWD7C7s+zRvHnOxu8X
FLR7weASzHQo+Fb863AkJ+5AUChmjOIcbppKA0H23kXYeXJHF8uPC+txYsbPrFOqP6bMnrqluFTz
U15KbnJWx1Rs+AXSjA73l5ffaRxm4eoiXMte6o2/k3Dldd2Q/05Ws9zqtkWxk+nDEdpW05ObUhBI
+JDKdeLXC9egdQOfvIERQ2hlk5E7N3WIZgeDC1tdHgJ7p9GRpcZYaFytpPeZ4m5CyXnyUaz26wtW
A8yCWGVDx9iVuG5BWdhW8H5048QwiIvxE8uLxhGzaN52B+X9zVuWXexwpwGLmRwmkLbrPpmxb826
N0skAOaEljsA2pCce+n96FA3nF2vxhk/3ka3nCVCyP1CdoQzMgj42dTguZhnhP35rK3dle3eHPdE
DaQt969uEv3qQclIHkIDfyhiRnp9SUhPabwBmP9u+or/tBu91ZMSi6eIZ6wUDFkd26E3bk00f9WY
x49YtxyeKJTg38d2rfQ+yOx+4u1BMPqPAQCpLVICp8EXrZUnqEpcq6ufAFehNFnASC5u3eR5Eo7E
JGACVSoaHQ0knewn5Lraxg27E6s6+F9PBtwXeWI14L6tbwRKVTXeU2GBLIUaLug+D3eQZ893e250
CIIMpuF3Lm4ACILMFmw3XdXSfDH0GhTjtTT7e+KQRF2ZyK/B4pUx+LnSRJ0YYBWgBXo+2iI4iJCn
z0POc/BJ8GsHX3/V6n65/X2zypwufssOqhXWLLODeWtRmlc3/PDVC1EOISeg2JkKfzJMsPXnTVfH
RIdQaZnSv+H5DC1j0fZPa13MXxLwRGlsU5bkBlcvdgBVuvhG8dGIcaEZVvuY63JuW99GzdlwO9ml
hOffP5L52LPrjPicIrgbN/EY1KV5Kbz9PrdOcsDNd9NNYj2U/73yLRefooq3RnMkKUH8A61DF97k
Ya9f7BtZg+2bxEb/cgh6T5VoEsfMFoSFQmFqaYOBwYMy/SqrRekIb001W2k2AMnzFnT8/kvnx0+D
qZBVNCInu5hwokvjcuTYc4a2gMZtLZ1tY/UIXQi3X1uc6VxKzbFUz5RV5MOkOc35kdVTn7k9Y4Oo
u9HCwjitknq0ECNYhksmCej+yevKUbx+DQIHNHC4ZDWbvNsT+cdpsYCtPZoq4+CUOakIiAkVAzCn
XZMWzZp3luYgNwJX38ZAgUg0ApJEAsnUkEsge6I5eAFclmn8113mbDA2e1ClAd0ZBUL8XHlVbNJN
l2lMVTBD3G8Y9RH8qS5TJvf9mVnzYKo2Ox0Zbd/I+BNE9ZX+Vgdjo7VJNkNPDR7Rtao7BO9htLS9
r+021MdbHWQ7GSykfplXxwKOEYHVw6nwe+R8hv280JTZD/+h8jEmDfgMegnaJp4ybi3cI3cVhUCZ
OVMEu/9LHe6dXF+8DdeGEyzrbHhqzrUO3Xh1+kpRH2lkxdG6Z/jfzKlJH5zeWOzRKJHbcYt1q3bI
fj1s/8AZIbJ7Jx2dd8l0IHHZsDJx78qVm0yhd7TJaDWZN9q7SFnNrBb9iYDDUb9CnARpGY9Suky+
jEufj1o67KZr0ZjFamk2iVUgj1IgJcQ3cgsqKDDDyF/KjqT2h4ZGYQ+GGRtmIgywheatCvmUlN6m
Jahlvm1mOa2Ok/c5g1QxEmajZUI/q6jmd2oRNrjITp9Mjg2xeQuLDlmadCefMjT2lElhOQKH8Rs4
rAMGOLl7ckjHvZ4WZYgL/YijKEa5hhlxbeolYCGrs5kKf/dP7Vo2AnCO6vXlg3zKkp0L30+c29WX
aGTkWEFtLwZUd0px7XvcCiDDZrsLbR7K+v5XGyFHQb5sY2lrburQjSBQDlo5eHrY8OiNNVnmBtH2
wC/VLSxG+cLrfa6oz4+RpkKLkJH386GLAzvsUVJklhTPGkHT/G2YbxjxLgJRnIff1FldZQmWhIr1
eCKm71Urxp3yb5Gd0T3xplL2ceHGrB7UYn2Ln0ikh27Mof0x4MHQgSVBp0uAa3fKkPh1eBEeKQzy
ap0YYg1dJazQz6ianyXLkUrK5hjyekFLBeTZ0yzvEDDDAzRAqzt/dIesvNBZkoIE2ZEjpQdJFxnI
HtC+DkbTzAW1XHuR0fUSJETbbmJ2b9rLJZs1a3fMJJJX8XIwozVmcS2gFOE4Ml1JZXOSuIuTS2nZ
HLjC4B42UpmRSwjPfL4rAB0uZCiV1JyjMHzt6OUeofkvNFzyXZnjj++XTiXc/CVV0cTVnTuLT9jj
AgBkep6FYDBQZIYISD6rYiiDrcp9AQ0n8JqmXVXyayI80OqVSUvF/jt4hU9Qhx1s2hZd1vutiyu8
Mc0WgtyZ3g2UAQxR4v4y/g02zwUdbf/AFx+1ZsD0+eJ+BSoZJy94ZeU9CMmeyCHNoZMVa4BgcXC4
bFVhUTCr3tTS0HOO+bDZdEGO1aBTqaOU9vBTq9STGm6K9DQRg5R2WHCg8QgF6IXjcUEQkkHR3YtX
4GclJjP+T/E5k61cxUaYwyxPnTXDiJj5p+/RYW0gbdY9KEjuIThq/D+/KdL2tQ1WoJzUOGNS4gxF
8K380ky7qo9zhQoNoykXfcOXRUEn4l1ly65zF9J6fDgYyfbV8tRGnmEm4FlQpRavehYy5+/b3T/r
mZFDU9JlIZlH/y8ohVLq0n2SyUZkKP8gVV7eU/72rpFvesk6tGGS+j6Zbm0q2gOqvRMTS0Kche/x
iuK98AvCShWTTm+bSUo6XXhH3vxw6MIFgbgjQH4lSIZEpmNpBxXE1GGh31MnhRi4Vs+tD2r8yDS5
4wyq4IN0C+IHV0k9iU0mMfy3mkDVg77K6Lug2PNOO+AJhkQBuB799pEoJ8MCNmFtEK34yDmAVgkt
T9gTW6EC5GjxcA60wP946G1uHqyjZuUZ4uviSYpqxU/+bNwVSFHCUQe/UmhKvVwQh2A/umlegWEp
Nn3AhyU90Pbj4AwtZvrEOZLTA1kL6rxThZptotusod13hhqVmjb/NGcE6A/5s66aSd2cTCVMJ83i
b5oCIt8Nq7pmlWz+JeiryY6ZV7V63TvkiWv86zMhLh05lwmic5UEA9y8WIHP+4J0dTIFQdplxY6k
Sn2WvuCC8VbQPno/tqMkC+cF/+vBicefnhOYh8WsrCBim2XlVA/qas01u5hIlUT2rIhnTWmBCQQS
UBXl4IWYtLPRi3ov6Qlp4WjjasDCdExEjMWDk6cBgB+FHdxPBxdp8ZlgxpecmqCPKyCJb8awJq8/
cnh2yXhll4zBJ0q7JgvXOzchAKJW10noaRPx/B7pZHzhH0cUQ5pYNh+ja40q0q7Zb6trM0SV68QB
hHsHQGMJAQISyMrjyW5qGKB61O0PQ3/VwA7gxV0l/8pb8H2Uv/j90iGGXT93LhduEeZR2/3tsp4X
sN/JBN7ZWbWxXNeQJTtekV7J3Xh2vgD+PLEnSoKintFR1nHXlCSVXoZagxuCxFELyPq0n0oAeqXi
5+4juy6G1mgdqjXoKdi5FmyoE91XTK91YVuGfosF2SY+1XAhHumvgSOFX1Vl91iMHWATjalyVVRw
zVuN64XSbQmhLE6eSd7up9d1d+v1RXeGevkGbGd9+qPq2HlbCviJfD+L+PwJ8Bt7dibLPSTjIVH6
vZ08Qg/VIP6KSN5KPVY/IKdT5Jj0FFvInfr9HB403ZhZEjzavnJooYGfz76TsuEOlsUuzXN1pggg
DGmC7p7ipIAg4UYhB/sItUGQE8oK/ThCoXY1vYg+cppAEwGNZDRC75t9vqJ/PNVL+5ueSTvkJODg
CxnD1nB0iitMJMfo20ArJNLG0449avKaMi9FyvdGEkWexlIKOYSY+k+nmcOM82WP3CYiM25dS8y7
A1bBtYYdWgiO4MEpTW+O/AZpK4rILihg2cu664AqAg5SwWZ/j2d1kOulQo6FbmV2w6Wt4vNGCWzJ
5KTaram5sUmuBW1lw4RbGFq3kbXPr2+4O5kLec3erUGuOy4Wln2XicjZQXl8KCoUj5t2ZcRAMrcD
3r5GoDhwrSoVxuuzL31kgkuyZaOcXSOi6EBl8AFxO6EJsoxYpLLuPU+Dl+YF9yucSyJYHPfeoVKp
qGvY3QB4+4wWdORlCjs4EYvEc/lE5vSJQR6faochZP1jUI8k989AkX1qwJMQLA/KiQlN/NQY8ljW
RscHBD+LdNaEQU8auaCINW6tv3sBsU/6wtAWXpiMtThhPwLDg+Ej2ddlBsEisfWdGWEpq4QdW798
hsAYqAHBkhL5YJTIkpfLwGgfdlxzIdRDuRQM3OS22+FlouIOj2NekjYdC4oEZsrlxQm1QoS25liX
2aO2sPCAOa+vQXJLOBMdCJ5E+F2T5brINdkzJhYvf8eNorUCjudsIOmZPZzoPLfchJWA9hhTetxs
IsShYrB/YDlKzWSEPWYTmZO3R3uA+hUCzqSfQRu6W65HHrMMDuV9vGMibDwVF0AphH9Vb80lDWd8
HZ06UeFP5AxJUs1KKUn0PxlmZYZ5pLCrX6jQW71IhXDZQvp79XrPiNHwH17v/QGUVzxoz8BJ+cip
CD0+tJqenQ8VIkivhKY5U3VPO1O/tn3tFveoI4Nrwaw5D8gT2/344fZiMmTQGP2ElELbR1Jw9sh8
4MNn20jrDGp4ifi0TL9SDqrRytoqGDN14f+QyFHeNdMW18dnKGncjwUTybdh8R4mx+fzEOV0UtgK
/lWq1o/YXTW7ECmaHazt23lDcH8vyrfUts5stRS8HSzbKhlwkg09D1qEZ4l42M0XnSodZO1P9ZDs
VNdA+/WRRLRfmvkZV1KCggb784McgxDE/3czZ7j2pYHcyMugdLVr+DigYgGqEUj/3xAmJa7lz2nG
JKotrsSiz9/ArH2eLUcrWqrUPHbYyFgxP8zuA3EMSiWQ+9ZTrqY74oneKLo2VN8mI6P3nCC7bqQx
wPFO8epLXHIF14xAGkmwYyZxo58zHD5xJnYzsXLkF+1GfRgw/CbtXGK45MrggEM1+m4lrjB+zJIP
1FbZDXQ5KbudLWIFL70R4I3b9IcLtSw60xFF9eoreHA73prmzUCNiLMn0Gii7D8Yafdm3sDfvMyI
/ynvZZIjA5/mHYy0FF+rcn3q90bQ3KDWs/vYoRjDdqCngsrTNhdV035sDd40/KwnW43FLd0sQ2kR
te6TdT08OeO9Hp6g/PWk2/GBUBdQZ+MedMLDpz9XUtFrfk1bV++uz5ziCQ4j4y2oymMBKpsqdSaa
YVzPgLYGoXogeFU86nUr1fKR9NG3VvzHQH2FRdSAs9xZ+g76GgPXzFFpMx9xlu+ApNDdC97b06c1
/hD1mdNINBdSHIGm7kysC9rUKtH0LDkUloDxMajiTw5YJKKesHoow32QrkPaSP/W08+BmvMvx9A6
btfXiwhmgbJOsxQAhpM/tD3k+oBjsAIzilhkuYK9eJq5Y72lWSlUqOMutzJmlfbMLsOo+cbkBdxV
NP3NlESnReBHG9M780MEzQNqjqHLsRErka82VSF6eSo4NANDyq439tkiKV0zkhwOE6XsrfnBjxaC
geIcts0wAQh8Vu3nUrdk4Ek8Hm5UmORZpCLNF5CKPE0uLiHuP1GywekP1zsDOxiRCDMYkWhmPgzY
/e0eJGNul7Fhmfs/n9YENWoM+Ulr9s11uL7/rOL8naDtiHFb9+StLu7f3D0srR1XHb3Is8//NDAN
V4XxjmAfWyCxNETi/Tx8CVPxk8/gu+rasc85V7hV9xxAd5JvxbUxzW7qfFZUgXvAVZjwHZMph1dN
BPBFjCBNFpCEvvaCrXuf8Wl+T6ezD9p3BmcIBmLX2i3WWDyhRBm+gMHqaYOPAqP+5O1+Tj/ede4K
F519SPjdaiDNH9ofcv08/zOeuUBJjw+sdoOZQoXrqu5n8QswjLeSFEn1NVWYNiUsuRsXHPvvcM/y
hWS4u/1/fg09ByA+/C4a6m1ghewb3G2tCcBVc95uWVKG2cCDMtsikT29gq9Ha9siYT2DWMbbyWTd
wlyD3mj7yK/iL8MSdDcdUFSEST6xLhnvWT4+N1rhdHmw8ukfJbVLTvOiw1Qu5bQHvycsKPnSZa6i
4K4Avq4GD6dIrYcrcUcpMcuUwr7ib5sOKLHaZqq7lT2gk2bYX/1rgw3V0/wAazaAKeAzrubJE+YR
aNV2/Wvmd45Zn951h455v5DCLpQ55akz9/6M5mGmC3vGWnh2DoglEAtqjQtJJ/m/sEIEcoxnuLEF
nUscUBLHYFEBkMWe/M6mp5dKYQCQRXY5R2L7UqGDwrMyyy3g+3Qp3U3MTwyzuXGMUFXjDY4uiOV5
XdD/pXhODoO2Um9v6NA4ILvCGWdL0Ce308/lSVUX5qkFNJaifZwiubBd2GQP4XWVJHieEMEMs2Gs
N4p5CgMLjl9vELa6BmPSlNTaRGcGCLJoFEBeSaHqu1N4YPzrf+APlSSOF+za4D+l2yKUcQFNLIuQ
Rx/vM0lkM5m0m6xjsDl1qD8Q4BGfdQc82NcgkP4S3g1MgL23+0szY1mCizRXwXE0uPjHmPaio89n
zHx1jSddOopSEK2QNvQ+vDIL+CYmY7kWK9ME6bo+jSTAFZB/IPX3NsyBSfsRDS08CbC+ZWVTo0Cl
buxbbil+AN65H1aFg0iXW5g3N27JRVSd5WTPtjrpMABPpDBO9r6Qi/Ypp0/LImVIrhqlDIBcIK1X
X8IYG90JB4TeuchzM+2rsWZqxtcXLw37TLf3Uv11uuhLzZSRdK1PVYcevQ6k9BhQdiNGz9V3nP2M
aRSeo71jI1DL1wuFTwxSQ6sgPFxjeAeu9svj6x1NtcsQIZExJ8YHRsyB9hDaOBco8xzZCWqr2Wv5
h/jLJODAsjSqzTzQxbkPDPYf6Ij1uVmM7z6JVVeRSJhNkuU05IvkqFlVsZRF1bS15K8MUYT3h57w
RGg/A3CuX3fKNiYWR4TuAYoqSKkTQ51qcBMmcn/5gg2GjCos+VvvYer0JbNmPwm22pZewiAHq+i6
lys5tGdCL5nicVKNCDol6sARX70GBoZKnXRDLll5ghpbJgmA/vinE5xTRDRqfkFr3GXhVDWLXqp0
KujZ5FjrOH2BiwAsMDVSDxIycm0OPXcFeNmclIb4q+jDVHWQ8iKPy1VsYu0kqqSOfMYBplBfPDyQ
6tUe9PcTNzUIhRov0AGfxySZjUuHrCehQpYOwIpLRp4qf/gwyr6EHYFEkoG28+O2IhPojMO5ArYy
XFDXqlUR6MntO2jf4rcksECdVk60mDnbheN9ztsQNYlqXMTNerMZ2qMzDH/AzpAvGJTs7P2CwykR
lOfnbWoHu5ODq7Ae0KL5oOIuQE/azYXP+W5nzZE0+UKi1rL8GbmsNdpp3iCH6XDegUUPjdif4zb9
2U/Y4JZYH9yYUwJEerwwvevq/rvSIEJ2KNKzjUp7Uqa01V3PpPp/IVx6TvDiLDVGZXnX+X8dLGIu
GL8ZBv3gszv9xbGdkwbCU0v0M90dG8Qi4TTr7Q0uUscqmrl7Flx0bnA6mm1626LuGt4jekevd3Ju
gGLkZN4BZ59vi5eRLM48TLnpe+mkakUfV1rF9GhRlP2aT+rbd4gJXz3jHYUhCU3Whc34BT+3iWrb
Kqp6fucE9q2ktpWyXIeGtqOQyWpYWteSV5Lc10j2N5Y8FIBPaRF7Lz4Bd18pYXB1FsrOaadB32Mx
nGvtNXDzfRy12wSl3NzhIfI/j2o3yQeBieAbueHzLnboOjmgWvLKYbUPnALwILGmX/+29f4u6J8u
H31KOAFtXTcmp990C5/+IA9aNPIzjLZOgPgx2gO6o74MLtb5QUDs3cjktHOzk4TeUcGMVHjnamiW
/d03aBrlI1g7M1B4aIoFuwPlXE8dnNDj8joRixoI16JBtsTcz5Rp5ic3h3NTjqCM49kko7uVQNtm
DCdRbkwOdB07n3tBhibfPRxb0p5Fk+oJlb2Fj9sPl7iBht02gAgBc1pEoHPfVb7Ld39E+2rDcvST
tp+lSNyDJindVYv9V2uej9w0MyU9DkLicDr6wFrGSxjLnyQdm8aGt0Usni0xNj9wuMxs6lsEqYAZ
KMZHM9HNsRzfaDYSWak/3miTQ+0X7JDSwSSDFSGttxFtziZQvD2xsUpmtO5KiePRPwT1/ha8e51d
huP9Bz6B1fPWcefXnXe37WseAAKgnbs1XdHrlUC1SYiP/VNzRqb6WECbX8RFcOtejZvxVHchyLa1
SI5bu3EH5rByi6CPo0Q+KCYRqOhACGhWmfhIId0gMlkxT/P9LpwLD+I5Ynx6Z0eWD6AC2HBC6BgU
pbepKzXXdHW6Vpa1tissbYKboQ95Yp1dCVLeCAYS+xtLIy2WfXscPEE6DLL7ckNhNKGDxGDzxhIL
RONaY/4NFAzAENQPTyxw/Jt3XgaBK8NDt6HYOL8qf66Lx/VpZu5m/pciQiUypWQNScGWhhfhLp3W
fuglkcMu4A8MYJHwrM0ENHfzNgRnkTsRLp9tHGsU4EBLHBdc1u62Te2X+hLyazcu1LJGNRkldQgp
afG9nnpOAUIyttoIeR1YOXLEtsUOt6ntelAL/RwnBxKM0qk1m7T3yFlyndbv/ZAlNvcqa1/Ht32D
izGMduD12DXJF6uT+yTqrhxaCAQkk4ZO9qDLKvclmihxxMP+h1SLmvo+eZ8Cc26aM44V50gh7vb3
Zx6W+lU2/0KQmIhpXAcuXq8Ye2N29my7v7O+jEs3bM47Gn6qJFZrwaHUf1PqiKKhA9NAvUX0WoKE
A0M7h6JT9uazFBGU0iN79IBPKaIcLCpODyhbYcCvd4wDhQ0NWln+aXoBAkdNme6Ay/y5JZk55JUX
WioPAiM3/47OiMMhP2QlgKUyreG1clWgMeTy5piXU/Sql4/uejRcOo1vi9SH3Pw3S2SxURWVLh43
odMaj1TtfDhNU6CLicvL+bPwFcDYKXyOLNH5HrFtSWbS6iKtkD+uu4A+XE7KniBlyw6aYK86J/IW
zDNitHJqn+LiQUb1gU1G5IfmkDX8+ExF6Rz7SjLrDfcdwT/01Sd0JgJ84UDwVKma+YVJJe4IdkNb
88iU1fM=
`protect end_protected
