`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BAdbOnoWehP3HU/IbOS7NRO86297cdnjJXc1YcgEHKnr0Pig9veGWHWM5ppDzshH3n3ER+AX7au6
kwbODn7mnA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
go51lATApq3afPT//Ni+nP/C+T0O4/zAIaHf7MF2oLwsGxFENFylSrhA1BY+NzM+lIYh8gqgHbbH
IAO9aO2YdzXfRvhpP0UULy9Q6BwUvvvuKHZLwkNlZatsuUQNiVPddhkJNUl43H+/ivQGDNRCDEg8
GnH/1e1Cslrivw1ibaQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AU8q8w3VGM/NEPCMcmK9ClE+ewraadhLrDHTxPD0Cp0TF7Eipm1loXD1OZ62CNZfaiTohORe/J76
jU+At9F/JTkv1SISXQ9EqWlq/NNPvaYGtwut744IEv/5zJJOSwl/9vQ5QLbbtelf31JLuH2xIxE5
Es5DDzjjabRodc2Y71TYIDkRnEUm6CbVkkPUUakU9WBfeek3ooZ1WwIIGKEQvGnoELcxmWNNxXOg
qB5Kr5HggSkoQpdOspx7Jzs6d4KQqNen8611yWCVDUzbl7OJmFfPj5hNx3AcOM9/MXvfLeE+A+5U
0odSu/x+hxRtidZ37y1G18jwG9G6y5aNx46dzg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
IejuVJehXqZlVy90ooaZgdNtDo3LUJ8HinDzbnyEqcA6vVVu2Tos+7OA3yX5qeFZ9AbQdEDXqpQw
BhCq2lauao3B5DAbs/t2Y33UUF4jgzt7m98rkZverR9nyGWD+0UEcUKvoo8XPTDI94Iz5S770VeU
1PxM7B8dbI7zActXQzk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W/aio5uiTI6uIiP14NlEw0yRMNPLKDFpxdBKGJxQC9oxIjblYS2cJjYe/AZJ7aYkNq82f77fyEQM
ZlieSB2aW2GtOCgrluX9dGpmC0SdkMh4fSOtfdEWM1rz+mrAjfZ2FJRALK2yloUGbhQENITKZfoS
3l8echX4/Y2aVUrXWMOQJrZvRJPcUBBceVyzEwDke791rAD6W93z1VQUbMLGkTRHoeOLjjYjVo5U
Kyi97iAvPLb1EbUINkJHJmwB/6GYqVpj929Ej9NMsK0SgejihRor7zxsgP3GZAvHQr3rMY1IcGnK
5H0tekrSCAeYgHZRMMu3rN3OHjZEWr3CIS5zyQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5328)
`protect data_block
rLngGfIMLTymAZoGb2VDfxYhRt2Sg6XbojZyGWIfmSUDqT+w2/pshzFon22h85OHOVql9uIS00oB
xNaJ1CTsh2bWuDa9r9bY9Z7RUN2SzypBekGFctOG7BBLE8eFN+FqQNXZFMnxku+qxfLmvcLErFpf
N6ygpNT8a86n6Rjp9SvEYcITkfLXLHSOBCI1/P+/jWfpvNOD99tfKnktQ0j6dSNz2UqguDNvnDKX
RfKtYXpbqLBUIBlS79RvzKfLjqcci435yH/LkXaIdealY1/qdVnN07Pxu+15CzxRtAKOXhuuJc2y
iwF7Jrlu1npBN11NqxpxSDkVQG5rCZNYW+GiCZiu8eOcVWUJaLi4JUR9kDJPdt1Hb3KPLnKFszOO
vaxh/tZSTz7kRJy4SWdQm9mY76RqCjokBP0i6eR/OE0Lzdd5fNIPosD0+00CowhihNLW6NcAQ1Qb
ZR1/cVjQVqqYQVSH6MkJjeBGXeLsWjGGw2TM2XkRCGUN+QcGEc8DuVvxd7cvHkuH2eIkqPn0hNl3
Q1XgZ2b6CxK/bvhsHHiOaRET3FKTaBSn9XhR6kouGxdRI7O+/CMm757MvhSgXydCsEKyC5NRbyt3
FcgPeD0FdiYG/PqMMB21rHxdd7M8FMigDS3inzzwT5Uous+zBn8ym1inmHWvuwutCy1JPhdT0mhZ
xg98NiZeOx8yM6ZspwYXEtrN8wb2i+cFQ6ucG8JykJSrdtoqJ6A702DlnQMnjFLPBnTTqwUplm4T
+GUkWPhXawriCQE/B93I0/0XikBZjQoB06YXokS0+bqrPLmbCXnn4sOCUFUUnLsktU+owUSqN6D0
ph2AESy3LNVPCC0+ojGosLQd3khHM5GYsxAhAsqmjZYf/U5og0QnttFjQrsyvaY0FqENC65WsJOV
2hzh1BqNYMjFmm1oP4pLZOYz86KV5xH6ahrbwj2SJg5ieWnJELR4eaqVI+SAXJmCFg3SsPvIYyET
+weiQu9Mq1DKaoQESDoTo6PNKL2SIc7myPSlAxtOIUbroY+m8x1IN2VuC4ihlL/p2OC2OozggnqB
vqtNxTUNHUIrc+mb3u43eYL6zQAT3JKZEeYxzyJ10q0XBDD1ei2KGYWg0SL8mWVSbYGfRvrKu52z
i5uJPCApv5477v5CfYDIjCaKyMG/fs2k7mXoSkkfLfujHK1LcEDBo6Wbl4DpkG+coVCozyDZXE/M
OIwZ/65y74j+8LPlogywyyeIRtMeC5TBKnTbRfLRvO2dRD8D/tfJ73mxZxKu0s/IGviTDqmuxmP9
ZyAbEKQklBSig5sK6swpqw6/HwsHz2CC0Ut8NhIl8rWRk9couSqMbbDn03/2s3XaIgHyb7gQHHWW
mMLg3Lm83JTpgbqrXOYfrqj7ilApgnx8Yzip4Sru7WCPIoAJ66ix+1aUSLxLDO5Cm6CFhnwvWMh5
gt5KlRBlVSHPSmg7RjKT4DIZU54wUtplcbXSl4pOJCCTLfY8gL9NPWPi14G2uWYg+DtWsEXo1VsO
ySJ27Y3wm6wNdyilsO2L5Fk0AZb96MYMGEuweA4EgcPuHo7OgfmnYf4JEZuzTD3ln8Jq9HgUvRXR
aX0e+/OPK5SmIyrZ1CM9/trfeqGf0PW/zyEkd/Pjl0kccrl+r9Zap0Oux+lh04TYOZuJIt0KxlKQ
mMCr8UMNUlJ5PFrRejpUNl6219mOyOC7eUzHY0IqR+8Q8+X3RRY9mICshmSP9KTz5uJ+xjvBXFtD
4uRScvLF0h88hw6tMaZj/6K+1ui63MGCpf930Q2unNna0qXdFP51ddVAF3kgow2hNWVuCvjhGCWx
Eess3/TaGiiBjsUdKMNBQU2dUfnK/HOORDUqVnn44y5Nu1n4h/0RW9+Va9TX4BRD1RWGX9Q/TBaF
8iw1gEJB7vJp7aXwb1/FXggRys9/w8m4mvstVk/qkf9HokXyuwEm1Seb5OPBuPiJSJiunNHWehCA
hwyqG11Zx7ZgTSBKEuz5KRmNEBJu1mWghTESWcGOwIabI4vY0IJHRtsfwhCiUWWPbgJYqdJz5hvU
X0Y17VUgsHGbFlmxxkKUXpw25aBb/UZSsRspD4iZy+6N5IJsLyXt9aysXsLCGorMqw0xz8TmurYl
ubw71adrfoNI7+Nmpa/vuGQKilv79gTAicaTl+7SArnNg7bG1cucl3cGWAdKSreiIBENOf/oNv9F
K7mv8c+QJRK2i8gI3bZqVhHAuwY2RsaFaqWj14C1ksTChWKyPcnNX4+fr96rW7UwWwaTkphKZDYJ
oRbepvo1mMQh4r0n03qhJ4R89lxlQhZDd25OmMtmhzsdSi8Uo6y5wBvh42TN6/U4gEyckCgr9I+h
5QBirVUkYTeraw6/A01zgiNLb+MVxIwgW9Fw6h5+EfnLrAoJQB5vl/C3yc5J497cgBlgjW/0Mzoy
2V7DaArlGrBf2HntezzHaCjgCiDSOSMocBvvMwP/g01Gt0Ghlto/rnhAw2iN9HDAyNcWLiX2qxXe
knzcJdIAj5NgmLPPNvvuAHZcDaCGfW6iYSiXcX/YYAaWG0n2pfLCxdSanNb2209cYsKqlTy6XfwA
1EvvUUeFu1pDAVV53jtlpo2m7+9YRoRKrYLTS+aOksEmUf7ynWhb0+roSDjvl1XjZifC3N9TR3Ra
ciWKigCR8LBzopwCgDaroaCJqPZD9Tb+fkZ5j7mcBBajUMI5nRg/iAIPlFJgn3/gaIGOGIgL+Bz7
D8mCLcegDX/P8JGUEDqVysahR2tn/6NVZQ5pEtPQ4s4URn23+TCvDxFm4JZvAvf8kbhzN8jzvmuV
brDTCUVYhQdaO5TxKRRQJF4w6j/eqFhYh4cg/SRAvd0nUmdZTZZ+UR1HxCEMQL+layXongn4x5Sq
27b2psylVbrwT55ncH+6RYJwGEMqCJd+o4OOnLmjqtQu+Qh/krPNjG9C9kPrEDRqggYutN3mgBRc
q9e3iPxf4btz6XTp+LVgfls3tM9eJTOZ/ZDnE/XMvZrIdQFJButHGDsuVoz87Y0isGAvQar3RxHP
Bt/x+NSdWLMYfr0h4DpWWeb/4Iv10daOyEZyhW7+kuO9aLd+sNzq5pHqlmvousdfnUJJYN0wJ3bM
tp6B+1FRIucVVFXH/LI3+dJZ8cO4Gtpdm8OB054CaDUkOj7tPQwsud3wOR8j0xK3GTUb8EO8eHdP
VqBwkZQOvfpAPY3QAktX3bbaye+z1J44WoBYkeyPIL3F/v4ff63qXI7+jBa1U18NujoPr455F1b6
vfikLRNL4kzJ1/y0MvEYy92lHu8V1laTvYcVvlIr7yDi7QiNQtbhyBJQJuNSFJMeyTQYY2q1oaqp
fSQdAJWiOtvAjlVTckCszYZlu2kgr6XPKlXTf5Ntj02bIl0ZFr+rJH/PXO0eDz9J7fgR14khr73I
nSnoE17nIG4Oeppp3JsA9ADY2lTyhB4IZJUAoj4NUrIamfZtIDsXw8CW0EDgriE/NYsyxE079q9A
dRNDwuhRNzElXYRqnKngUtsiFivJCEXmSKtJMSaM/4mlSQFGKJ2La7lGUN/susTt+Q6B3Z8W3Wcg
C/tfuC+JtiRL2edYD/eRVh7Vyz093uSnSt+VFHiVUQKv0PEANpBS7st03lEE0Ub5StXr+3ZjGaC1
QlKBq1g0OK6pp/g7Sy/3jfoC7VbMYwGzATavtiChaYh6qc1cgH7KQQ83PEr128e5Uo0IqNGiyLVI
d8LempeA+CtOPBPOnjM3PsqTy84hvFn4wMBC54kpexyNq/lAxOXjfn/LuSOTnF4p2W8xhaZj79aK
3PFPZQOIRfkRXMMidUtvpO/GNsiceNXCyn6LPga0IDZm+GmUAvMnXRYaPGw72sYq521Te6QoUsdg
pq+L5e+E2tsk/3l8Qan+Wxeil6o+SjhUavwt1s0ddEAAMEdqi1bVF9DbjyyXq2QlhUp1gd4c9Rbh
UwLrRGBktfFZXS19sSrnRuPoJ+4xEgjS0aFHLNApa2OFMI353Cxm8S1+0hDfWyxHmVbNQ9PYXB6o
w/Y88L0salf5F1LSRitqergr89r7mKqC3tNrE61I8ddZyEC65tr8RyP5+96hdlkGwfaDH61IjFEv
O9B/YdHiS8N9BH3BLTcEJrircTqteE/jvnG0EA1gClGxHnzo/wjlCVslpP2Q+w1GEC8P/8AJTnmA
D7598SpQyCh6u6X7WvtUPa3nAqQNoM4l/iv3Qf1ebvZshPu/0VEvcejj+kTZqAqZyR0hu7bQQWks
bGU4llZEA7RWUac93VBMylfK41HJELbx6VyWeibJ4paF4wxdZmyIfoh/vBzd26y+0CpQL/+H9PGz
95prkYQvmH5vUdSbxvh/rQbDQNUDIjeeSEaWqlVWCicvpFic4rky+wT7DQ34fHX8Y/gNSSFDi8QR
yO3nsulfL4w13AuqNIQTFwrcNOUdyLn9N5nAVDovLBarTWH38j0LwbxkZEGpote9aK9nl331tk98
7daN5rLQywKGCNiM8wcjXwuSKHKPFInDb/tSQEWu6eIKfWfjrksOnEx+QrnuE3X97d72Q27bcsgg
JtzV62MxkDN7fPWvau1ezC0kbplTISj/0y66WO5WcCQO26WsXhTckZrIaJ9ToizUrdnwf1XuZQzK
9PQM35aQZhBAP8sViB7L4rgjHAnAIX6VV2wpmwm78vwr4oPhxClPdNJxhLVsW4iaoZnmb+UQ2/Yv
rZW2hCr+Qg50BIr1jgTH9CPG/cpc5KxZYvU5iGJNmaOmEYGIA2FPF85XZ8BqMsHi8VGFWASKUqxH
iNTSzQAxZTknFls/Xnw8DZ7zHypNtVNMSAr5Yatz3lCa8B0agCfPwPjYr8qFK83JViik7JDobyXo
rqmCFIvh5XdeBkkrmbM2T3f9jM5IP53smyKkepeAG1/hn+7mFCSdDDNnlr7JUHKHxPHebiuK15B6
XmkyXDjbtZ6Dd0jaLFsRHShhNBdDXgnv3iDFodxGIw05hUwY3ya+apzDwJwlcvobHVsCYZQ0SmH8
B/9W++jn849Tmj+3WorkAxrtCUvmDGSI/IGanhhfxrLOCWzNO30eo7FRtr9BqiKwZREEHeK8I8pm
OgoJMdaFWKAWxRlhC9qbr6+6uuig0kt32PCWH1Rk76b/1cXfZ0JAyzfNRtop/ctr2OcpKUKEAIMr
OONfs7cBIOIkDTNWrGL7pLbOzr0o3UyjWJ54CdU40lQlQdtlQ4RERalYDWkfxU6p9g3zAMpgY5LP
P6d3vIlDcjymyuyBnGPdVEieChBHWlRoLqJTMzgg44NKbQK/sefVxRRSMQrkR3irTu/8Vd3lZq9M
+LyFs4KVLe2KOi64+0CQTA+S1x75mYR5KfsfXhB4ijbsmctPHHqhJG/I5F6HsL2mTqlNc3CDBfZ/
RrBZw/mSIFSyzqWejqsIW2GZ8ayA7IAZVmHhVvlruXCbi/Fhi00RNPh1yqonXkMuC3d+Mhe7m9wM
tSWFACNnN42cLuEhGk92hcdh54At/FKO17qoEc+WWdu/Y8EJ7yBTPdNiOdMD4a/9c4oQE78Ggtyh
D4T0xIAaJJWzqS/bEEPIU+vdsGmPi4uC6A0tc6kzUlssQC+iU07R+7pTDZJ2ndr0vqxIdvkzQicK
AWEXEnifYDHI/RQwTmgxJGIPJ2zGWbQb2RSUv8wUpgV6sTwxN4p7Q2oUHjOaEMl7oxMFyglXLxbg
yyAhsqcJxep1kERoK1Fxlwj7i0kWNrR9L8oTh3jhsADAggZTFvZF4gdemjx937YIFoWOITifVzDg
M0ap48PtiC1U+3VbvNMsaFK1Rt3J3TY5/YGHCQ4LX4UN7c89QSxJKqRoSl0hgUs7fSLy4LLI9AAB
alJ4Z5IGCOQA0o2+Ox0oRESYEKCD5wA4AHgUQA5T/of4V/d1I3pHx8KuSEcJsE0DwIFzJQ6CUpZZ
wy74zQrANZEcL7I8KAuotwm5O14srMlEccVA5qCi+/X4lBdQWflC2eHzo5IFei91ljAxdm4UFWoL
WKD3yosZj+Osbeaz1gjB8dDbzEuAUndFjMj2u3y7oj0dnoQbNBY47+g19xwRYxKWEE5KmvEpejHc
dtYZlZRAyHfIx6XxX9wjgn2VFqekVp1UUyZto/PO0+qyZ9p5VZ5o5BmSjjQj9zllj76qBo89+qyp
5iF72aQjT4fMuYKqDtjkkZkCmZe4+tYe8PTbBBaCf560jQm9j5pFMCP6mAnY7NORTmcRPeQ1RatX
Fznidr8xPcRBT8/Sn1zNazPeyO6NE5wqKyt0ZkqJHbbSgxjkA1PMdtYnfs3oIff1+VAG3BJaLc2A
0u76Gdw1Juue6bdw8OWP3kMpI30L0prx40OJYQ966FBMcvEV/UBeWwPK+5TeJSNZcr1DowxtldrT
mO0NsnNrQPFSwLwgBq1qeI1jslgTEIu7KaQiBJU++yJ3IV5+e+2bawB+pXnC+8xIxMwghaHgBhLw
IbN4xmKUpIig/y7woQkiYklOuj6p4llfUi0Yp9ZopMF1cRLgai6UAcAKmk17vbR9fINlqk2QPVQt
r+Yz9SKKqI9D2ZiThngjOYFrR5rOt3AMKKF+aGgyN6Ju21J+TCwlIHBEF+6lVUSnYwDoSP2FSLZY
W7190C1hFA9Lo3y5MmzCxmR5SvUZfjJMvi0fzysu/tOkXEmUZMglbJ40Wy5XVxtJMFzNnCJQeRD4
J4RDXEmxg1KL6tE2Ka8OWrgz8HEUXSJkl5KaH0N6eZAsSBSHFslHad9aUlB9WpnBo7Y6Otb1t1L6
78G0y9xPZPV6LfHyKVX9OHIv3jtTr5bQU8ZJEwT3upSS+po3v2DnfujLXXX2x1LXuIdoTjO6O3J3
o5FPUIVwtnmm173fLnOvRmxjsqrG5M1PUGz6R3mtqtmyjJrACF/tPmshRd0rqgzJgFzvKXYOn+ZK
tsV/pw7FAbNlY5vKBejXMxoTfM3/6b9XLv3sMcq1VKYxT2CNNG3rNLB5XwcXd/SNrVzbJxZycBWz
XjdWE+Dk4iFFgARH6AIMszJIPJYDEMUH8PLPvJQeQ8j/4XJfI3zDWczvUfi/c/N1NU3glmYCUbDs
ATzkmzEPEKqN7sLqNiDkRHVCe8BfaHk6uJdq
`protect end_protected
