`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P1ZpzFBJ2GGs+/66/mIJyM6UqRrN8O0htEasQ03blbqDymy+SalwoKpTAiMLO6SkLvL7F4gmdbzr
1BHML+1NWA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Pzrpwr4owCQQKfrYKFnnZisYDCIg7Ar9Zd/U9Eq++FLY1DYC7vuxEvlKpYTkxTj4sT+3fA9+BHvC
+AQBNAGThT6cQEluOgz/QdNqTdWmQlTs33WqLNquer71PcZMbow4oWjZk6UjoAoWdYf8PTPFWBTv
T2xVzOBC0AlTuv1s8kE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RDBX5MPc9fZMG4sNxFN2fm68q45RoKq6E7BLz+rK/uacaz4ipjDoTMzHYXJCno18xWjNs3fAoLQA
qu1KLis5XHC4T4ZWR4bPGw1CoE/CdpkouDqYQRcAgoMSBIl+1toFKTaZ+A8Dg0QZukNaBVDxPiRS
3Fu5AVrSYJeCSy7sbZgOGprp54e8MVXcgQKv4MuDMz76vTSo22+dd/ATDWnXqYFczUQiGSOpMCSR
1nuxHpAJiJqiaB04WXzeRaI1/VxIfjhiBlJVCc6SPjN0DctliCzTtZiAk17nQtN/jhDF2oui4y5n
A5NrzgjZ1ny4wt4Jn/k1A2FRAaJvW8GE4TV5mA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
K8qr5qYixpzOGqWtk8FoZ+7PlZbUzgLtqOtudPp8SbkkaR7Zp1qCehWWudxXAlyBo14Pa9LWcGgA
bdI1bLsovc2Dr/EOjuOytKzvdJ08R+zNXSxcnY8OgbIy8x0SvqIkjcNDMdVjGsC9O3ypP9d6C8qO
AbpsqbeNbvNQK5aPRVc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pcR7+8W3Dh32LE71lXylaDvDaougnfKYdtQPsgZ5cdnHUhGEIskWT8EF4quhlwPYbaCZXVRDHGw4
Khrw9Khuf30z15nz1ZpbjBsh2uVF+YdHF/ywdP5QOx61f1YLaMoNT+LNMhAadmiieAtfnkW9q8sW
w7fW3coyOmjWv9P+sxMoVHzZMQdY5VIAL9JBPuTDDhe3TQBx/rkhhIVXIo1K4sX6nV462nlzhspo
TaUhBLjgFUjViWO8Cc8zOoAxfkH5kUIve05b58FV9ecVkPFr5hFUSMCMsU5XQa7XYIC49fOtdADc
dGPj5OOHCz2pcHXEfx8EiaH52mGSeI40qZd2og==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 31872)
`protect data_block
LePSP+XnkFidLkyMOvf4BllOrgIhYT4sF8wJDRUMRRK0xA6SmUKVtHQH5VlH1VX6KjwkN8chiI0q
3qMQ64VgpDByWwnzIZMAZcAYi4vL9pOEeWrcz+vJZKGcE5MzNSK6hC9yKfHWee4l5e0WHW38zT7/
7sZ7REnxLr10HGmeS7+36uJ9uPld3tiZUoAUSVdqEJURGGj6LaanzsWBYQBkClq2avYzcWhbw51G
oYWQUt1wgK80FQUd2KK37tfimUj+zNlaoC6Yjuw2Q5N5jNseiRcOF4R6N5P3UyZ9IaZzOn7B9WdA
Ja7VngyftFHqiER6peFQDerrEXf/WAlumX+ThX8U2qpWs+aULXWml4hT9vnOVQra6QFp6AnFWkgV
kkq3YeCPWrP/0yOvOm9vxMvxObO/HGiZafxpsMsl0ayuOqUBzgZc51A0PUog0E5LDInbEIPdpCAL
mG8Nz8khkhrc+gHK4RX/IONoJ1wAijvY8SYI0Qv5miidVMjNTY/N1ZPZXfdwy2hiWcGBapWfw4/g
3q/8rVTb3rHjuLtdR/lZ9XxT2XzoOkLXYAFbu1OWO9WCGGfqHag3d3aGh7GIPK3tBuJJih7VzkTg
Pa41l1E0roSx/oQ8FsQPlcOkFTfGn8wVc38Vm0Iv0rjjpiN935moIYGCWNPit5/xSMh73iNsHbuu
JSiLlWdNbnI3FNi3GAj+9Ngl3L9sc19SjqM4kSKcTXda3xvcmPozJ1ocqvbqTNiLcbIjk7Z30/Am
kUFvoEvWEdiC2bafscA8vfS55A0QDqPuLeR8AZhEIJQ8GkVlJK40tU6Tj/hNh4ARKHYwiAkv/7h5
xB1Yo3pcSAHZg4auSe7HaTTF8THT87anZBGRyb+hshxYfvqzobzuc/Mr4LMiUn3R3h+01rFwdoSi
hyZrW6ACrF4XcMGGLGtnDe0EuiB84eLwgQT8byAaS3QlndEJ4/sFTnh1u6x9X/RGAOjMRPwwH4yc
cwlvIRqcWuO3lqH4cjXrSvOAcPfw2rK5UsKDwfx9u8lPFu/3OEXISftMu80e74c5G4oXiZeF2LaJ
bhA/RU2U00rPHFLAuDd2ilLNfjyroUdJ/WamzIAADJHB0Cc+A6Odf9XhdKXr+MPcvQXAjLzVLOLc
s9djaCRCDbUmLaRkN2JtoQBxG0CMR6hafA/tmByRtP9WHPKtIU4p8UYzx1rl6NNQOwG04E7hZvcL
5X1iaWQ583QqtFKyqydLd3zB1bgGP/eURrN0m9/gy3Ac+LsFZJwdrQ43zZUsc7fJwfU7gUSy9Ruv
ieLwIC7yBouat3Zp1EZJW+4kDVTmAecw9mZNGpqNEGaTfSwubeSYfiF73UeyAhHq2V/n7fV5xfov
NE/sZyyleIEpzcicR+fdT5MzQxTPk++P/fVEg1V5bD+kRBucbCy36V9mvF5o1w2m6r98InRWK2g/
dHXVziMRhAX0qpkFc3pZFCWbiuK8M1BgvNVq3hRQs9TH4oaDau1pP/njKhwB3WQJsWgZlObRWm/y
BlrvIps97YKDTASajrtsknDEaxRQCOn4XNpK38DYhBxV18EjjAOdji0Rt0PQ0uA+O3rqLQb4omTD
h5u0sI92K2+OjvhIjyaHZsIH9/ODponvn3+uqrR7W4s/ag9gUMxV2ZmzJrqv0jQjdss1ne1JIktY
SD4Qhx2YNe4Z536uY6Zf7SjFcUB/4h4Rx0H443FUfdcB1IimeXKnK/kiXSFxtN7C2a/w0HJ1+wTW
/eUOlaIU6NtOWPgS9cPPW4HGC3SaWYOTteVDDSd/GNtA1pyCeXojakrSJCvWm1O3bcQAkF1ylvc9
jWyFJihcWJfV1EiOwm4V2T4oZsh8RyawPF+07fz5GJuncU74w6RcDsNCV7tZFO0yEXFIAnu1ODNW
hb11S0yTOeTpHgnDgZ5lbrdbBbMd32SUtqQlj/xTwvYz4DRGliZRSMzlowt0bh5MKorYodLUyynQ
WLPjLHkWwMerHx+WfeIV9Z6Be29UQBrvh999vdEqXVSUp4bZbkO9JFO4X7oVVW4KA6qt/TEya8eq
A7WEscoWpgT3rb/gjZTkF95ONqKaSeNbaAUEMpPD+OI8irlLBAsrrarM01rItXHe3l4dGW99MbDi
pHn7VrNaIMLLbjTEe8dbk05dcslpvZGRAyjU7sXrZYQ+PDQt4oEJ1F6mBVPVdoDJUUW0auPZE1BZ
m0ehDn8Qd6aGD7lOF4GZNTbr9YuQJdKG1ahvTZ7bsTPuqbxOGBJNDu017BubGSuYDMVPBEj1V72U
BZ/vXtULuuzVx34vwjc/kCuqh0cv5FXvpSLSHfPKLzPeB7LT/jPj0mvzdqS1E/+Lw29ChXPPVg1Z
ZWdPIBmxQf9+9gIuZ7KqvIv7qPFN6oPoQF0nHik13v/wxSIP4EVoOc0Px098i0Jr2NOu3b8vMo0r
thMegm5RDaXB3hEDoRuTBpTDilgfzFI5ErAMJgqQdNBe9+NZKN0Uul/O5JJjULahh/SyEtmAcuwV
XLa7I+pP+kqd9nytX/I9JY9fB600V5WDnCM9iJdF3u3894XEJaB8+Ow1QQCk4pAqqfm5IoyfzPZH
WOZ3bqE8LlPuuGx9KTvCH7B4P5joQ84+lsCV2UI9F004Xqsdc9VspfYhcD3y47Wjb0hoCUJwkJA5
DreJsEaWsfBfRiUK5Rx7VNkY8ZeM9PpvWV0Xa4dPZceo8UOQroBvJn4pSLySsl5mSDWvqvIMnwXb
zMO/Yz+Lwf6td1rnP4rzOJ7OueIR6h0A8LljcAWwH2uNq771Dh9g1i91ZIqMfevbeZFzo8c/6JTX
93qHLzA0rH+B5uYeUJQtxyOMuB1nKBZSw0r9E06ZMrvJexpffAYIYfHLcUvd2zUOCoMrMsu4StKM
YZxu24FfLs6Wj7RK+NDlg7eErF4ykYHjIfpoKerkG2yl009DNS2U4VJjQE2D1mixheXI2ee3MWPp
CfAJd1AT1ZHHZR1pu19tIXBzp84imdNFkqDjLhTNZqzAEEYUEvntCEWpufQWLsEKl0yl15MwwHA3
HKA1GjgUPlqgNqsPPpqVVHarVQjPStazjfOnvkdm+vkqh33ggSKriPAvMKsnyl6IEOB41L86lusA
LK2lDQS2843cMpNRu8lkwMHlEtB4Z2XgRnvIEyhOA7Rng5uoT9CeqAf+R+OfWKeMBC8ePmcHib12
s4MvKSxIGS6DxydE1G+0BmjLu883va2EGxeEyCj4sPeSe4dzkYDVhdaZICElsQouHPCN+K76OSxg
9iZgaUMAZk65RpRboTn9BtLIe5zzopknzo2kjI80yFJY5IOFKBuL1+dyv/rRVwidxgGhb93jSVJU
MRjUmtV6xq2hYriWu9g0krY/2jzITx/xd0DwxijVWBRGi0pvtZXzQXCnu0R5ecJavM0t8EjPBiYq
42A2EVk9wTlKNqwjA1wTh35GozsR7TWr+qzNBYHsxKsHEV5enyXQs41PV46mSXQSz0dGMmIVqlxk
oEEiHWF0ZNiU6kTJwZNrq6NGTvgLV7uBfI5sKU5zI5fWKHlTyOEhOl/s3cWF3hFW1zZhiKN8qZ8j
a3WfVOOZ9pCOofW4yLASKWZPKPssMUTjv29SHOszt+jpq5BtwRMspd39gKgwmNDFm+tmqGFzDaNS
zZEwkNONQk+RXkxchX/M5boks9qjyA2Px41CKpvOEttGEdHEjfxHdIEHMT+iqAzEV2caOL9jsQ0x
misAPqMKt9lY9DH6APmk+n6Z0UPLtwLwQjrdk5sZgmyWpJPrPjd1A3lNB6rGc8Ro8cStSTt320BF
jXsyvkjjQrPuA7zrU/4Ej0YEp/nZ+EY/u0YaN61bgBFYgpvuRtCQtCGMeZg9jW294CaZ6vMjrYGg
jvZVjwBg2KxilQKOBIh4BKnmA59X7PZqYzb3dr8FfEksPpCeEygleumdT8UWuMJyf3B9tYzwJRfz
VBX45Pt8EDqHVflv2nJI9/EXCunAPUVwD4TMDdAMTNHNVxOhjparldlM/J/QDpDWn7gPf/8Cgj+j
1nmyHHq5mdGbK/OaWgx2ItKCFM6QzoUL/PXiY8iSMknAnCOQfWRWZa8x1haqDZQupuk8ZWTzHUWL
NudW7ehPO+3TlWTT513Tzbd7H+yvacuyTsHh7AweGCWtrHivSq09s03mzfRhjuxzOFHbeky6BXiT
rbg0h+QbXdcPGEXmumwAgQAfYtk2X3VbAeKAi0ywpIQWjxrEUqyNkR4hYD1opKKSrfQ2TJjR7hvR
PmYzES4eqx1mDGiMwqH8iCKHbDcbgs69PWKe3Os98918eSOZaHhgCKDkYH+KdJTop1NQzX6xmfEy
AHvj+zQ7TR1Tqt7W5U/WIBZd6IW8KyZLB5pbSmQwM7JRIGOBCgpBT0fD/QgfBBNI4qyF9kwmsYo1
aTwXPm2Piy/IZdSkpS1E7x/SyLEJlxa/q+KY00OoxeEaN889hymNaQOS5w4oNn0wvXzhKGNbZEvB
fW2Cr8awd6I8BkwTQR6GUmuy2mO0AN96NaRtdSZDdkNygOqw9azolMQrHpfWQbXmDY9njLRoAnoT
ybaEGS3WoP44d1YtURpjIarSD0ScuqLdN+at5IG702KtkfKerVOfwf7vvePev4wiHQFDzyihyJ6J
KA0wK6kAoP6QGPSy2o94+7Cs5zvE/RUOQlHCFoBam6RPEOuN/lFVl56QVxky9aKllKcm7PEZqLGp
nKs9joajfriajY48al8LCLXVj1d0lOHKqI7be7QbliYhKrGJtFed8NlwFTLmKhdh4+EP7infYOku
ZtKpm9VGvZpLRi1bNnYoNvD3P6VpKjKamA7y6PfMk8FSqmbOq3lHkizUDXVo4FO/B2Qoo7pmj0ll
X1xUjgf1Joruyo0cvv8+3uKeG79186tg04iFoyqU76LP5SZufukyKQdSwY3+fQ8pB/5ryKpQjdWb
kc62yUJ3FEnH2QT7GRl1BZTl+bpRGHxQATJKsBUdd7cK6vRJNbprcvoqKrVHoK3NpJvtUVXs6wsV
LZoJ56Ua2GFog8kd48+bE0vLGXcPEfVWyOmBpqMV48PCY5stMofYzkTdiqUsj6Qiqu1MTG8FBuEv
1TOqwx7stQkpRQ4UGWgAT5cvq73f/1vXdiGMAcKOgX1vmADlWlxyzAIpINSZgrDlKL3nQPsxdS0o
GJ+5dhCqdYsj7NM8v5GNFvT94dSG8S2O1nLWbfD/hErSEtvaJe66gKc3B+You93nHxGXgdij9oWt
/YsNmd+utqFc/qiFGJ+9tern2jppk1uvBpgE56+zZnFHxXgwcLqTvANnSuz6X/b/972hqATunT3Z
lzTFjBHOBA77JYlDlR06aRLXj1lR9qXZvlaHM+YJfSyy/8hleJmo/gtxVjszHfJxtY79UVG9ZQSY
tO+SXDQG/pwIM3OkxCXlVeNAhELJ29QvIHAltK7iq4u37p55uir1t/GDcaSUilXqf66345Gs6nOR
+Y72i/WZ5n7uTrLh/QuLsPStrnoBvDBMBZzIs/VDnzj5Jju/ZkAfIcYm+bd++x4YlYYvwEesGYYH
H61PPbT2Pos/KvlBmbkDRdKthYmta41FBC6zP8jLOMqf+52I9y/019UWPt+t9DCkeiTE0c4/gCJP
kjLrXJ5GPvHxV87fZpGi/85Oisvw+Nk6kfPI6WMm50UdwN9lA7sV+SqP4h93upYZYdzYSTfNvavc
KQz+jlKuhz30BHJb1BNjh8U3Y0GiTo0RR7N49L5vqGmjBk3v/FkoJuPAYbM0VbFziVHZiAkTokJ4
j7fWS+EJCVEIZd2O1B6XLb7vH863VVOhVSU9WdM0eGeVv6QcspooUlSw57FBF6cFTEEwRSFFlvEb
JQsfyONBqMLXx626MHa5J50AKJBzqZHoF19hOUtpWeOrZ3LkFB9jV+9F4cc3b6QIsSE1ExrElMU0
tv79f7eaJC/UtcAY/ozQYiAuPn1YTuQ1cxdJFXl6YV+xX5AoOwU7ZPe9IY1DScZtHm0Ll/Q1Qxw7
nG7qG6BQ4+CebljvQ570mm47LRJmHEuYkb3AdXEtcuaKeD5wkgZlpwGVrvkMUv8132LuAPTYc7RN
VZ0A8WvPl8Vxxo/FrOH3X6k7ATKTP05gPcdujAEW1PXNvQctfZcpazcs+z2aF0PJYFY3u+jIVu/X
cmYM59fEW3S6LHWV03fIi/3Iqww8CY2u3GpepwR22goZT4MCEorR3Yc2zC0dsdsaKFIEKfWN46/w
is+GsC089KNzvni4n+GqhIlTYTctwTWYjZMxFpRG7rZW3mpRocH9vZ8JOApGYcuotzOVK8/FRN2x
DC4WisnHwHyjowa+pgFp0yz6aOcVnFqLa6SSoPRNskqDB8LkQNk4063TqapKZV+MkvmaO10qoo4C
rwuVOzab1JiVzARkZzV2djbnfHZ88K+hAUWksr4MHurSJipia1k2MT+0jVCbRqEydXa9E/jCXGRb
Az+hq02NUTbvBmEUTFr72x6XI8zlS8mwoA+olmGGGge62U5ohw9HWFBisLeu2brviCYt4tqge+ZQ
02OAcP2Oc/+6Jxdcv3cTSwuVtOY5Q1OyZHtsFkZQgQktCQAG0SMbJuodcUmiUS3stxQS1ZjPpqqe
tm/5mtz/9MK1mg+r6MPvR1tdf3LnJbHPe20cXOteQAevx2uOOg6kNOY4NG3nILcPBoCCqb7vjc2c
t4SWftZg4K1ZDpU9zLA0ETqMaCqa/DnraDa3Used5UTwrDqz8bufbjSiZrZq54YREwfAzH8MiWqH
+pC+p7rr6WoOEg3PYGNKNqrv9+/5YteFf+KBgZMFX6JlndnctEyHGSA6J+9QlNRYVljGI8cGhVis
dXLyeP6Fz+sOBefgtTC+ZuVwgyeMS++KOzOkjz3iLZ4ul0OovV5bCWT5KuVtk5Crg7KUuV0Sn4wk
ZYzIpVVfPoz9j5o67hdGspwNIyPnHgWJU7G01i7SBHS5LGHSmy4Kbbc4YM0XWnCQy32e+uknlr+m
cyog3J21UV7f1doq07G1TPjyv+6a/oBqRJJScf2+BhpTd8shbCFxwAYSu40fCcRNGhNRJkDqvqfZ
vfRnV31lktERrihJ4rhPKvU+y2Bkeo/a8BD/XE6Zh7aAwddJUZPeyUJMYpfQ6SS+lZs6Pt6/Ozoq
BGi0/VBK2K8tuIUUlScoqCsHC9KpqT2BRbO2gn2b5wvc3cMMZfFNiFnjpLke3DDxoFjKPdYlGKzO
5Bw7O82nehr3cq6toYH0CadJ/LXtc4VLPk4DGQNMGPizuy58dvjPTtjQDgrsMaOnY2uyqR5BCxn4
lmEg5qzACq+90xuKIrvBU3OXk+5EPBZ8HBiwahMyGeHEDTVhLPZ6MpnvkQJO2bfVkcA0vA2uu/0I
RaQ86/hpWKQxEAUlMogsOSwtRqryGNfD+ukbzqCrnZyRmon24jsnLG0vjZml0HBXP84gb+cRn0Ly
SK/SKQP3l9AgblrpZ8voQu2/n6qXFCqJlNlQ7z9RSJsYCal0gwMOQwSOocGXT785qhbKe6wBpC5t
wTC4Wryv8x8BczEUJ8kZAnh7k8gKS6Pq+AJfbf3C29rH/e/jmIaH3AjQLMb3iWLTUVykWVIVww7e
0H/Vc7XlJjzudKOmeks4/LZ85M/s6LhC4+qZqWLA+pp63irxjCvhm90BTMuTQSQTrlZd7Vk9doh1
OEOdGCb/Syp/FUUnUVbqympi4KLEcDVt27eLkd/ag7HeGSovKp5ppvXb7iv/bZO6FbqgrdHn+Epx
gdabVSU23oxU+LxRdrZgIADxvnWM4RwC9APK6STzXQH3V0Eh0NNonbXVnKBNKUXlZVIhPBR3V8Nx
O1oF/obfun/+Rzc6EHuTTV3PIyYWR+M8lGB88r02FiJ4UZatdkWyKCDmTsc/CLAqqUQyJj6UZsWg
ht96ioIN9PdWUgduuSMNMzVb8IeWbAy4vJG0VIY3hFz+F/RTXhhAbPLvZQdfP9hsPKMgZulK1LdL
xICHOhYK9WO3s265A/+dntsebN719wkilS8IT9BfOHXM1bjaW1eRXxjm3+zi4M2k2/n4zMBdesUR
b0BK0dh2RlaQFdxt4xQSbRxotFYBYtaG44A5AmMi56+o9Bp4mOv9hn7PdWUTsa2ZSAADSnp6TfZh
iAD/wQQMb0eLZiudQ/GsKc+5gPX8hNE/7K70TazaI/lm+vwmjWXOIR42KuHvGiVJt3w02OkWzkjb
ZxAxcq+ANP5j7TAJkNvWXTJyYfifaiNZvjaX07ZisuNj5GEQR7Yv4NERPF51v0ZRWL6+/6yJQ8ue
sv3Vw9CyteiIDFL7qT0pPOcLc68jrNVATaQ6jQ+FdPNdr9QIcA3vgGfl0/AsDIcjtTsiYaeML4I7
c9VHSJ5UYBDrNgRqcyDC7Ke8ZhY1K/uLerfNnuS71GleEgb/zAFSyU7SkhGMOanBbH7hOcte2qC+
oePqkHtb+9DkKlylOeA8qh9UZQ6aRse0qL5e3evUBuqhiz2l3zmVHdJC4Yu814/LjukjAvoXpWgO
j0j6ue2+DmUoB1c1z6DEne2tjw2xbYX/nDj0uZNRm0bs0ud5chuVVNZkjn5JhzORPVKUFzcC3Bct
Dkn/xTZVv5QXYLiDCtENBOJBTwzwfkyTwYI1eblQ78lxpxzdzPnvZC/jUFNqr2+oLSoJ9FlnlYyz
67ti17F9qmgpHYEfyPv7/ITXjm6uzFhOaeYrWXv2Bm5MlCeUr7rYBNAOvDXLRoM8ZL+xw9HZWW24
+F2hmgGXeAL5XszZOk/7oixTEtCWibdcefjmAZ+O/altgoIp/RYbdJazfpmJ8WVPHnkt3KSfJXgw
qwPbpASFjTuGWCCTv7Z4tyah7zqzAxxK1PBjGL1iceUTiyc9Ji+tv/srJ0d5oKrxVZ2+tSkStgeP
7O+XNwHBVtHXxDlxlFrGRipBDD9ka9sW8mUVVYnO6KP7vpGcqehBCR85vwkfYAEWXJQPjMkejSid
4mOiMYhrT4sF2nDUyl2mchk8wQbNIyBoY379Ux/1tMt2adyhOH+oBcak7Hfa3tFSpH5fY5sD7Kbh
DjJL9c4/YZ+tXEPrm45UKwLc4W+n9XY+/uPH0dZ6SRriyDkkori1GwjBSrqrkfD6WzD8FnlvL8pJ
v2DR2Ob/Gf2X4Pa1RDZ7ruLdMLa/OqwcQVmIT+NqC+ABfwMlhs7v59kd5DEF+H2HENTmutnproTo
1Vajr4aByx7dLwUQqfxjRLwH8ySCE7mO/cjzdumOUuK4qX42noVThuke2/yo5O2EuMmCJE2u9e68
vtorrLpnuJOp1hvzMlDXABRr6bELqvSOwer8e3S6c8wfsw2xlwN628j5G8Vv1HpMa9nXIRzOA1gh
O1p8pYmG5jTjYFGlun0kIxaqZfZupGvgEgJsKfN1prjE+nIWD3zwD0nLv0C8j45DBi4N8VLLU99z
MK9noEY6qxFHCdZhz8nqL5Vj938z0hXEyYKvstd3xTEq02m1ots7+L07g+9TGh+RqaY+6eiiPYvv
Fjx80Ft7A+hMSQU/cxLotkk/sXn5zslS69KINqxhbk6OsBQy8PQPRGAYcfe/1r50lH43E5t3oO6z
ZrGmVA4j7gepne94lsaYfoWoEFBWCqcN4f/NYIGVIq73MGYnDVp6Xgog3KzdGha7lsiQfTXNJJ1P
DC55Q9AURwb22uzgrfomi4ey1qNL442llsX/BKAKq69Ifd2rIgWSmHPde4jDp2VYPOSBeC8Iymjw
vmqel/7T9gxm5W6AB5DDSxQXSeGJl368ykd/7UZ3NScm/QocuRnn49cfY7jCOQNoyVQIWRHXYena
2Kj+YvYuDA+X8nh8KFArMbEWgH9ZOb5IPZiNCPNjVs4sZtGAtJzRk0rjR6jqOrN6f3tN/A4wp4FB
OZPZCorUy4+pGJBBzCDfR21FgSu2J9tKW56SG0ymHArBDHvsjoVT5qp9AW9fIliijazpjPiS5r7X
y2s2y2eAC0OnsCc/LBIH3Q+BZ9qLQEpaVevREKWzhSOBuH+x6+e5azbvoj+kZNeiejDuB9XBVtQH
xepDazx9eZcrv2kOAkyi3QilSNmnnZF/qfYyNclKFIGRDb6e1KXuT0rs+IG2Ttqt83vPVYMUOOpe
tj12Sj3RZ8b0Ok4BAJY9EIlROTXWgj/P2iT5GLgNg5LVrhHuJ/pkuskl2KrDhbzuTW3r8TekjqFN
aUU32aYIGYYVnUWJ6h2mnvkda3K/HnBFYKuoE23vsyaMLQjX0/JVGsQVDv/XMwm7ADZT7TLjGCRc
QEkv4V9TCQTyrU1pD4njkKUTueYt3BgRqGnDqASXnYAQ6JxA7doDfaBJMLyN5cWXIL1dJBRVTSI2
42amlfDvpuLl5f8E9Mh8MRqqYNEgE7ODcuUzhnJu3chsJU3UOhMAg64G4yxx1mgoOH3bpsdAzhZh
ee4EJuVJHFBK8iN7kKRY/JjOk+8nUXLCRRRUFvT6ofncHqSsklIRHhmfmHcFb9xpTyzaEFQdQFpi
nJFJwSfE9gTwZyHMCWpnQo/qaczSBdl09zxYudu2JCMkK9aBzST9/N4SxD3qI15XUgcnDNII4IGV
Oim6BjySe4w6Fwopudxc9SqRfs6BISFhSQSsn0aZQa9f/lsJNjoihRkoKjTi3OFVC2xOB8vA1BwH
0mixxJ7OuDxLJskWTbFg5YWt/HcYCrgP18PMZ8ODB0VCnkSeFEPq99/vZZNLKAJX2qMzkkAakYjI
WMI276lPUht2pbksttN2CokbwoxmkWq86IUWm465abSA1lXec9IJF2rXdEmAYaTvJZ7VXefwAZ12
0bIUF0v/W5QXJI2mBFZotr4JBJ9LdKTjUb4y/FSJEdyPWA9aVo+nRudQC0tJSDRRaBV/YkqmADqE
D/Ix0lKkR53I/nHf90S0h5F4PCv1x0zf7d1Id+2uZ242SQwznyAQ+VH2xnerLjyu07lUqESfwgMq
UClUAcml5X3il42P+iZHOAMFpYu0TKDVM5jhIwIO+KUA0Jb0aQsXPhsIKrdn31zCENJVRMh8962t
6lKMRNBCPqFeT/7P2v4bZ+6DqK4XacK3F3ngvnpg002TtMGKxVf0MbvRDGo6GWp9kgz7UWJn8UwR
jMw24uNdHu03izcteQSx9gK0alLIWLQdeb7LHUsD9GuvzhdLgjsjde44W0GcJGwmTi6iXwN2JK9O
rkm9Q2ymFhRnUQbVU52MJixUECyb6G2eGz+hYHlM3Ic+Go5E1hJVyXvPg68htOGYTTyLJmtfcfgW
7QuUzGUCbtemBFo3jpEm9WMizsZ8uyDiqpVV2Mz34NVOUrr9Td+GzpvVRhTbZdOwClPUm3zOnmlV
74VBl1Enw3IohNfiSU8YKiTxYMfTNIvQHkwOlZA7+zolV1ep88i2sApLtn6c5MUhBUcscY6KF9yp
oP0vfM9O+4pTln45/+8L4laAMOvzDIhAep90w2Q9IVnNSZ/AYiRmz1Crb7N1Bzicibuj5/OyIKdW
CuHP9Uo4uF1bWSn60pjbt1sAIGqtZWJBpe8rJWuNtrKwNqB+xDYYCewh6gUBHklE9GVWcxJU5dw+
3NSTJkCAsCqJCrhu5V7S8ksoPZXGNo54O3ABiI4Q7YsrXTnwnONVXePtXCGKfjc4HedkibCs184H
TWnb+irVBFYG5PAT9zWSzzkCasO8N/BGMHQ7akfN9Fkf49ZObbPJhfsD7MZEWmGZAClel7XNG+57
obV8UA2X0axRZ6SuSpdJFsRZCzWPklAcvrwZcYE7Wj1Tw38Bv6gBBHdfdSYSRuCOc2jSfJVs7Vs2
9wVLeopGBR1+G5/OgaPHIfgNauH6uhDYP8C1x83KLdW91KUpL5sQley1nuQKrvaYCtQcOjXQUWLQ
TVWcUOFvYsi5uj+5P5BMScLD1h8FrOwYcT556whp/HX7hxZ5Eqh5c5W7Mo9JcIccO7CNawyaYHVw
JJQ0ULa9RpLa1OEzUINlqex4lBA/qbbjk4G+KTlOLUU2O00rvyK0GF3vkZkhmgqutzLKwBqR6mie
KH6JXRwvzRTUUJYQRtcBb7Ld2eG3ORreNHH7k/0DKW+tskBVF1l+KDxwO93pDKMlrfQbw/UgvLjy
k7kRBam3GYEgOcMTrdu5vbsAVRFfvAeZODMIyw5KmSUDc7RQzRF+dG8NPdCyOdt5M7ocuexc8mV3
ngmwX5c/o8tXsq2lv0Qw7VOLSVbFrJ66f0U6xvW8esOss8wZAZbxaDvBCX3R6Jo13m+xTLsMktwf
OsvLdcswNlRrKnnJw/knh+FhHPTJLr6oElInTc0BwHyV9rcW/htfCeWC0JC3dJF1bf/4ncrocDZ2
zkdM4WP55wvllbrD3fX+xaWC2WmbtJgda8yuM5pEFFlKuRkzkySMMown7znVF0ticV7FOlVn/P27
E69Q0lf8TWbwPnQ2UVy+B0Nov5wNP+KPZne7qqVAPE4ldNziS5v24xotW0XpenL1xfzsTPvHAuhu
or78DG/bw8hnlxes3VjgQIeDnoge0o9Xh96DkWETJ3Er3/gM9GnBAJEWr19KjDwY4cnGZsxLm7AZ
/vOsjPGWkvxrbevslBiRG34DnZfKjXBN15Rg/+Xf9wIhI2fclO9erU4uatNitzkl+KwLtCDR4g8Z
KdZPJSRy8dYcVIZzQe6sBwChIVTGQx5PU0BuRzLBvCO2+LpifYMZZvGwhddFwIije3kJNgQWHSYq
x/9dCVRpgQOJCvdfxM2EIbzM7uNYl96tz3+/Lt9eoLXYQOnWB1j/ncRNI4bC3u3CQ7xvXygGU8ie
55zcGHNh4ZdghsKzI77cy5lZ44TstaVaDverMR1sjAQ1k4O+4Wy8SwmCxtni4iU3V0i+OuuRMkjj
PQcFNOx9zq0r1yFpAIg8tZ8yAxCT3YzPlE/0ZZzx5yS/Y/+s/RO4Ava8fcb4OEa5626aDlwKqU/6
YciZh6XVV4ZyVSyvQrim8D2gI1TvMYKFchHZ1LGzASok+xH3uJ9A74dmGOW6pbiov4CJBwe+sf/C
S7+MpFdpdp4wkTfRb700EH+5OebZqyiV/Aqu6yrGqq4WmGxb8HW+Cje7xnXunxdERzLVTdwrKSdt
CXP+B9XXC6bRg2n5/EH/4l1cA17goRp0bK4Zpa0Mc5gS+uZQfi7OjWlHBQg4NNcGQ9iRdH/uqFLs
oNe9jADAcuqs5Fw/u/CGm7UpXA1NhDrNAtW3Puefnvf7oCSS+lWQ2KmQLy3Fz8vfBi2f7AwAdU+1
8MLyPvMjg4NxcW9iaOLSwn/H80q/UTycxLKRTxL59c4VWNVLuX5T18wQBkEut5nBWx6h0IBr6FrZ
NtwwosnxsiSeKst33Rf1zeJnGMVxDq1+hAfKWYi3cOHkb1bIcmNwItDYQGXWkzXK9LXMhLmXQqqa
zSL0AyxKunBUi/mRKBb1z9CdrVgHuuO+hVut010xXvfuP8pWiWC+cbswWhsjhSL9r5szZ1N+HHKu
7/XGiztvh0L0KAv9pwyq2eljC8IRivBOY9TMsSi2EI8YXmaj093DcpYbOVfwBfi3dse+z3tEmABy
AbJMq50yYGWGSxLQbEzo5AbMHkk7vh60sbRpTDnUq+n4tcVZLVuIazmc44SAuHi57D3MXn4UoxV4
y5tnspANmBo2xIawdQ60Znx8czZxnwbLj7iJt4K6/XPXZRiALamFHGM1KxWG8mUbEZNdxX0/r7Bz
K29wPV8xzryMM2OpitYfByzDg3c/wXxG2QjJP9aXaJ20NKh2OB4pUJvp83HAZkNuf7bRKQzJ0CK3
qCPX4ODlV5+CKbhewXHARcSeqECvlGlJniCgqRUIeYvx+E1VYxohaE0sVII97lgUSS7KzEcall0F
poQ91t7qdkaA/I809cxhyOkZAH+dTZq9J3jCTBlIug21i7i8yxAOHcESloYGuJ1E6xLbkljREdHd
g0c37QFjKL+W5xUJblcPcmwe/F1uheCQ4PaUIt2ECOgaPsWE8oJtnUi8iNmbq1K/uuj3GeoKbFD9
sIuURPjrJyZfx47R6Uvf5Q8E3IYqs2DQkQOjSA1P3dgNs9w0PjhyOl4IjOGDXovYkUXZvJoH+jWa
bVOJ9fdYii2RG+vfn9YNP0PQFY7nBhabxDtrIqsbzNmSkO7IqgO5y/W3Ba3XrYAU6TpQa4wRUR2l
gTOHfLSVwGkdIVVG7rwwgfTexcUO12cgI3QrZZriV51nCtXXhDb+zdofxbJ3woUCmdHmTvUq0Q4Q
1ITRb/y0Cfhss7XjXnOiAdmcNEpy52MLIZIMeF9+ODM2HT229vQ/qzlF4nn2qA5PtMWYBrhh2m1c
JnjSft+x9eTzdFcBHLT9eRMOLaxyqxgpEYY5kBnfBTg8qwNEL87AHISWvX+2OTnSSqlI95RuORUK
8a9HBPU8jucKJh3L2pcyamEnwAw7/6HSo2Zygf84hLN1LJzSeEw2JmR1dvx8QaHaJ63SIVPF7xEQ
AqozRw2q5oLXv+twvEILAqkWP0aC6QaI1TRqiOMD0LvHNpIulJKfRZILRkLexF2oi2fpPoKs0xmz
cAlWdwWUgL5F0rXOm/s/KDHtLEtnWQGiupYK0Ydna8AL0zJFRJe2AYsxNU8NGaY7Fmm1lggXRkOU
xEyXnLIlekpceloN91vcF8dd02/COEWKmE/W6AWZLZwLiLCFhs8CpZO6Pk2flYaQbmHFSEUypTyx
JyNn6/ryuVeHsgqu+Jny+BwPeZHGVt/RaMLsiJwRArzBr6wlI4ngnhPiPdd5NN45LjWKBReR6/OS
fJWkyCxBPBleReqgWmScMWJiXGreIFBh3j5hWRLdrFn4P43UZpfI8oumOLhS3xes/ISsl9JL0ogp
1ST+82fmcXy2UJv8ZgaEkqIXW1oXotifzC9tvzobiQ23X/VInAJTyVBlD/Zi/FXkiVWcEFbuTbT9
PxBa2FQq/0kV/dUjBidVVU2W28gd+XiWMLw8NnQApr6rwZWkqOMhVlRJlSKTpL6wr7pp7dCkwEzu
04+yPi0WOTN1Hj7VsrG//mudIKjcoaKWsxQGELbdPjhfHAEKLv3qiCSLramWC8u4qv0xAObFqu9Q
HbRY10uhQ+mUviZum23bYh3EPkCCLdpIkz4c2VsAz0UbOAv/U9uDJaR7n7VOYOzGettcs0Nf17D+
VtoHXAuj9CLiK6FfOAYnXlJrgw/lodBLiA7R4lqCBoC1xntryHKBNbu+NWW8XViRB/uN+w3CW+Kp
pZaXsUq9I6xnnhKdiMiu60SNyGsLZy/aWBWzwQglUPCYSxmM2xpjvjKcL9vY73OtGn19gXrSAKsg
CnR6eqzHzayQ4PYgpa9NU2VvKLTE/1DbzS3O4IKNEd1FWe6YA7tmT5QZ1ySvt8alSAWS3mpMvpxy
PKZSj+sUbwzTJwMGEUnj/pWlPiPnc0n8KQntjUBL4YO5RMb3kEaa+8P6+/30tZXaalE8m9Oe+dmM
LuQGUF0wI/bFjDrbUWAV0bU/zNSzoNLsA9Qit61P1Hi0of8yCntyvOic1ImihC//96pixDqyEVnk
7R0iVXyG5c4J4ufsjqO10YM33mDcrn0XayEoLPLDQae58BAfQbCSgUTlUp8q3/QfS7ncU4kkC6Zh
Rcvnh66WvditbD5Ya36thzUgBQEpIV9pRuisQkfzbQlE23UhwpSRaiPaquYy8nkr6i0D6iPn3Zed
RMoKrMpytHmDJJgCN91hQXG7qBCN3Akm/MytaEQ1V+b6+yDjOyKwiXU+GhO84D9JkoKGHW6ePVzt
lFY1b1BSwd5wFXl797wS7eqhokvn8JVHV0IoViSpNkbaGDyvyxvt0Q+XkBf3wUZalvIoFrZAmbiU
oLrhBrzt5EAgv/kO13M32+rCK1SrGzOKkI//xhlrN1yQQkaxCSXD35F0WPfXuF3dkcAGbxY6Fx8S
sF6SYBEoPN3qYBKWre/fXt1KyQBC6Qt4VHexfiXepznQBP0UlHFCeGIJKqDPsDrjmJoJiHf0Kvil
j6KojziQRYGhhORvk5SSHoZDlJFkXyIG4tgVMWwJPYecABRuwrIYmgisXA2K0hqC2Bf1AvGwIuBu
ydjggXB1KuiMga0EaC7UjEFQHNdxDcaApGaWH/kvGcRfi3XxkeAhcA1TcnM4sjb4MMWyOjBvWDLa
v3KzG9yJQx4dR2O9Cr2lJb9WkT6+A806xmDQfMZlg0KBmyGwzZVWvRFBJc5NluDQkAetOKcZcv86
NAXAyp89h6e4AF/h5FhQ3f2c7obGHvurrZe0UBz1pHRTEv633pskjb6gdnPFUW+JBKg9T1mUp42l
YoldjGjBd26PlroLvbDj+OwYk7tJTizCecOdF4Bx0GfW86hjTmMJ+oeV70f+OnFZO7NnuDA1BTQH
EHf5cNoGYm7d0Y/bomo9wYxlwHEhOysRDVHMvGQmOy65mCjHRAUivSdvKt8b/syD2+R7bO6bY5jX
S3OBw6wehOGxeDQsvKrUskF7EFmUlXMa9X99JafQ0iX+XDLxFHs+pWWbz2M78LT/NwTRWKYp3SRQ
QbRB0SxaroJoB/36gbR33KwrRBhF7KnEispEDKMhuhOM3dA5dg2Yi4Vj0jZKg0tWElfObSfP/dzh
KtNSd6PgjzAI8ua+ie+ZYgzgLn3PqeQqmYaVmpOSnH0oxYqEcDllGB43HDjHwqD65oy7M0wtkYhp
seoS04jO3dqvF2JkjpVZMFT6uH1c5q8O0hFeCYCfA7T1wD2h9qO9ruXRffWj1v6NFGOQOiPFf5lG
m+2td9nL1OlzcMQ9PDSLhKMsAaL4QhMKQ44KprDBY6JvUb0q7vjNmgvJvIMabRF+hn39Ci7wJsQC
Zvr95fK2xDiYxd1qbwTfxQHGaE1R16pqJIll3EmiZWwEO6bQxInnmGCGeIzU+KNxoTZMukq0sdwi
2h7wTgknzOI81xOfzTPg49ufgmn8cPbSL877iC6HuRLNvJc8tcDLhdMbkGEZa9FUdYdb5EfF6DML
EzIVL3JDO3q9925wyFt/PrYvmYWn4EavMEFHvXvG8y3RyKlI6rl7C2wCGqTeSruIXTmdQh8AVJxh
EVkWGBaMGH3pYxt2bap6Ai0na0IheJqA/qds+3GAc0C79o9mFSfNfeX09lK5brkyy3OA232ym6eM
YWRl0pXLFavOb0zzCOSDmu4aVw+NIzrX34Fbj/P5zXDWNynQ3MzLlPmEWGbnTByCFTTfLJBNf0gL
MrFYe2ZzzFzOdnJA1d7VU6cg5dekGSwa/9AKNhiXBNz4MFONIDGIUQGHct9HHbBpV+ykIZRwKVoQ
dYUuJxl6St/o1A05buuTLwkrCUrEe8PV393pL2fEg7jqad26MaylG++gF730y4a/Zcdve4E+720z
znt/T9Shh3VT7U8fL2AnrVz5+f2Ih9kfiIX7vpoPqoxj1R39qboV3KEinQplF0upoqciMJKc4RXK
heixfo17v7aURQAn8BPXGVRuK+nJ8Do/veX78W4OfRtF0IgZbOjmacG+fnQaIpg/vvW/aQtFNkdR
KYYoMJsVADe2DWeDWUblHaswPW6ThvumDbdPzgcCPqblB64yP3I3uFYeohfal7ZJ6qZhWF8x1EcV
CWy3iPC+/Z3XW/QQET3vLxoULt1DL+5tC1f9AOghU4QrnHW8zpd+AYL3VV+hF+pwFHrHBhTdDeQV
LqZWVUtEpTteHLS14T0weGXGOKwYTT4qUE0H4FNxiQXfo7A/K68hNerTUDGJuOuHD1vr8lRdHMwo
nxpuvRergkBNPrvjzbxk68mrAXr6Mg+rYbEhDO3lfVHFMyu1u/kKz9I+FJEHdgHUlQqXMYeOmwPS
+kRP6Nd4aJvVSOSae576WxvjJ1Yz9CPPtulCBNlz8BguYixsKpy9FVZsJTf3I6oL1lWrF/CAJbAD
QKli0zFv3PTx4W5RTXa4YMRvEfF4q4S4LkjcFdMRzend04a7fHwoijIYtsom2HfGiasckLzKAwLi
vzTb4h/+3dYIHp9X6hPReeHD1nfP1zIn5D4Cz155Cif2pvEk9s7pXDYgp/gMxgZBmOeGQRoBB5r0
IIbQBwsg9MyStTPiWvT+teKwrAY/fMgVzPHpZAOvxVHhSaWqL40e39gSAwwG5gL0ffIFVto8IV6w
mN1CJh4/lbQwF1jGARpISsI4FR3MJBvpipjIVijGoxV0FPWan4gWWVhvQFnF7KFM3WcD4MGMergQ
+ceV4Dcw6Jxv3pcjF6lBOCu3niH/AhAU9MiYqK238ZJOfrx3z+DgQktiSjdplsulFZjYnqBK2uKP
oxfLghIDFczd/Slg8Jl2K4AJTeSCPgjJehCm0gaVjyss5BAxy5IaLI0vb0mVuv56a3v+U/18dN7H
FxLWMRODHVmcl3Fi3x7JvtSmUfKyCtqmIuHgjVc8448eZ3CrCkTrIlxR8dzF0vxh/mDetoGDxe7A
zwq7CtJ4bKeC+h3F864F9DNV6vn++R+fYFeKJuOpNrxJywXvg5Og7C0Zq003tiAD8CdjbbqCaYs5
E3hLSw3aBZdVGJJMH9HvmKXQj7Q6QDQ4XPsbJBzymzwFC77D4WyRsciGZqCcn0HOR1fwasCuc1fJ
c0OZPUJykzSLRS/ot3bmkQpkro+2RT8XRxh+aCZjKSQ2T/0pHOdTD+301hWsr6sDCH1wRyNxFIQ/
7cGwy+b3Z72zYcmqY96M41dUeJQlQgjijyE7VYfB58mlRdqjltnC9nZcuO4ofbCkxWS5eQRnmCRl
hfYqq9E3U4Bs81w0R3mEUI0p+pyfRK99NYTar2dRDYaGIevr6OicJu2kwt3wq3pEKAjMlEeECQ+G
itFYb3ekK04wPL0qBpRKJhBROi5sxgFEgtEd808aIc5PXiRpaMZm39FLzIlSB7bBUTgclFo38jzH
DYzdEJG9YTIQs+1xv67vYd7mSCfz1zluGH60wZHo2YWuyOaZ48x4Ee4T/YsEAsS0ny8RIJ0PJRWy
H/3eRwA90VoS0YoHxcZ3ELFUmBUJLhSisygk8ZFNpyS59wFZTLtDZuCEiGehGWFyB6OpsL+VRnHk
y0L6WIOiyzg5l/CrWKOajEShMtAoz9+SfwaHdP2xs3oqMH6KINjGbWvdO8Wg+6Y7Pun3sQ0Zb8cx
DFdgLhDClx2l+7ClfCv1mkfw1L/MvSQ+tJyTiGIA9ZsumWJudnrbsW4lxdfuozdIKrdk9RL/aJkH
J1+Kcm2ErakGO0Md8DOyPxleKGlWIeKL7ZWjegSNIt8ssu0tIDu4dW/nmvQlglhjL2gh7wu6DeZo
RDNLJ3upC9h7lYHxTIITHzqvaeHbFubZ39jqQzERyx6nC/9mjUrorZnROg2wkGSKF3XNu8Of14FL
rPnTi8mGyGUaqEImkbMnfkN01OoWbZ4OyQglMP7uN5YkdziBHUD0haex44VuwjTTECaX5EfrysMu
4aI7NSKTzo82IElI1m6ObqWVWmtWESUmZBqe3ZlUR9U6krqJOaaNBRZAZ9yA5saIFjZvUbQPrslq
gOOG+2E19b8zhyU6oPN7RJ74cB6vehLD3mjoZVEOTT23rkuKLALVFYKsx6d6DqFHEc5yhPI/aV9k
JXZu1J7vWZXbN2rsMGpzTbJTQ/w3N5KKcXnUxC0oGvMj+HirFsL0E5ExKWbtpBIk0gCGvwgT0Eu6
g1DjkakO/tAG+OwIq/KyHpdu2vUg8LvzAoRNbjHc0E1+XP19EVLvA08ZoRyu17Y/73G+07VsPq0r
edhCqHT9/yEOdK4QlWr1xS4Qg01G9eg1P7MKbG0TY0rCAIAZ4ffwNou50vACMCw6cqvFu6dfFI3J
mhrGK9z9H2ALj820Cy1MAGydPWOGpgUHBKbtxd0btxMeGHYpRYjfwq8yybCFM4MMRV5tfZeRgT5v
XPQde6dmkvdtZFleXHMiPIu4wC8L0vcysMX5/8aDVNTe8iZT6pR8Ug71KqsvKWk5BGAimHmbCUQs
GVNschEPVdFKpYTYBF4CNYcgnb+QF3HiwaI1KWWB6pquWUJYB0GQqbCzwPBLk0UCnyHl5BTgF6kc
Y9bLvvTOfzNd5IMuhoX6ogSjM1mJiPyctQ/j2J4RiipLnBq+M/Y3mPzIjew9eER1FLaIt9F8EOcb
Byvt++91pmNRykC0ev1+ZSxXYeL4yJRAvQ0mlzQsxlNE195tBr7UsSp4PXT8xiY2tyDCEun6aO1l
tw4zPhM9Ddu7Pfa5WmUMQnt6zoBXrhaCHofm95oLzzH1fqJAi/nKHM4mEMKazU5YBHAj4OioIdgf
/m2/iwINO61j1+hu9WTXz4LZGutBXJRq83n+Ay6740i4bNJsERINtYJRs1QP8lZREa3GsFGPwt/7
I2pQy4hwylEmGcC5M1VYiklOgw0c6FNs7/fTbxuqPh63+rxYdwDy6hEHXx87xBOwabu5XEiIhHuS
3G/4m9lf5i9cxzRjlPrXDB7N2RJrz4AJg0HY/+eUotEcAt7YJBTItLNE/gKLpi4jc8qtA4wcoqqf
KEFCcKdaXeFiRIEe9Lr4UdW7FDOgKuzjqyEKrzG4akGA/SiSX7So9ig7SZc6W1uO72WnJwT8UkIe
oHs1s0PWVxA1YzIHm8ZjwkvI78cIyZ8oELki3Q0HdhBE+l5rTXMArDSCgzfRyfJVFRqgZxsl3+2+
VVVKe/uVCznK8MxoHg780Wh7Tq5PGhDqBcf5sKtmdLfIYrV+9INS32iyH74tTv0zHNJozHUW9Y7f
/7XqJh9hRNC4Fpj4j43czndEqGUAPyqa2qzeqYDM/IFaGO8be4DhqI3EocQTv0AAqX8KiyyJogzA
s13qMRDR4TLKTacahas9rp7P1WPi0p13hE4Fjqh09bY2SHlc/rWYu6z1WKeQ4mwstrPGZXNlLK1d
ZNnDi6G0uxDJq1c6BZLTzN3jc+bg7f9ATOgNB/A7AIFQSxc9MG2X5eML0FHdMpCCmRFdg83Ruehy
mjCY1uf0WxzTvzDN/3oTaulmnjYzsGDyoy+p1mvauY0PCvtVvDLpNuzF4sX6Sd0jwI1Ry5yjUtrp
vKYuG90Kb0k4KUPpzld1ZZ5xe0yzXEgGh6ke4DfAyx8DFleZA9ZNHCwasnVhEkYoMKjQRLHEWhsu
Pwv1l42cOj5dEqy+UaLuvjPdTDf5nS9AmTslYnjOGzGTiHLT701t3H1B+dFHIH5UV6dZzLRSuvre
1lXSC4jtX5bGrM7HReypYvjW+rW/1/aI9Jwl4kiKckf0Y6/ig/LjMaKNnTndg5Xu9yfSr+p5+WOb
HTEhg+wso4U+9ZCp2PkefDHPl+EFVKbC0LdT29cTdYHMYlu0ums0MkILMLsFaXo/0VIgYWxA+DL1
Pgjx0QCvY3GwHK7+p2aG4yhuNy1g3eWNd2H+qiDEuvYmmrFQAKWbaW/ZWpqNkcCnx8aBlBSrEohX
hQraxew3PSS3aXTv46AlasY7cYWpq6DWEytkR48uapbMubH2rwYjpD7arP/YbVo9gutgSH+s4KYt
u8aXbPM5s9XcnOt/U6Ji/gmJdKOAO2xKkv8+/oxO0H+aGka+HQjJJVKhrLhXBXatdubezfMXiL+n
YX4ZrlOWymKUT0ljfQgcUMKd7IHYyNWd2XMpBAnzK4256QauSpx0/KFWUY0pPwyF4fZRfKy8w3BG
ERgocCvAvxMVp64Wxk1lbhYd+ifApi8BVxkuvaxM11D5tmFWa/98GTg6MigApk0/WjrxvnVOiCJh
M2OHvo3fVSJVShJGClSaCgdQusUu9n9J/w0TkQbkFFuI3B94dtxYQmsAcQqacSgsHVVo4z7lyIU9
fqnsIiHVgl/0SoQVQzJXKwifOXz+R3k+nScZFWNF4cSfkT0oW91UBoTBjjuRrKyy/k7ehgC3lLMF
YKG3pi2mKsNJHlUBPfz0qjrj5Tmn6QOJlY91KzT+j86cAagjyscTQtV6anQ7M/WokC7vBvMbFbcB
QD752tFglURFr8c5aa6gn0TMIU5BwT/skf9c29R8mMXAEumkQApV+i26A1nFiJvqC0QCP+Z8tI7p
d/XxenX/BRQ17faemTYjdlU6dOWBpb9NkgMzWEHHPiy33AEXK+Cx8OeSm5k/4arXoQqQmHHT2tLG
seGSvwQPm/Lf2Jb869p2YMaCIeSyFvJgqpPWKJ9GIv7l6wXe1j6witMCnx+C0iTb/4ZEzda5tXr3
YP/0rQyQOlJnf5Ld3SW1aIPZEb3cFOV16pqWw+tHx/oTcMF9fPrIFAVcreWKGXFDCQKErE0a038j
5xK83JMsw9unapi4FIi2vgIZkj6GiwNIEdZNUfwMwzQ7jgN9jMB3UgxMR1/4NhTdYG61uR51M+9P
yzindw1cjch9kWZ4YqnAZ401hQ7P1CsXbhYQOuFr15ueZBO79UBYQm7cpxVJeqVmnITVlUsmROzy
iJYdPg03yZKPYA0QrGuLiQYtXpzK/TZEgOBBBqA3VCsjhJKiCyCiwRPjwJbBR3TBMQm1dE6T0zZl
qMgIl5H7P8KikmhshUv3Meq0t62pzSLOXZl61Qrm0Bi6JAMWGoyggef7ZSSVh9k+qLznxCr46pr9
VHe9eN7x+CfwmQre3dVKDDSEyJLWa1Am046ZQkw53bFypeB9RlQLj2FtISWvjudLoOZ3YcoEUipA
rCFpUH0jmbUzJ0AipGVx1ABf0mPUv6RsLHzUwe+MvmxD03Rwh9838HMN4ED0IrkQ/tPf37Xb8nnu
xqu63W8T6VmZkgg+jt9lN/XKNN6g0E+wKBK9ItPKtnIom58uZTOeENaVDPJc7jDXWiPoDC3dGZkE
xh9Dxse7jYJZDjGhjJVGKUcV5hG5tCh8mZqeNNefcngny+yLDrcFb+XD7df4nfPdeeQpdiGjik7r
jZXsoJUlTtDjH3y+fi2uEN6QMdwnTaMcBgZX36nCTALRSazSK16/X7Fv8cQFwo2liVUyVc6tT5rd
sjc/t+fQZvPlNcfvqjZNY7Q/RW7xUvuH1SOxW1sGlMahJd/aUCw51GapvjxEpTwog+BmwWCEebn1
8ZbVGd+oZxp+lgdy3RZATRZAnNbN3zRtu1k/iQNDhMvubj8bN7WXNBq+dY1SGzgbWD9fp8BQ/kpG
fmBAIPOjeoxz8mJNvy6kGcqTt344LZOf9zJRXY1GDN4Pt8FWUi0ZUdBOlUFOdXWizfTKypDRHaZw
aSth1VTBqoZ5KYVCya+8MNRjcM7z/wjdDjcXH1BRk058q0AcE80XST/9zp/HrJgZZG/jJSsLVu0+
5sOfXi8cqXoU7vHVdG145RsIMyIJYXbCUwYhagVC6pQ+hZEIOV7VBOQyTsnnwnW7rGgV/b4EI9Dz
l+gTEUX0N5oOgb32zamShudwebllF4kYZOrQeRfKT+sfCu4TtjeMP05dcmIFHpSKw25QocAlLi5F
qn/oDBT8XiC5o31U2qjCIFVHmpbhT99/N2H5hxPaOIDi7mh4r/p1ZYB9lbGh1Xd+iuepLntjACgt
weMHPglwVOJ3woNKNW1R+/O2KC+M+fCLntoMfz8o365HGnJhpCVk17aLt54HHwSD2EoyBMPNmiaa
yK9XgQoQ1RQDxtwUgiq49EqXjt5OaKUHJyEkMEDqcWYhZ1K4uhBhtP0Iqo/HVyV5ME/hMnd++gya
fVBPJcJQGZpJF4mTWBIe5Kgqrgg/U7pAAwLjLU5IUd2scENT5AZF3wFeTrIoSxRXaVCccThMPmOE
qduxkaYtJIYXiy3djm7dgLLIuyz+rh3QR+W6iZpcdQ5FDvrgdvM0xr6r1oXkGfkEFa7na89HGqBI
TmVv4XRrsEquPXriq9LHFSUZJ3YsXxJnpyp29tcVDl0lIvCPwlqn4OFnYf0Bajco1m9BdHYTF17o
k9oTnS9krNBAQlYJ+F3apMZV1mQn4MP7Ab+zNNTsbuH8vKMNG9bsRLd6senpxvLLqc77ji508Xf+
5Nut4gIOGsEDv3dEYXt4HcllJNttkJd/Q6X5NFByWax0LiABtTq6hJmjefUbWUhnBONEjDaRqAXE
oPmz5fgyTLMUOzrJEahZQI1Ho5d3ydxVFGK2corRbsjaTtrtpc1a8KZSiI1rkX1uYxrRlrEsOK4s
2+hmq1qljSquMeepoOyvwP3sIC7AEtN2uvqcAg4LCjhveKY0N0C0a3fzgdPXITEdx/m3W8J6cqEX
LsiSBbcRykf9XTT2o2DbIHBwhc3+/3BRGqRWX3x8oBZwEYoF3HRGoinAXmbRrU8ojiq7ZehtrGDb
jJgaC5wrHW9uEukxPfwcoAyt3mtwG85uJMNjV5VJeq/nx4HXVmqBqwdrTSEWosARkmWnnAF5/RE3
gKi5HWZVqnv2qbGlWwFIlCq0HvvZhVdC6PoVj9iH+PfjDwxk6pJ2eN57PTUoUhzT33qoy6/V3l13
w258/yP/0ARutVVd2u3HMQx2YM+abKiLEXEdp71vOksZ3kLx0HTjXx3SsxZcVOX+PdRAPGR2gYBT
OSO5tPQ2Udk1udjo3RZZ7DBaMWqTffbOGu6QcGWWNLpKyJdA5IdYgxApo/4rUmXTh9jk+nrC4KUu
ny+Nnp9qhxX4SubmrncgeMVKYO8nh7YF2uKqAiggL0keP7BEJaL4dL3WIc/02BTaZbg6iKu4+4+U
F4ZG46DO38L5UNMNFqqWbuSd2yksz7k2hJxPzgiyCUKKlzz4RMd2Ia30BR85Fx1kKeCJv2xzdgti
4l8yg0KqZcRLu4+hSCFZXF25M3FR5YmBZxMCtAuW22lySgrWBXfsuUdkGcdbzYSXK2H7yU0dSDhR
9iluyejPHQ+gqYXjzyLDba4+ydTviREX5zzR7rHGg2akYQAC8aPx78KlZHEoiF9CTYrQviE0tepp
Wke14wx+inHyzVJFkMXYtMfJAWmgbkJN4QM9R0zt8KiQ2pdiXOFnXRyXj5RSr3+RcM+efNlDMYPe
vDfHJexNzPVH1wypK7HI8+CMSqiHtoW+tc5xHwbnIl3M6fqfuM+5Lt9WGeCuWEiF+O0sjSJCCpvd
gCMczNEQYfv7IQxMZxpThgx/LAPAFlyjyVXcNerN2nBFqCOB1ZhLj7noWJBeCflOGAiyDTlDNCAi
rzxx7jFHa+TN/MuxnW8egx057VZy9gA0Kr/dMEsdn4Z6asYm8xV60RTRSb1oZ/hunx5TruIkz4z9
E7u87yZBolv2gEBMH+d2BAKv2t4i3wG7I2/5fg2dEce9+y7TqiOW8qh/yhlIx4Aj3z6eLJqOY5BK
f0V8+ZmFJYK+dvivJRcU68R525bfPBwYn2FDcfGB9q8dFO7LbaNu8oOz6aNsZtDY1WfputBZrKOE
aMd37XY+e6aN9wnFcubz/UmJMPVXN5FHrDwsrpIb3TGFnoZ92AHm6JJ71dBQhWi2tLTfit26w/t4
R/KlJmq8GIvhkJdswULvcwtbUSwC/6qsTYMh2efywpbpUHC7urBvsdu8CJ3UoNGmdXIJ9PvSnbGT
x0GCKQZwcz9rVYacA8byo5yq3KO2v05IQpB0sPnNndq/xcNpxd5WneFa/L8P8bUWR4cKKNuIyHw5
ojsROR3jXypKmoE9obJdFfYVwATYYPlCE+btgrpMcvgAs5b/i1E8cpkFEh0fjvFpzAHbXn3ueGnv
d8Vh3NoBsC/ej2Yd1gf2PdUs2dLvmaByU3z08RgJmkelbLo0vqaToAqMHTXFHc43Jk1tuB2NdhkH
OWgCdUr8z3Pest1dC8nlkczGzucI6y6hKzJBBjy2nA8DUWP5rgZEv1ja/q/njKFY15M1CwYla0cM
9z6JG4x49R4rTy9FzcicXzcrlWW8O8Bhd9xvqfm8KYWSzYRR/l5ILP9MFoHNBHzqYjYkWwT5WF8B
7tg3AGE14sGUcdeXjclEtz8aONVwdx6ZGVNj8ZFWh/46SQT/GowcdnkNp+W5MtJaPM4N8SAVrgt2
y/GSwgXBCs66vnKvkJshLSa8jTMbwxGdAS78lhwDSL9UGIsowBKcaHrcQjoxZoeqorF6eLwywaDI
4ZwyC4Zlzhmni6W0D69iTCuBTn+vNBHAwD+Hp/ufMIRqwiQUdKXxzlpFadsoVNkvId8lK+axdS4/
ZW9Qy+8cMJxgF7AWoCr1hidhB2GFCjh/gbL4HG/1UM4Ee0VOIQGJmZTc9vD+hTAb++7HIVo4vkBV
y22t1wfXZqaR/qQPQ+8Wz1t+gMTRHtLTVN38DRue0uEWe6xtti/okIJNf8AybMtGB37Pl+QxavbT
WOkJs6l/HvShQKr//9nY8KkLyVUfoRIU2+6zrxBUhqa2SAGYlwexAM3fwCTx68K2PgOHskPtx/q7
3u//J1Lq/xIhNNsKwLAYlFiWWTjrqaLDu8Sp+jnoy2ilrtvrllhSbxvIPShP3Pp6IeIUxfigttfU
IzkHtFycAnnFvVWe8vGy+GQjNSuxLqjqQ/PEIETdO7dh7udGWlePJbYNVDSZb61qUmv2tWjBeRY0
r0V76Ahf/zzUKWLaqC7lrUAMU846RPiY4c1oUoPW2FEimu9jFq/iPC62aF6EIYtHnDzT1KMInCvE
tVdFC41vsdWM0P3tFHVfpVI8ClyEV+2bYqsz6yU/dMqA4W1BsVh5YVsZn73wnmD69lZTBvJMyuLa
Xnojbv8/flf+Pz8iP4bt/RDMtiibS74svoTYTWqrdhen4p2lhe/xnYsTTP7tUj28+UQxobHk/gRp
bJNpDTD7SXXuxiMXAFRg9Lam5hQpcOHaisXtpfStIepy5O7zyPzrS27Xw+UsAspju+kU/mQ5icvl
qwyV1Q9UIiRHME8boh2wjEiBFwPh8ePOsrre4wGfu/Ea+C9qK/yZ3vWwCUJxeOSLbbFFezbr2e3T
7dVkGeRnFCstMtdUtIqy4mY+uZmVk+MYlj4O6l3/i7PK/8GvdRm67srse1CPMs9I+OrjcSO3o/Kg
TST8qSbglhWaSnqqutoWnnG4vowVAXtCnH+rz108OTqoxxqopkT24Xj8NWfuLZjRQ+amFj3MVfSV
5BBoLC9ARXz953pQp5C5xVzukJNtT80CzZXw2ULDa1r9vIVPEbRi0yXfQ3F1sahptjO8u7W6+uRc
7w1sjcOTj/lfXKBOBcmIcgtsNlPMMWiSAo6uq2Pby5GhphY7ZDc933uoBhEtkPPAGXdq6i0Iphc1
ujz4U3oZfaHcaNEeIwS0wE1r89derTEBG68iXZFfKlOFgcehf0INc9mQtkcsHea+8HpWJlOpbIPJ
eufF7O1qMHTpeFyNN7+kefy+ZogxpREgwCUCnaYypwgr5ueUpalrMkbx2/N5m+I0Zn4OMkTPniGR
CYlsAG/rfs+SoHd4NNtkrMpN907m5mgXxybTYT757mHTE2hiL9ecC6DMtM8gBf78j87Yjk8sOJEj
Y8ohg4yzWUKA7BUu7Ck0FtKmjZbAk7Qa4F3k6y5IlagQTLt1xnqctGcu0w+A8CVXRC9jdS5qaUVi
v3VrJ5rnh3I7TUw2ZfRtXpCROXgA1nRQRRjJ6Y9S9l2vHA7kw5PFnnE7xq/TvAkMXqWE0q2YaOIm
VIqV5agWTuonYPjrJglyzv3VL+zSoanHvHT2FXXbxLmnifZM5Q5uG5+G2QlEJGndo20k77kv92DY
GahrrXmOJvXUkxdNtn+oyAJPirZcYWcv9W4iNAm4VTqy83EUdk3YZzZydygxe4Krv6GvhsWH1trB
9L5hx+PpdcfAcaXmUnbHsaQGfdYQq408neJzaEWoih5Um9j1/VwQhURbDF4khd7gGEc54kB3b1OX
MlbKxXIZ4bke+qxH3BBl3uZoJ6lBfsirUVWwI3epFvLhaKSEvKSn4GfXQQRgtWQDPPLPAGB+hTPU
zE/2DOfF0fGoMk+GrHScA9vqVY1KvrVgQglKeT+V2yezL6BHaGdqArGxRdhW0JHARtlRtT5OIDJO
gV8xIh9lc1lclcmpWdWh96CwJqv4ONxBMI2QkR7/Br+IkUJMVRebPIz3zQuguv0pIk31JfOsvGTj
NRkOoCLRRhPfCgbk2v9ky/NOX7KT6Lco4G03es9nX3+mh2dyKwnYawfDvyzI34gwbOOKCSnywlBJ
c7445GwzOjmbrgPzcSt4DS6OXxwmxZYgHkHm2gWCxNeW5K8JmaYOmphgMdyP77D023d/HtwXaER/
KfcROmB/1zDzoXa4lZEcOtfVILMOpYU8n/oyT9MNzC5QoWluAvskyVxwgbf8pKAVjbaIDT6IDB6G
71XWRVVarDQidS0OLGGw7KJzgEHjh1b0QLNh0I03diRKNQ7ER2I9JjUAG3ZYBIrT1KeSHFFoalxr
V+tg5Qtp7gp42QPVcxrhDppPi5J40skMf1rWueGE8hJKMP6rq4NzzP2VHKGypTgbya5g/l3A/dMw
gKRTuoWoYzeL6H3FCIUN06hxX0jNmTTCdQjIP/t93LpMJ9TyHfmAkD4mehbo11bx/W6s9YBi4LU8
EV53QNIPpkVfuGTdPj3lz5SuzQr+Ij+pZ6tRMrGAC0H4G0sGsUb62QnoYDnIK3UZvNTcOUodLbES
lcp8k0HW7SEBah1xioHrrUmqx6R+El+c3LnOaqQk3/8Ef3s4xF9B1eA2Gl7M6OEg1hn0aCNaOIHn
MNbrkG3OZq6uXcE6a+dDh1ALqiEEdtV4DUVJPOUTE/bODH3hQF4qlo74SQPh9WVMsCjlyB9qZKjL
NDubYh03nnneU9pw8nQz+t7Eu7JekdgqhqpVocWWkajCgzI91n53A78Ip3F539bsDyCUJ/46HPzK
Rvm88DfQEIhIMKUKH3h7s0ZooFT88KpkoNTEo7s4zVC7TbK/vu4i+IPo/Mw5mcFIA2X3vq6+1Z0b
EYNQEcqJplqZGC3GCmNX5JIxpoSmWQU1zaAfSSMvKRqqdTsb48NvSZrJIOnxU0C2X6LesIi41ZtV
s/tGdLl2zK/4WCaTVR3BPApws8QvEsv6NdRV86npTtdusvvjlwJ3V5tSNSi1hzme1aiPqijMpSWb
43KtQ+bp0rv99ffj1LuuUEtMWOYMXqGg0mO/1OjBK4Fdlp6JqAf1Vz0qEBvliMN9U0HBf9bVNMT+
E5IWv/C9KMS8nSBxEmrv5alWNQ+ETLq8Fg4JhqVM/XYavYNOhmb2oNiwCpRVS5yQyLZxIzZfDg74
EhPOmx6iOWjf2fJLAdfWBVd27NQCf7WUSq5nr7RwhFBlePF/3DsFs5gdzrn9KlaKMe+yeIo92eiw
La6KUWwzDy66LlGVwNvfqYXvY6+tqUxcC8QpDCMU6KhonrgxXl3DycGX0CH4mbijoDDEW7zkUt9H
cTZUnfbWuDEss+v6cvm++lawhmQgl4j4RRDibflMwW+BoqZQvyP9aiOLmLP9+NaxyyuEECUjPlc3
HmUTdZ6B/vDqsWoqQnYaK4lKqhVtQgrhY5HF2JjGiYV1QQDdaO+nG1+gTfsuuuUfEVFKzv0OG1v2
mmAZEL1rf5ZQElqMJc6snx3A7CR4uk0bC3fpX8W+s+B8zmn+Hbg2yVVRmVS3lN7IFHln+uTlEaHF
06WtLfEQK+UmRAUiC1IzprzpPYclPYPMiLM2RiFYpYXmftN5/Sbf0HDhnBKAWPu9Q6FlkBelP091
kgyUUjeuDeM+CjhSXAstUTyNG9+g/PwjiBagVTUYOxjsfprkJARdg97hdk/AfjuPe6OkSdBnYvMn
lYiFAG3yFJWNLvC0WTP9AW+35YPfl4k9hAOm/pd28xifI70ctFkECnPvc4vxfvqXxFGOAAvr4naK
BIbRkmS0Ww45hg/BgCzALbNZNHEyP5Ib7jo2jTc1LqLvoPId6szqh2ufGtn0ljc/9DOGbXIw9AMt
kiPTovGw82LQ7ng11iXgrXA230uG3tNvMLieTldNLVs5pAQTPYEDQTnjDCSKCNfY+HM2XdpBHysZ
ONgbEH01LhZ+Rn/6fKkrc4UWG+STJNBuGamU+UB+/pY045CNX5mksJSH/N4QH9JMEvSypDZOxh9O
CW1ojhIutoR1IKP7Peyu+o4kYxqaV3TUpQndtWKUavt+1DfRvxcFkzbzxrRp0GsL5fWlb0qqZB1j
pypDTPhu60IS3P/Za1h/A6CX79XiLi6tOE0dbB2DVpYx+C7MC2mxLKg3qAqjan9HynPce3EIia0M
ZkpvW0XkFmdC8JGaIDZ0XomHA18UWvyZK4CmTkX7BXbvr0fxTwfNiclxPzT5AjNeNt4a3L99ZNNI
nbjv+6tVq9hQNHR0noJlayDH74pUStk5pwUMUrTt8v6mffPOpBehXNLLhacG7u6Rv0hG/77JSGX8
7cEOT8M7eoSiQtDP9DAlV+LFqJESUcm/YlvJm5DciqXoGJdni72gn2IGY6ofWYNOk4kPKdM3whNW
8ywi9lYmfgHzvmmcgtvSN7TJs7HXBoIPmebzNqh00H8W3Jx0iymuPLjhAtcc5gScIeUFzkjK2K/1
WqG8X7gpbiUK8xwFrUFZ6Z+eC7WvMATJkTAQh7qDDxzv+sz+5tJ6tttDt+U7QvnOYJ0jEIR+zoOZ
AR/19EC1VZwW5NSd+3bKqcefqeOROCi+s6Il892dlon5maRqhqX0fCe3kUxzzMwSBxzOsVgJTZT7
/SCVm0o2/9ynuCIX+UwkB+QlnVqFqLMbk0t+f348IWIRltvUN9ZrQVgxGICwgig5NYpgGSywdWuH
WFi+9ofi010Zi33WxH88sm9dbaEoAEM6KGcvSvUj4ieIOcFmx/gRXmBdddHDgqFtFng4XQP5LUWe
CHLy4X0rPi2vqsrgOiusJJ0tEzYMEvQr8DENIZly0dic/eVWBuq/3ZXfleGtSuYFY+j/FVvMDxMy
eCV3JQ9leDme9tWPfeRvIgRL+v4rlDbaIt4etl1Ntd9ZwP2/4uyB6xX/ujlJAZmJ/AW6wBoK0rOR
2rKesaS7uhWMYtg8T7Qli56MFZt4inxxddJ607Thsh3fK2CBmGhjDO7spSA4F/zVenBKWzgCwLBp
ucHBn3ZuGzTcxlrhpPvsXA3w0k7pbDk2Y7OJ91Jh6P3nbIM05ccf+9YZ57XG6BF5FGsah6/7K/CL
uIAOQvTE4833AO+FXO+dBejAN2bcOof3CYus44AqeqaXYwtCGGEMTNnNQ2nEMKYNs5U1bvkjarud
Yy618Td5b/drTtSbYBIU3poRy3UFAHH5dvN1bHwNB56o7THHwwbRfPrktc9DYOncO1ZmxNaJT5Hn
AMCru5ZGOIqdM3H7BHjMsMimDuW+PMAnvF5xCASKow9g4LoHhEvCTK0klMv95UudkurVNQ4eTySc
IJ2OgVgzP1/Z04RFkPXrjlTCT/CnRMzAMg/ik59HYnnVMG/JdJ6TaJ2dAe5/K9AxJaZ2hX4+13w+
imQtOZ8D+//EGluPtkpHSx4Gvac+uVWhuIqTuSCQxR12qtNn31iUZtUxRqMNFgLtaWXB3cBGSm28
HmRm02Z++Vxtz5IysePCc0XFUEKT0ev3p7lxsAoGD/9HxlFfphtJLZxsFClEFHHVIHvULbzLp7VF
gxEoyGiXbSblYvKBmtTGWG9YJbdy39s4i7G2X3deBSJY8ae+hKXNG4iLqrXOPX16a2ny4LHWl39D
1C6Set79uPkl80mdiH74qgZ0/uyXucjLXFjG9V0hwXzt3UrXQpZcIfx5SZa99PfkXPEiwk4ujNa1
pTa5n2TudP5Abfcq4jQoZretrMme/WDiK3hcJFF5Z49R+XcSPXMoHpgleg2r2pEmN0Tm6sIV54BB
OWhK/aBNLM+IPIjf9SpDPccF+vP58LlTPIH/f7bwxJEGF0/dK8p4oBLPYFIDfLTYaH8+dHVeaCYu
+RNBoGx0H2APdD66MYeQm1ny1ZEL5TGK35ZnqD+ejP/Zf+BnXTkUAqzxeC39jkuPn5fQoP21aEDx
BYUjyYQSE7/WKCDR5CIdmydvrnkgzbDyRF4jNxOffT27O7qucMAA10LRfPRcLHzUbDpv8hpywT/f
OCRVxthH0KjpSn23Dmttv+Uq5BGJTp57d55FsYYElZD4dlbPf+uI/6MAZjwR+4JRrdTYAbxw7hcS
WeOkYgqr+vVMHYoTxvliaqUjjofWjRPcXvEBt3yF1fQ+s0XpPB4gyZLf7jvFRCkcc4cx2ffTkUeY
/ZklP8RlHfvO+DO7ta06jLJoy0VLuasrWOIV7NZu7RFSARFNdbmsq8UeJxkaq8EHHtyUvJvRAJ6c
/GgHMQ/3MFO2IktVmyXerrX8FVPUzvIiiEC2VlgT8n6Hw3SezNBMyTI0P9WzOVIPafVthLkVJrq5
CxV7SX5NdWlJmZpBj7yHXuRpVTKon/b7kxuCOf2Uf61dhwe+G4nLSne5q/f5+hmQ/7uVsRaixhyB
nCrypCV5wmi060xj5965GeiKwvd6oU8U4bX3DdjNmNbQAqjXwPcNUksM2wRGepnU3DV5G3SUeJDS
NaLJimBWLR72tGB4qa9qQFCAVSQflrRne4YNOELGrjfy1AIXcyl1KwfueY4wYGpM6TDm9/3QckkD
aXcVrpjKFLewDEu5GSIs/TJ6JDbqMLxflQDkHvNbjgZJeF07PulbREuvrB6AKBuhM5WvGHYS+4/b
GdmoYxJEABMXYr6odv06faka0iYEtEm5o3faDGFIZDBUgdkx9CA/16yunobzAvWWQ8Nv3tDAjLZU
HVI7oGzDFu/I3o0UqAqGESmiiCIOOD/0WbiVPxhOT0nZgS1GRsE3M/QQs3PRegELb6nG2l53qxPX
tVs0eQQSeDMzBINNo80OHdiRiYymhFFrPssj086iNF4SQPEvafn10OW7Z86Ue22cOuxBCvzqGGiP
/+dwZkpVi5xI2G8Wx8FnToT1fd9GtcJiKfv/j836AwZPm37kOsubeyO1PT+TJAe8jd3xVTtTd+xF
DYemNATubjThukPXrdN9J9BOlfJ5cTnNn45QBwHiuM7s9WyELZxMFt/iVk7zct8eKxlqaTqQWg5R
BBZmnRE3Np0ZOnS660eIBHTQrxHGrQlF1vonKNe1oSRVA3zffKz6Sk7qS23iuo4DOK5UOtTMvHJ1
vpls3zVur8x4cgAIYWwsqu9ugB15cg1+wxqrRWsEjAXfF3Rc/Zz2907yG+pVP3bHytpVYFQv/Y4T
pOLhLbWLzzcqY1Sqs59YvxMrDiVC2rZwaahmOBJERK6l4AhcDP/+l3PTLeKqyEp0TBZ7AnABIdny
lNxhcXPCaDY+DgVOWGUgRgyv6P0eq0cQNw1/Qt07pukL7QJNC8ewT9o2vaAyQ3P1rs3XAZo1wjm1
3Ha9Oah1KAHSFYWV+770DrTws7stLnhbf1hcEyL9Zb1PyNFMpvtdFp1bs73t/eE5ne8jyj2sTRQM
p69jcmvccTWKoXqxyvm6picjxFWbDQlUR+zCJS3+Qs6N+gnpyWTQraOJzk8izX+Jw5vlwoUWhXDR
IOEqcRnHTkI8mqZIORDL33ORT8Ha5FREyfvhaORo3/apHsEoEg62Xu/xcelrDwo3sD25yO3ivDbm
vkoWwLCQoXYIOQ5diN3v9RwyiFB+j6SRvd7ozIKg338ib+iNsNWXaG5i9Vz3G3OTFSBGl5oq5cS2
owuR2wPTHldPkHyWqIE9yJGcov71Jepgf7c4Xc0pt4T8Wckwu94coipPvgfLrIaejqDOf95gOiwH
ZLj1/4gPAJbwXwBPqeETthtDBxeUZPdnMLQ2GawYE0/N/ZsuV7WpHB8a94WXJkqBThFtB5NZjakQ
D1IJHtf6KF9+PbgK8d/fWmoT4lDt+MODbldAIIqx0js85Tp50gJSEN0yHK6t2WIfRnjXweJR7xkO
AdnwnB62C6U8mh4N/03j70UAdfUkxo6607mgVzJ3SEjDrxDurdz8A62Dfd8yHEP9GaNxFFbPeMVd
5J20dHSKTD0H2D8c1riGE8lO5gKgNhhRCxdTJBRv9mGRXkz7EKoqvT1+u1J4y1BQ9fLlM+9Qw9da
eJSWZ7vnnY6ZfFka9RmOmSOeDpQ08MKsv+kFhFRiCLd5vG2/qNd6gvgolqnvw2OO57iddoSLbfqx
J3Dwhdi7RaoX5v/pdy2fVr0SRBu+8M7GJoj+NtbXq4ibRxO67KrD83vqfO/+SO3z/U88Hzy1RuIY
Ung5jtZ2lLvisoGzzocjHDJ5PUIawN+eyzesvN9i6UMm78tPcwM6lbXp8ocKL+SxJpi4S/YQZTwS
EOApDBUr+i7m6sHSlcdzO5BgSltJ/zntSBfDXefW86mBx5quu0Vkh9nTIDDyaji7hmgaM9kPBNCa
1YiyvNuVgg3jKHT1H4/oA3QhNccthreQdk30LclgQapONtutcOOzyXZTM0J9MhdHvrC8V83gQbuI
uZxGU+BsYGimkFArSYlCSGBFpGtorZYSJjshqMmOtV41VFuPhhgGUzAgyHndfETS5UfFQ9CHyNd4
gFdTpeLqDH0hQgoqI/YdxVOzLrn8DceTbGm7NK4XlcSIb7aqe6tMtanDNd+WP6DszrkjTI8PC9pm
nRzbKmPVNVi/Sh8CDwEX8vzTfZaJrmKjwCIIkXK9XuXFRLS+kVUJw29NecOQrGcmN6yw3aA19KzX
5qoXoI3Az5ARcLmlCeA0GqZBAKAwCWLs/HO9J/8n3GE6cm2vNXlPXS/nr0vscrSZ8l8bY9m7GWCi
qFjHdF90gza3cT4lMC1EYI4Q6QuXtUnfuhNOxFZH/Ki04x2bHZbf81gF2kK92yLZZ9pRVxKp4f9I
j6jONV94EDr29chCeTbIOWrNh4wTqI6As6+cYUwPfUTSACDxM8cp/fmIgp0QfvggHyMzQxT81K04
dKBjSkDBy4hZ5Nitsrixm53A0SuvkDGW/Qqym0HZbB4Pp3Mi6MINw3/i1QXt2qpml5ijJ2nIwhct
f85aPqhiktPP0yQOfzwrB4QQ26Q3kZji1uIaO9iOmA0027Wq4QZmpsk+dgaxNSmTfKARk/MlgCY5
bm87ttuaxkd+JEIZ1CV0eVqf7tiQ2Fmhz/5d4Sfvb1PM1ZWXaTMsTvpzoZWq+7rAj4eGkh456EFn
C+lU69HqYCbopd1CtEaO41eQuHPXxlMRE+2oN0h7hcmX3DqutOiwaHfxQw1voS0NGElCBC1GLAZ/
O676cgog3dxzhXZFCpnu//mQH9nk1q3+ua+EUAtXy1KvDCltT1ykqaAdwQugFzBi/+2isbGj55as
IqxfmFCyxb5LuDKCX8nPc0v06k6uErS3fEqN7D8Jpd7U/eYOiwA5DDKlca0sFrw4l86M2sPpxlnk
u6SvHcIIPwTIbJ1AQ6uf+QP9T0Zk242W0045SujYYsXT3jAS8uZVUsVf9DO2Zco3ceyXoz5+h6zx
P0e2lVgzroSaYZxyzPQPmVe/CPTjRo1DyYAO0JMaBVpyu0cbeZRbvGMp9CkE+C1OrIc38AC0/sdp
nGAstcPAVpewh65rU4C7BTEOpFo7fCk91QqAIpKVsnDUHA1jy9hYTHcQ8TZ1sVj0dkga6abkLaqA
imulzWPmca0vh0I6uQXbQlS/A5CC/Sp9lmc3REvwVL3xYpF/VRak8fJ69qG+yCcbfmfgYr305pvl
xgaVkTQZ6RETYab21KE5C//0pVQpWrlpCzVsCrWEAPg2wi03iGBZKHaadKSeaclFB1HDHQMFIXh0
4OkBH+w09UKkbhcSSnq1IlnyUBC/+E7oDfNFfJ/iRcybwtulSiviu/JgcFEWNb6aJeMCsc0SXJfS
TDNDWHqOdWWE4ubFKGjIm6Berx3ReTD89qKt+b+xKRwrvpT0xWC5tfRh5F/jeuyt9iFbhZaRoXPp
gtYFQ6rv/tVRGXYJvPXWHskkKmjWQDIT8p1flbtSSxEPHnqKQCdvkirlFzEMFSp7rnkUrHxVoEy4
mOQkND45LuhrSpX8tx8umBx02DlbTjQw0uJuSkM4IOvz0mgOAvDkeeQRxsXbPE9hJNxngOUqysc1
eYmAdiCV5M70dFyWE/u+0E/867vAfeLU36uH7QbWBg2RVbL8FKIRCZTJEPqYbCTAVhey35eq6GaT
KaTtEUI9kyXjQm/y1t95/oioe3WPFo3G8+YUXzYo5ONVWjdFPOzWLFauaXtayLRRwgB4qiBdQCN4
JcsD5R6TXQMU00Hp38/u1aVgAYU4dByBiq1F7bMMQAk6jaf9g6SkVhBPbknyzol5/29SXfGSTjxr
CnYn5gcgJVCSNMVx4p5y0Cr6CDJunRaPJZ2mWf/16CF9cEb0U/+SY6G60RbuDpOjOOYcQeUUt3XV
y6IwCiYVbUteT9ofZaSh88tD0SRUHuFmqLdf0tAaoGOJGMnUhuOi2LoPFfNaBSLtb4VYFrbCF4Y/
vL66kKndL+jWrzqyOQzmOPjtaCd+akD1J2AHXYyHpY4j+wPHluTlTU6Uwnw8o9g4kHkmXsaZcGiK
TYmmsHfc57hROxh/wuRrl72Ax4tMo2U2VQ7WBlUiAbtSoPZ/QnNymrKLcbRoeH2g97Uwh0Lhss0N
or1oTO4f2Gjgkhf5Ph8RoytWH03NM0rPuf/xBJmtoJqBP+WSw47XYZg2ijusC6/toHnLd5h59Wsr
bj8yDARHNd0Hj2FnGex+IjjNJW6pI0c2SBeb97KfUbf9E9D4viXjyav1CtzeEbCPajJ5J7b+W0o/
WIX3V2TDwyi/cCVS2oT1WI/GaA2oE+3JcDB8ZFWzFAQq2hkmx1hh3Uv3akm3qjmCybBMVOXuvopm
4juwRXbtBJKYN6MOskCkyIuZ6rVYSvM48gS8xKCF1EPzxCTk2Ox/E3iVrpdNc8NzudEvqChEOp/C
OWxsVn5mmCD+P21i8PmtaQl9UspZUJLghbH4PeoO/oOxEh0MnK+Kr1r0YFgfPOsFPn5lAbs/7rtP
tyZv59ITKPyYdm6r5bx4VhCeNJ4lQ5Qde5r78+FW9UrE7crKXAuxZKE1IIEt6/rB1UCuk7QMS4wg
1qPOMHVQ41FNz90fjD2Fpw2FaLRMkclbdFt31+S0SaF8yDZ2rwMhv91yPTS5i4fHhN7TNykk3lCd
c4WirEXgR9nffKDRj9522cUUfOw9BQocCjClcZKuGwzcE02rFNxTfwSMizgAS+7yX549K8SDgAlc
gTJvEE3XO4mH5nj0O6qs2TjAYw7H73nHlm/DUSXrVNddcl5hIgk+6JtDXKrwOOsN6Uh6bn62XLkT
80ZvojhqzqgWgi09znIgChKJ+/UWEDdWycxjAiKffVpx60Z6yfSQJDRxiVj3uUPhRCj1vCDk8RNa
cqMB7ZLdf+E8A0IMfSprHb5BxyrDXTJjMKs03prjzox/wemVic8f2OoneAZIucdF+BmXRl0ZCknI
DZMSn2lAY76l01INMYi5TF4vdU4est7GZvHyupnf4zgOr64v0eFFyxNSoDBLS+VWnlDxA42viTph
CHOpl+uJ7Tz7TM+A53ICuaP/L1gJ0CV3NvT0vU3xaAPThOAjU8pZqxhyJmzUWDSSO+z/UsLiWomm
nDUbrOWh1pAwL5i4pg+LtSd0yAONdXSPZQ7yxOLcqVEjnTv+mbPnErcN2z+UK44LnkeXqXDeU3QG
9NwT+97/JeZzkNOlgAcmWCchyIlZtpJzZmSrba6Qowe6l0FSncgce9zruq3FrdaDKSNMq2ptRlqL
dx+auWVX9l9FkjHeN5pxVvmla++KBB1RHErUzQTNA9ZIQFKvmuDrqihzm5eAl6B/QDAmeYsced8b
6BLr6qOYYpe5NvJiR+lBPSHbpA9mO+IxE1M6g1v03RGGPnRgqAZWdrzHH8BqBeT5MxCNks8M5MCY
T4dQoFJoAWO++9+k4VJybUvKiwOwsOumv6pdnv8qBhUBHfNTGtUAf0pVD0cXtIaGgImSZCUzvwZO
MgnZj1Dmk8Tea+WgOZY/wFIKGg5t0sPh1K8VigemLAeGkBih9haDO5MsNCIkB8fUbHCFMxqSu1W7
9lcHtt5VAfOWkKoxig5VLPLbcOhRnEmkixFimEQWYykfaXOv3mdkqw1nR866qRHwVEJOphxYmOBu
wk+pn15eiuJXSIAk8uU698jhgVRPjLTrAVtRDdQJkG8NtieawKP795DFVD8hDPjE3b4O+NQevK/F
9NLFTPG20ntl49xribEsK3ark94fDf3+iw8e7V0AKdFmVLb9Yn/GBJ+AUl0H/waVv5DCG9dfnTr8
mguYsvDiSeOgKKI7i+oSJInUgxg4WrShKrhForpYmnGCdGRObRSFYGHrCn3d4SLTQpGCdrUHFdgi
pUz9zAMBlYgg2SjF35Ey5sUfZ1JvZFL2RWCoubui/KoDYSZST1C/+zPhbthYLs5L/mWsN6nCoYwt
Cpxh05m52tmaRNGp5/8OlDr0N+dnz8ucYvYqH8jqA7BSc0IKrNCi8238HY02+uOU2KEJuix0+O/A
AHSUc38b3J161UadFjnnLhrXTIE3LLqo0pxui1vi3h/VUTyhTRmHkB/unmYMfY6ncUOj8bZBUOJn
dNR7acKUx66L//1icko8hUa21bxX2Gd+KJWhwSa4PGDKzFRP580vdTcrEsidrqahvGKUr3rs0iHK
baVgXnul6F/F6CSUCpXvHELL3CCZWFZr8aT8I55e7xMIW90V0xNFR33Y9O99GPRL8rb263Aq11w6
Elna2reicpp7Kc94tLgR9h3fHjf6fECR1Euidd1qz5BYZDlQehY48Rr6kQVBUw8/IcsN9QFVmQ4m
OW53BRc3RhBZB4MsqiVu8DCrPOqQug7I2Iqa3ZAaQVPmaymiSP4blWvEXnVvOeAx8u5vXFn9ApLi
B9XmTqEKV1xeqYecGu3pRiukyU3EzcQArgjP3TSI64IC0wIW3wLlEgZHeuPTjvabjALVNFZ/7Pgd
L9jtR7egL56J9SKvcSdrNomwJrXs+ZP/GZ0EwNhupJFyNUZjKV3+kLYsk2igo6bx9JUMthAj6yzy
CYGvI9hfB7BfdHZ4AOVLUctrYODx4hu8Lk7Z6cbCu8loQer+ZvBHswTHhrgBOfOqNG4iuSQa3DTM
59DZjjz45nOIg77CT7oyFR9e9ZphtoBHr1ht19gfXj1u+PbDeUNM17frzaanIPcvGR1eBcrSWeJW
+Ihhq6IBA3Uw5Ef2w1znHRBYmzTrHnWzvjVLnZ+yfJEKuCgjETBbkQQhEghBHJyc0zTi2O2mMM3f
QpBNldNcws/jFK9AWzzgX/udRktGjuIOqup2yu441/fXPzL6g2jcnC9g+w5FoNU2H/lyO0TPjQHv
kJf05smSeE4mImq/RVfxfy58n0V/qhLG/ieK3872Q8FU/xXdYb5gtfiAnY7PxvzXDEMfpLnQYaGz
RUk8CpInrh4FOkVktbhanpcKikIhB+EEy/qEwsz2AkvlK3IVZC5q3nyHsteyMMg9GfJJLJo/DOMh
1Vt4j6T049XxEvVaXSWnfKzJztfB6yNMjxS8lQKWfp7VgkrRX3ek3csdaaSGiDiM2qjiHG7wUEz+
C2rcXqAi4WyN3wuJ3z0w+XfDK/X48urDgmQ7u6Ad3FJtL1u4usfkv+Le6jxc7IztQ51yGIP0q2nD
9vvgaFflUPUkU9Q4/yZJKYQdhkWqPxXPy+x9XakWeu9YLNU4OSH/64JPPSJmWC21IQzpaqvlt1dg
Yi5r81ryEG1P3E1D19r6Tdup+ceYAJye030nGPbHxfF0WlRjVlKQFKTgmZe/gfaqdJUx0gmbEV36
B/A+zKkUQQsQTqAzRsn6//Ri86pLPyXwWR4CdRlDc4teMGZhYmQP4g34SVSbimdVHuSVQdoW+PiU
R1nZ8HcRekIZGJRYpIJU1CWgH5r1KBROhoqpgrOMq41S4S0myXj38dmhiy9zWgzWIkxG7i6ArA2G
f5n6cFi4/coql4vWcKazXFFsMcm6BTUWte1SsBdtrDGolgeCBfbB6LYZ+DxwA8O5bkqYn6ftWfkI
9zvspfIqs+7rJHTIPkaedUw44HGvN9VxiIuQS0EmAB213vEyYohDt55GnmQ2Cjscl/1VJEh4Htv3
f+2JaDpevbhghBuZr0TmYuffM2mVQbZpuSww/n7YuBeewiNsnEKEfLIZkpxP6h1XSqeMnmQIjFrV
egeMgAPQ8zcrM0jH7l2v0gj7D91mFLvE26cBdnkfLhPzjAdGY8nJuAEmsZJ4wkbqSC87HLNUVXz+
+KVGB4tY3gujmgnF28s7GjQkR6SqbHmV4RACz2dUaalWWJJ/FMYjv3JUiTqqXH8ROlp1jsr13zCF
B0KJo1IrgqYx58sJUTk0JcmzPSTdzcQ6ko7B0H8jazisMViXTby1PdeZztLpXcZykjxer10dnDHM
ZtOW3UaDlRy6tyh6taQQFd6fcpMmKtKFCFW5zJkGbC6HnAoklSMQu2102ATtoJfXdtugr0N4Upzh
AoxIIReQRjQ7dWeS6KGtUyzKHBb7Gzk9ceiDF3hl+m0PTyZYDxnZaM8f56rFEYbtldWpVacnGC6R
H4SsDaxgE93EgtJ7jky5OLjHGo84fGps8iPKIUZB+FqLql554E38WvCMgJw5ucXsBnqpDIdDqztO
RmOKXcQ3oM8faqEoR0naujfMlshJkOtW1lOYN6JDq1qUdTwCYFCyAnTl1uIoeurp1cLpWxodbVP2
qU+QWdl2bNYa0jtKDi+rUK19uJY5sSe3/WfscckAXM5iUrzlrF0E8l78xmBYcpepIa3dSQ5d8tky
A7UgjEVvjCISBxO+l9cZe7AFgGXSl1M+Gk6vBtj7oLgSk8Vy1C6syGDH0b3KvO9DiOHRIhEcHnuX
XK0cvJqFEWW5Sx+ZhpKGXuU5ec+Xb+3m9OCD6TFzirEKWdAafLBiO/wX6njVEOcn8fIDWJigi6Ho
CT8Hse9AtQ/JLLMeh4q2Y4CJKoPv+CiiJ+i/Iomg2LgErEhFInvH7Ho22Lin3uafIux4OoFq43H2
Psj9Kh1C4i3BN4yitkPOtyyxY722C9zTSH0ysB1h15LB4uaOg7dmW7Ihne3DFH81ecfeh98WD8rt
UQM8Hbs7x9eF21IGVZIYAzwCRrLAaW48NcFdCXxztyXlUoZ/i6YEZ7b5chyMeXLZP+qxZ04+IcTP
1yfBs8ezwFOuoTd5Jbqy7ZoQuB7bkN1LMrwdkGVJ7xprBpW1smL7ht9K8IChuhNMhndWFdIFaseo
R69joSksgfGyicrKDYo1kJ2Oy13wgaDrRfCFeqEnNg+JKHxiy0Sjtz/7kdizXhzggm3yhZBGdMHW
4U2ss8V9faaS0BA/h0goY7JCALsPOhHZkX0T54j+A6osAHfpI6o2DAR0aNRD71jMY+c98qtbEKen
B8CVU8DYr+bUypuD5WAHuVBsr9rgekei2a/HnAZPHl2xuXfNckxzHmUtCqXsJyaYHPNER7T4diqX
ZxJCdJkGSmXsF6buITug0z4tdrsxhjtfzO6AqotOK8svs6HIBHEHknlwnn0R4+7V1PTB7T58pusw
BcMMr3E6BOkjTauDc1oTtia5EqLga9yZLC9N18EQrE69ks2wvkVHvxLgxUd86542COqpTjaKddIk
a1M5PYs0jJAW3wEL8+0AmiC135mDIPPhfykSY+Mp60DYR94TaHND8+XYQgUyc9RuSS2F2JP1aU5W
yyaANp+i6fYPhV/0M17AlrreEL7MbqVmLENg3nEktSOp1UNIks6uFxcnlzMh+LqdWJIxnwg3gHlr
jkLrTAGDV9xRCZRMNvtM9STOTzlhccYMhzO4yaUuIenzQjRIFzUW4U0kiHIpPcU7IMuV6Wx7mmee
ojOFikfEWrJBKbo/J1ipPDZXKN3CCkeA/YFckO+LRsRglg2sxlAiG8DqXS0P8sAtONml90gsZPEm
jXBYz7/gBW39rx5VMNFn6zQGNydWMaB+Zg7AOZtE2zIEt4e5cBq3GfwKAqyyjNsQQjbypgNUevMp
f2E3WzPdErBL5ct69KqXhjUiPfOaimrzGyPfEUzXmZtK96QIzs4tKvd98/f6BQHvlOwwgFm2/Z24
b+xOXBwSyWA73te8fwoQpGVTliiimvujYqocUZw3wKyrXJFEsrmmjbmioonpvXJmKCLxQDdtrn6Q
1orqhPyHoX8wEKE4asZ6CVzbH/Y8KKDxtcucyImC0A4uKIVLGGpFG/sfAotKpf4avlByPlbTEDiJ
qiQxOyoq0WWZiMZjSd9vm6WzQ6qWGO5P9D9SF534kx1S9YuzNJMf+RNlKqxLy6SNGYZXaG64kNhr
nXtwgpNz9gj1w7JOkOxeJnXcoFALDP3TjiQD5uL/B6O0cKOuj/W3GdD295BD+UFUcg5fX32o7BJt
xDwxuPY6JER86qLbmLtTTshIigUbaloH2FmzsvDAxINBKCjhceJ1UmOt45Yf8Ag471V6UnC1mOmM
S9xbM0fL4VBEck1qDAKUFyCIAHNBImq0zE0qByi14vSfy7YC1JF12zokwtlQY1nO+LRTr91bK9Se
yTgMjZBj8hkbNzhl2obEze4K4TVkPe6VJqMggGuWl5I9Zb2LLTbjGxnyv7BE62RgoqpKRRSJopK7
WI5N0cG4kBRbnT0506FEu8d1FuG+D68idmgp4hBhBCxeesZ9BaztnxwvFBj2iHGZNT7ftlD++InG
kL0vuaA+1h3HgYWxLuP9hrAOUHF1wC8KvhIzzp/2j7AaCaPoZQvs4ZOC2wCloekVepbJ40/8uzgR
7gsQScq9JCPR
`protect end_protected
