`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
d8KecUg0FZEzu8MBudooHG+vUyDDoN1W0Km/75lw4i8STC1I1resSSflIbbY9cfp86z04dVAPIrx
5CAJFomaLg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XSLbD/2+SqGDNEh5LP9LEpPae/btogITkLC4aSgQx5/fZ92RCtplSGBUhD13mpqpRdK81bxPGV0Q
/hygGnD06q/40rJLFbruFmXLj6WM41nITGY8V9GJ6Yef1YkoYFieWpzbK6pNljoubRJFF+B5gyrn
NopediIKolm0Ec9BYNM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M3FYtESaf4Ci7BzhD3g8A7Jj9n8rUn3DARC9J1NBqX4NE30bm7+paG3FmSYehbT2J0oDiJKa9Zm0
Et0A9fU8bycECfc2sfr0VUqwVRcY25ud8p6n+boW9z7Icw4oOBDTq67kZ1zwY5qqDjEhFemYuwP4
TkEkJnDHCYqhCTBN26xZSTi0y/sDMe9tUzAwI+Ng3dKbgjbSg2Lics9b/8YeGpG/NafN0cjBpQCg
1F33k4YymjnSQlZ4rMZfzUsM99WOH8byFnwMpOiKqzXg+JhhpD6psvWQ0PM9aUCBp65FzBIA/GsC
z/oEBShPIP6MdbVgs6AgeT+kfmGbEYuNLpYFww==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sAxnvUapeCYUALVokFqBnCqY7B5/gYCBFaZ4mfnL6u3nFEzjFy+f6L2p9THiQMmWoj9i6rqziPJc
dCXfOPEXQlOUJUuJeAB8U0dUN82t3qjLWTm4FQ7vTj+ge9OQusUELDid26m6x4RGgKbIia4SrpNG
i9QCTWcrnD17+3IkVOc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lm+vp7IXDizEFo4j+wq3u8SAcrBoUccgbOzKIUy9Z1IOdCDJ61oNqwoVKN7Lwhq+lDrhvGsx3E55
KSqrw85KDcpUXUy9PL8GUjHFMXJbtw9E8NfiN3anR7nV/4UViEMaTbo+Ak2VQtUhBDYpSFmIFro0
bjwmLkgeF6fbu9jsU/jA8HD2NyDjZVCPfdwG+6hq8Ks+C9oyDf1JQ0LjopkLLvP3eeeLovkIzlKh
pPUtOjkkFIUuNd1cHJZxukvz7umMexhwOmlYSPUcNCXkvJ/QMEPyz9y1/5eT+d4/1oHUc3H4LJzI
Av6IK1rrTSy5QSdBAQ9XhmmCmv2dGvskb2NKnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`protect data_block
3BEC1WGFwO/8r3XdObluV28H+D2bD9qs2ANRNhPzFY5JXVp2KJmRu3Tu1WtqR1AxMl8Wpi8/sPk4
5hs0rHPpGs7wFqkRaOokHgIf5M44/EmA6DhcvnUo9dHzP3gE4S9WXXagHixa0481w0Y+wY3xTN8N
2KQEmAumieDZDgzb9X5+pVp2uxvPAw/lsgJ7pLmNiwfPln1cC0TogDkunpTez39bVxxuoRIfOohe
cBWAD1ON6MtFk5tazXvRHUARMU6/hQxB3Wm9oCRQ6GC8At5GQyg2PN1Baf28gj5cPzq/+k/cqEy8
//cVo80/a2Zc4W1R0XWadg0OO9xmceQZP+HM4NWDFWqMuZJuvMeXvXaQZw7KEGG+ixgrb/wCRrx0
aZUhv9BRFzIxYVYsWEvq0hZFNXw8c32qR5ZcX/3jTH3jVAwSZOyohSbubDiKa5ApiCgipKQpbr0X
kt7odNfnUkYimkQ/hoZ9EuKL+q4uj4/TQ5F1VCD58rABjpiJ1uE18XCYeNJ9dE4+DLVah35MZwZ7
VynycKVsa7pctKW46itVzeP+rsKVC/cchxUCFTtAn8ELjV3I+85VHGClTEJmJin7UF6LltbDwCAH
d5iksmDvqVdcJaFdfr3/dh9pd3UGOdt4LXm7SOE0cINByA3Kswd96e3ntISCk9VKDLrekFQ4zM3b
WwgQkLlzlg13jTGWFoOKIZuJ8YhD8WkVS7tp30mEIx1xRWp4gGYvnBdmSpjOpnWsRxfRWfex2ey4
1ISEEN2gu21nK7MHKcnV9mmGBhbo+iwaW46rjY0kMXo7xONuqcEX356aTA3JSmtocTZ2Aw7qMxGB
g2vxPhFsuhEIARNMZMl528Fo3OWcQdcnT+Tdnr7q4n5tIc+gV3Q+DWZ9yxo1eFTdBtTqzYsN80Gw
MDKrpZZeHpco54tHUv1E7WU+c1GySXmnilxez0HgVqSfY+I5RBkLUe6T0WPzezD+PwyCXcVl1snS
CRmNUj1WKy2WQH0mgB2tlXbbJekSDH32FS7KkhdBUx4c2c3SNMvJuVffbTlresf+RMkNd7g1yI/a
GTYDvP1+40ko5Hr8zJsGfC1eYID43CT0zfirFQdwBarySJseXcauPX+rKX0TdRvgSw+KnAk+9bnO
311HQQYx0rnI97mzikW8rQxmqeV9HtxyE+zRREtHY2gzEXhgOw5hxb3PIwDKAfeX5OUQ6cIYl6i8
kEnH/CPi4kUA5dDCdpeaDqzAINaOcEcTagDmUCGfdKCmTPaTP5GxU/DfHLnEuUbNMJUd4m1TK+VX
ZS5lo25gEn57kWgWk68hqGJEA6UuOkV8zr4F4dHTuM8J8bD6b+fWD2MjY5ZLT+/eZHQzJ8wLvnX8
1HbGSdsOyCcivQ5VnPmBXDSMP/xkW8yo+uGLkhfqP6thIQzL15DEfFsA1qvJA4+NjnXH5INO9rQD
8C32XiQ8T3DJ3Q4FTOkg5g5GdFf5x4vUI6t5ylqVdRje88Q+IQl2j+Bc83Rd+hc4hELQWpE+LOPF
w4XQQV/7o7X+uRwCMpzQqqrLGitEOGR1ULEHvJsZG5giNExWSaDp2YFNj8qZ2UjmJ+vgwX6sOfYP
TmRQVMsc4p0K/HpspGcyn196BvFECtsmaxuPYgOfyS0/juiXTmh7slJasUPUM0lcnUgUOxVBrFwa
adUk52JiD+vMOIxNd7DYe8SUnwnRvVy8PasmHcI70gpeHTQap24UZJr3DWJzSrWtWTJRGcbmgojk
503gndggZi1TLFHf/RaR1RLxLdlGmblWWyL+y8J5zJzAYDUCjVgG+JGk07X8qhbgIGe7BXIMA7c5
ppPK4CeQg9bstXsUN12ErC1bt4VJXwiTV4DsbHjducCpiZYUk2egtG3JHg88+q39822i8wHz1ioe
VnNQUNVp1GzjFTgX9g3TKFFv1EQHoiprVs1/g1K7wR3RfK01Wd705SAoz+iiIb/+NHKMHH2JXBIF
IJwL0thJP0wJQmjU5dK9p1NyvDq8s7I4h8A63P3cBj64nQGsRwZ30hMJpElVwSVMvW+wsxWfMwLB
IbkNbeF0EtCOX4Vc3xpELbM8Dtj4XGI3srh8Pc0TxY53azGuQR0gancfMQkAwhV3J8smZyyVuEyX
BU+ygpNp5+IDKAiTjfCgmN8htceBKW8usG03OfbReyiNJIUylj2b/K77vSCcoj5QF94h4t+wJ/Hn
huI7NChuBKwIGlN8oL4FxuHqg1xG23M/X7EL46d4Za7VAAhuSPe8B0+7oDHCPLLsDOHaittGpee7
ZXoZ2et1SqosSSNr+6StHh3TCEgsttahhMYl9YpH+IsWPoTwC1p3ctwz1jmV+pDPCqYeDCgqb5tN
kF3p3CniupzuVffbbDUbZXmIl0LZty1zqvh+tIcKghX9EHoBc1/7EPreP3KLj5JxlLW4jAriZ+Oj
S+t0PSp64yRzhZqECjL8SLti44lBE0SQLnXmJdS3u8d54e5gsrNOAHch7kE/HhyuJ8gaN+42sIJH
N8jvWpgnTRSaGQoAnrgHX+S6ONTLOKlgo84H9cDwUbS+eo3a/F0Bwz7pZe6C0lHV9bbjhXOXOveJ
c/r8ioL+PJYyabegMUYRAiu/YOrJSHpf+Owj4XMHoQBhJ413e6UlBu0baZ2CgVacy5T7y6goZt/e
C6a1NXQGR+mGBJYU9EncFFVi9/9lsMlhvdOO5r+9TX6hv2bVdUkc5PS/u/O3Ps19OXU2LRRzbkTf
7CuKX6IZVzWwWLMaMFt9x2IjCHaMcpwj02PZ8mWipa6c5priTyNEPW/Lbe46wOSehxA6yZMTDYUv
drRvaeqZXc/+65x5lCBEcnVVKO5GRIf8Kda0KsO8HxJ01B8GvZsbw8DZhvrURQMGCPseIVZjML3s
rBujlJye4NGRtzKAVuu03pojXnmcxYBjdL8sLfASgi0pzP+Y9SHir1QgvVdCy1+pWivLX9LsdBm2
epwzsRtf04lgeKxtNNGkLgnidwS+6N9qW3cDKE0qHnsbJh3vy2OWaL5FYE49ZN9bALAqUtVUnfkM
iLLWi4LGa1975/HnKmZ+kZ9RyqUJh1HvrqtIwZ54JSBe9rQJGLwK+R4DQby2si7z6UEPe284sl6A
tAKURvIeYzuqSiIxsWy2ZV3uS5vyJmzO7riGuwUsqYoHQgMzd/TQm/QD7tL9Ky7vitbhxqU1Xlmn
Vy8VPJ4A0dhG7QN/9SIs/YdGHqvFBueIgLQ5pVicG6muaK/RUh3Mlk9298x2uICP9S4TcvWcDJ96
YAqeT4BsXApto5D44YFJWiNIHoUm6/kk8RYAm3zqbuaG1YYee3yD9IAJmSoRND+8LUQz0LbFVgCH
nn1imCw7OfuiIvYXehABOljqcuCVwtiQ74fBgywgiO4DpEdqAfThpVQJSH71D9wh9vKaS8kki0on
ztT07JYgWudCvNpLxEbaP9W0aM4ipsqsffMekOiLIi0gbDXRwZTMwAGTcyWjVsbV7/Rq4Al9NtFz
Nj1WLAegQDjCXtt8+vquD7EhrPvZb608U8k9LzMydghsRmpAE31r78XzcJjHjWOoiEmmgHgKomCU
YUNMq3M/Mc4myo7oncMwG0kTzf7GPl0GVJRgJXS2pOzF/oJUX/nyBg95+/oS2q8hWH+O7N5PJttx
sNVrfWrwY1plBMItHIm0rdy6m0yvEEmxQtdwUCFXGq9foXk4Z0o/mf94ifLy06FrR5/4V0guwLCY
fQPrrVxy2pVCK56e8qAy8zcXlxZboNlt2k7m0K1rsay3Rw/TNdAAIaTiIF9I5o9yc1tkeEmbSEPm
ZUPMcgezgzZc/ZpzeKh5nRZHbLtPq6UpVryFMh1irYsqybZiif/8EEvddSdB3HOiudU//Hb3+Aof
PZjiaez6yXXJCSA5dwCYLbo2um5B9qynsbA+kfNyrRt735Q2/16845TePFmiyIwVixVeebV96muO
CDPg6EmDtAmY1JmCtj6MQ4yoPoMMxD6QOypJzGguL3GlaszY511ROSTy1GfCR0h7PSlGefYl2Fwi
jWgfMzKtx43EpP/YY/N2HymNRuA/Iy/SJwLkb9SGvmjSRdK8Ud0qfb6TcU4MbIbb9TzenDj+ijDY
kGoWdxzMom+IMOw1Pkp74oJrT1094xTauhk4xE5S2MPVI4mnCNvev1Wqi0yD0JpwFdWAa1UIHQMw
W4O6FrxqFVlkcJOmt0IeT8HCXg4IZL9YOpCYhpLg4akeUAI14lyD+CBwQk4weFPFaMXxBvTLwUQK
tEPfKjxrwOl8W55VhT5z44+gwxZdD0Mesu6OlGsptTYzYNPnibMQWbNg+vm2/JsBqwLwmZSf1MT/
4NFr0dqTmooh9Kc0D7Hg0Pwp1blfV80hCGFG+C/7NB0qKdiQVqEuOCmGtqQtcCHds1+5DqurP2NJ
eCJgxcJPQr5hGVDP/7xFh5cLbd4WmsYhSz+hUdUB9Ql6bVK+q3boevjh1h21YZVSHNAKORuT6ogT
ShGG90ErDarcgpuuouRU/ppAUR7eG/H3tuKkCbkzCUJTqmtq6JamH7Q5VnvoC2/OP4DoaXM7rK76
JDbZYi0GowCU2M0J3J6dDyoFK1fvWsj0zMMipFx3e57pg/+X4nrQCRF9xh3hgWynewriurfsMoEc
1DaeOs0i8AYQ8682/0msf/gHMwWxgXLnkWP7OAKcFjA/U6b20ALa5fqIdVChYuuIg9gtAQjAvGVe
jHVf4oNcCwi3i6bzh1FNzvJFn41F0QDUVFTRmKU9W5lLJh4tiprDW4JRcWKYJ6tS0rOzGIlQs/3J
+z9uYWSB8lRobT1U9DyCrqUN1lI6LBqUpT9SDDVs5p2UZlU0xWZ6FmZ/SFXv+v1eCFnj+Z1t4rFN
7IF7yCuG/2gqBxPzWmDHYkTLAGgrUrwg/VbSq8iKVlTXCCippQ/qmYnzWfZo42IZRHWVkkugQ3/x
373RW5Las1/YGXk4N4SsKYcXQ8WkEezSurOHHjo5s/6RPVWnFeW2a/0pAsDPtAWW/4mt9cxiQR6J
BpglxRi4JKlnfVE1KXsYilGbhxJjoowin8gZSrb4eBHHp/7/1kzVF6VgpmiksksoCcVQF4nICb/q
hA8zeq7+zw0n20iG9qsrmfoiB0GkC2luVCP2tswIv3Of7q2WP8QVpDHove/jYcB5UoqetZt8n2vE
/c7Cyx/oFDwJOhVQiWiC7aNArtszIWdsPIRicO2MlGFUw3OsVFBFj16rHZTM6aNUBpCS1ALu7DI3
JapddQdg6HrmlKNawjQnFr6pQVKLdQyvu4x1wWurMflESk2tQszk8j/8eRwHy0PfJUrGhTDnDS7J
GFIof9uOky1Sf4BEiWubqiftLOE0AgIEjG05b9scbuiWXZ8x2iQ5CXJFxwWQiNvCYalsfK2vhLze
DgBx3RexhF+/ysYq80hct4a0G1OlmZPW9C0QsULo3wPcy5s8640XC1WpmR3etg1qlphpTWPeR8fl
tuFKJGb1vRPtzphiifw4zL46Wo9AdSIZ1tEPuQdS56PbTeUidz/QqZNworxNHVLuEV1dZfxBE1oC
4epV7E1I/ftowE8tcVw9aAuuAYHjngGmGt5Up9AS2JduMvTOfL1Dr6tFy6ZJ6sMGICF3AsXND7+D
Xnsh8pn8gIKnJZqp/rrHTOAmVR8G3SlckSYiXTkyY4kS7HAPv2/eBuEGF82R9SU2oeXCgJVABs6u
6fMFXtnRM70lZqQCkdHaVlY+Dwlfc1hf4Qy6lNUij/cHKjjwFkp8Oygy5j+FnU8E3SRdUC/4wrWG
6hoqf+DffJ0eM1o70AprZRKORRyo7GsGt2q6zrA8d4qDlHFvtsr/Y1d4XFFBRN4mWx2pfNeh3I0j
spNJIYmz8nyG9VnkAiGONayGIOKdEK5zPbOVdb7fTPFyNeaVyUkn1ubgBk3/XElUUQdlcYPRDSUS
pGnOlJQoT5onPEbOP6Zbra/sYlWWFpW/5gOOrm7CcAWDHzK7yLCXhZugqrEs06WMgaIy6TGsUZPh
jklT1oNOG5JmRPF1cO7mvECK2pL2mkJ60n+0MENiVblFnrJpfkJnwn0qQPV+PFy7Nore4NuGY42P
gINSdmcGEgh24EhAm7PdtHtLo+EodfS268TSpvaZwsiHktT5d/QrlW/RsV2wucnhG//tFc1HA5sz
JkAIWuTSKXaC+3vfyoTAnQchTeaCoCVXTz7lqm5iiiL1zPS/LUjdxx8UXuJZhakhABYgd2ZgAap9
YWFJBGuvpB5sYPPPCImQn5uPbKTHDNxnPlFel6OTvM5aTr7HJAGNKVfm5W6w1NMOZ1DviUhoRjfi
PZJ1YzGVIOBTu0hr6qkrcem3lpxzvoEeIkmubzS6dofWU6Rbex/p+CB5Vrk1VQC2+U4yb7EptvAD
sC3gsIlELVYgdwppn94qfLK3DVP3OazM+yavDPCBkpJ0pPyCGO38HSxSPj/ZrJD96SHklyBc1NVP
DrjlzPS1R2nll8kMUZL4566dNOpkJrD4/UsIzzULCRcCO17kGbPpAOwl9Abb1nWrTxUneHeFv0Ur
e5LIkIXTwmOUBB6y5jNhQpa2D0p3heU89M6oDe9wXwczhw2kUdYK5GKhheeBaZkjJZL33iyVHinN
J+k50+2v2EMFQd47MBWQPvCEcOEL+66wYaU1/zjk/i0B4KdnDUaDJQYzBszhXW9FkG6b4AAc2Vt1
7wMgcKzMdlbRE2O1wdsZ5NoftOcVsPN6Ub34Ut4+0HjfWGHJ9WLpQhNjnJRdZKgTn1WIvGwMY7w6
KfQW4tDVo63xJQgRZDOdcRthZ4MMaaV5CiyMN0G3fe1j29EUV+cnHa1nKHhnTDozyFLgNVF8nPB4
efezZKoYkbL45zalOhTsfv4V3VYBia0u2v3diuTSe6vPvaXhp3QeZQwEnpDJUNjqzDOuNhTxrj0d
Nf2LEz2e+tazd72ni+vMVXMDz2JGpd6QOw25EcyFf/H5hpZvNrxvt7S8L7BmNWsWPHC0786cyNin
R3wJPuY59OTQMrHgyeb0TrTrJ/S1KWLWmp4F0SAS9mxOy34HVt9KKxyIN07GmwswSH8Hn7Qz+zKk
fFmKmtDdeAJBHtxXmQROxm5bnZh2N75K5g13nifLuVs94xBHMFg1P4Nd9w8TvOz9NArK1aqupmU4
LW4lVCKb0LRzGAPzh9gwi+4HRrBzor1MNGpV8RbJzHS2h3D1ApqgmG685T5oPTQAZj2r2b97gm/h
yES5t3frRM/RbFUDb4o+X3FMCPdxpOv0FDVd3m/bxDgtMJhAZTuD7A2ClhvivaMWV5uKEkHQyFNn
n9mVR8yWhGtkwtdzNA9XK7bdetcXkg7MoZ8ccDHqQZKqGW2dSrrSw1T372AGZe9s5zzT+ON/wnTQ
YL6ejbCzdrW3cUfEvJkkuZ306mByLspn6a4EA08zfjY3KB3XYV0K8NmSra+mHYp62kNO/czHtAPJ
qGGuUt8pMQyO+yTcvUavbjkYt+WNcPyHdQn7x/ycG1S6RsaW1B9mZ4vsaKO6WX3fOaTlwkFlEtVh
tJgAGgWDAFodDlAt+ejKMve2eKGA4vidCToPTP1feD5LF/DInswAyY2bImJOSVgZJGJ5cZtEzlgI
/y+LSQmOiyzILPiqv3esnSE1cZV5fpJjRxNYuP/CLHg/ArUwanlkTIXhEH3CoWXKhhc2mkPSUB5t
XYlXZ3UDSoNyNDti2PoHDOaLNOzFwTiMDsB1HaEOMqKC5mQ+DOrvWMDFgEO8+EutJykj8m7h0ni4
8QsvDhjwo4h0dw==
`protect end_protected
