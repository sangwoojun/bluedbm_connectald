`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
lpxzCh8oh6z8liD+PlJK2jR/wrfrCQjZwTuk/GDi2FBTcWnBuMt1bG/PWWbt0LUtK7p3GTKbQdOy
W3TaAaUjaQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G28AvPC/fi9ig1WH+Cm52NPcfgfqLUHlJyb98SpHA0ZgGDuPDpwTpawBjCl04NeMz/VjLjqF3eEc
1We607cvMurzaIUv2PsscX49Su+smdjUJftFSqCcCcSDKsuJFKxzxK1a7vT+n8l0VX0opmrThRYX
rP6uMZMixF+EJlui97I=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VxW4dfToEN5cq6lISW4Yh74zQ3AKh6yFW0bvAB5APDCfTgnfApshgoJq7QoO4cVUIwhYJ39Bntjc
A3yFcjPaSvsYvHu2mRu0Xb4K3B7n2Zmi+dLGu+YCygWfG0almLNK+iyEdtR33iOmufvDuw/rzpTh
Ycn4vzbCVvvXLDMGTF+5ATnOWUJxp47dwQbSqzHsfLvG1copclgL++a+5kyoeX7R/bWHClXYhm65
KMvhddNN2S1a/dyCPwQPVRKR3ZriLvlau/P9N0fKFVbGhg418PMnouJ/9FqV2UVxCqLh71jEG5Im
8MuL8Lfae21plimd8lUjcuHylwLdi8W/j40lbw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KTxSQQOCOy1g/CMzQ1VhmHLMU37MauEVWWWFJeCk1U4RYKVobc/3BNnW7UsAvgg2EM3gW9N2aSxz
O1wBUFmC4mdHhIr6MOobVZEQr5YcwUl2wkjy/lJPDHyxITe2/AS8BvtEqcc6HDqhW5r/0x7X0LoJ
OufH4R60MeE9PAP/W38=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
S4ffMg8+ru9k+LStiieah3VYPx2FiuWFVDgDs8+yvUNDGu0ZknB3jaGy0cLmnDsgCoT1Qq52PPSa
MT+8C88hIhPam7zh2RrD4XT/Mu7sduv+zr1nAUNRsYTFw/iMxswdQ6v7yBi4mQr1FaQt38PD1QI+
v5LQLXwQghVlsGsK65rY8f5g49xUPvGSTXTM0leeALZIIj/vgzjf8Ctph2ns5q1dkdVJXRWuG3V6
7+GOcxymAPdEe1TUNUMXI4MWXQdWgC8h/nxz52DpUC5g79hnWbNe4gZbMZj8d8Lygnk/nUDu52QO
IbW3lkXJxkKGjdpBc8MyHRYagHPksB+mHDmsUw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13296)
`protect data_block
RQ1baw/dXRd9j5dJH6LV7CMSsATEXvFDyB3cgi47Um6qVjz1QUpo304IIQsIHUTiu3accEowqQ89
Y7RSvKYxuiaQTbV9mlUGKcfxpwwBTX0GSBY61wr69cSO3PFnHKMofmidUKpLscLCsm07gjtEkqr3
lnZskk8E/jE13mDP67qWIKiexDQRFSk6TF2p9nzVgNxN2TOHJaBVnULXC/5wmxccHGtDSuRjuygG
hxcrVRVpuFamj25eo6jIxsXu5A2Gt5uF87NdWQP84WleDiBNA1J1T/j3rT9+xEOc/pXCYR19MvAH
6I2YNrSfE2b6q1fwBEOMIfK0SeYOAuLt+KZhD3HQRjyH5PEXIpJBj+p/grIJxh3S4e1bpjtBBS8x
oV/BuzL2bbKhRl8t3/iOpLIAEWLJVAh6mebk4cnY59gxgSOsNBAIDHaghjdWfalNKnI4grh0/jXe
pL6epTqwwFLJPlVGfnmQOLiyCBlCTsy0pNOCIOrzaicVA5ztPijCMKpAgnuh1EpoMTkcHdy6xXb2
Lj8iwE4yzb8P8nl+/ZAR0zDFVb0FFI2UrKPWFpCUPFLHtWnJNpfqilR3l32aWFYfHIg3l/uLOyIH
pCqRlDAPDPjAae9m10LdCzP5Ov/KPHOsxJrY5lwYNQJDSNor0o+5y/A6uIPX/hBw2um1ZiAMr6Ts
vtxwQ8k7CRUSTqLKriOKNx6SJaKurqiotz2zR5VoBlUlaRAv3gDHvUL9DrcakKSa0oRiMlGxaFmN
KLFeL8FMBJfzYZpEFat7tX/LuYDwBwSW4pvV8QClIv0ox4FgzwVo0UJVFDAKSyL48HGGy4Lyq7Cg
A4DRWS8imUpGlUjDfWucfA2xOxJF96Iu2Dp0ekALzkqiaJuOI7qh0oDkXPYVQeRjt1pkulmVZuSQ
cOCEr9kvVtIUhEPZj4lk4oaNyYRz/IMOiLPuqC4wiWZGhVGBa9dBmJQkIZ/jIY0LNZmuDwMcQwtK
IERHD13xnJhiSi0o9qLPJ8xWNcBsdpK03LTEVNE74smDv0AWKrJdFDoJLYBETLsy5LPGvhltjdaA
sgitPaZVpfosq6ytQBK0Gc7c2h9hpRqzMHHE50dov9r1Msth/49ljxoTu2qAlS48nfIFPkwzmKI/
pH01v/SD5quZD2Z3L8sfYpEIA/DTo11qSqehhtNh990z4H4o7QWBtfBjdM8k2e3HeFBpJgi3OFhS
Qgw3TtFReESLCOE/ocyzGHU8iegVt4MJxD0VErD9MorjE6BWVRjXBxmznjTH180RdcJt6XGCIUde
vBw3pCrPps5CZ7JmLkslIO9CkKu/1MNVRjtuECwYbuIO8a97gv5sAeZkODXYEsyMYj6aW4xGwH7e
ST08LDMZ2koGvivoFj9RQ0LzfaY5a2gbaHc7iLBBN5iukTOqS5a3EUPqOZIbcIRP6OEF06Ttv4f8
BFhFQKVWwBzbZRVGIx+ms4juM0SJF0iO47fnETYExR+3T+/OOhnvRu7yNsROgo3z+CVHarM1b9We
mM5LFdhxKDDBi+bzjEoIwmI/US4jaVlTcYncU5rbFzh+fpLMk8NRmXHObeXB9l458GdQmfzW/GvX
3UFN6wFi2UpRh1IF7G/hVwsp2YGvJh1KfvwudYNwktjLhhmpWbZv0VahSyn2pnB+0NuwadOcZKso
N52FKrXIhHX+ngZ4K/GvmiJ/FkEpMwD879WxbiIXAkVwCn8exnirYSs2CN3g7PhG/+YEe4tywVhI
De2L5Y/V1Sa1bWWluauk5iJFaNQIWmejmlrgN6T8u23cc3y40+hTmyIxjgQpq7mWEU+MEUhnmOJc
T4UUCfFRfUbc3kW7LeW+GcoXAQCGn6xWoOvCxG9GGl85xS6gkgqiNI8AA4pVl/UtxNqNl2P89aGG
qy06dAzM52p5YAVFzaiC8A78xNxTvn5+xrfFq6dtHTspAnJeTzEt9X48shuIZz/+b9fOYdpLSpxo
JbhH8M/0HT2wyFWfsrGqoXnkIf9ZbsakblqYlU3qYHQH/cb6P+FJ2GN1pBOYlkqERwUlRaPaMVVL
2DIkRIbHQCZpix6vYJIo4ssuvS+uKPQWY3jTv6k9NjnBtUik3eXASJ3KjlS75OGUz6VHV1Dw2+IG
coO8uB1U5UfD4HtCCjVl0xcdnWIgkt/PNmiX3JUi+UEP0DlDwc9VslwcsqbeY4zhjIv3MH5NKWpA
T7sKT//TxmB1CplBCDNJp9rfAx3oLGL3on+ppDxZyK/DkU7t9TjnEUpwJ65NW4ofVnEWJj3l8lSi
mXvL0ZjFEb8xYm/+b7GOjcla5UMNhhR7DGdXrwP7Kh+2LblBc7Y1K482MVfl0L/Xb8nHH9XZKaP7
pjfg/lfBbra2vpBpIx3LW1pRnnHkoyedDaCq4PGS3bL5ZsRQhW43xYyfG3cGPkiJ8du44mbwkrpK
/MrHz/h0z7AAW6NiL12g7H9Y+xqLcBfLAlENAgAbrP6mT3e1r1i4Yeykxb75zrYY4CxtsdEgDMkM
FBegtEjvw/QiLFlfmk3Wn51aXnOQOYqbqwB4XPDamv1Eut/0SnJR5Q7YUYrHP970VuLfaZjhe26I
F/gwaWHRrAr+ZBgJMF8C1dajuss8Riv0L987FD2/FSlzuWXZPwjPrnMo5yv17u/aHrIqwMvAPHlV
mK2WWfTHe2OW/y2dbKs8Nl5xjjKozr9gky/lCHPRnr8+wktNnrXT6uF6rgH7bCb39oExza/191vq
Sxn7VChyX7tJ3uoFfNHTUo/uWl5Ud8Q2kNUS2+Bs/tLoIEQ2r+o7vuPVeEuhosEzyM4DdXrgVzTv
gBd6lOkCacrxNPlQWiprljyr4ngM3zaDqtjsogfmWCysVSHd4fhTTxxHoS+qb68LJ5mw5zYm39Rk
ZUKaQ1gRqYOWaWJqfdTdVdoV2S9cvxP0tDL/SxMShTtVdPBWiLzv6ws+euoG5Q71R0DS3Taxsj3v
MENV9SeVfBH0/maZQjeQm4qp4P2jqXYgtxpV/68no4HBf5ZKnHiftmXwW0u3068J+mp//cHPcusS
1aGhNGbdLX+8b8zenlZlEjVeLHoMRAIjZNJpStg2tC0S79qYhp4tE+FkpH50CKd4U/U/7SZT8xXy
48QJfZMvb1Gk4VNTHLgLRtcph9pJ/YYhjYmyJhOPqoFaRZTGbLiwOIpTBczZz+EpMxzucx95N01e
SlRoh1JnQrTkT543ZOsFGraU0T7noqS18gYQcy3/jYwDVXnQrJrotYIpT77tvFU4xhFBUs9TeZUi
q66W+5YTY8lmpY/TRS1z8CKuRchnYci9+gla5AAWVwFO62uUsgZQehYiRvsvJaYqM+t5+p6PW3zg
HRT1TDMFLK1NU91ezKBYButRbiT8/5r2yT1pENUIxi/bVRBnuNlmsq5XR+ufOj9VnqCa6I7ZLtkd
2CtKBmIS2RpUKkBqrMPD+Bd1B3uLKymsx1TTok66nACYLH38zkaTdtAAiKmbeehb5zUUtUgu3eKx
URv7qxMrl6AveLXM9yBbBu1pqPBssJ/CUdK65dKd4uXC56IqS4E4tmwm6WUWUmHUnFk1W1GExYCU
3zvCuB1UOlvzxsJzY6kuEr7AvVY8FSVosnVRYokWdPotxr9BFJsp/VW5UEaHQ7XenKZtS+U84I50
mtyJTerSPW+Mweas9TbM+DVXV+gr8RoxbhqM9GZRars4PnOV2DVYiMyh+YLdIu+5d6odE7nvfOQi
FyIl5ALqODhahI2mKKz7pVxJgLoWyJadYiXxhRRCXFNEzJDui6fy3w3mWYEaFVaZ4eGs2B3XQONs
enKPJ3kq6bsqho5zcsxIgmpO005gO4tKdec1HC1UZarnc2P8CtGLBwp30B3h4MTANI19B3mZzi1K
8my5m05dTHcusId62R8OUxmP6tQa97vWeF7kN8jX0M48aqDheHd01NP+ZoAHeTCZeE0QTrjO7dQb
fIetr4+qOGYnSc3ZThrCo/BxkZpeQzj/uuux8KuiKVsKmBLFsu69ZgHtZz8VsDlcGd6Kdd0QQGf4
iljg+AhJKy0Z5lpwdaWGjXapFrHxQU/FsjfY2qeeoZa4M0Z6hd+BUz4CvelT1sOTTR9z/ACCTsiO
V1NkhEPMCeSEiw6EuEEHLnE5gnqvFBhJkFMJvtMF83+zlS1ko1OzkbSOjRFbz2Xlet68oFKJQ8il
+8KPXaCLr4rTjM6kM7kk0YuHIrYiFmLFUPq6Yjpjv1X9plJFr9qzm7YQ8QNW2Boi+cXGO8ZQtFR5
Q5MtUneGuCAPhw2g+BkaDitOMyg6kU9KhH2E3Ab4DQNXcL9fagZ7/L1TEdkyiVIhCIO2aKCgAU+P
+H9ARlHEOK3ZYrRbSkbbHhARqF3L7qgaXTTwhhFP1jFaPMoUXGTX/SBLHEgrxQMTCJn8avALTsqq
Pz3D8KP9/QutNnZxBHpASxjDrCPxOmMtPfPmM2ua86VbXb46LexaIXcCAhh475Ve37iXxNveWZ2E
u0VYzpnNEgVaT7M2saMhYXemh7H4ZNZ/TOse+cTvDeGMOPrAhViap1m/TxhS1CBTL53Wxob5r0Nk
WEdgpjRkm7PmYZ5q1AzilWzQnDut2r138wDmAkBEcK9PklU4vDL3LaDYnUT6i3Ngu2pAIyPlbIjA
rgon17q7boVsvauQpu0Urb/CC/rAp/SKnNE27tte5J0lnfon2jtwZwHSsKUpSB9Ary/418jVbLvQ
aeET+SQ++zAbhAZ97slkqL2J47hJvmZbhfNIUePFv9UXwEJkjOHM4JFCf7jh7cbcNlpbRC8uuvLP
FADpyCSAznEqkQBT91d14kB+rZzNIJ0HuNKsKqgXCqSwRqOSuryclhDXha0CqruKdIxjCC/tr8UQ
XFwV9y9D9Bt1e8Pcy5hKxEK+g5RFFExVUaPiwdh3j209XHNsX5iocSeFPs6clodY091QsHH7If2Q
PvK8DeE4Ra3BGoDWbfBCdSWzIKBjvlo7wkiUBjTUl0KVWPitL7pNCzxyJJoDOP9y2lOOiUpogr9u
jqXlqO371JfakOT/adVBpM6kgoG81iZSxM99Ldo8080L+0H0D/DrCI2B3oMURmnWHbr5TuysJHDy
akIeAhC8d0qGC+Z9CRi0Y83zELJlDWF+rkUyrDlVbTFZ/cGEj51gkCyHWUYpbQ75gj+kflYas0Xm
G2iITB9gMWoc4tgly7xs5gCkKLUChaQ+4V7OhO0q5GZIa1fePffjx67ng50zS8P0Hvy0IMcYH3Ys
SprnZgGuSByHmxD6ey8G/XVURJ1VUPn0sVLQ31kiVamES5LDSNzxjApHkbJCssgynTOfmzkNG8r5
XEkam64tukbM/Dx+mCdmO1Qkvi2zrhXHTp0Ln/cENUAbRkhAGqTzNMGLqFg1rJhlCwy/NJO0bBJj
E+obv3V7IhBzavFz/pnkTy+sRDWP2ILVA5X1+Tp+rzhl+Jxfd8lxGZnyvqQ2FcHfieNLBatTsIij
IyfmuVTLM7kDAQyNv76odgRJZdHTgY/n1bdh9JieYrksJTmZHKF0+Yl6+aByiTAUCYcBAfdQQ07J
Kepe1Jqs85tlarNEOsTNVRCy2QqSlZoJ9JYBrgurBOmV0i7XOjKlFZ/PaRmvFem7gd1msW/78oj+
3Zr2GeYt7/k3SWHgVT4a4yeAIett4HQdu0ALKKaJaHtNuoL9vO+MuvN1UpAm3I5vlpCJP9ioPnDa
Fj2bOZN705aSzwgTqkGCtuRupxBEwLQTGXedSQ6yIoHS37Al5JAH3rxIlGQak78aSzhfsXbDGX/k
pL+DYOs+32RRUxh9vcZ2fzWftD20F0PCLc0vW4sEjcO6Rqrk+bkFn+kjk7lpS3CT+eiH/MOdHWTm
usMPv/4vBthJXH5Po11US8eZlxfl4TP7GpiKtEtpAduCZorh/D8Le+c2KJfj1YyPMpBi5Gz/GyYj
Ir2tyVudTNQhUYnWgoi1VzciWqIZSXd22JOZp1xv9KbeLcHveCvoY9HtpLXeC0e7zd6WLzW0X9Eq
G/5yBITul7yrUC8u7dqlE/iN/IkjKMcC4jCaBMSY1FlVtGpHIqUfgVubdn14tNc5F6ltZ17uA+7m
wvipmdAOkTLZnZNSBxpTfJbqFBuyLoSU6iEGNrk94RAL/kON5A3SUrcDSvibQb29VNqXFbs3ZNVQ
7QzOicRERpW5mtiqdgovnpfncm16ACQPSOrPlyUsc1I+H46E35lkruQJMwcdSk4ic9YA5EhKkoIM
IE4CcbjxNw9Ror/WET7tybsIsrmQ988kuYvQX6XUFMISZI3RLj5Cf5gPQ8cBSNDAlO7lhUZVrYCR
HAC8rg8ktOtvn1Fj4rFCimORB2h+YuGUSAqm8W2lADos7PFBsQ5pvclttfiMslPHtv8Go+KxOJFy
vBNpZ16PCrdUEcFTPmAs6pQHFWTU95aiz2JrR8/aR81eIxUZsprpKhzhdu+kBiPYnqI1+Merzxnq
ZInls4F9t3EO7FgXbWvpZXD3Wt75Pkrb1FhTNohfQL5YevfI4k5unaKa3pl858iiSkBxEfyEDiE2
O32ssg7Nj7cxMLqpmvdHZ9Rx8IKHiKND7qQfYMTL+mi0V8jBYa841X2FY29xVch5akRV6mFoMoZo
4JRPtwui0G6XZFxFL5oB5KfmIZnQdU0MsWnP/jfVgK5hXfH0VcHGUTBhxN25bhcZcRilcGRHWg2D
b/Rmx1MuOs4xqZiwgaqphb4/dZ4Njy756NS01SWXOAoDEM+UXpd60XGNBSJk1LXWI5YZBnNYAwWU
bPBkJL3gpet8mxzfyt2AXqtsqnmkYHVtYl4PhYjQoH2z4XMT5dVQ4dD9OoJ+xpGfzpIppevDT5WB
71IOMv00dA4UbpZS+TJb7D2lRMdsPMiZIBvFftkhy+3rHHJsHA4i99z+mjDyxcoy6g8mXWRoDUiN
Bkm5bfLeAh2+WuEV5ts0T1A5UT4Y5tF1NN6Q6lbWA2cv3HHhR/rtRdlg6WkVgYSIkCey/NxLGaWT
hVI/GDw9cVOAXsMe7SVwHjadvthfgRc8cBaFW9ngZQRWrEZpmjkPVCrw4rj/GfX3a+QQUECRARpz
4o47xWGJ3PA4eobDI+CGUJ7+40mePYco6zRMNMbBjNt3Stb0NWu8noIklyAyeK/eefqh6LKjTKeG
qET3dHDwE2xNIfpupnMs1RvHX+UIn9t9rWcCtK3Xtr0uiJLI9ESoHtKkZlqFufEYUoSzSPSiKwWM
asleiSJAK13aofLXErNbij39m8iaPcGnkcFudXUKZAHZI57kCoIPA75vAeM29hxoQ6evdfJi2PXT
HTX1o2NbfiaAZKxbyZxVUwB89WkPaC8SvvR1TO6L5a8yBTbIDwnMz8NsDTlKYin4PSkZzMy8SkQk
tRwHjlcCa9BTY6iQ6JGpOofGD/dNeYGIgNcx0rXnA7srSqGchc0ajAsmm+yz0A66Buvnd2fMZ87x
bFc+zhT6RcZlXCZjJiN5JK4bOXzhYsomQyIJbjJvi/fAEdRC/zIkL0yc9jIggxVyAgyO8cmXgroN
w8960EKnwqGscPwzadhlgc4hQhDdJlUyuOTTWZ1fQ9jw/jV8M9tiCbUosXo3lf2eJKNZhxwSiYje
jr4W7rZlm9y0K7CzGPa+IJz3v7J7bJZ2sCxUPaW5BNkl2WLLOuCIqYG17es4akSfuar94ssUEFXf
d6pm97w1TtU/gA4UPiSuwb1r8NPHVEipUtF4m1CDHuuoprkzWAkc4/0cKghFO+OdYEnG1Py3LroF
FDaWKxUacO6mKxhqQZlx4krzM26EaoMvpOHuDQjEJ7pbWASbGmeAdsgkHXuLvyWsrIgU0TjP1ix1
5GH/JFuFcL11ZviI9Kw3P/PbrFUtlY4EAN36HHtcV4/BdKMiGBO6pq7jEbGnUOvELq0YfrSj7TqF
7BU9LzNYUsk0s1t/ARO0DFf9uv3b7riqC6ebzoC/ZVHjeNwUFatKoyE1pLTO7PzSDGj2kIwDU5Ks
NQbXIm276tosHwJL8iF3R2UYm0c0oj51mvzLxWqRPowIuA6cwwRNr3acYF7dtF90cm10CvNgUQui
LD+Z4OUfqHM7l+rnwmfmSjtyuTIK5l/BZP8FmZRr2jrJU7gIClW435rn5+M+KXGn6coFZluKpgQr
WETmCPseQBO0vBMZDkx+oKVD0z4Q41V1y9FIXo5aXLEJOSM2NfMYrlUdQhNMx37AEN+qMOuljIMH
JDJypqnOZekaWZJkVoF9ukJFZIjxpWrsQMvrw/QFMHqCmb2zDyDWISU1X6Ms7AOQAABKo/55gpYl
wNqXi0LbeE5PDTK7rgCEpdq3FmUOsyUXP4naBK06WvWTDmyYXzdGCHJzY708UKvNrbausNaqEpV6
0gNjsBSWp442rPpRUAOA/XD22+qxHt8vhT04hs+xXHsJ6cDn3xJN+kMC2UsV8RqX7K0Jz4tnqT4S
pavU89hqbrzvJ8n1SU07VAoQpy9K2yP2E+3i+9TefrSil0dQDKJ9xwEUydNC2hTxU8rLD3tnPuHp
t/KDDubGdYbdRjArI5IZLVQ2Re4+epBvVW0EFMciyewY4BALGl/MugNf1pfS8O49gZq3bilvHjts
hes2lLp6unha+WDuwrHwCgAPFtrkhv4gJdWFY5LNqaDNK1g9ApC4eqQQZdVDFU5suLYztG0w9005
imWvAs3UZbN5Qins1LVN3BLUJQPBzgbIN30mmGOuzE3BE0PrfEGRZRAp6BLdDrt4P3fAvVwGXQbY
m+uB1QTgHt7w/jsgF7Cg9hC1B6z1U/jZg9nZi5MQpXND49AYTcwpGZNP6dwyVcP+NTtv9MSe1zG+
VanuRw/o4HJyKx0/oUWMWcnCHGAKha1zREf/QuEbSHIM9woew0Emaf6gIQ7VBNabI4JdT7sM+Gr1
Jbc8mXq0FL3GREfxB1/vX6E8I45V/avjPMJn2Ap33eNFOAGrOruq5Q0OdGKYVnF9Cb8JKr88G+st
pCa1Bl+Q6fftmTGHTeGVDi/h/xH20vj3hdoMGXnWyciz+qM+CJBu1XDxbFvDUG481dPl66PI86mj
8crupnzplq1u4efs+KJBozHyiAUzAIhzYdmrC3g267wrGNGtmVbM8D6MRBveo6iKiU5e2eFGXysp
c5F5JTnOyI6O1YmOkgEyL4Hnw4tgldm6FKRcpuRk7y5ANFYlwq4CA0vUW72/lhV70PojDBJyKe6S
spEFZCP8HsCGgNxx1Ahf/8AKuuxxripCKxBFGNzslJjMfWJZ2/PKSv/sCXX3b1H8dNCHktzsrniJ
SkaEHUY6DzvygKWN9VC9vtMeJzRAoo/x5SVA66/G6Z9RRay2hQ8xuaqddP+q2LH7NR9nOY+KkJSo
clcMK5UNjeG7J49INdjx6PoLoG7yfg5WPPwUNlKlSREHH5GTr4DB3ImOkCPQeMpPSFoWhE9B+awr
GzxI2m/IasMo/uo+keAuJsuM9HdzUDtqCUwlguhNlLCwhOhOSqhW1IlvbS1Obn16k2mXjyztnjzr
UFp+qLBUNMOOUG0XkcP+kQZqk1crqcvcJ1QFiIV1GSeyfLq5yALPGHJ6sO1gQRX51n7o4LKc4RkC
eRzUivWuxnQMN723/aIcB7FSWkZnHM1NM3lz0S7AgXnLqhCVJsS0zjkGLBYjHJyw1hTcuj1cfMSP
wiXIV+gcgZFF1PfxZB5k+/oyB9LvkOGeIraF9mrkUPO9QE1NTFrLgLpP9oyqua/BLEAgJJN7MkME
sTUJeAGVz3tnEdRpWbPGhyaswANDEvaC4HdrQWzyU8WidYJIjb7P+v0dL5/1UxVZm7fSbTgWA91N
KfR0QfafbMWmmcpHA+I8kOdGT0vqGupbbQV3Nt/MNCkYdYDtqyiB9gLsXcO8v9h14CQJefMIJ45Z
MRouhToIAnR0bjQRZ+W0YwPlzrRc6EgGX1gzt3fwAIn0LFCx+JYYsekn9BcYAE0JAOH7NQ7UiTmA
+Sn51eNAA31QmKVT30K8LetOD0OSQpLKYt8wq+t5I/tlhrTvwRU8Banlq0w6m8araVpMsVxTcNu7
8Atdol+k46Jh6Usxtut3f48C9qqySnFYxFjwDc8/37WzNjJvl4fvPN3eGPFI14rpe+zF/7MSWnoN
pA6u2XWtrZLLAUlT7kjNi5HSOO1uSk+p8ntzqZLwqQNSk0A4IHMcbOqPVASrgTvQjdozDmd3M3fs
ry8NdgIl5zv3L2wRhJELNWyRYisDeV96nfWt5fHxYAcQyXWzdJZXmkCwhLwxFK1o3DZIhLG9tD1n
vHF9C0AFkG7uBnbKWzDZyJSFGP62URysVEeTFMdHFdZ9WYzBVSZZjI019zn/qxOczC7dgnJQG0QB
R5kRI0rkUQZ6CdnHPKR8bCJzSGUmo4JpXQxZwvdM/dhQaszgYT51TKsT55UovIFBGP4hsuwWXAro
hvQ37NvT8m0+6/pXogXDSU3EfKdXNwgtEP/Q5XpVIWc3V3nSYqqmJKO1+GKAHkODGKZ+Jju4euH9
duj9bDjqJ0yCK669T50C5tCvuW9rQi0FhHzgcEVcq4xxgt3QxkPtEKKVeBdyJJydsxcb9G+OBPDx
kBuBeQHbPYvDFANFM19Nh7pC0r0vc4OjZLeR87a8lgGZ7lz+0SscJw+97N7pY38ssS/9CffhUS3s
ZRGSDAJ3Jm/ckQju+y05Ig6K/+hGYM920KEqELt/W403lomKOg6tQOey+MOSklbYTGmD/83p83hI
2XH6HQzyYO/ssJkBuXq26ZhhcxbeMSCMhT/tFkxSZNPeyGW5NRmIwO3tf6t71gZ9rpptrLfUi81W
La+xVs7dhpHv7p/tBruKkC6P1gmfasJNt3rVk0oK1jZqEXGTVrQYoXFtfSKWVT6RwVxiHKrqtV0k
Qvdy+10wJrr40wIg5XAFy1zy1NFkyhf1/IR/4r1bqS9qox2/vTijj4Y5FsSTFaCYUgAZoISwcmmA
eL5svPvy0q3rSRSSRZmMpy//QoaG1ILfQItzqn9jfWakPkEY5z/DFTw91dDIbVrFZNtcAbPvHfFO
uFNODpGilkdRsYozEvEjzSEHiWcAtq5mQ4duxAYM8pvy6n/270GmVEzvXRv/v6i0ZJd7XWFe9P8t
mzIKSXKoPMdeM6Gwh4n0C/L4KwuSWMj+KowrBrEJYZyaXHi2s13xlWAA2CUoiygLTebXQM8RoOpU
wLZpwlyx4qXqn4qs2w1IWzIYRGK+3XG5Zhb6qWkts0Gksb+UO8B3sGD3yl+NGY+WHIU6G0QSBMzR
v6POOed6GYATOzcHP6QojO4/IWOA6d1r8bEwYI12r9v7pBnw2hyPyHdmUp+UhEoIPIJfxcABneLT
uQbrYXBv0HIl79ZNT31+l62IzQ//K3lV91oEwYUSDICSFC5c/PfcnofeAC8Y/Sx6DhFlIA//nhT6
DMiZZiJpmTQSGqL1nQbnvDIadgWLxhNtsTpZoFXHKvyAN71rAMDCllzFiOpDVMCFYNybj0DfusHo
wqO9iYAAFaPOVv35E2D64lOkpgfpUwATZ0a5zxKE0nX/6Oj7QfggXdvzdmbI+Sk30r96OsiGHUS2
SAMfRDkI8wCyqqKMIGNoMXiDXSfLV8AiRzRVBo6A2QH9L8wdyKkRgNTduYci37wnSMPfYUB/JcqP
bsxV+d2EHkZ1a4QCG2noD7+Yf4LYqtv7XvfsD2XBB/IYc2K3Sp+xON7NYJ0ed/uZ8qyrOMl8xan/
pRZEEIzjrwnTT6PQ07Y99mR0aAgMHN0d5ksD05+O4vziiNgWvV10jFclH9LRsL8IEQ1+AyOAFIzD
pvj751TVWws5RW3iXP1v4OBQE2mvvbQcsbctlAW/St5/6L3H/qRGWh5HEX09uhfw6UqGH/uCSi9V
rYhuoCDQ2o/QZGlnh8X7d2yhMMzdXZZxJCf39sfYNi0rkbzY7AjXkatoteDo2h/RNeLkxK5X2Rgp
zYdqZGRrUHnee8vB63yDCZolY4PxliguatIrQp6g2TwfSIKo7/gmsFJr9tw83lk+UUkl5wID6bYr
w/Wbi280cB75qrYhglEVCgruAYGh1D8QSDC6rvKIUgN5GPtnbdbT4XoNAzYqT5ZfVGBqYANYK2gZ
xleXUeECiOdSIlXaT2hIPm1gdPBVa3JgEVToj9KL7dnQdFEdb6xVcH0/+8xdIQPKSjWnwQnOqSjn
PJ26/XDnm4hOU3r5JoJMJlvuWSXHWxmpJJXsw9J3U/3kTYDHWVRY5vrHLDQrZFZM5YJjNuvmg/kS
LOFKdPCQDVl2q+O2XhM0rqr7P8LOBovqE0DUa3l3hK6Cj7HAnR/LTYF7kDRYalOvXipa3H1BK+Yv
LoJVmhby2OKNJx3f51k5OImVuZY3P2juSoPhHEMU96AaJXjBZQCUHajZNyIpiGYLO1xbIZsOMapC
4nR26CgWc3t4KmPZz7wzuVrqrfSNbYSgECzm3LoYh9I2W51PHMHfXnkBjLwC3xuWHSQfNYL2OYnz
lWuzqxxnN899LInxOLx2giiltaRc2khvdrzIi03iYu5t0phmdyPh089WyC0coE0xI/eghFmSY9iX
o2WYPv0KNSetgwuKQjQ/G08cQc/Y5DvsivbR6a8dnJyksQ7SXvcZZ2bL8CBkUBlQ0y4PhmZEXxLU
76NIgD2gebRRVHrmboSzsznjIZe8EhMSJmTNk0ig8m97ANs/k7sQWv2hrxi8Hp68qzOMVUtDEj9W
5av+UFvZzIl255vIyS7zqLkNLqngVSzS3HQ8jJDNSHClJgKwvfsDHUaA0oGH9Tdc29sDEBsrAZ8j
xnPZYkGr8Ui5gNwga7dLCOHNiYolWSqBKYPiFDLhxRtzZ0sRpgdfjYnQTmv/QxPBDP+9hvoLlLP3
qGdkyQ/a4VTApg+QkKpT7QpH8MCj4NHC6/xJMOq3D2ycG0xJNvUK+1kc78okaknIgSzwoHDlXave
+/5und9RZfDUVMb9cP1Card+57+KK/SlCvUTff7DkImbeMKvfkTnDIZyvV6/Pfhz6Kk9wrhnnhOe
fyQd1jR2km6imXpF3P5KNQcygkATdIahWFetosKJjk0hCBDNPwVtOwL6eDE5g1+mrL7yROia6oU+
uV4w7g45oVeKJSqdCL6hfvDeGlu3hPk409ATBHK1/6GephSf96UWS6t0nFZ49tnlihz3/1ThRd8D
Er6UkEToquVTjHLhX+8kanHTWp3wDJf/yBvbJvaO60na0/ntaZZSynL+0lndvuyRif91WVx+8xWD
j8xAuoR/x61E3GovG0IgLCENoabdnkv4LsSfPNor2Qt/MED2LX4RnqVQUngPA7flBTilNcngdemd
0FzavdAz4LYEOu3vjQ4DX6QFaOEml7VYOgWsseNSxSukVKM8WnqJPYMinlxz2xQls2XA+gV4FIFO
26T2cfvZXyIfJwObPSIGMn68wWu84evE3MnsgPAPScOvlYxJM2kkq1elr1jU3+Gp3wg7LuFqXziX
zO+FZQcrufp5U0byRLL1M/VQweSP4++LU+zl+hA9ko7erJvu3GrVwhpIK1w6NwGHet13esIzpFp/
wOKAE0UTG/sUC5jnxYtlOpFGhvg+WruDbpbzvTYDyNXPONCsX5FlTs8Q7PVLLd8aN8RKe7Gpyn/x
+NuDC0NDpSk/yna2WO1xYBv981iNrDq+FKoLMP/yYktI+DZ53hmkB6zItKLYDkWVtaQh2SNwtk3X
/+SsUCp/0NhfwK18fZFLzkgsWQ+/PQRytci/+P2aDfTB9YvPJ3h3jSOjhl9lRZ+PGArwuLuxWZHU
yi3w90cN3MVjfm4WGFirOsxb50AvaLqQwbhzad/MGMlle0FqCujc9FuDdFMqIp7J3yh2N1wN+5pr
G4YRiuk1321WaZbv+W+T5qJ6U9QlxM8uhfdoqkQcC+0KYK+rXgFuABocLgRbtYtwMhoaNFGT7cnw
35D/4M0LlvmgJ0mnZ2OMrgB1tlJRSPJGhfLvXbwp8i+bKgwx2rZD/2fLLqrfkorWFKwF3KPiME6k
GbmPlp7RisfebXofdr+ANXWMFhRS3F0avzYfLDVR02E05ZdflhplZ8+QBkWHHQTPj3EwRATtKBdD
s4r6OHXY2rVvuAMjru/Q1cM2ccFbOTlPX3JGeoMEsPzKjWhJP4xdj8PKU1+4ijHtdw9cjwpgxoFJ
QqhNV2BxF6+ZwXzX6yOBAY+KGsanwNFWSZ5CNxHb8c6IkxU5Otw0k292VcBDWcy94PJsXv0tFcVe
/OuauAQ3d/Q3V9EOBh5y7KssmekMxquaAGf6nlmgLjaFq28RnOA2DnKtkOx+SZlbsbdwIrlRIaif
c8nz7ZiEohNdIdVxQE2o95o+CUYThgLsUxTOI5EyqgB9hLavOukLT/nGxeYw0u6qoL6PNJX+VQ6S
Tdg2UbHeSDShoqK92UPkxTKDIdctWUyDjf006OFgyHxdPctWfwkM8QQSBkSEpkY1okzmo9yYqETh
D5zvH8PZ+VU4fhvKe2FyAELaXSxdAObderb0N0YNogzrsa+pgWag1s01BWS8ixKTWLfrOHo31KfT
XTaTzY6X8QXJgNM/nWvS3Wz0yl6/GWMw8mcko/O/aX0oyTARicBsvykkauGFUhsOTmEhnop9R/WX
UeBnSv0bwUM2lXajYSrEFEA6MtSsz9G15JIA4+keBH55ffLI72STfgw/pAlbbqWFpAuyjesENINW
2z3S6AyDY3hwndMzSego8jFZIBsUbnjGoXNJttXaSnqsRPy2Z8SZRx7eeEe90j3g72CJGWsOou6C
xAZzisPWfKiF2x0+T9W0RVgK8DlyyfgNgZFW+3DwsTGho95fGVJybL5+0dGvWGhLAzuEQv0NgFKg
gbM4QuYH14c+/pUaQNP9Jrd9RmW79pydCgIesjpPwTF8SEPVh7dQMTmJYQSADrud0pjI3Dslhyvu
VMHjAR0os+AN8RKx/S8Ye3GXIXqJ+FohC/JakkeTaSC9rORUnJ9Wvhwa7HhpdUsL/7eU9UHQxpKo
Vkzc0R2YUeshe0LV/2IRhSJVkdn/mv6HPq7rG0OT203tLarVwu0yn66DYwsEhgBrRxhQCDwRJI7r
wpxZoTdPlWAyobD3c/L8AHDJ2lrOIN4QWBeWFCsxONY1a8yC/U87teSRm9T6r74d9AEyXHrGO8yq
5RdGzetgHnk1P3BeVWN0alC3ueVfsselA6pFDch84fa1THiuZh1DYbJWxrKLtXwyN5RujN45dQoo
PC7clTiaHFTJtYzkCu58M8V6C1p/JKysosPPe3J7tCJwaFrM7IerDjL31t4jRm2TuVBneXi24UN9
qKFtMHodHgae/++Yti0CKWPByGFzVuIzUMcnGFYhdXUA5rclqVi6RBIyHxLuQM7XnPMePSTz5Wu9
DvxgiCc0V/RKPB319v5K4wDMFTKmnaE5XbqSRYXmPeSz3TRqjpV+7NHndTCvJ6LBix6/fT5FziEH
IylVQJdtbD7hcyI5f9PCFEYNGvdavaPg7j/EhmjSbZ+lPy6I8Ya1fQz1GyrTPDQf5SnN8fe+ekJe
1zw16M6/VHd75ALtVf4TlJ7r/BKVrzu8T98wExcGOL9IOj7uJ/SbHQ83z/K8YzhboZYmmwwNHJyt
WXGz1xZJRqP11jQMqTjTCrj0bp2mAp1uJDr8ngrWEr/2INEx/mXEGoaS9ARBG3GeJudoEP86asWr
Gfs/x0tb5g/YxhY4GWo25gk1B+ukO0ZOCz3cdolbzirUS/ZbJiGHZ8UCWof+qtfBkIKX9ugISF+V
d4WQXMeF5uO+x8pJ9n69NA+7iMOhdJFVCkzCEB2ffEpabAG13ym1oKchqd6vFdt04AymKWz1+C6e
Rp6NDGZUXRtz7Fny5LSEGVfkUT8R7KnceAF0fnQ03CnDGJCPwm0nTLND6oiUZvnK+sym5zVYgPW0
JgVPJlAwv0D9/OMNwVye6rMXe5CsgDJmh7o18PEzw1BpOxjd1zJknoJoKCsvcii7tumSf+UPD0oa
6fWrc5Hmf1z1A7MV5sE5jY5fZ4veXIpHccIyHGIGkLflqlTWDqN7FWaOvwQ4aVzCngItb2wjFotu
0mTFEbaIWJlVP8z+c/8Mu6+wIw/rJ5ttYLz57kmi0Tths5CShi/xWoew19VGbxnp1GIR/FdVpPY1
ycCMMzO1h3oVdlRdcrKoUib+AL+AFDpDQ62zwuepRRNNPfbAEZBRy4xdHm5aPrypYSE6ENsdhraa
3bHfU1LRrtNAEFpIGHz1pjmCFhsh36s6AEwU0AEo9UBM3VSZEgHYc1pVhSYlzp6RoPSMuqHXTMbg
4p6iBHjAYnfeJGyIKAUhgKI0Cq8BKCHyubeQNGEsG8n7J1y6DxSUWOfyvTAbk5IUkVKwaneuRGm0
tMbz7LgS+fICnp+YpBHnzCYOS0BBmY8rHbuWeahYkGSMXbnXpV0qejzd5G3HQh+zxt9ivUQCjA/+
31Kqkt7bUwqy2Kmaw/YE5jyk5N36AERDP0vNAoio+HjBN1XQzotOG13Q1dgwCdecl7ZsyvpVteWA
lc27oYh73aGvzyykIuW9aems6XK/R0kToLVeIku/6/3N9Ko99XV33bB2gLOpHDd/wkClnlpSa/mN
dl6avyFGEeYhHLgylup7OpT/A8YYvN9hAFLzcln/PnMmHf2/7o8GgR5MUGMZNYUKc2h0prYbF4Ns
m2mPaNBFUTItvsN2tdrayg5fwxkCH+i5S7rUi+JwWfPGmOrzaPl1VpFzC2rAAqnxPbg79Zgq4LmM
1z+rrpVjK3YqC3P180Iamsp5uUoagx4mUDiJmuSGxaTgM1nN3Qp5Lxq7x7yzEIRgOaqSC5LZHS4n
q9cf82UdfmanYRFwwyjyeN3lrIN/ypqEcpc4d0qKdXeQkunb51YZoun4xGJuuzyGB17lIiqHAp6k
QtVyanbc/yMRmpE5dKypB125dEqwdHLeMPvjU/Qyp4y/l0SFfDiNWEnR73BKoqW4zY9flUzMRuYO
OzLujGzwEFOl49Q1hBlGFSKPFoFyV1dt2DjIBqlYxBl/zS6eZNqqVo3+X2X8rCxOJy9ubPgP56Z0
xQGH32KeBQxPd/0V7FlcxGbQW0t81iUHFSRU0OmxrHZGIUbso4r0gFjuxubdldgKrXJnYO6iSNGw
hJP6ZvON6zBf4SxiK4lGHAkg/hEs2igKRynresJ16+T8LMJfivnByaI5FumBQMMRSS9SKZtZfWc0
fI8Een2qWl4GpQM/bkXbTEDszFKhTjSu9kQ3kVfHd6IpOk0bewphETIpj3xIX11GRUHJtIXcHE1T
dKyB1BRPHBoqWLfbCkxQJKUegMRWsw6/AYeVw2/7S04463FCun7jOYJBid/LXgaeeyUwq+ZXuU0e
I6aZoofPhq+b2czFz+iIdNl9QvI7d4xp12mfz6L7J9LiTBiOOohWgnHBHaqbilHUFFXGEqIUQvqu
jhiRIFE9AEqUdZ2Qlt/m0FHTmwywvXbkhaW82h3ZWU63h1q59eMQ7PWpu3s7aJS3A/Uei7rNPGEG
Ba5ry8wpqlAD9PoMtKzw7H2Rq/9WM7gvctKXxCVvHV+pKbGFGDx/O3F/7ZuQhTecrOflsiovxfLt
qNcqHKJiG6n5FKw0iG+yRvpfMjt0twTDxugPKkcfOLCdldACwrP74Z2+9ZBAn/XmTXtiae3GmD3r
4DzdEBRVXGXllrQyn5+cGc/XbE0DbTvs2/AB773GmJ5O28Jlq3ctewLu2xlCcqf+RW3mQScygcwI
OP7Rq7vPEO3cl1i2FUf6
`protect end_protected
