`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MTXJFkLYrcGmstIwGuQ+K9WdUBu0OUSMPAPq/gdGV2wnT63hu2YRIVMl3u63iXp/aWfSuXjTLQ+y
K9ga24MOyA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Up1PDKC5Up4jIFrFPo4ewB0Lo7MpU+rkTWqxDYZijvYi8/UgFE6A0l8k0zuw+2bcRz+qKriMg5Pr
3lnOczKZcNmYc0s64pz1daiXX9lkAL8e+vdFzjKs5jLqZc7Y7xDtTvCVROUdkwLsHiKefUqakpuD
CVNebf1Wc9+Uyv7Fp9c=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sK46zLhuakSuyi5tm+555VwQoJHjmnKWK2sz6wa5owubC74ynXGnIzRCHDSnNwKk+D22wWjhmZ6G
hyT4iLVy3TzqtEgszwnYBytxpeo4Z9KspKywkAk+fpqfDMc6Kngo+mnGlfQKBD6VmKIMmj8R6qAc
1efRzwOU8KJekQa7idY7e7OwByGnuaMSKjCQC/rZlM8c7GdYlv3hb82Sy/AQadY/zOkjMMfuNG7a
5S7te1qZWIp3tBToc5WYAvyKYwPRtQv2x2brGdCzQuZ7BxrULERIPB2Xq04Zu+Diz5/Xzr8+ljko
jw2qRK/R1OY03Pcfr2fEJL4JwsWi4x265ll4Ng==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fS+yN7PKOfDz9iOtUWcTY8I1LI74c+fses04RnIoZw5q7CEUTAEmIomHLAQV4+qI7Y6pqXzcQSDP
oYJ8//FXYLkv1lthj51C3Mi0DJmyvqNWDZoA289DySY7igXc/ORPDHMu8bb9odStvvoVheaWKaWr
fW4DNsV+TiW/x+fMsOA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B9mZfPoI7twY47fXG2Vg7P8ls1IjL4LrbSFr+wtRcqVO/K0JgZV92XgB8iraqlyi84mUoXNvQHHz
DEfAPsiNZXfK589i1sJ5XmuY65sDQmjd5eyyqMTMNzSJNLgXbH/eZzKPwDA47Cz5VTHoQ/TWl6Lz
eWC3BBJRfYQ1EkYyoH1/qcMfXebToX1luSKBF0v0oaNV7TexEekRQyUxDC5SDXPrQCcA+iNAhX1b
5xT//g9xuYP4Df7M8ZM9G9iApwgxHgCdex3A2yluTpuqOGEBkifnkaW74YSAzRQXKkw0P6viyP0+
swtUZuXIfIJI7ZE1QayXouNrN2hoebRqIR+6+w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16672)
`protect data_block
xWByLvllaDx4yQaG8ZGz4o3o6c50HP/0uHGDyTDsg5gsAnQdZ9ZgVJTeyz39a4GnsGbAuiOzC57S
55GP/SPOSNji2n5q2L6nzSKK5Gj+tUEhzCNn21yVmxaflztU3LgdI5u/F9L4S5V2w9kaNBtkADVK
2IYKNh0sirNfyfw6h9G4uk9NNpnCVI2vGW8MMXdX2QTQHYudD5OGfKaLDi6Yz67mzS7c/0uMRVON
jnPo+Y7njNvwfwpXNClKqJKh51cAITZA9vAKw8Efj5j3Q7fKhxY5PcGroa8yzuFm88pOqkdxU56s
TklggypEzli5Ux7aAJ4sjz9vCOff+br15bMswUA5f98b3zbU0kIpZbfqGQql5HRtzylspZgJJNzA
hzqDLCJEXC+dfgTUioIQAtp/cYZSvi/RYTPgt+4xn8WUlJ8Pf1T5RB1kIYIBThlC83pVobf5Oxsz
ZTw5PYC2BIGGG+Ngn2VbLmoOAADUe2uoixeOdOUbqb4EyyeIZ6z3/aZ0B8sVwwvaZWjaktMA6oEs
ioTgbQdNjfsrR3luKkNlh5doatDLs8sd+BGgkkpzmtoytbcssxJXiyGz88UxZSN4kXURhkRsvSMo
LHKyTqxPTX/M0rSPiyuFVf4gklJjLIJv/xijy1CUzv7GX+zIi9WQPlsbJCVlekCIcP9Hv3ZG02Os
fyOGE2teayiOnXt7SeYgpBUeHYlH9ZF2cOa69PdOU4moZ9gzgudDo1UBA5SP/UfP/+glu8cDQ0dp
ORFWwoeVksEV2AHTCv4QZDKFFx1NEwr3DgMnnFe48JGClQPtMKRmDkS9qBioYnt/+sn/lcoZUCL+
pxsx7F75K7Nl3ZMKpX5LiR7lUMrG4KH8J27eP2Ac4GWSnsT3yJCDiEyIV7qVcNPItlUSEAuZtPrR
ZxlOpmLKzZmX9E8L7TAThtDfND5zX4bzA7capw3/zf/4Z1iBhLWPAyO8FujcmbQY2T8qAYahGBwc
AYgzbuRsmxzLyy2ERYn1upEk49fYWCwF7RjWRgA7y7WQDwJqiYrABevFtqwy27lKZM5r941jc/lB
uVargQI30BWl9bNDZwoXME4PwsopWOWyPk8Zng0SNNj2pQpRr7sM47m5qVKsfVv7r+4q6I6Kzb9W
4jEFsN+Jpfw3V6SrNIHA96AtMOcsvESiQvYSNmCPBj1vQer51TXffO/IU45sghGlYNSxn8hDHDSr
8J7cKYFwQPhojrEsNn/hhpUGR371fVJ2UtJyxbb5Z4MEfFwEKuOfYmRcdSB5pw1fRanIb3zgCaf8
Ee1wzocxTy4HqUTaX4dvdkM6RCwMDozzqKxqDRgSft/XrUhVj3A/QmYeEPU0zvDmzQ6R4uvivlFg
KhtoIH0PhV/yHh6JRv2j9xFPkl5HBFKpdXfH6FaluxUhA6Y0x4DRWgmrQ4U4zRuuLniQY3xQzOY7
v2M6k2ccFRoT3AZmapzL2e7Iv+txY5CjXJHcShAo5DSmj+wCqBodc/ed3tan7NorVq6+p1T9lCK0
rjKZ0G0+OeFpNEyAZmQ/+5F3KsIMU0MIjsnSddXYfabiXmZlM8DuIJdMj1lDbxFzpbqG13UK4ugy
K/EEMxKysKcwpgczZ2gP1AH/JtMT7R9bWPLE3kJfsLteIfENqWHWGG6vM8e+JIVT1UK6pqOxYlUt
hyaP5AGkNE9YgQkEJrTqtpNtznrrtG+wHy5SGW+qRTLasgjt+bhIg6cYFRZ7oF2CIby5I6E8ve5d
Tua/l9rGoNMn6XV9rmh456l1kNXmkX5p/kD9KShpjuMhG2x7vGMCzY0kI7Mh5SK17i/Mz60040aF
g35Vq5B28cPyts3iP5u466zBKiL+Ul8c3ElgJmH1jrL0dmhS008WL1j3qUh6wsTK8FrKnbzAEiD6
bHlhjpRASqDM2gAaH3ogjTzsH1NdnL4LQLfDQ56ST1yNStXflRbtHa7VDQT9ohhHbCufNw6W5O4g
5rcy26SDBj0+4glP5oIDHYWSNNgvH3ps41IjWkiLBiKcxCgdELpSKqZ0LU3mtD1b770VgHf/h6B+
eIdURtBv59OQZwhXVSH0255FTK3KQsOjwUOEEIWrILq/b7aashr/Z3hMR+UT1OHJKA1MhmRx510M
/xsOC1BwJn/KZDnkYbuOhSKNCRHasWr+AXRaw0XunKxxnR/9z0wYZ90WzxVLX5KhUyW0dbP71dBp
T4hfIWtJzwWCBWD4W1K7dHSxylLa32P/304BSA+nGZHFacwP+Rsn9PiPv2CAeYALdEfQSf8ssjRU
CzkcCGl7QYTrph/YMABWZ01U7h4oy8BQ9ifTLORJtikbWCL2TPVpsINOseTiNkkcsXjay1gSd+Kp
ha5kHCSvEFB/+NgkGlaDHL8peS8FZlsA0/i7RiF4weR3AlNudALyCsUekEzamMSy90y8sp2Vjbz3
HEDRBBGPhovb9xKfAvNq1FGFUGHvFAKdgRvPOjxKfPAFkKmfkM0F4JtmzglvcSzbbSC8VGOIYgJb
XBC5C5tzRzODrOpg7NYQEt8zeoJUenvNvFL9bI0+6R6jhE6MB69ccm1GfDSRCmcTlnm+29EKLP9t
5LXhSlsqV0Gp0ioIEtWUP/IZh6UClDHsR4+XWhOZ2UjxidRmeKJg+OJbNNsvR9GzIKWW/QdZXLbK
Mr2xKpjhCQ1OQ+8tGySAFcC/N8qihtv9j56nia1WmiDuOp0LLunNd4oULzcLmcQvpboSJh6A54nr
kHpsJJqI2mVchlefUCOSoKHXRsHElCVAT0XDoaPyEXoEHUQ7nFyV968Jr92dPCxzxR0i1RR85AbS
qsmhSN9A8Gac2IEhfw4ebtvD3jMrrKw8EJd08CIEE9+Ieqhzm0VHWxzkDcBIKnXBc82Lb1xYxWUg
ywaqC1I93GwQDeRR0gXIUOVc/4h8rC1/XUij3zmj8PIHEPI6ZNA2F/ptqMV60n4TrXqUB2P3aaDt
/vK5mS9FKXjOK5XCzGFvRtxX/PVcnWfrLqqXKlWda6bSgfaEER6hP87Vt+TUiPVjmuEZ69yNFHi7
LkL7DD5k7HxF8lzt71oQMUMX8PuSR+0GeiPDNqcPHOaBPmr6yphCq4g1MQ5E8Hq5n/Jq/X4ZaXM3
g1S4tPqEy70Sz4xCXvApcQBw5enkwQIhx/OdzIr2dM4RACXasKQ2rq0qAwXahPevUbD18ZqNgOH+
8RrxWOv7wX3LJguxZfGSVHM4fQLTCR5hAe1GDpDvXryWSBlASXIiswDyADRFSjjOAmRSB1Zh58gn
PFTilsqsbddbUdYMo7F3euL3PwmJDmyGn9kVRguOS97rCA+zFW1NEIf/XgDYmTPMchNFyxOuHuDn
Qk4EPh9eMzjJGud60Q9VxZDMySYDJMz2Td5yizXHJpb+kq9M4ITtXuTCDJ/vjC6xMSHdVBvzd7Uq
t3pcsVUxpstHHiF/tPItmcHoEuZ0VdEB6DTq5lXSGz5OZPoK7XYo89rc4PQKo28p9ZEc5NjDsHkJ
j21+cvAChJd/BVeKcu3c7zRfOP5gqbyBYVCgzh6ApltP7UxKhZjzWDyVN53kazZL3k5o20I2gixc
CiMPkZtGefGFNayXhqpQ9GmzeqlHHBhAJVNOezlem+6fOCx76yJsLFL5Twep6tDGftVYlCvcP9Bv
rvo8fBtsRxwvcw0Gl4jOWPFEbsQYgz4WSUuvk7sRRJ99XCZhQxj3b5ZQ6pWszW4kv/X68OfiEZRi
GzG6YcSEZyREt/31w/A7Vz49ED81iQKj3T+IDWcq1IzszIjO1CDkk701Le4/Xe507acxvrnKI4p7
zj73ibhV+HpJjK4WQLx0BCLcByj4WALyOH/fs7bSexSyvgkkNMKczqC1EVIrMAfCEdXgeFeOb+bF
9QM3iYTGhUxGszDbPT8xsPdbvfRQbWGm76mxmOVjEUfYR/4pPlf3mLonLJGIbxbJ0etot/dtP7KI
E39h0UXHSBVuK09iCXXTC5fLA3PYXkNFuTxVc0oP62otksDV/QNauEo0b2hTRK+lSvTOrAHqN8KW
tX2MooWb7kSOj8xfpuevfe+HV/mCucYbf7UnUhxVskEsLYqj7p+nTmpZ/i2/apmNSKNHZWRhmRsl
cEHy+urq4b63Z4FiCKiA/cXGvmb0SejlObwreBAfcLH5ybhjldf0A12LiwQlm+9C4Gcba/Cif+kP
YCM3BfGMkQtXHHkq8QzfNRMnB+zo5WXy0WcDJL4I0W6h6hMczYSQ4ktgqK9gtssHkOwRAhVCFpyT
OkiKfhK+mPsm/fvWGsnBE2r0toRpXJUs0ASZLfT8sEKgnDB32wTb8wWdXSOOnQaGGhzuhL8NwCjc
lUHYmVZezOBZWMg4fB7JU9ajy7NbZbw95gnbpp+5WeN3ViKKgORXYHw1InfSrdjaealYeNxHfvSi
sJ2Y+24Q3ILGyL+dkOd2zAopKWFtyOF2mj1raG+uSyB1CbIV5Y842ds8RXUbYyAq49u5JRDTNUJA
j/dPPZENzk9LDnaYCRW4xsxaNFh+lXjQHRD8a/l/y9mBxsw69p4XXxxOr/bGlZLwF90CE6AVaVdD
WU0tug289Crs4mPE/iG9c/tU4SI4UiFoW9Rq4cOg0596/A7OP23LVuAe8ltqjrq8U84ELnfccEpK
ytEIInx8zpSX2h/rJXysW63jzi4X9Al5udvoSbrgbZD0C6iYlgJZdP8JXyDPHhtvy2aePM4H3Bv1
WvZw0cdTjAtEVtK+EllS9I3T7oXK2Kw9LOlutD6AhzsGXwgS3sEOIZ+CKckX9bdWL/KT5PDyw3VM
LbUY5AeeX4brED/jcACE01dyn72JNUIBfz2ppJLi70z4HAt/0u4MCD4xwAW9UQ9O6PZFB9Vz6z8C
mPLB510zBL/4M/guvCKl0foLf+b5HF0W9bZ3KiWUaoOsSrecaxYK1HCOlMtRWwT9fYvi4fhXb0re
1/Of51gUWSxLh9ylMpOSTFOAxZKS89XLMK0LwfTc/BUEFrw53J1D6ush+6iuChVoV2giUOcKexnB
YpLqGGzW7w8tfdQ5o1oDUKdF9k85QA4YnykzsIq4Kp5pJuC0FSahmgE6AA2G0a3bGLU7dVdZRSE3
50aBqA+RUQe3AtjPDdEjQi0NRJU/wl8DWl6cx5W6wJryNfYUk4+08Lp8M6Wky71iK274BD3w1AHj
YaycFJsPFeeCoPbJ82FCztTlRGwuRhxkr3A8rKznoeiKe9z/JvJGODPX5l7Vh34PKXZ4nyw2tHp9
8T53931tCxxwVHApn098ucTxP5raWk6+yu3NOmorow8B2IpZ9v5JWh+sZ08XFkj5YXx/1YryAfqq
gzHMdUzkfAyLj0/C0cJ1PGKlEsxNvRP/fWYG5WG85uoTg1HBkKRXA0xaeM+v2BydHtltHaEYGAj+
iIBqDo1Vz0h74duA/QXKxqG9hfJce/bS/F6+jbmY5qENNH6nwCRJ5G281b2H93jhOUHrf46M4rXj
EIZV7orDPUBWqwD8tXL/AIWOb8lDYsvVDgCyTLcs3cTz8Ev+A1eWzai/7qk27MbYEXKxKHxOwLrC
eTEJxPVXQ4bcuqQPmBfKY79j9QJ7+4JF7itrpS2uAp2do3isc4d0snUFHd0bdbdkDWUPi4ym988g
8A259VD9ik3OfqlKeKrrUB9qVTjyhgLsLeaiGjCJv5oQ1Lz7Knngn/9F+/GTIWaumN8TUPpS6vEE
JwzVZbuEOuKjoekq7hu+NHwounBzzQp5xoXOXE52Uqg7anHTs8QFWqeLp+somUl74i0DWXe5bUiE
RPfaYas6BJwstqZ84x+qsvNNJ/b79QX8Bv9W1iPH/Azw2Xo99IjqBgeJm7txCjdoqRfLTYkcP01I
8x/c0tNz71BJ+VzTHf78P31BJdFryFIAn8y+Q1eKEvw9VeuXP8Axhy5ETua46frXmklpTq3Vh0h/
Axnzml2JNm9Mvu4TikipYp0mwPHmne4Zda729H2siKt4WTo6ydErJpUiOKeDhnk0nFgYDeHNPlzT
CXHKOgcA6B5UZMrWkRc9bYOEGc+AfFlpuFQycdrbeonpDjn7B094QXSN8pkh2ONjrvfCgvIXZKLw
T/A3Itb2QyzyaKrZsqXBAO4MZdG2ZHSXz8VkVzussfXLA1KhTG0YIKmixAfrYuGrKg0dQ3SfbDkI
GMyXNCrhE+ZC+R/TaTjEOTdc13U84Wrwdpp/b4Freb33s5HJlCHcMuvAkFMqsx8aiGJ/SdLtCppe
HeuXUVCURVUZ6AcJ+yTY81SXo0kBtyAuTkJHsUBGY4kjAQRSdDOIhKvzf6IrNK/WSxfQAqDK+lKI
O5wjDUFfoxPyT+88Hw4FZyIdTp9egC8ymN3+i6xeZWas3sXj/xAmZMqzqgIAbFO00Ylnp2YnDkZO
aUqsab8sweG4r5d/xYwJvL0rS9jzZxhsk8DJeY0M79IIPasJs8XA8C3MsLLKIHxChq+qRVO3uZAv
gFTegKIZ4I8OlaiaYCdoEH73Wpfm7Z/CkxI+0CoXVxkS8Wr6/0XTK9aQdpRUX2/DgLflhcMrz2Tm
068g8qjiWrUYB0c1Hws3TPLBUhtxulyx+SjfvJ1bWgRcID1MaRPg0MDcGITy7QCHoIBm4hM3kWdG
9lTT02yKhtWoewB3F3rUltvsllccpYAqVWsLcZjZIBwyfxNIs3ThoNk7boyNOA9XAtq+XN6fLfXv
/m84jYe1ZQQbDQSy62QkCbTlkFGcrRvPYJd5L0Oa0bYUV0sm7Jr+EbNzT4kBaAA6khJIEMPw1Uyg
tnalDWRjSyFNWVTDJp0FmCCBhW4WSUEx2tnJQP3f+aXYCCZpQt2ZaUMfcUrgxKhJsx10CfFhDw3k
oB6Gb0md4ptgRzXIbCE+Lq9XpwNmuvSk7awc5Q8iXTo5GujeZL/tDfch75xYic2i8Y0ORKOi3G5y
3HOC2vew2nCUHrf4bL8K+J1orAMHsf364xaG6Mn2+QsFKZDeL8rBycE1avfqpnWE+M6mEobunJ5V
yPayjTgZ7oMYao6N+e9+aNhafzY5ucGvdZE81PvGfsJUi8Y/Gwfxkfc7vj8cw4LPjXYwlMW940dv
PB2mkdFf17Y0+dHsgfGif6SpmfbplMcW9OgZpylxgywQ7beTBOu1b2THHDSjbCVR8X0/BxVO5Cmg
iJluMnoBwGN743J7ic7Y+FLUFOPZ7e9GUjPhEDKYipQ55ipbxF5m/as656QyvwglpzjnGC7YGX5/
1eY2Ezs9Jq63Uj/yL0DpcMiH61HjVjjCXbFkE7K0lAPcPAdSnmiYIpddqqMlJrD5PIEpVsDcSQTr
D72r1+jR56H8tisOpgn2fSTu0JcjZMygiloK8+OwZAN+5hhlMCbX01YPoYChHlei+PXn+x02e0Zl
ZKZ7ue0mWWp1t7fH8T7LyhTWBCQfQbFiYDWJX/Fpt8cWN1BzQ/3eiDg67CVSpdjQzvuE9SyjFzZw
MSAjAozhH1NJAOajs/f0T7aZ1JX3mNxaZkYDL/RqlPIqSz3XTVWQaCXM5sU895LZcmYF61vpS2zX
HCs/UU9KU/K9RYTE7jo4sVTMskQoVkHxNN3Rm/QNd8F52HxMjPAz58rvt7BREqSYoDKHMSNdPQsP
+soLy32ya5Nki3NFhRPYSCDJAEWJXfy575pNB/UWI+9FowIK0MtaJTZdLOPxMzndSrimuY2H0osw
59PKimVyXezlz2zCUi0mq2mR3ykzF6AAYSZmeOvbpNGy/A6GXnQftlc7A3l9Jy9Uy+RbUdJlEoL0
7sJJhxUQClf6TLvzmwc+pw2/yb0J6RTz+rr6PlY4p02lDuwN7cxdTH7Y33oOi/nTkYNLjieFH37S
2DvyYh65GaeSEo1dsCJOO/vYKWH861GstdBeSjbRgnkoungYsnJ8ZIJC4vOUKJuRrVXaefxy18zH
7ZP5C+KW5G5sT7mWvM5Hu++CS994+q31lfRt5HsdcQIFzN7AxzRuf9OxIP/rJee1FwV3euFhR8pn
ztI28Xx5YzkJcDd5DjQtkfDfJxoTlV6QsvpGhf49j4R8VwAZ9LHarvnPcHBUiyjkwE9KSSvwx43h
h2roTTWL/DnlVJ52lRq7/k4E2v7IMPbX8O8tv+HFybrsCevwWBRShQ93kj8GMRZuVlzAS3YSAwSy
niBXLpmvCTWMBl4wTYo3vFjTPv0lvri537+iV+bG0YpAxQYoCZnL7GJ7MyriFj9bRoN4Wpn7FAdq
P4l47QZovbKrkjVYO3OYrdaWPDlfYdu+81vr6bg6FMY0/li750b2Drw2yeAZt0wu9lflkoo6Bv06
6DS+0wvLaO4OIburJHorX0pHPe3QoCha4V+BFwerAgRifDmHSWc6xPHOD0dPa2woQHcU42tAsBGD
uPNMRpFC5C7Wc8v4Z2d3bx6K8mNq7qihvQy11lfpwNiEK+L9OiPzGbZr0crdIOqq//tSZ887QCRm
VEaZ2yJHouzeXjI5gfBDjGFIEFnYpRHPszwJK/8QAZIMgL+dZlNVBBDUzGkF2w852jzBUI5zTpay
X9IIXBWtr5GdaG9l2QCEZamG4x3tlfxbOP7XcqmgttR1t90tGEJlQB88gvZoJaKJqCI64z6ZDWY8
OOAGzcPF64Ll121l+eMyixphzPh0SYn0ucx+8zyQdTHuXt/np59X37Oeajkv6MesyyqWCbnYFLUT
lKUT8TcEyiz0wECwqwBfMMtGHLUEbasC/AEMN65dcItOXmRs87d6AMEloNlEs0UWX36USnbi7mlM
1sSP3YFT/m+9uYTathZXlUAnWdTv6ukAzp5d47ib3nvntylKbcnAgX4iUZgvi4k0FuxpYgxb4cEL
4c1AWa1Re7x14RsrFw/8zqaI9tyvH23bUBgMgM3yZvmOA+scOGddrKcrf4vS+D1JHSEnKB4Hr1gN
uYcvy6oUTH7MaJuk7M9wSfIxLcwTUB57xK+nxKUE0mK319T0Omsqe9sabG6bEelxj+e4COumofeF
mqxfFxBxFuoK4cQveWYqebHFjRWK7VCmUgrrPuCmEMsaMdSY0VAJfsG0EI8xqzT8sqyMGLI6JviI
aasFdSp9k80Jsy82llwq+BaCph3MiEIeg1v1v2ZYjfPA8z+4CuavdkFSztGbP/gPQ04wy1OZBo/c
aNWauG45u5aRQUpn8gOaW/Lf/E/a0ZckUXSb07inDVO2YFxIhi9HgJyOVo52RM+LhmtATdEgytCa
wnRMTtXYsWCTJeCHSlgnH5J7g9AmRTvyQA26Zu/Xhdu37iVUOBtrXMUHhAeGrNK4vsYehfnc2eO4
7dZWpJOW1xheoUKXa3wvd35vCFluiC7z1+86Cx+DlYTDF0o+YeE4hu1UVvSM0IOa9I0RNZl9J0UH
EWJ1L9RQQOaBARt0DnCzsZBpG74aJYhWozJSq9bpc7ViDCSly/gLnnZE5DLujjvlnyStJ3ly/aKN
rE7Z3YZI2qcVRqRIuo3S50h8s8EfTx1ZyOVevXFuakE8SSvhM2t2YO87sXVsnEP8ODlYpJ59B25M
SpkQUCG5CzUA52IjibvDOtWxi3l1vXASvD/Os1nxUhtpCgo1XPDlQq5jPjr/4iDmNMieiK3vDQ2m
mdTwkdsLFvE6XZ9gANb2alEII7xf7prXxmaMFyj31dzT91UrjCsFbK5fcnPdB2c0zr+dsnv+qUTR
HAV1nbB2li+YHFMXGkUrehhhkc7V/eOFyR3ITZCzB9OPeyjVLZYYSw9or3DV+jGZ0wNWUiOV+Ub1
Vf6Ohit4oT2n3k/GhGDsrhE7vut27LXXxd2wHt0llW8/4pqIKd9HtxjtdPOXNfn9skv18ILZVm3K
4QSgszhr+3O94+w8xjwgSRCrf32rEVOsm4mvp1vwmA/JU2IIRCFppEzVb4E4IikxnBoU4oI0s+Qo
OAj32MT+2pFLxj6Vw+rk7SbNxpsMzHeLQg9j9ODDkfv+IKEUqoBRYlmvsYGj7VsVBfA97cpJi4C9
riurF3GlXRkh4WsyUHp7DAUKcgSijiOAbv+qZzJifO747n82wnCM9bb1hhTP5Rck/vHF/YF8Z2UH
GUSQoIbUIMiQzzrucvTRxGuNIiL0OANh8Qjz8J2U2DCYVy3z1d4Npf5a+XYiHqgWMxMa+O9pEzws
l2EhN7oXbiye7UKdASsek43ODTUPmYQWnJy0eF3tF/CuoZ6eVSznTN342pak/b8rxETWAFHyaPiw
1+D7WIROorpsu4TlS53J9ln6aZMpPgHCa1KOd2tWGObv+og1xmg3G/koEo4nrh6HhY3GjBen5dVQ
FVIn8+80P3nl/UDGfCBLhf6Ij5epsmibQkx8BtokVSIaa5B2msR/CfSZib1XhUKdJw0SvuQgmZI7
aUd8mB925affv5ETfQo3MptlBzgCrHvp1AOM2HJCN/nW/t8uvkwHO4JgP4t8bMEDrqbMjP4G2qHx
/Txtp+n6d2FX0EhOpqUrpLcyR0QWaqEW27cpZUSMrL4V5qP/CG2KRj6Kum0/3iCMBnNDBi+GsYdp
iR00V/D0fgDhMpgXV3Kg7tTbCyNZ9Xf3+JgJAAQcA0EC6A5C3ifPNyXAA7Yi7Vzlxdb9DnpA9XOm
+xGVJCSZ7pyyKbBOh6RueSicrZ6ugikIwyfrcYG9NKIINyV2EYt+O2ZjVWOKlECHzVZniNZk5TGF
pxo/VsbIW2cmL26ag3TXioVCk8t3iVaBX0qkltAFSHkOQJXdEkKMgeDuYutuN+fquj4rmkmBNd8u
pg0OdAve3B0yibhvUfHwAxFGjDQqFUm9Zb1RcNDzJ6GM5CM84+nH6DY5aKBEuxf46IB9Or56wXbB
tFAGRNsig+7wbxbEwmZhEDIr4CxZF4w75PvdtMJwHomzigr6ESpN6bs2Yy8Cn5ZlfWwKcQU0Nrs4
UCwXrHRU1xQoGZgJn3dPV4YwpfEUB+wrina8ZRy6YsV/CRa6ZOOdD2gBw8VWtZJ1b810O6/Bq4AZ
o7YFMMcPLa8P3S8TrHPO8TBDhBc9VetEc/BYUaY47P3QACwgu9hXZNkfTqG5yvvWDeCLs0f5/ant
3jAVHON0j690jWCZL2QCl71Sl3WjUFkGKCmjsf8kD/Nmfa/4rOzsxMy8Q3kThQPxJkHG9VNMBUo2
BukfG/OGz/m9LpozCv11gTbHxSC8tlUKgUl6loaWsGwThx4a3rrpF3Ndt3SINFTqfTqTs5a57aht
z11d0wbuwNuKKQekqsBpX4Q6D7vzPIFUTrqBEIvya2nb7xGXm5nUzKWjVOGb9QHWzjh+RT/Otihr
P2skSVHzt23nidFCfRpnXonKZOElTNflv8+n7wXi6FuSmF2QfMlbQVJ8kG9MUjnxqnZZ/1axz2l8
+uWS2ZpT0Ix6PjdYWXuS+w2V2PcpAsvEM9BmexH7rIA0GtuE4iOaXJm78LjRbf6+/sOYwm3g/Q3e
5/SxuBN3jnPqZQJG8inyuIOsTgm1E0CJLqlQDll9VTJtjLLo74Mj0gamYDlR/KsdSGuwngXJ+3YD
R8DJZGtsKQ6/v13/DmIlGkWOMj1v/h+nm2Y0dW1cuBe3Nn6L5iqfJO4uGbpdVlQyzHFZlzqR24NQ
oq4zVg+1ZRnek8KvFHvIPd1rSShonl245OrEArdXPhOcF8rQQyct0XW/iZQlRAlvxLa9UlXnVAC6
DO54zEPt68Oi+FgadGxc2XKT6lFfGtZeJWfLDPXzT7y8fXWSOp1HbUKGyWfvnXlb8a03LNNa6H0l
KT301vuhaEwoZHwhmHjKoNuGKP3U0QhE129y1KHXHi1QqFtjphuxf9tFyZHrD6xuThVk46//dMPe
+kKQizZEIf3IlA+RT3rMAjruaGWkb5ga9isH+ud9HiBJLmc702krolFHm7Pz4FbKo+hA73PFDF1U
iM7M6jMVPigw0f0ZlYUna4Xd5UkjxUXScpd/PtWqu3ugA7o4+9RUeyyx+B7bVKliQEJ1cOWw5syP
dNO4eoM3HpiOwGeNwle1XQ5Tg53kR2wxN0HsDiaeKKcyG+v2wpASuojHTOwJDqk6yIGZUf/NTvrZ
YFqv5aUBvKjtCjtc5ds45UflsqdQC4kbi2CrWXs6JVlYXLgeJnSuRXh3W2DMGF3HAEnKqc3F/Ofg
HOyROA340UZn9RfHYw6Rwh7RmHaSLFIaQaQ1T1tOBttaUY5GaiEoqH+AMlLDLtytEcp5zNLe1fI4
d4/QfvtkspHow+iSpL0vPQNWbnrSX2osdHYu7sp7bdHXDUVbpKOymsrKP16GIvfHzXqjJL+wHXSJ
MuqD+a9bBcknSToafxYNgKPlX07Dt0mhhCGhChnkta7Lt7KtbQPBxwinLQ6bbkTVCdsdtWS8Q6BW
1j6ow4ddC1r12e2HM7RYORyNbkoZtkvkMadOCKGlC6PVKgXo6UDtlYtVnwiQVy3mzMpqU54krZlJ
5PBXFD/A0ZiI/2X5JeDKAomotPwB3Hu1/j/dkow7KzqGizYhC96s6MeEOKzd3ZTnbCggJoI4Y1sz
Zl0n8+fKBmFBlD3WHc9qOjfBhd3cApZeSPsgkpOMCcBv4Km7rxs+amscgA3qbC6rBzXGq5Z5Dc03
Dvo9PEzSivNGV2SqZRDt+cMoyqUUF/Plq4c/R7bfnZkPE1B1W8/26Ax7GMd1agvyoR6u2ld4H66P
P5LTqtZvT3TvNRgAMStEVQ9sL4y5ukuGZNOSxjZI23WqwBNwzLtFfyumQEqHgtyopByE+P52D93c
MrPKex5vUBMRTNTHFqDBguRB20gHUxWlfNMheyBmteUP7Z1asGV8oJdpCS8A1OghtTvQqzb0wvz/
xigx2JALTMg9S3t7pA/CE12mJ0j5rwyb1u9sAyo9SfhEIzRpBZCF0tsmLiIAUbLOFlZON364py5z
24QXDdU3MH6y7PWerB7cNBg8vaWrG7/uKRyMcrpL7m9GTIQ1uTRP+eqND/qsd6zvpV15G6cEql+8
YbjY6Y8gGyjGviTI1bRgJ65mofs6ZbksYwMCEnDlYjFUlt+o6ZvAiLBT8armWsW+UzPbDd9qRRvG
rxCSkBBfngCv7v4iPcsxbJWRi9+ieD7zw0fhOl3vOOLrbMw90fEPMHr8LSu2pGA1xXMzjK2RJSkV
yqfBudj/06Lm9aWTEnrmoHkPGtnYPTR1MnpfzpCq/MSY0D1bAXYlO8uieIjhwcV8V9GALd8n4DyE
pebu6VjJTWIcGUPCtJ/6iFnpaFDThX7Qu++3QF2CjNGEzZ1OmMiWbThG4J0760dc+7zU7igcsWuh
1LyLl6Qwwp+fi+cjH8v4D9mcQKx30woozSNpPBJlJceXIVy9JZ6U2vh+lajqjPGX8MVPudHMLCiC
up3vPi77XRU4Gu0g2KytSkYsHxSHo41dbC78M422Nq0CDHM9kHIPa0ZkvKxZVsXKbb9VGaOHnB5i
4AZl+gpsF6aZYm6YpYHtpq+kwqDm+oWXzxv+6EpmXFRsla2Y91vIcqA8VtFy4ETRPOgQSD0aOYF6
1sKiFTet+eOWa/Q6QxqAcCnI/0ZsBjK+p248v4BB9p7UO9dlYZ8g4uShrxP+1NELye79XCrrgtQp
ozGMhW6nMlYZHKnKAv3QSJt/2xfe3/x5bU6s78wAX8NafGIHzyqNs8pi5MTDQ8qLq51sXdG3mKds
iXKXuHLrlUAXrmoa2PPFBHkAoYX7h3szZaFwwdcFJYWUzLRYdMZzjcey40H5L5xHCtZ/yCBBhTzj
XnaMzJZfIRDwHOR6HPVFbbW+WsivubPPDpBsg5LuZBumUAxHziS2s2Vri1/bPSPiJbqmnehNoYvM
rHVJTVpYWzAYjQDA4XpcdbZ1pXAUi5wMq+0VpILSNANRUKkpekRYy0SGZmvL+cxaNzWwFzb7OT49
2/L0VfmPgp6uMhv/8g+wHMQ8yiazYFX8WNqTeNxqSa/LVO5M6449PoL7jdhMe2dtD5HgA4xqyHow
LzPIZrJSD6CeYAzfxa0s/Wud4UDHlaicR+UQM209CDJRLa7lM+rL9oA35KXhisM+Fgr2p2oy03rD
1knZgUwX73Iiu3d7ZQzzI+hrOWSFavSO7EymGMfQo84Ed8q6moBynDZM8q9teSLS6q2cvrDM3Qdu
LsphPfhdTSBh+I27RwU3tFNGIN4I4vpzk5TuMO/qQ5ttsf82G2wHnWXhx9XvNfdyp9DbdFYLd+Tj
sdif/krcmc8pkNJtUXcVYuxvGEBeernRM1YrRZ2xw/QyivxyEMvVtjZupG1LgtAZMSC7He2NAy63
Zhn55271wi3re42hNAtI3QPeLUQP13UMZgKsdPRuG35Zs0C1RhhgKhdT14PFidv4qJttO1pA9Rla
6SSDLhEXSsAYdNnwF4QhiPcCkr3M3OEQbbH5ja4M3RYS5h5nBXTNYPiZ7Y0D+4fQos7EF9FNdLju
MgkxUG1bb8h3x3oaEyFOxLvKi9ZRWT0cfzxOHxQjHXi+S027/ZXP6Ju8e8NB66ulfcYtMPALzHsu
nsPqPzPZLY8gv06oYaS32Ne5XV1XlShG+g65Xmw3wKlmfx8frcG5LoFiwEDExcONEJX9/qGQUalh
RSt1MEO4FB6oaif6G5HCc4cnjFNjL9G54zzfwgHSw7yDCVqIWrZUmYrYs9Bhycb19J9jgChJYr5S
uKRgwvpOpHR2/cr44S4btLUvMIabregRd2wYm1NlForIb0xXPxw9/SReBn7P+/v3YxPN3yEap1qj
6qgsjXmNTKM8p2H23uZS5y2XLGwRuTDtTlPRgS1Kac9WxDXgXq1rYTuXoBdQovZkqnIroOBNrfTs
ABRSOg7xuRpMMeQyQm5UmwP5F7oSTrjcl2SrNlb8Hc8rBeHFO/AVXPCAgze8YGKp2cwzC7kneNRY
SbDBHr9bLl/Liw0DnJBbE/+07IMbsu/2anyWD23xcaEuasIIe0SLfgRh6s9GSL7Jcr9h7TnFq+J6
eVBd7CpAqi5sz2XKDSa1H04uzdI4T6Wyhu34ayZxCPUSDOZCC+wjaTwxWIGMqz2Qa1kPvweyKAx8
llF00qPmNfwA0gyn6tyVDDoNZ6VwVsWzxtsyj19upmI5Pu3tRSv7LC7iRFLoSjxAm3ep9nnKYZBK
vNw3Q4Es7DmE0yBGKvaMU7nmFfROk0KbBb/bFglA5VORrhxoMxG5oIjG/2YLOQc6YC7TxzOpnkzR
HjLRsrzMUtuWhPh/a5PSeNEDngIIVuGzCOI4uKtcmmfltWyuMnqcX3Hmc+AfHJQSV3hko4YYJo1z
p0yCh+8SbbgyKVR88quZZADYZ5or+aqJxEcv/XBVbYb1y1iEU/qn3V7iV5E/JuxGO2ljBwWPTB0o
M5hAQX1Mkt9Oi5+L0KbKImNlrcq2rhdEm/5H+pXZ1XQt/uCjTeVu8uPJfKh/ks8Afj6FmfQavZiq
y44xZIOtCjoT9VQX7FMbSGhIiGQi2QdB4w3izqSOW8QYEDyHaV0QkOkLEkb5zQf0rHU2MAlo1aAl
CFzucVJJ9MjcPH/h8CVDErN8RYyWj30oZY4BdC4dw4ut7rbXzf7fTmXVOmzbyRHNIbN9djuor2KU
D3Uol44e72/GEQalhkm0PW+hbWNjrOe0qT6VfGYPczPapjIqUb5kAYo4PjqqDwPDj1ZNpPcLBsiA
imiTe3kHvNlra9KGnrbT4kSnRSi+a5JW/AqXLhi/Mmfg9EndyWkwJgrp1+9CcJFvKNFhpxRBMq7J
waoUSNyv0t32VKwgWYLE8SoBWT30nfzAUCt/w2cGq4kUgCvpE9l8aylFW/P+cfysRzakyg6InQxv
8s83mZJMeBAZZ+gFjPNEh2kxwphrg/ntLbO1Zp3DjCB1MwaRHtwkkZc6lUzW6p3bgi0BV58N0ic6
GaRG7Shh4B4r8FUJh6kW8BKnwa92qwBMslvzlAIr/MrebYlcvr3sCWTwoHgVK71CLRPLAY221ij9
tTvRHRLVWYEQeQwNtBEUP131JB1M1NtOleD55Vrk1bX4twlMVLI+o1SEQIXUNcJuM1f3fDGbiJlm
lNXiEdA7w5SHqfrjE7CaF3f1dK8lWlv0YkTkI3SMIENltvOjkCjTuDpPigNH6NzgSREgc44bsNdX
cmquMkbBIv4MZtTZvpcTmm9A18Bm0/BzdbQylzvxtAvhWTgkkwpbdsR9J6xbSo2DpyXcC5Z94RFj
jna0G5pE/c94P0HJVOXvvdabjuP9o+wWSaDIjZyvXtAjSjJB4Zx6GEMVFszUXcm5Y7xmLoBRc5RE
dGfpZlaMVL1eui5JVkfoGti6Ux4EIiI5AqRlc/4dGJkasaYbUpqTRYQAvZypRWz0t8gWvmkHrjQD
Hy59vERnTbjdEoToVsou6JMCL+c1ZNqLKzqKVEOTKuuHxZrjlHR0vS8mi3nkV3G2F7tQrUJzByjM
nhmbL/xZX567wyXxucYG2T0PHYbaEa68FqCaF/xI9WNtBipuIamVcp3UWzfVBmOsQbUsbC5zIM3F
epApXsCDkhWd6AvRDFIq+b4//DRdwTuXc3Qy4y86xfTjrYNUUgXeyEaFjcsRa+Npw6vcpriCREan
nbk532W5+HGRyQGsQCS3xA2SSGsxRLWRKtpS8nHetFAQvePfBbV9M3oC/sAlaixh7ilMg5ub8ot8
ySXvrFpfkS4OTdp8O2ZQBJUXVEF06+DfVo4YlT1GNZmjz8CPLzuFvuJQEiTbj6gkt7X24icQNUN9
jFtnKVd5l7BgrkMUdG+u5InnoQmFi/6YZUEjB5q+bKCapol7CqGOCy6td04JN12vvkogyVWZ+6pd
cEDu95SXHpzWWkF6tbCY3ghiBrgG8+imZJbG1rEWTCSRn0XhEa7wlDmYVYvccpPvCjQ71Fo7gL+4
DYINOT9BizK69ruEmZHI9Wx+zJ2EY94fU9NDTz5zkSb7Ew4xMpbnAjSOYdswYQrMl+HUqaw2tfx2
/xVuJTARv7f791UoZ7ecf5C5v7naqMg+z7ZUJO09WYbWmhKQ0y6Sak/9Mw7PsFeeAUbxkTfU9AD7
2g3Im62j2jhbZ+SIs+SNZDCX6VUMdaiFXBpAu8rcjHMCv+ac4iqrfAcwC3nbqP+djEAwjCK/Ukg6
KVgq4hOb46jOgprcFOWljVK1XIS1rASG9bV4Anyx44jaw0DryUkDq/Zd4+7ILESoarfOcRXCh0Ta
08wuEjpJycn57XM1O/+NtbQOmzFmyb8k9Wi8ayIVXiThO+Ox1MXwD1cgyFpNRp8dE5UZdSN7cng8
iaRTFu/3tEFBdP9pP9A15NSZahnHEL7PLhpSDgtDcRUCKicf/VQ+OOhB2d9qbddeF3ES4hReHuiV
N5vg/26nmrmfI58jLFHvXISy8xqNmIHIs1zSx6t2jGhiE9L9MTbRaE6Z4YSRqbdsHpTqi/KeiVlc
eKJYzLTO3CzeMDru3losy60VANM28nLrcn8CKUSeN39PRb4+a2PliLx7jewSfBAP50qn5XEzHdG8
JYun1Ckw/6lh6EbVR9v1eyVAuFbRWbF0ljdsFXjMXiLPlOoirViLmVg53NrcpRWOGcc39k+0hxRu
3g/+smNeOGTubrHgBda+tKZvojh9ouH+aNzGFBpMOAG2NEzKQcGFvNRnmiwfGEm4jNHTgLofvPa4
2DgmeLmMewNivEOsSond9c2sXo2rvkCU5HXnUIr8t8gn9eT2zMfXONQyiNQhBXpqsR3RQcQhU4or
jbawWWpoKv29VgGcyyvdQnM5Rj7yfoo9qL9tNWQFRcX6MCKYpbua3A6SVeXhyeQTliWZ7MqytGoW
jN3b0MAm4gOmcRUDSeOk/1jTLkhIKvnKc6PSHuCdVzdqLQV/l3OIuWkWtp5UkyFpVBAefWzn+ygM
Vc2ITybVsSuWX3581Of6nyNlZ+NoYWybnoJ9rjLLDff8eQuu5C3LpSi/mTX/eEg2sJoYPwrVDyMT
QV0vg1FQ8KNYi7FluDQXg27dvKt9iRjvwVSNyNl3m1+uPPJc3UrbSMpdJi2G6v6X9fZjkdZM9R2A
qjx2CPd3pfxJ3dbTtND0BK6KtAiSVTfuFLpx2gRwhFqoXLbW6QyFJtHKRTeTyOkRdwLxGwUjOSxM
icTxtnCc0nejdZBnR4mAA71+h9RXoJmAkQ5xyIreVXFV35uQQF5GvxmMcBGlmkQLypgjQmXpe+p6
wveL9r76hLWRM3CxMXIERwGnQ+APZCqo29YYw8VNTl3DJWkI9cTMB23BLP4deBWRY1zwrGNR5Q18
SZkrg12vG7DmN2NcGhUaim94ZcSO1JkmKM9qfEbdZEtOWafYv1MzCPt/CjmlTlg7jCme2+6UlyLf
moi7dwxgG3oiVPAR3bcQ6cNL6C1e1GLJrFPt8YORxSX/WtlIfcWk6x6O0M6U97VZCCC/CEMp6Dct
igNTQJT5zSrJqD/3BYhLeQVAEHuhHVIjUEDnodz8UlfTHO805Nxtx+wC/1NapKh2zB9nWNKwwRXr
xGaDdviIUIeSoQfXqe8mwfJv6JT+1XMR3KiwA2W4vhi492aPjYVrmRkun9BHr+YdAA6Y4+opTqHu
O9iiF6sXpQDrTGpYoxSixA5J3X6/4xqoySjIBDYMlOC02VvYN2hqHDyCi7bBNe76ssdQxJklAzbR
EEsW2zXl/vTbWvyMRGEih642qrQVsnxs0g8G/AyXv8dJb9pBi8KAH+ZCPZSbnVBFfInLJgLYyr6R
Qxu8kpuflAd3L6tXbLhAC0jED+RuuKuJL7wc9xcY4K3ZAWoUFZEP4CVAmnNVn3nL5BFSbA06Yzh3
AstjAi2ml9vadNBDwyZt2Yk6iErwdidxHZqmsl+fT4x7gndvG5WkAZr7v9KJ5kQDXBXZzjE9Yiae
iHuseay2+H0uJiLpGc7DxlSJKCYbxW0Pk3iUYkHS3VnaNahTri0nFPyupsdhFFBBF/B7s1/btP8E
VoSux7G3SOAZEqvP7jSMslLLNC7HCZlONWKHAaOn2yOoWeyI+Xusp19QoHTRhq03Fo4QM6WCPSXZ
2YlTB5sql1CjrNYG4vK3uvM1jz5TTvbBlNREt9Rh3/Dp+39Q9wSFGrs9eFTbTRpDb+CAtBeusTyM
BaszM5/14EMEAf2WNinj94cSgforv5dHgjDB0pgQJIYoPD9b9YIoatkKXNaj1MXhaXuKJNpP79Sn
/JhEtevkChiYwZSIa3OQs9IGSdHUzh3gyvtn3NQ1Vs5Mfyx+g2x2Zzo10twDYIyGOHRGEKPIowB6
zmtjpChp5g7o8ina1YhquEZclIfZcR35UBjMvRnm0XB8pbnd2YCzAIa9oT6pZ2K2jGMzzHg6kb27
O5rN11iX0QHOASAcelV2zw0P9BJuwSlR7Gl39dZJdCthyZU4/2puiF5c7qL5ERSqCIO72cxNrJi4
5fFwtOwuRBwxvUdW3NuKDlMW+NUSMOc6EOEDUQJRfM9fr6TRrEWtS1LWQUh7wALy46BvkyXjtNp1
fRjftuL6AFNsCuHgzqPsY6A/J6J9pIMIk7IcRM0K6AL2Y3Ojb3kx2BmxGMwa03f0eVBIDoiHmgPJ
95GrWRbj6WnDcG8gTCDasYnt5WF/QXDZvJKNyywfL5F8+ddCupt7cIGG24yL9wSJ6+khBTeqEozy
0letgBLjZKqGduBK4pYSrJ2MXJ3ZztZGGSMcG4veXf2vZ3Pce/qVDvisZmImxnDAx2QYbtk5HAnw
v2V90e/eHZQloh4U46h7DaqrnQwPSVBvJDp4/EFXnuKhUEPLHov0P5OXjfCRFUPcCRWIMvXKMSbN
A9mCb5yRyQ0QCDSy/a2ktHazqj5qqSw8LHeWhVhk2BoBWqsCREvjcS1FlpxKz4SZqOQfsLqU5NAt
OPJWBT/fNcJ3HmUi690TsbXPNhJSu+OIW3oZTrtNOXHiyFbUXSTNYVNUBW89PdVQFbj1n8dIiLew
NACpuS+lTaUMvSHjREf9C5KSsV7jXUuo73cr4Lq8gXnnIgezYVYSN7XFXj9UphiaXvbKV/bQY0a1
aF6GwipE7RZlDT7f/vR/f1I+BqkGTNme1bWHPwPM9Q7r6KKW8xqD0u4nQ6UD4txC/BCLGEC/h8kb
fLYbsEXhLUpCt9gOJpotx34F96ThxMlsHcBx48zN7ZTo6plkn5zkFkl0XIjcQab4cpwei6FWj6MV
nSFj4jiq3LN2niTVLMAJXQLaGdPGDiUWsivSi+SOsLGBzMDAlrE/f5pWBfUdcd3xbmXpbu9Z09Gn
LKx2AMH9rfDuz78mxMaRiHJKfzYWAUw99eSkiBCbYaQxcN8P4sLynbxNOrhaww4WMkO3ZrNbMJyA
MqW623VCZtPVaaUJsXB8RDBoSeFoKFtm5gWOo0X985zJlJeiWCaLa8XnZqwMJR3UWEvgndnBjYiX
ky5BwUGnYKMO4Z7dIu7e2cW7ErekVHqYtBUEJG5JYdGuG6qamvHmdhLUEvzTPIH9ex4QhMfxu1W3
EAr1gwq8/xO/nvLGO2vJwObg18zwQbGEld3OKdZBjT/34CCwhIx41PHizNqmKwqYB5M74dZA/j0g
WGTBbX3kQ5gcbgS25F2X5+dfTEFhqUFhIxLNdiHleQSOspWmnX69YfAzXnfeYudIKvfJXuQRss7C
jRzSqf2HkT93ZuMc5RmYCuuHHtf71uPA0znfA29FW9hJxKX+DXtv34EQMebk9Ih82DzS/JHvfR0e
pQikSI9dNm8Tn0FKSzdgNtFI0Rjw/bLXfDi2B33x8y5xsFILiSppJgJXEcJ8OpBuwtfqlDFC5Ab1
4Y9wfIWvYaQNyMAoNHYk9VJdwrdhV3KBxt3Bnry36vBGQsGsQuAtxcaBUOUlhcnCb6qdaBiGl23W
nXFl+WC0g/KiQjWvFmJEs8+yTA28mjtf2q5E0gIJtKe3xNIMzDupjUwF2yHgiHdLItqc9avjTHoD
khNCN5OKTN8MjldpqUr+jeO4Egk3pAB14jv/FF71TlRue0fqpkQcvSc32YyQmTmKmZsd8eQdCKC6
I7ztEHAl+v9mRsLw/pufm/kh0ZF4kBT56Gjb1kVB8qOBRfJ+rlI1/EmG0xUF3e7+0CpiuJCyS2O+
WQ2mBxGXkr/qmBYat9iih8tI0x8grswmbzeNgFAFiEyUp3U6Me4NMbIZ5NTB+U+zDninHOyeSpIa
l5rcc2GSm/IpOu9fEFBnUmKVoaSVu9Gtr0/Y9gV/Rlxw68P1r/NKlLPO2ZECWyhtgDIdbbd/nkXA
k/w3B6fgNPGE0IbBkcvsm0nSZXqlD+A3gBFyKpmkNa3Po5p35Lix/PW0UuHd3gSmepieXjnPptWm
FWawmOdp5ybTc4hePHt5oP9aK4ZFvnayXPvBcAF9m/AUylALHfapmFSbKJqqUB3Of8Nsj7Ip/yTh
DvQ6IvTtWlFxYCUlnSR1fB5l84SkSx2MNDCwZIltJxpmX9raaN98vPIJU6fMub0qD/Ln+ACl26/l
Yjof70x59AsImw04iDEuqt0n5MHB76iGdt2AGO4LlxL/ktMbOiGosZa4dsnMZWaUyZnINUY+p73M
mUpC/4MZsjr1YT+pckLjRhjwHwF0IYI6XOKe0X55lfJuisGz2SLFw5GMK6oSJZxktKM3W9VrA+hR
FKyFI4m9TeDQYvzHw06bnUrSJvvpRA6hScHHGqZAtx1/XtElqH1MEnnC7PNxRWcx3Qbyw2OVb9te
dFb8uQr/MFtZypTqcweb3Sa3fzd/VXF8LXUHoMbbpgngJ9rUt4QZsaGR8vdzpIVGdNE2utnEy1Y3
5hFIdAHkSNRQyLINO5/RyeDOPGclqIC9QXwxk6ZZ7cUICLs2E3ZyyaTG9VVAt+lRheR+ir8GNR4u
Wro8Fg/rIwDK24pZsZxdn6RhqU7KH5t+wGSoeK8X8+u7fYwcFfLnS6VhHTaCUUz2wM/i329xddAm
DVEuGvKjLOkhs2uG0XAO0IDaqiRra+SLQ9pIkBjjpFq15iG5vG1a9LDlFAS7wIBiVvpdgZ7aarp2
gIlE8+dRt06ffUn0Kvx2ohDg5PC7yy4MSN7uZas68vrN8n3Osx6MdNgH+M864zx9x+yWNUelokP0
v/hZ86rj5a/dhZYxag3CxiyK8HqJW5vjDNBx2sO5IuWlC/HLukvMh782Uqr9U3QHeZtu19IQqWdF
GVunIf7GjhzQB+hSEk7fSvlWg9xkhbQTZz8gz/y50BZZLQEZHtqql9enotKX0xSL+8dJdhMyGaY4
vcBhv6ud/0wADhykE2wCPssGCdQMf5XkawJONnveAgJXaB1nwmjY3w64L33XRjf2/1LPKWmGtJXD
RMS2UVnWdldcgINl/LX2Yl5ZeIzKvrIk48Mz4w==
`protect end_protected
