`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BIkOYTQQJ3S/pgAtRdTaDU7YlCnll1e2gss8C4h0Ia+6M/R/aWbvgbdVBVPdiLAgI1yMsFS1ZNmb
VFrXeFQxXA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gksw9Pu0Fhkmgh5VyQzElsTTU7aoPhuAmt+2errmBFSicX7yhlv71ZQHp4/I5JpApWeH/6FFw5D6
b7b40oKkEUtggaqJnqHiJhjcQF2TYS32ghLkLvbIH585hJJzu0kIi+LkV9Z55VjgCMWVkAVfz+Eo
glrtfQLo5OC9eEkUlSI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j+u4GtaADVWJUaqtrPd/w/jiHJYMpeLS6xFVWXRn4hd8zIOucRBlSvM3xmnVjcEAsYtmKdKYGQfL
Bq1Qq4BwaiPCSXtWasXx59aVgla1Qu8ziLNMcbTH7z1hGvfE8gOb8pTCMdKv0cuasviEXFPaBIyF
n+F0Z94kEF74M5lQq0kJQbQw0GHU1drSR5ScYorkOqiDKrTBAQnzYWNL6aWDzAFR7loL1ohqwyxf
VEQZPuYQiFgf7l83x/wAnQ3S7tMSIfSrej/ly86xQ+jRF+LnKUHdEJUjYOSzzcmKm8ieBiXbcNL3
2CGZcy21wxYnPNFC2uJbyRqMzpdeTKLRvTPkkw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dhCIl6NIF7D9YeGF5BTG99xCVebE4c1ugGsJijjceXDLdE7S22j0eFnsTufYIVg7gfbLPnzdZcUU
Zizc2buFV2us71VpNF4qrOrInJBBzngOjfJ1fTNJUK9xYsSbYZSTs1TSyJpGo9PZ8chlBn2bZy+G
2pTd90gW6oV3Rxxdzbg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sWfEbE+FP0UJh3N6Cb8BpO+Y86VRcazogKX5612005R0lWrS3h4d9fw0K1gBeclv9u3BTSs65C64
ICyBEkroR9COVl8TZTq8OnxhNAOUStdY0ldCcAYdR1jf8oCzy2NSVW4l4dvjOw7rax8QD0ip29F5
SZgdzT7r2u1q5lzvC0+Z2a4aeCsx2smNkQvE6otVSGNa+5j5WZ18rqOwHk835ELoF7fFlCDQF59h
WpPqONdl8jKbKmKeTUeEyR+MNe3ii33k8fRed0A2krr5+JoIHmfSTeHhVaA5fNqu8BJCN6jNjWGd
mWtCA28dc4zYppTcA18mJI5PL9DWbHyAa2UXxg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87504)
`protect data_block
RoSnmiM7Trom+0ffqQiEgyrN0kpfnN4zSQ7rFrKph9i1YAs7EpIFh88P5OWq/9CsOi/E5R5TVPsJ
Xr8sd08eyjry3qNb9LRwIlczEdagGbQ1OcgyxfNC8h8e1uq4Aj0FuiPWbRxRQmKHPT4Acn9Zu+0q
+uYpIxcMSHoj1RGkxBQaRdeWO7xY4LE9zdGWuGl9kVboolntrPNu0XdOTtxbrWMHnS8Y8jBDNq3D
SXgSSwbduAVAEAmGv3UA3QCnzHWhsu4JQYYbFQDaeXodvXcRJdmQNGqjfsj4DNy8Gqs+gWtGv3wa
vjRmfjl8SmB0NHeInDRzaa6DAXuSqPI86mSozlRfgnYPj+m2dgEr1p0C+d2J26Tvhi5BdvODNKe4
rna+2Ou3ZlwCmHnKmILWJxS4C64em4erG0mNpry2812hoV0WAWIuvygAxrlTiibG+HiSAiOCE+fM
wPzddjzTqux6Fr7qCoF0imQnfUwem1GTPWQAL0asz8IUIPs7mH3migiRLJAYViHomqt9IYucPgMv
/xx69k1b/5XaIs1dm6QRnpzbqSkHVWl05uRbuvvL1K0uXY1KFtEixW5RWnbCxDoZvYPYoJXii309
IeWhuznPzDybGpEji4gzUPuIArdLayX0VtZvtSjFlKJiJmhUcIzP0Z/ydIFmcUh9I34uZ3+GVIIw
X7RsTtKhfOMuDa8KNbGKAkcq8L8sMw0sM7Tf7a1TOIW1JsdOUoMGUxjHjaD8gdBh4D32+KYigH8j
8nM3Qieg32IZQ804TlxU2NrlYAPD0VplQtjYPI++KxyV52FhSzHY7Ae2NvNBTetkrMQNb7xRHnuZ
J5ZmocPDUkYQScQ93+tXhjUoo50siCEI4iNGQEzjWO6PRVYpaMbucYlJkD6Zg9PVINygTyMax3Be
cJhIufBBMcV9SX1uBK14tQEdjttpTC9msNJaD1Wd34rJ4OV2O4oTUQY2w8scHbC58MxmjAMnSGRd
94fa4g7FfCxDqeCJWd4g2AULBVVf2hE3nu1+xvND2dHb4fAqr3j5f+PirVILyV8WgA4tybTzbTqj
jphRjPwuKyYYUsF8QfROF7vHbid0qs02oFBRVHDQu1AtWWNDzh6TT7XpHXYYob5AinVZrZF79ixP
s6fTYVvx+1C6ji7yHDVoyHxiNJYSWh8sgu26oqs5kqpHAU6OMBhQB7ektaHjOfz7IfCHqThiZ4r7
h+WGNRo1RsC2VCPRVFBLUZinablsVrB/Ff0stytv2v0am5D1k571E7R8UA/4plcyP4m+eK7Tyasn
5lQMIKDwi2qwVPcyPBn7MVkc+KEuH+aG82/vPAVns84QHpyMhP/wBCUzZLrhT+Zs2Tfv/7PWj3d9
zb5i+OPaCX5ZkASPA7/YwFRdZKjrgtX3jR1hUHbfQnsTVl2K04yPOwpSiP/VTJfZrrer35mCu8xk
XxixIdkEpiPpW7FGRtRaeV2276VGqZPnmNZGzfIm8hCGHWmFkaavX5gBJiLuGAc+S0JfJnx3ZpH1
EaHBI1dB8djdHq8hu+y3ttndWwMXZwAFHxkxy2em1rj6rh0JmlvqGNFbfib86yWgfvzkcnE7yQze
YXO4Y2GuZ2VTnMrZ97OxgLixwMyxCkJ5xTCLA9jF6WciKxjHZkerXVpXZMEF0sOGhVsY8wrqyK6Y
f9RY+RGHpvTfqY+CSIKrb9/2/t64C11ail8gjNrvBO+P0TLOu8/CDhFT2ruQDWZ6Sm/YF/ULuqmn
52BZjeButwomuONo2cn8MQS9NhuLqQlBA4V2oVBQmmk5APF0Q+WC7w46Rz2u7s9uVi5ICZ0tJM5Z
EOWGEdNUj8LRZZsWr5oB4nH6pnzcw0euaCPSMaZKStIN6p6mjhdrF3pjwa7WkazUv+BZLvH38oCB
ys7vhW2qoWp7nkZouHaeIJpWdMo/Oljxc8RULvFjaedPdMrQ6ndfPj/hw62Lk6y8FAP0Lv0OwHNy
xISk9+lhNI/Z31BsdqxSycjD4oyVMiSH1j0PYBizcQon4kLibV9PiKKZfA1L6G8ojoaaQ6Adx97z
H44hxSrQPd80MRbdOJykGctty6617ubUc7qAw73FZ3GlbhJwcQPaSediIM0wU1kD3zohFbBfa192
+tF+KoWA7M0c867HIGUmODSilUYtQrMS1v3rRMboAZGTRp1q5ZpZttBoX1oTtw89INPhk5RuGZs0
yPIFQ7Dn5iPvvWj2EOZZ1GhKQDZjRp6jjY0+x6JHg7CSaapGxXBxVBe5dKFUpOIVC+7pKSJ2X9bX
FetgiJ4ahi8ziJ9YfmhZulq/Hq56GHDh017YENoncvQDAksAVg56YqmYKPMA2eZu3ZyV5yEuaAS2
ahu6IAhVpHWon//4cJt2TwDRaWG8NpFbS4BG0FMinwU2M8ESnu/PF9cqralR4cEja39R7OulKwJI
xajRxa5IoBO1t7daMAsDNCuOEWxNGntjVZKCMqjTuJdyjiXQqQvD8N/swbnh6cAFhkUCNHVpL3La
8aP6vieczAmUXNyTta4ev2o2fCBM41KFrbeKqSb1bcHHl7hlyIePXxgh1tffY6f3Z0Fz33Xbqk2o
sv87QoqYyUoKDZqehz90UxHBkbIhjoa44PtTWEU35rUF/CwSujRi1e8XfBtyg8H1w3a4rf/6znCU
QyDPVR85Eew/jGW4BxBtb3w1Nm9HMAhcoG0U7gELCW9A/hTmJI9RQQEr3v79J2zqrLBC/T5dNuTC
gJVrQsAmmE7OJljb0vOcWStjPrmphUmmED4KglML9c9ya6yTQw0IdxSFS38NYbQIQ8qx4G1uTn47
DKPEHjvmInxixhL+4huzstRhTSH6jBtrdv8rXCTBCOV5hK3Gl7HzrMQqK4ECz3TE8AgJ6sRW1o60
i75z+SrM/e7pGuBhA1ohb/2nM0IdRvEmJiMQ+JNPrf3niuG8mYb4iPpxcHThhOTAhSpq4RlumO/N
o4Cr3q0S6NfdLmbiP5nPQNnznsRwml4alyu3229g/BaXpTxLq5NimjN41G43WQtQ47ugqvBnoNwf
CauUM40bBaYTfiqI3XgXLjaBepxU4QtITWY0kFR2KkTdS8KdVS3YtDQwADSkhb5tfm0RqSiOv9gy
sLo46idW0+IxvOiXx/GRhr8WeASrXjevILTWJ1ba/0YEXlngm3rg518LotZ8KDMOVVX8bc5aG5Z7
yVXK7fDX42b0tFrXdqu0z55SOJa2o/gL6jSREkUYkfOP3cD1m419Y0bzM407CTelScHGRtUsgsPB
lbiku7apUAg4hIhDmo9A4zvHyIXpptA29icSE16UXY6/5GkeE/mZFxJNXuaiZO0yn3GJJPA792QA
7xawFuKTG4xYzr9W7vkkXu8XcG2lghPIPhN5z37QsGbaiFw65REbeSQkDWpxq2sgMH2M/tZ8PWND
YbuWK4g/E5fAs6gvsPCTKxx6i2ZxsQz4a400nYhsCHi8tYLILU/wkd1EpNDdi5zz0gnMJDz7Fry7
i2+QTrO0yFuM4PV1oTh9OfYkoaU/fwlKuyouj+dNo+2nPJfKdMUKpa+8gwPfZrK5cNGkA22b1AHj
q96SgIGsBQrDDs37udC6bz92q+BBz/RoOmisv/BNzQxUsJtGNVXOAbtaMBehQjyOCNCLUUv8e9/3
VJzgvR3ck9L/s+JjAi8S+P7KXo0FCXfYEUbgp+t1pEVSHrIfacU1Q5lEGCAcGJQcEAQD9LdYDIP+
gQlXDXojh0J0uuAk6gkGRDuDHKx4CvGlEO6l4FexVzVbNYZtQrLnwWcgjusRxbcwnORcTuaot+Ej
uiMvSTRAPxWfqxsjYrC2bsVhXPW6hn8/VpWYg8js4yVtuE/gBhXD1xe37kIooAL6+KGflbT8eo80
PyTa188rcJ6XaNhUgdTrtKjrsT+6fpj0FubCnIiiJqLtdx5gRPLvESdMAp5kZEt9wGVFYen8Tt2I
y4LG6zKD5FYk3ZMFPj9hRse8ZMAz5kS1LaVgt/h5WMTIel44XUdZ3syLYgwGXGhY/agd6BicR5d2
UzcIeLKeGmHNQYVkEFxyhZRi+swFr/QUfJ5N5igAJZu88pEPJlOXwrfKwPecZz8zrcdAJyXeS3Bn
PUAoVQf74Dls6Sq4KFnsVrYnqyQ6MwWBYRarxQ1y9cVRcME+whvYdGVoAG+xh0dokfmWPxLzjMIj
wbil29nR1MTtvjpXU4L9FO/iSajgC7dcaqSSYEDWMW2vRJrzGx4lWYIR8SzFDY+Xk3YaOu9F2Ffa
ir/HiqPUY3xnRAb9mpRLhTbjLw2AKflXSmS/qrlQSbveNwVhVGdmdtRQ1NZp/KmT0bYKaT3ys+9j
w4Vs0BnBd4u5Hxib3WePlSejkntpKCn+TZcyD4705sX4rhXuVZNgokfCE7v/zegp4yk/TeWGsPMq
Yq+lCrLqlS9Oh/DE8mHc/xM5fqjcUA3V+PUiTQZyLU6nnMKnDGgxVinV2QgZS2Sr8l/M4gudsLrL
COqis/UN+iSXNK7cXdgpJYtxBgAukR1692qO5XsDrLbwph33BykAsD0m2RB6UPE4NHy99cMxCj6L
jqxbOGRWlyoM+ZA5xo6Soswr6f3QiRjCMtTm25YxmGcJeU/1eHKLsIQILsGC0BohGsVgqy+hmGb1
SyRtYVm1idA6uKwmYapuV9X3Qz/I6Qvm6ng0FQvcFQT0e0RZxULEBtuSCcKknkNi9HZ975T/9HW5
vDvicdTEgbXz54zcEzN4k9g3reN8GV9msMoZHgngrW25K8D6n6bQZwS1aqqOgi/50Ekn0BDtHYYv
sidtRXUCIDS6TLTfJ0rTqzqWxk/EYjuObxvIwK+GGqZLb3huenQosSR63vCpF/ydvdt6xergJsjL
nEEB9h7cey5gWYJR1kOVeWrGtnqRCap9OsSTwcX3wrh+RlEoFGRR9lMJmK/qpHexnCVT7VHGspLM
1eCu1Z6BCmooC8zIEz6XaOsJBmsAMa5bVTTQYY1PHYxhWK/qWnSC3LUN9O2b/iOmnZdJDhVMQeyo
y8+/vOmoAhewvdAuDHRVZKgYjc058E96Y+WrPygqmlQZw0+MBx39Jw6ZUO/5TMjq6C/qeEWaPiIN
7L0EU/pG7y3hTiR3o/VaNXHBm2Xd8FBWD3Yz3VyWN7HBHV15ghA+6D1onrjj4f505Zq2nzxwmvXk
SB5TNYrcT2OND0dtkf+bLWbfdQ8iD6DSJ4W6pMlwqcS+ivWqU7cudTYvwijuKkH7/Tv2OzsJiCel
abbZbGODCxWiu4VT66DOXDPpclQ2aC+S8an96drrYDwF3JrxonI3zJVuPD6UYs41v1L319Bk1vUI
balc0cfzYkVPyMFPEaGvPW4F17IrqZ5lcNHTXPX08h7fo6r642IteQlouYvNft2yMSfztHeijLi7
c5UQ3uXrNdh0CD6E3SorrmyDrKvn7lLIJ8tpNOEEbM+tsRPLieszuqMcxV0xRVFV57/7vprPz9eq
C+CMtx0+16/id25712nCJfS+q8EYQFWHxVOZ9P5wSk/IaJW1YUP4sd6PTDEHx/F5TVzYNsxk0DZa
WSvX3uSCYWvdwgagbJvfdpPaOkBPv9NneUhbwEnF8M6zZ4+mNTyqZrH/rCZeDdq4gwMuN3hEHGzg
Z6H7Y3bQ1LYVHM2BkTdWIDaAL6bgqi65EGfuAebPG43ycq2UunYe+4kL6Lp8zYzLC41hnQkzG/z/
zvxsxNEehylfeB0Ez9pwFk7Ey6ZTgfzB24je3vvPsiziHCgXsbm3Zksy/Oe7ZUWg/BSJ+LV8+ytE
AJFgh+Z1DDFlS0p3xzVPI/3qhUpRjSdqisxC6hM1EGBZPLmT5HvyNERfRVD+K+rRJRYV0W7Enyfg
6LPCQK1E2FrXjZz2ClGk84O8cTXs5tiAFmYgqB1grbDS3M1P6ivm1fechGRkLbVI+o+bIqBNfFuY
TBOPf4gC9mzYQTmtOFFBFYeRZJEvI+FtN3ErxlojpOdJkVBbQEiFIV5gY/Sxl8bLRFTiuOU/eKpE
OBE+21P05snXZO9epj71fLVTtmuwWmgk1E5kQg9JQ0tCeT+YzNCzYpxIG2J1xnFg9+27/M8dAxu/
+NeGoL+rJxJFKpsGUS2Ug6BNPkHy8UYKQKi0ZXRu/KqZmJhaf72/bB5YOO0aDNCitRSQ98hWVoy5
M2flDfsWWTuOMVLhiNeHDeU3D0eGOh9OZpPNMIKxNO6CmpzmeBx8jnCf0Tr7zl4txHXGLcKnT8WB
bMZhn86ftWNTUtgmds3jQCVmBudw+Cb+b3GQzwQ+P4OYv1t3gLH52om16XYwgK9bJulSzJtoBY87
Zrb3gNE7f4HPfFIxYYdlr+yeqT5srjTTuwNqV09dQpjGOP/J22HyD/xRqdt+gy4FTkgOfyR6I7cW
TyiiG8btLK6O+Pa+dSSkaog2co7qwV2qJUs3ppvbOAbv7bYmTsTGw++P1kh50XWxyYfkLomddZli
zmTm0qYNtJZ4t0gXFRrzcgNyJXIEV2e0+DE9ipS3rW/YV10YMolEmkybjXH/Kc7hs8WoQtVz2AQp
NYQYLC1SYYtdel3eFuWpk4dTfRNfyL3fEzxLSL8RG9yn0EOtI2H7BwlzKFNFRDIA9BCZOXs8OkG2
Jj8KTzr7awvN6AgwOz4MO2xOOrS6nG7IdEsdyeUq/n+0omFLwr2y8qQev/yUvTqJd+DZCgh6k7an
oQuWfYboF0kLdyE5tU27/ZW6PcZH6KAEB2pIK+CLAUaXPKN1QhfW2CqojldOxlfqpL4IPkVr1x9f
JKZ8YKzL2X8nXEqFR2BZT3SdTuve+r4q7e4gIxBKpWoZNm9YCOlHoT2+rwqK7aNSY/oIaygqtq6y
b/DesArD/TKvz14xeAeVN5msU/ZhsD/MBu7LfHzVQDnJxaR5yt9Pb2Ovpe99Y2Yna4hDu80VwOTp
el8hqOtEkphm6kK1i0PJNCu2lJvbwOA9jaG1EZKjCc73DujdHTgCikE/bM3xPlkaqgMuqlQ+9qFM
Dgft1qY5SLuVM5edQifiYaTjQ49JHVpX2QVxosxN+i/MZ38mQPCnorlTZKC+kpH6ihe95uVDW3F5
TUGpcsN3KZ1nFXXSDqnS7GDp5Khp0wg+XF6UEh/6298h0HzJd3Wf0yK6CI/z8NvjBkVuYvpFYCn/
BfSdyTjBqXE7mRpuNohSdZKlOsqd458hWs9LkWbWTEK6JDAVFf29Q/Gobrnuoh4Y1+W19PLsjQyC
wtCfhS8j6A2K4AQHlqKWBolfMdhd9eXS+tolgfFWJK2xvVXW+IvuxTpmZwDw/EP6lV/LxeLhhxoQ
v4Iwmytvo4zg5kMIWDtA9to7tZwAgW4IbXU6IYtsllgOBQNatimumyJaJkb6veinW9cWxtUJZSp1
8E6lG5/bWev4PqNoG5jWDOtv+xSSgZppVhHuRHEiiKrh4Nsk8WwoGHEq21jkgKDCGQPuXUc0nw1x
YFiCn+Yzqx5dmeaaTqn8ubQGLKrsiBd/352lCkbhF7E8oY/bW3+cyqnegqomcU1dJwP/y1bDV137
0Ie7aZ0kohHg5RPLrlDsFucl4XYWhthU2MfGcysEJQrXhIThmH7Yfs7JmaG7fMJ00/9y5sKh9OgU
mU7lvuvyCOG8SH8Ep/PlDraIjPXJaTD4V7TrXduQYmftOW/skF2WUafkGlb5zMC3wy01zgsA1LmJ
G0AvNcbPgQNHzgxhyJBpeYb6cznrRyO/qFkQpI8omvk+yBRpD0SatxHUlhovFWzyrnr8mZOKSBjU
6retCosrd2pM4tt19toNS3mNM9zlyZGoPcR9M+K58TT8ImU7rS9ld26ydzZOzYXrSFXOCLsfRiEE
OxXXwcxXIHaZOrhW1iJbZ7gdGM+SLPAPMOAme9m7f9g1N5QAoIgyF197GCCtBOgArmpOuX6riKmC
5IqrlxJqxAz0z0yGwd0H1eCpm46AIgtNDUEwEpopMhqmea0AYQV+cKEcQefr8vMMGsubJc9cyKle
AFlBJCAeBHD/1OqYqwKWN2rTN14M1H+4Eg63QrLSVoWp3KgmHB65GFIQ/KD3NqBJSl/YGzJLg83Q
LvIubm2dhO/o/i5ZT1ZiY3O9TuwY/V9lGf98/df9nbmlOWVHPPgBsD9cucMAWcD4PYA7/omgHc9H
2Z6Ty+wLaIH3+yPgMmeebEs+uBkFfuOKsAzsSJwGAz5hAw2LVYRDoSJoly9/i1GGXnbbF0Iv33De
PDI4KeESZTWaDsCC9BoYhMbdojXkqoGL6WX4bdybk3mGcpHJTaFEBggEZouES0g9qsBi51QTsdGk
DapjyWXmJx+72+IxWq6PoAGL/+Ta7giTzIlf+GghZgf6zwjRi6jSontLZ1z46j7O4SvCuwmkLgCb
nl5sv+WhkU1gmQo3FjyiSUb787QkoF3n5mZYGq4BN9255i+sm4uqcDYM7UTPDhGB5Dv5oJQvhE/J
cjA/GQUMN6fCOsDW+2IfESQzgtnBacO+5mWaDuX1SkDkDymksQG/Z1BFX+IOUjqLnIv+INd3rQ1y
wY6CeIGHx6BMqXbb/OQgw/hVOfPrHRYcXDlhkiWv2duePNtfG48frxLZ9KXmayNwcy8+P45jT32+
UcKDjXZEDpnUFDgRmx38GhpavE3Cr4LaENPdNzTiFRNq8beU0QapctlBi2mgApkASp9BcaxMNYST
crxYDfbCILcaheU9UTL1vBzbpCnTGyt8EpC/AT14qKYDP5st/g7u84IdstPk46BHTLgH9mF28MgK
uz59y7phjkfNiQnraAvmkEXa9wPIfQ6SMXBPFVx99eZJdX3IlYUL+TN7bl8XpcgPDxupDCHgLADZ
zjbyXBWg+6a9oguyux3LR48B/865elt1a1pyejKGHdO3LlAzFKUX+BWFMeG8NCvzo1P12LGe8LUZ
WNASR3cpQMRZHh0zt/Zp7QH7unQzlpcm5SbIon+3j8OuoUn360JPi5Srkjmt/0pn4sOGePKZGHmp
xx+St1BobXnPMwuPlhTgEIjt3roIMtNY5lHUn7Hr5U1JFVZc7EiXj/e0/ggC2JoT0Vitq/HbtHdh
cLAJZG6Yr4KstJSJLzeQvx3aw74OBpQ6TmETTew55sCInA/EgC3ZtB3iPs+VmNNxXTevvKyGDHLD
JWeuRsLjs/f6hnMM/sbc4mqWMD+nj813LP6MCoo6kK1sl0Q3t1JcEbHtMYy0EPFpn332+dRrCrwV
AsCi6OS+KcHqONbra2tpmSYZKs14dmKZnYvHwfwzeJqe6QKMuncq6BeTN60YZ+7pfm8AG/vZPCmk
yzRyC10HRLfSg1oleHgLHmuBM8g2cnScCsK6jJ9GB1x5AnfONHVPSWeUh4GVK5d4FbBi44qgEDnT
U03Gn7+W3pMou1azb6GwRePjoJEkyOgYR9alPRdr9wtqICddabiG9IR1hGiCbbo40yl0ILXjGWc8
WPhD8LxmQ1i/usfqcVd+4kJf0JRi2Ee4t64AMQTGoKYtKtdNC1jZytk2FxW8kGoATScb3QzdfQYp
K4ClLX3z4USaLZvk8oxGVHa/RSZHYmiCmKzWi3XAGuQzpAQMG2Oxc0HuBgpysUpgply+ReMbXYcP
Ns0q7CfQzqU7hTKVQVo1MOdfbjrhhL182Q3qYxD4R6T5V2Mpc9T4Y+DRKx6gDXERgFfvgnGCrghZ
FcwCMD1KlqU79U45NUo9w6ANDpNlLlG3vH9CnDy33dv+e+6u6fHPrfCgGxMafZZ8YTkFdaJtFZWT
Q1pQ+4GEz+NHQsRjph5u8e+N/Vm+xDQfcBGKCT/Z2GI9gVRaBCrL0cfB0NqD3za8QAtBS9hunj0W
neejBngevzI3BCfSWjTmT0mOhGZmpRELl4nVeiD4OADpPQvXA8fbTfpJvn+O5kK9aI7GTeRh6uOI
iGhh86efa9fA3nNCtArfjL3bUKjpC1TyMGljqF7Q3JV8oG0jwz6M5/Bb/GixixyoSghodDVqKXUN
Mbm61OpAWTh86j5CYSu9fEvgVfrtihSPkWDwHmgepxd+otsaPNXG4dKoOa9ubm/m7vYI4ek3I3ab
LVkwb/iG+eI/juQWBCUlDKI/wvhnp1x9e5vok4gl60mLznq9jRwOzn4dSzLuVfzJiBmQIxnaHq08
UcCjgNDdEBIiP6rngBX5pmJuLjH0gQxiN5hIrYiJMj5Xp1i1CDhd50cMOaG3OGg4bTYVy/2/3Pz7
IffURci+YcaWzfZ3NT6wqSveYQMoOM19bQ8T9ydQjwwFpBTfDciYvgMXP8Adk6FprfBQNbH41u67
nZ0yKGAhgPYUh3nognCPnCRCVxVgWWG2PXfhJ0+6p9tk2Puf6LxcddXEx2ui3NNzZD11gq59PIgz
UsEZTQ6jhdMJ9auAIc2rPcA15UdbfhojSMOPLWqLxF+sGo8t5kaGVJPOixvHOPv0wdroUjhHSlS5
hp21oOGGI8T/UuCxx8BB3RmBgYLXQBwdWUaLzZYSKLRwfJEEksdJtF/uXEWM2PsVjCePyTtPWSoo
K+z5CKzF4p/Rb7SjoMp35+5t+NEdzNUKFIxamPrY3UKHOKEX41nZ2m6DtyPzVMGQ+BzWFJdWfw79
QsYN12zFn4smFMw6XVsnyzHWsi9R9//ji/1J7AV+Ln+Ua5/HDnQleIaM8dra9Zvcan3XhlAIYMFU
Bl2Q8OFiHH+ztLnNJUGVK+hPH8R6QGgCFF+R7ZmtxxbGjkARdP4zDPt8BVByosTCHyGUelTSk/ve
GpKg1r3JfToLZJ2Qmg5aMjNzGMUpZKsO43QUq4syAj0z4/3x/kv4FZYJS969+anB8FO00FkwI+jg
Bcx9Zjv2QxT91ttiRPsNIPfczXdzdac1QjYkZgPVc1bv9iPUBSERPmSJ606w/ytadWetHjKLwMS2
5FCBWRjG3qFnFfFkHiR94YltUa0nZHOZwDqnHQqZDMaMkIw0jp4T9ouzLFxrdwewpgTmUMVebmu5
2j8XIKhjSsxu6oFRfHSuThvMhVUv/mXRsNy608XX4GraCloko7fb1o0OeGo3vG+/NhUpsfeQ/H8T
oM6WZznfCErWf3kwD6eye05ql601ii7kEpaZl1kNY2fpwRlFRk/TdR/PlUFuanUrRokR2WAob2xo
lox7yAXCBRlGsI3kwBZu1H2I4fnwxoPtAhdVau6p9WyHN2aE1Q6KBZFtBzuOP3z+CO0RKvmK/pLL
50/bmL++ZHY7ZFp1/BIJWb0qtIaoQRVZM5LDjWQjRetdHXHDJndWE8cpyygEZ3Hr6CdVqpvWxoux
3ADNijxZeth74ZCRoOMKLX8ObDOYOZ44nNBuDYy5yYSh2KYV1apj2vSywInPOJFafwzGCrt2Tl9z
GHehjb4Fl72TN6qVVS1+xrDhM7d9JDYZpo7pjSzxreQ75+LgVOiaV810KrGh6UIIKvGkRJqShmd3
TVxKuNEuzfAEHCeD7VDiE7gW70y9n4MzwxoNHyqCeC6NVoibWvIePe9LkTFswH9LVJ9292eLKe3S
N7uVcepINnT7u0zYRS2WV8/qFtQsKCh/HtKR02HJTu3EtcG19JMw/7vqEp1c2+irky3LJjjIlI2M
h5ayBDZ/P8vVTuLHjUjdnxOTB6a4z46WpuLF1ycPV2+XxnYCCSjbaDtusbE7b256ySENSFK8079A
N0/SqNRnBR+oAX9NDl/AFDchUIfnu+6YltpJm1Tey3vNI4a3LIGNOAipI9QrgXn/HJEOSjRpPFEJ
CpC/Noz+lPMbmlQUOd1+Ch/G1mcJmDs4WxlyXp0HCmfvQuQp9oAO8O7h7VRnJk5i9sry9Tg4oUru
Ab9oW8ZiXBFR0G/JizQNrIUUvmut3y40/V68zmhCu2igUqmgA9epkBYba6mpE9g0KYo4yfFB+BMz
cKpIXXQUotTBonEpPktuGm1y4uFxLR1LVs7LBJ4K6bn5aVgP14gy/3K9EYoZ+htuerMZ2/OgXWEC
0PjUlx0Qm7r6Xip0E7mJK23gJsG7tLLoRD92QF88D0wBeiwWn5SJpSdp0a0cLBJlpnD/2oCHV+Hr
CsutmCnh1SfVUDw7Tf0dzxeStJcwlQysTrjr9VydyCSXtmy+U/nxwUqBN5EtxZ+LmUqPjdgJizzb
TAjf7aFn3rABKq2E2xp4uBM5ivH8OHbQvmkWPxq2P0aRD5sJDiCcd9AaXXbxG3fViRdVUhQyVHJ7
OGGr25w5Uja+jG7aVwpayGd4sGNxGZ6pmVBNp8L7lbKRGXRQ19WCz6thuDE4SOuf1r1CptXyBEkp
GPhWd/muN9bryfdyR0Ywx7MfKqf89pIZ8GEbc5QPXkSFYV/YfTZCp+kCHpc/6kUBC1hC5ry305Gx
HEBlNuFzAK9cY6xETiEJszM+KellaHnnfWFEi7yLEseFtRwlMMPH8XAk6cpVwXwmZfb/otwBzVag
FTr7bR7P5o+kEFeMq1CKJMeg/qzppY/1Jv5ZD/UXqZMxE9XFY91sbXl1F2yuqsfMi9TAJ8gsDHU8
XmVou9EVB5PB2ptlKMcFq4LJoWaV5adluKBGQoCvK+JxkUl66LI4NbMiUvUEXiU+ytILN1Ypqm1a
cj7zlGBl3YQJzy13hiflokavA6t5cmYlFP7ZTF5HxvefVz0prGd+zqiAINbhzul3prN6RMDWpsgD
yJFRfJ3iij2UHN9UeAj/L8PDB0jN/RF5IoXpMEKLlDzKhA/pj9aDk7gQV6esrjEEzr8pzfF6vchX
14OIUMSSPRvjhI9qAQPOG//qqAEjVvEwLLf3zibaA3lYhu0wf6xF/CdPMGv74zhf0m2HQQxZXSIw
iphizVpmlWdhWehEYLC6SSjENLKtWJhFaVhLgReGFHdE8q0VxKkAD0aGCJvxYGA074thw1qIBgIT
uMbdf4lLSX2JFsrHQMhOPTg/aIRtGtIf8j2fLSfR8Lv5guu4/CNa0AXaSgvxTzDtoNuww8MGPo0X
ivsqe3ryLS7P8UbwxTPfvrjRmj3uQ+XkE6k5uvMmyMm+8YdcepgqkPkCttfpiSgGtC5uhPVuVJ1b
Iai4eSeFy3EvDhyvRo41RhLnpbFBBaE/Vh6j03ukz1m+tkoFmpQZe2vd4moCbv2llW+jU/smoVqj
xzlzV1DECMXrnvJkfJEf6aj8/b0BIoKPwCveEmSOjZkXa4MSSN7oocKrfDmVj/Yg61HEotugcWyS
t+MASANPpewk6126SWm+PfPsA0u5fLc8NArd2Ge7x0k+Ibkas3lVJn34K2Zv7Q/SlfMK0uG3kf2q
Q7PJ6T/KxpRmNyUoQF1d8H/c66u8jSnAfPEJRUPnhNf0jEpbl83HVJ/TptSwjNvY4sBuZQnQuAIn
TKPZcyJ1mVRLDCkFoJE2X5XxM0WLcyowUZTEiOiwmCZWsM55WHzPhT0h87b0gusWnFYU7yRZO7K1
EaGcBDoqxrcBKLVBRCrqTQEegw1JXRIGX2ERbf8LuOWeLkOVrR83YQ5vJ7A6rPktyQJUu4yajR8H
ocOqeyQYPIvzTk6cInFEBbi7DDC2buw6VJhcR0KMVyPPC2PjbqaI0l+DpkC57AvV9pTgxGRAtX1j
1WmtaS2gsYsOWjLaNcZoYXHyCFn9kI9ubwwUQpIfhpsZUZAqgTWT56uOC1M0nUip30y1CWDjP1BM
/x4M+ihCfBlFay9q+A55vIYZWvFjwdtTaQAAjU85H7nh3l2xz26k/o2fwbkCEwFbZYLOJdR9IjmO
sMk5whedTcD/lZLPKnUlptvbV5ZFL0ryn67Ll0pNHccimZmqZH9Mx7vMJk7WomXO9nv9gjxbUc5C
IfzvOjLwtphXQ4twMoI4ROQtdjwiSvYI9X0UUS4hqMMLnjgke4v8E6/QE1bs7Ha1rlOawkmoMBLO
zHyn3oVv0YRon+xWYorP0bbqSMZ5ow9vUJSH5TjBLh8vH23fKFYgNiUulCPtnmiIpAX4bNvWxAUR
CPIhCMQtalg34wqrDPo+w1bb0hDz+8Z+xkDJOaUwNq62A7+6oXvl9WCvnS4iJG/OW4pG23KYFv3H
c297/xgUsiomlqrqKzatK7rInPei8UuN+i9QVbItG8YfMTwRAFLJGTk3iuSvGjZmXH/p2xgo2hZQ
t2TCIhS82Wk8+ZcKKgMCZpql2lJNGAJRvZ/RLTy9EyO+1t2wCENFC3ViuveZl7cEYff8q0AgI+OT
RrbR7mFjgX014RZPL/xxgjO2/YHZ41UZ2jo5HPIVjqcYQt7nAT4Js9fmsUVbGsKbKMU9dm9IgXqB
wlOE2obbGzyGYpSD5F9SoixDLTlD+Zhe5gvKfjj3OG5CLChlrbJIkkABAj3lhiNJbqivBPA33HQb
zVki8q0IcSa1fTvbB5NqWXn3HX48LWqRsAAmxiwSPPAFiPoQjxsVlwfH76e7tHhQfoofDGM9B2uq
W8JLMiyuUvhL7D81KpB2+lNCPx5WFoUWdabryb/NyIReXXAc8T+ADGkafxc+wsi+dYxo8GSNEksC
HdQ/af1GvJpS8zsKNWotCAxEGURagGir1HWMf+oDqrJVQXbN8k6tNMlRudPJHAuzzUAg8II3Xsh9
tyXGNytVuyiHSqeXQQms1rPK/I30f05mYqgbsl0M/7cne8xPTH6/HZ9m6M1vPdKtuER3Ha75jJZF
SNd+UkGsvF6KRFVU1bjIrYBZ8JjMupcmpF3VThlJWWbzdLsbnLrPNkjjm3MV5WMR6AjP7n8gwpX4
9eo0v4uRcSZcrK5RwCSjfUQyLiRWB/j1nbx5NXr/Zk2S6bp8mZ1w9dz8l6RVXB6IzgXKiz3RVKSt
cfUnOK1ch878V9OctV7Lg5YxkvwCEnM6iMx8aTedkUnJkJTtwPoQmPbO9AcaU8Tfb8Fp8Rm71XTK
OwbG+el+lbok0lfPrvFItmcdf0DW8QvMPNvTHa0lcyXJ6ToQRlxo6tXFtodfdSd/DXm2j9qKQT55
1f+9R1hms7W6584N7ejSG4JbDGN/A5CxXsSzz7jv8d0KfE9okqV1JhtxX/wHV4UAjeOZr/rRp1hP
e3UpAugIj8OxpaeSoEFhwiTohZH3ukCmfkL0yfyAbS/FahXxumQeAcAYd33YRaxUmX1WKlQ0fTQt
OBAdvkZmMx0GQ2anUwuh2eC8gCmrB9HOodGSE7Zu5l0KPXMWI5IN4PcbIOktf4F3i5l4nev5U7p9
xiFhaVyWSh3RYxIdYZdsNAJLdkJ9D6Jo9WZthwGc+N3qdmvYnXCSEMe2qGrgppx6VG48Viw/oedz
/0mewvc1efSihldAccCUbaa2iIqnfrJe8h5Lp3iQBalRqXhyrwbrtJizW24bPfeeg5M6TiT8XukC
fQqQmdI1D3NYMnSZmcXBexl10EoyPHGLqQNumkT0IiezCQ00VUXvIHrhvJbgTGmNkREjDq53aA5U
Aju/vT0lch3ZnApzC07+1dkqyNeKeevrPfhKMfmAWX65gaAJ7pB3XLvCi4QHbNfDlw7e53lOD1Ev
vRdgl8aFMLQHb6LoslbCqAC2vnErLDT29h4cYC/5UnFN/5abuV/CoFy/lkdPEmG6U8bXyCrjHrEU
HxoGBg67NMHpt2yDIF/Sd9saykPOR+LxVjxMxd8G0IDvVrDy1D4JbZpQds/8MLE4xqT1N6EX0cGn
4ydT893S0e5KBWvndrEuHuw+JDDNhN9OV3W/MynqY9P1CxUulAsEHgUsBOZETei97uikVbslybr7
meW6uOMqJ1u1POCSGA6ayGLHsOqLpwU3vIiobeA58qilnHaAI6otI7N+aKlaraQbituRKPc0NefW
q2joamRFETTOR6YMaxwtJWVQQPEsWO9EXfpNrWCUFsAoM9mbg7tkiDp18BIE80jUg2c6PLieF5j2
G8LYop1ETknGKkDTa+RWPZM1CAUK3UaDTkNlrP1DlRlNAf5NmG2sWdBCyAjpCSSTUCwBiPud4Kmw
z3teHVZtmxeYdzW5eG19X4ayhZJOyrIwpO1h3EYmPZgOtn06dsmsEBMdGuUxQaXZ2vr4WAVKGx/Q
U1s9Y+LrZMLYQQa8Ag3WvekBqgMl6uvL4dPW+P6xzlE0tMMO3DrDUrCvHueNF4DK/6SgjntFV4Bd
bUQVYMZcCCHTpaNWZcf3eK7wav5a3y7T3bF1lWWQbJt+ISv5U39jXdlrKF+MDH7kk++MpTH8KV5z
HwSsMXfDuq9E15Dqg63vq5tu8Usb+9PvrG09gO7xoLGL2HOVox1GVDLY8ac42G/i/URIC49paMCX
8H/azxKDduPY05PE20s6qKeSmtCSlVA4Ux57+nnG3A6+T6OHoHrtj9tfYav/OMpPGK8FrV/zp9E9
Zv/vM80I4hlpRprAxiVD9W8DAobaQ6VV3fqS01bkJZo4NCa/bg3veF8AX3AiKlV65bpy9o2laLwh
oAMvzTL43Y3vtdvCC/NmS23XcVVNZisbNEPSWNN9YZsm90+Pa1h84Bbt+9u12jd4L7ygXfz8k5mr
FLnjSbmC/iLvp25ZawIgCfl2nlnZulAsjqEsRLPiaINe/T4WahJLWXmE3V22ijVl53ZcxliAEcgp
xT49Le59lWXQNecJ1GoY2KAFRqATrGJ7KoKMYlUk3/b8mxiT+Zi6tmjUmKeyiOf6Ymrnz16Q83Ar
HMq0TwNYoJo8T+bbRNDG3GwukP8+euzvIILPd3B1iJ1EpF2N3oJc2I3a0LetsWY1z7aPvR6qrjYK
jz+ZuYHS9hD0bXU47XVfRalgtcl2ueTy3VKUO5u4h/ZkORqgVwPv0NAs7tFo0H288T8l1FErCtPz
ugvppHgk3xWeOG2nA+E+50L+9bqGDU834sVKSMdOCxBNVmnE/XhMlDkNQ1+MO6neKsuUJlVUjuLv
9+pGnUjsGRyXNJGIEqhFcQTuyuhUgrZQk64+mYY93CnDnc0u9RewMqkAomh3P9N94LjI+ytmcQyw
zUMsEQOSwfP668SAkdOVRW80ULyGxblCouyOLoTR2OCC+INFaXDncmkl2PR45QB5jlMTXL4sU8IX
St/bxJziXcM/ru1SJLBtdcgA5POXLvsxQuxsEQn5TpJXrtk4DJat+gImnsTryY77aUbO7stDUwQf
QfkPEUYUyzbEUqKxIz2M5r198C7HaCkHAhIb34iv7iFAWh8PEIlVgzx88V3PpERWiBuy11BcR4Ws
X2zpI0gnSIRr6FbJZiop6mk00AMvMYbbO3QCoB2e7qpfa1bu1mLHYUwYe8odnL6Mko1APsvd4ULo
sbSst+bEUBpvG31q3C8lemYTn4MZwDECrlatdDJGpzo87jDJqM0bb2vsps0M9FILw25nf6fw6wBn
ZlrZVHVgN6d0OGVsHRh4H6NJubVtvCnKrqBALqOFmhjTAXW0HQdxr3Kiq7mOgW2F8Rp88ofeehvz
3ieHA4cqrAlNXWf4B6/Jxofm8j0F2jO6Q0gHJUG8i6ssURI5BSm21eRzjPIsUmdKQoV37UUefICS
sp/Zn64FMlFEa0v/SfGp1p5i0Rp26tjG3c+SJ+PRQ0pXCGUGl5i0TEbZTTeLZNK6b3Rbd+1cNSg9
LjzLyCX+bBB6zCGQi/1e5mvMIVfBp4T3JNo+fHlk/YNGVgCLbn8t+PFdf79IOpwIlNKGQTHxhmkT
2QAE5nQVAliHLCFz++v0ORV5Yh5VIA9aZ7bPA4KsgA63tIxCjATEtcMQ/HmzpZzAbxUp4pXLn1na
6JePQbU3KH39AYx+KYIaaPjyVg/20BSDKD1c2VyyOt5AamzNwFm5HCnnPDodMqvcpZvARbGjCMfp
57MVOh+uQUA9aiGizdjEGbmlYm/D/lVbLuw31qO3sbxpXWN9V0c0OZW0vEjlT2Dkv/03lDWfTnuh
mMIOb2RAe2eDLZJAcHgwxIjwnV3Cmepf0BcbNlcIpeeDpH8VU+9mun+2K7Yonkzd8v6AWlSCldeq
oVPf1tibfB1I/dlp06glwatFzIuTZPW64XzP2NpnvIcJ7/Xj4Bn1pqNKqcLKz182AAppXtzyQZf/
/BUd9yX2jbt03ydp7dqyhwnFvUJbIXOio395vowqkR+3KSvmweRy9gsHTpvTWPnkgZaynppzplY6
SdVArndfTotNR/Sn8fDUHaahpYnOxzfC8XoXp5uY9l2gEGrXF7oHa5L14T1X1+hMhBH7jrm06vQC
pDRjQKXe/Rqc3kY8voqv5Wy7P/yEg4g6AOyk0fhhwMtRxPnWw2k8+XHDt90hXS2udfhbWmGLMtHf
kjnm05A8mnBm66v3gN/u9h68eTbyvveyGwRZlzDD1wkObATeoret9ViXO3RO1DDxVD5hy5dC+ChP
SuiqJLq2Eyq68zNnpsDkpF/9+xBu3/O3LuVyrdiSYKw7yXMq8RqOioAGhEw3BQ+YUky29XZq/roO
laCY/SaRXTjtFYlo6Ez06JMxG0bPT3eOTAGe0nEEDJ68ZwkuuIYcIVZtZ5UA2+oMBTt0YakfTM5c
7VjBMJdyFbH3k57Z1vGDxXOAY7YojPW2hN+i3vGpy0u0vt7PbAaK/KrLURWxhUhcAF6W3c2wZxPh
RTow09xV8hVbqIJty/Mk9oMdnM3Em7IyzlaxGO4yOOei09erulbI+yGyHWbP7VaszmExUJ0NWy2V
HbHMWusNcxrxCQqyO4dIMYDyFUBJOVpUDjZ3U73tkcWdKF41mIKiEig+b2Sx4XpugZ3RfCZ0bbFI
DQraYEZhKiDZj6X6WV96M68jR3V5ONSd9v01SBNpoe90q02Vkgmn1XNnYzZ26F0MSFU0qg9HB0Ry
1QShg4NTFkn1eUXp+je3Ym4f0sJCHS+9tmc8hKCaeZlHJJSseuRECDwLlMc1Z3KKgMg3pkDl23KG
eCUdacz8QyqihBIW7jY9X4K07Vdtn2jxDMGvVpvqYPMYVrjfzrU6xzcpuHOfUB2IPX/thDJlDd1F
Ts9t6m8j6ChuxFoBn4frKrMZgK89S/DLKdqroHPbDZqwgWSN/BdfngVR8MASeUMxr/eLR2XWxPda
ylwaS7E6whFbOj1T6Y3IHxnPmYP/dVXLF1yGbGmjl3rsNwQQ+/NKUabr6/Jkt1DuJW20zrfOcd4u
S+KHuKCB2P5IjmBF2xkg9rihOya7L1hWCyNL4iYJMh2jN/3kL3tZ3wIPDYa3jpJdsilkUCghTARx
7CQ3jiUidw1IAJ2wBD+3JS65IF7WFrI/j7CNy2BpqnNSNOhoq4VP38NmmVzthQt7r5CvePblR270
VLWn0gOlZ2fMv/IFkNkutx9LR348Lg3HGFtqAOXaawHp71iB6BtbTJ1ZiYem9GRe/P+5gLN2a2eT
fN9ZvXSorSLyYXYds8+ZYWElYREa0kkYFUSyZZv+28tyd3FAN/mVfdt/2cuvzkA0BI5xJdrBp84z
4LfcF7HiEG8pbp+Fb9bZrHk3aL6iq8kbNKyIICfD36wMBITwWWF93zqwoLCO+c35cPUrXfZ5z2xD
j2Z58ZpCxOPqo4qg0yKqLdwo87UejFccrheFaRf2hQViZ5LqnwKFSkY5dvz69Kc245O8oCstmfY1
Mz8+dj5l+8hmXXv21Ikm1Os7FR0GF0Q354XmZMHwZd3k4/aGf3K7mI7POsXjMz0Wmn5zocVqGQtW
Q62XpzToBvGGn0T79HmAZ7XeU7Bet6CPMyhoEo4+/oyB7Pr9I1xW8ZU3a/XmDmObvNBX1OeM8qY/
KPxEy8xfVxC8BxUPIhgQsDpCrrc7j6Zbx88chTIGBhttM66wO8aLKsgAD0WtszceMLFgcB/mI6So
d2MOrwe7sRQ9BF0fcPHlWxDJfX7/2V4yRm5qb+NfV3Q8gKpe+nED7Csx8s2JjXJ7au8/jdNv4zuB
zgILPBkcr3itP3ULxmK7//jVl+1zMMlJck0K7rCMfQGx4XsrNMfXRfCph9Wj85fN9VK2Cr1/8XPz
yxX7LwRnBmhZkRL1fUW+fgjh3CWgFoGnr+6z6EG8cfAlKKXzaiSRRI5Zx2tfDHhp/leOd3sN3hJs
FYME85A+7317vtw2Oao/Y3Hek9Ul4dwJmoeoqhFUWHVxupW73tne02VOukeT562m/ACjfF6IjFdI
RUMDpAdOLKSrWR9/jc75GzYYptC0ejeNeVIufAbIQ7UW+llynJ1ahoomNz5XIjI0g9VXYhm7RzOB
22aO8OEfLnqjyqhnlpWo/3CG3VlBZ/FzQ69ZEiFJoskuHa5DpD3jyD2hqOEM36BW9xv+X6JFYzyr
DRvp60mKTWuiI51OlUVzj67AGcGn7d1zmiJjqtX6QCHs00zPEWRZ1K9QM+/rUM8V16laRsu25QjE
YlR1y/jRS8kMuQERxhDQLYpsakAD7urEfUQvvmSzAvLa6C9R5+zAXCIIZG2YmC2KOobtnbSAyKLX
QEFUDnSiK1NUC2c62/GAWvTXhuuSMO89uQm8AW3jiul4rsqnPXEeDkf/AsH7zMt6L6XREkci2Qnb
/XI0TOcAocnu8tSVC3VnI+j65aTzgzywgcwEz1XynYh0A/zXY1/RDpllZZW2B6MN4QhxNEguwgRP
sI72OMffH9RUdi7Yd8S6SYAryxPNblA+VWyJDRl9cteU4V32BLPF03+A9JnZ6PiX0eKA+dR4GXWs
/B7m1ImnUS7O3bDWkop2UqdbHI8zt2R5eHqOhftSP3PwgkoXB0YkDsshxL62jB1vSXtXwOqbgU+7
BzWUh46hosnJCqmQ0vVgIjywygPTEQQdyxMcchOB897jIEItyMpZKtHRTJrwJvJNmKp9b6lvAUGk
dNxLmuDCEAbx9fJohV731X9G6+zVy0icqVvpL2OrSrFYLSsXniL6ZUhGhBcMdz3aWHOuNJGl4m3b
2z0M5MVOuzooKxbXLBrPsEfiTC5XAPK9KCatCwAyCsqdL084/oHabaQcXdYAPNDa87Iy/+RVa8yh
awUGN8UcD1a+kcV3GQlaaZCvb9mPO8KeNa5xcBa9YoTyhOYtYPlcraheoU3OCmAZHDbRdfJUWDi/
CbHgCayC0nugbDnWZzRBXtVBYmvY+oprx1r7YAJZj5bGvriuRwLkIDOzzBj8J+udev8ICGwLc6x0
feeMWy3H9CXGd4AOiFWcQnQcnkWF7ZpM6C192YFQ1TUMTW6Dx+H+NxfdlBq7K4ynJVWutoFyLXiU
djQMogrs0bZG7xpM5qZY85XGxkzoS0XLfXTy6CAUhGhvzo0dJm/IU2nJLbXTyWHwMHmgKSWCw/lt
auVpIDDS8GS1/t5/FPfybuG/OHvq0ZT+AH7MxByVdCEYc3pcZXh2UPQipXyU9ovtNyel3HNrL8aF
9r8dZLaes2p6+eHLF01pM11K1abW55uGvOfENV6IsdyTxXTeHLDH9gTLyhJDvIgm5r2lVzRIH82d
rVjPRDPeQv44Qtb6yIAt3TzFiLsP99Fm1paIOOqiZpM2sD0p3i4yYxzJGcUjMS+HT9t/YI1zq4Ec
Z2tKfCExqDmtZl76GWQatpIX3Xc5XzDF5PbEG+kJmYDPC3qWCW3334P3/pDMzXGnst1ZxMuNz1p9
J7Px4r4YO59wOMFxTzQ5zfTBWWlPPPVd5X5vP6X3JJUA//5FHL82FJ/hD4WTepZ1+/Ze5r8hBPWP
ebwUo3ytu88MyFgmakEgIdix1aI9VEllyx6GMHDiYd3Tf91vabmsM9lg2Sv/ARYVSOu8rnFWKhgl
jVYzcU6N9C3F9f4wYoQfa+hjDnE51xAPSDlf36IpMBukLuxUawTmuD41f7wgTLHTJjg0ZB9FFWJD
Zpb9mATAETZObSIxNaUZqYl/GlNS2sDvB22XeYk7Kr0zFf8kcdki8ODjhPhaONv+vDt7iW6LCtmm
R3mh52kuf9/BNqZ7DtC+MDiKR9QqUb70alhE6UNultVc3Vm29fFKQEQtS4k0ZMmlIE3JQbd9RIRV
Nt3Mr8bfuLUTnWKaKmNyj8BMF1MrW2cZkTvdPZJvZPDyHvAt8fbn/cUsIbkUnIqHt0pFtNtDbQkn
wL5VnB+OOiYjxR/dbSHdsC13GOdMRsvr1gkpXOfYHNthXNzFZRuDIqrp/CaQRyOFqn3Ew5nE23xf
jew/JFqKcJ7BaGavVS33hM9kogWM4wEFXcdcj4GNBS7hquJvJEbRLpH1JnQv6w72//bA0m7+TII3
j24FaFeugPr7fk4acY7JalmvmMnz1AuGszBndU6aqgfvWVOP/shMCht5KtbH42qhXZEUNjkJnICJ
AcE8BSmRWcTg5Z13vDQx8/CTFN3Q9k1Onk75sRHQ0gCNVk6qocWn0Dmhfg7Tn/rxe9y9NXojh3RL
0F4NZR438WZr/MsgvxhUMPuI/KNO+/Fgax94c4yOzzdxeeV+IZYIDnCQ/qSh3fwgB7qs25RUT2+k
/O+uKOyFedXfMgn+H+WJpNL4gUHjrmF84XgwGmD0neFMxVfG2L+lFroUn+yMGq9RxmZ8ZsTpxdT7
MpSUUsQUBJKuGHZ/HXRf0GkTa7sSEJwu0dXt+IHuep9GsrXIvfBfaL771DbghXDHlqLQp3t+mfXX
M8aBz0cUIsevva2vAmsZWw5Hpt6+gpp3l8+NRToB/QyD8DA0vW86DFLtRwE4Fzknvm+WN8bZJ9ne
//LRGr0mrmHnAf9GFomnsgmGvOd5nzE46yFOO0agGRxaKqJrdtdIfwSSzlPR7haU3v+WslrWMfFV
yMC7dYMoWybUfQmhjpzqwjpYHai7QxMdUgsMSaHuoR71BX25eTkmGttasl3DLpKDf39b9x36sefk
VNGtgmU4ag9eiFUhzHhqdX9tRJ4O0siDnQX3iYg+ygjPE7MBZOy+3mn2m3NjKi3ZFZmcyrd1f9pu
tGY3cS4pHKMaffNVQ4ZVl5wlyey5J8xI0uKIoxIr7S2MVDIu4qVAUsVHP3gysf2OT2cf3k2wMqL4
mLVSonjm11c3Kvz25/jqk+vskVnoVunqsCipBLQm0+uBrznKh9pPVsVAQ0SxQm+XOBHPcBP5vejl
XZAVKsu3P2cBx61tSx+woTJ3REOGy+Oxjdi4ju8t00G+3iOjjQRc1cPRqzKhAC8bM2I/VHB0FIIW
G4oLUc14/w2xp/nBJckTxdZHbjELmyUudYUGzWXrsk2UR0cBpl4jZXQmZuvEP9TNmnMnHKxvK9Po
9rviDfiJtjbPV/kmTx+M9wh7yJmVvjAWROrwwCFeLQBgScbAYs34yXo23Q9zFg2WWfV9tMoIiban
yacgdA3HEG7H8NQVQDDcUo+nLdCSD/z6r3tzjubAodgWIS7Z7mTG2yvry0ZkReFOYj9H+LHbMIjS
l2xcEBSnSANM4lm51khR+L641eJEAoHuxEivpx4D1xmJsDXH44DRnoHduRIiUMJ/Os9KexLUmQnd
Ws/DSuN1dvZR3x5ps92nB+yv6ClgYq+znRiuWjcdhPdsc3c5YRnfGpQFmat7ghwsVhw9tDqjCWhF
cuHNoKYfDN4hLhHKTZErI1Ayy47N1KfyeZZB6XQhVgDOyjWPNJI74pU78XRjaOwuPBpBRxH5iUd0
vHWQUqbYLrkO6HGh1REdjtkqNmY9xob+upZINMCp5h2hJPktkXHwGAK2VYS2vDvlw91pQiB65oJ5
uuL23iM+d+tBlAKOfdbRZPE7GpDCjJWMiNFj25tqQnh4AV9kcig2INislA83JmpX5d13QuVt1VI8
0S3zBkVDTUFqO+rhXCoijcTdy9fmSTgRerrNbWR/CZeHVI51Fh5Em6isKtSq+P0Aan+7i+dTOJ8D
dt7GJguowVBfrOrWtcV4df0AC01YeBJyily2GA8F7AtA1brM/PBrIUk6p9RYbUe3jYzu4rwkjJAk
BvRH0DuRz9zopdf6Hyn1gmfxo4J+H+rTbC9HUIc+gVoDjln11JG3Da7xVtHaJ8l9/AcpmFQmgtVr
R/7N+dX5SqLQ4m8+ZptuxG2jA/Az8r/JbGQBxDB4TooFxRvN+1X8aZecOgVIQSMPbwLW9DrUo9W/
MTt+eTTp0KVnXce/4jmqrfAHN6hohZikFg5N7a+tAN0QStEDp8N58zgGeqZ7+RXLAZUwMHr8wiBd
k7BHmpd/iM0F3PvXOM0gjHW2VNeshfNHExhC/8tEXYp/pLa/SIEYf2zkbXbdjJzAvatggi4KmvAl
ysxZhMk/eyUIUjzLSGQaSkNKDLDZp4KWPfQklkizvW/VvDcxOazdpUJujlPKE0DZvWFa6qo0BF2S
iA5NJRNoZFfe1sKNEDLz2/tFgVYG40eA2tg7l+ENPvlTMn2Hbdfk2cXT+OIa08VqMjr+4kj0uRnq
uM7221nA4WdWRT4QRmNvn6VG2y5R+Gk4HO8ffpyMxoDai6OrhpHNXE67xXVw7BcbwD2wLIyhu8el
10EnFNb7zZANNKfhp9z2XAb5C8MfXsrZRgpwSpzcG2cOI2Yz1sMSGfLJe63BJRcNHjpn+/YRyoi2
YVLAmeS9iFcKVX+LPeURWLXYW37QtgiRcngGTXOZEG12NR+IjKZzllCwWVUozZ+Bb+xdYaLQYxqa
O52dYeWXZOPbnBg/Rv4Vq6NAyGWvxfJJ/jSZ6cHEUZXsxgxxiXk92qyLCprIZIdSOvYwtwUJBOAE
L87qCFlED1HuuIgfqXd3QwGUjH2NIIohW87+505936lY/UoEhJcD9/4FRHXfbbUusmM05X/zu77S
JZOVTpug+jfQ84hvsG8mFAyGLql4o+V4O1yvX1HHPJdNNMxRB/B5KSrJYlD+Lz85JExUoobho9yl
CMUY7bKSAuD1i6HHgGIuKzK5sl7MJC6Su69qnNccba4fnc7d1t6HXyej1JD4SuxkNqDf1sIlWvy5
9otNgGa0zVVfcKlMv79Di+wE/FRpD2cM4PEUGAAqhoFT+L+wnNYixp7XHH33wS/xEIltnQ43HSIW
+Mw670k1Wq2T/rImfjIbyb8SvpeqwWm6eZ964gdbbNnpcs8h11YMkf2Tf26cOo024w6kKqsixGtO
bsUFRiG6uROUjM7B7t3NDolQLZ4QJXItbywhmFr/MMQsBdPUSAQ2ZlDcJw7si1B0C2x94yzLtqCu
1l3y1GafQCv1/k+LMecpHiUFcCBCwg++eF54amhUG48mVBBf1gUVEghbJxsQjqWynVIbAU1CL3EC
nSTo8mbPM7LlHpLs0wBl1AU9rc2mVcJKkW3dLGUKnrIiuMOpMLBPIdwgMq27MRwSxKwZvTIqP1AN
t5NdANZxdL/1JmKLQycjv1+6ppFHzyVPygRcuhJh3RFaBeTabOpvAs8hOQ7hR+FlfZC6SR6IzCTh
7xHeThSBhMki/Y6domozkTBQU0IOZTlH7Zrdu6BSvsWVoEE5ePaU5pOzeFlu+Jc7XgV2LuXm2Jqz
1AwWGzvNfUwlzmorT7fhBIu28YOwBPxJ9po/o5ei0V2/mrblxfS023OC6nRwPDu1CPbf3pTl9WWW
wqnocqnarULVpc6jTS0C671oCquwzmw2HfNs+kTIa9DclEbjrg0FG7MoK8mPOXc9DbLQuQuH0VJ5
UQB7ahMiAU7B0+fMhNadSittp5TeRLZdJoQG3Lurz5cjHEIaQ5XAJvTvXOSfmi5w/a/HDcZwSXLo
yAuUNERHifkkyLXSXs3iGdTzMNDVGZJqn5FNIvoX3xEgHT05aE/R3fO4h376yunXcsA5QxIYs20/
RXU3au/0y/u3AYyv3ItaOsFoU5EKARi/Cj5oDBPQOMn/3pz1TEXcHr9RE4Or3ugAl1w5tAUnSOFD
OnTNRHIS0i8i1SG4JdOq5P0PxzcBN5/WH0C9slu+LKQ/k+miLiigBasuNloNp0ffnMoxT0+YM3LJ
cIxKbid2oVxypq5uQhFVM36qbeoclY1GxKdRMH58Rlfq3bub+l0TW8vsSSG1kUMaUTpUoiDVL2ap
gyAtSmzVRqPq9tGKMCqpDPJbQo/ETKrcIcB4Bv+quzKOj8dWUXYIpgsnh0/p/H7ooh8mEg2WvBxo
foX5ht4IRHCk44bIXjFKvbheVxXx/Uqh3t+683774JXib8BYutF+kU31oDPipxFSpC6ydTnMnFNM
KHNAhhz6Dlb+eKJZTdGPPrOF0j6WLcSaY6gVsCZofr5Ssm2IFvbgF3p6/wE5YrP9RiRhxj3N/kJ2
YfkhDKZkH8zfwiQEXRVfiDEwPOLXmpuOl/zswQCVSH3REY/ytbvpMYu4oQKAk6PVErkIMnJVpTJ9
1DsTXSguGRwLQ4YBhbLb6ngaDC2cQMmDYXcvLF5KGjkkJy6e2RwQdyNhms7FNDJ8iINzWXDrDgdE
mludDE+CdofN4/RwiIaZLY60uoMYS8OmCfxz1rPBckDPn6/lrx0arXkw9XCgKtJLgTuJAYgQ9OT9
bSdq+9sTj6/l+ydRNQ+w12/jaUxeXKQDVuhX/KGzpgSP30N67MiLcoPyXTgmh+FtYVtmCYvaYLNs
rmzbeIwPDuU789lDUXEVum8i500jIwRPxLd37zS2ow5gxiACQry1UYDl7NIDx/XvbiVPOAw0LfJM
1vYCyoh5oTNTGyrxOo92KVM6AgEY9At4pk0rEKK8TZ9T83sOjPEx7Ak1IFENxZrPRt5wc+6fLgBg
G6BEoChCjevanRfefgkEd+LVU9qc88+xGqHwbE7Qy3bZkbl6ehghWQt3yIJ+/L4cJEx4gJQv3462
P32VGruAOnBXkmtpeg/7Q1QY/t7bum+ZJJ1MTBiuLNW+RLKBoGitQijOQZu15vnlRiXEFFooPm0u
jDTc/WCc58MHL6tA2OQ+PFwsAg2yBgQPCbJSmI3nCf6FXYPKWFenlSg8H1RDrrVO9vvrv0r81p8h
2PBSOY5Zq50NpzX7HqiA1SsVrpFVp7VA6MSvbCGKYxdSJl/ghBrA0na75qmidmoUuTY+oPR3ZBZW
bkwOXV6SWWJrp0qVWQzS5jCvwyKP9fD1MpLNzb4oUYXgzKrkYe/sYzttCv/H7e4foXhzYq14kk3W
reemIk5KrEVB27BYKgDSyHAWPc7ckztW+hQdaUGkqoFZ9O8Axi885HHILyPq0R0GmZeJveigOh43
RcMqMGqC1JSWpHHn2utIAflPIirHcrbS43TWMowdg3iU0+EUwGAZe9HVzH6fyugX+e8SkfQFdgu9
ONWSWsTRpkArG8Wlxe/4cODIckNibsBjcEeDLoErk9UGM9pl74nSjfABazxmT6sf+YFGWGU0gUrr
89Q2lLOb5pBG8Uj3pkmBrPH8PfRmJx6nuv2DNmtskq1fFgK1wHwsqA6x984bcF/Z/7A1580Q1i0K
HNHeyBJY4jsKlEnRmRAQJ1h775eRVN3+tJ4fK823Xcyi5Pty3yTUzMEU4FuSso7iFTT1z22dOiBJ
lK4QVt8zJXaBQtEBlLg9L0FtptyUwDNloS7uX88FUc4NpoR07LEkFUF3YpbrCS44mQ+Pkafczk8E
/DrR7jMqs5yp3yc7mlSyMZjPvT5B/wfLNeMhkZ2UsiILSYvh+3FWKcjNVBIyM88P3QueYGKIwAUj
ZHrIPfzbGymVQR6AekQnA6N3ebRsl95/UNFRpCS5yw2GDbLJMUVBkOi+K3tz40yzaHk1HwxcZS12
sT/Uh6jrXafLc3cJJuu1YvIY62DUK+0avnZ3IAE/OV34pZ7hulyzu5MXE0zVbhsdxb0mtwNmhGDV
frr+nsLQPRKY5850GoBaHI22YsCjKn43o5Ztu4Sl91W5VrPP4qixWOCqH4K7Cp5G7W07YhaHFU4p
WVX4DvF33k65lfwThe3KxXPluI+87TOHwfHGDSUK3vY9YVKvyRi9zBV1QKbM+asT+WNMGd7ymcuQ
u/xyt8hSNHj0YEVCeLwBeQCmjFvG6ezP+OyNTn/kN8U1NDKc+tI1N1xzNWYIcVpbKkHwqjvZ8CpO
+oiPjckBcEO/XjfQwb4PDipzUTIr5RvlYZPjrLYcqgGX3RsUI+oOQ/XRanVgTt/39tAfAC4qT08h
BDb4Hw9+N4YvSyTEeEtmuydeUsTsJKgniswRwfC4V8EeZE3nT+nMxIVCOH8KReqms59k5DIQRrCb
Lep4ekZF+ppd4+K9UNxLxk9ejT/74fdoA6h6iOMk4Y2igwRJnc9kSnF3gWRGPbUjERKhoQ6odVVK
7vd7Y03l/03zPdf1cpOU8EWSw9jCXSgX265EuykZJJDCZj2T8vGGvWuJLxTsw7DAIPH+2BoL5uat
0UOlza6rXKXGcmbuJ4jFo0dRNZtztS7JKMdDmxOE4QWDKnNwn7U4ZghI7Bm6xr9yUvebGcu21RjV
bjoLnLQn0A9IPaWeVWKaxPFAIng/ND7MwuyKDkPipRC9juVIRj9kaJSUVrV42EXf9YdyfbnFQ+fF
NRjdVsqJjllUS0j9MTm1cs6bkPrCNm+8DJPnFhTFkB+aUvSVZUQrx5hytjsch1kY9zPiMd4dTDuS
xnyVwpqFYzODk5wpRuZTeJnE40ML+1W767XqN73oQYq9Kkf5mP0j0ldbnO9QUpfKtgmvZIIA1cY3
J0NqcUz/Mk2zCWp5n5GqYBr3MxAOYKP+2EfwmH462kVIe/7gAeUEWoKL5/OeLcLU3Gmrr5hjjrLa
17Sqxac0Ik2bvyDffv1jRCL8dLlugxWkL6gGMoSafOPkvO0Gjeet/KckGULsgdjTBos3BlLp2rac
6+7hLDtBvj37Mq4bXr8XKt1niCHfMm206sYHj40OgtKrQWZz9TQzafTQ2jnioem9IG6u4LQfy0yF
Rk3Zy0eEyYj4eleMZqxC391yn1FG+BZCq31XNDOH2DrM0cBO1wAQ3g9JO9ln8H001RR4FnfOVujw
ri11DmTfJJm5BX4Lx0QqE/f+sEcfKnCmNz5HjBq8WPGkpzZKj02dCtw28L4/vsFNYCVQUjagRV8x
rbOVc2KBDI6XKhBwBYhdEiHUKq09RdydnVrs88RjR5KkLOSMQNakLRGmdvng5RRBS6lyA6VBlrp8
3NAUZYRf4qqYfSKTgbgg1BBccH6skBB+k48z7KpzDZ0KGsrPzYLz2jVJYh1eKzJPJdptek6XhV9y
bg8wrF4ghziz67T0Sa/BV/bXbpadTrtWGxbbtRB/u28fFed8kW4lRPpjBkoaTNP3diBP9PNjaTtc
JgOtCgr/j9AbKpFhGHA1NZMB8drvlR3V4amarYvASPStDdqbtI0caR8NQR76ep3zw4ylv6E3Xfhv
reeLpeohWqda3nRcc1gqTLQtEVI7Ke815quLCbZatu5tzLPsACiA67K5LtqqpEjP2ef/NvhXdbIu
gBwGnFwRrb5TMZz7Ji5Jl3+QyP02TgrXSmUYlgVU3zfQL3NLkPUYU4wPLzlQ4xk+pLetse9onO15
2KyYn4nzdUI/D7gSp+9RUIKSjv7lEN2eA9LjBLRnhz2/XzAgaCGtD99ioHm7AI/RTw9uImESfD40
NdDhIb8Nt+ARQenvN27YpRcnC7/vZ+3TX8gGheI67Gnm1/gpmL7KxOj382AsdKH4sMSJzdVeKxzd
7rNW2f8PZR3OJ2s9X5lWYB99krYSqzRyZHqq/zujYlRZSrQxm+es4wihE7PBz1VjZpwxdhi/JkNy
5yvWBV1gyy8Oqp41pAEZFQh/E1cJLsE3IRwkPR5lXZ/njhwsd+I1pdSyVEXEaYqV3e1XVR3B3gL3
8aWJqxnH+yX9MucrITcIRbIdYlaP4v0O8QfpVd2SiIXg1CjUd+xgGi8lNlBhLJoq3ttLkVHIgrC7
NlLyyfV6fDHWbcaMIeIzqHUuYyvmDwmCWgZElyx4sOAmTo478nKtKJqbRy3fAYykm47sJGk5lRU6
Siu9UZhQZ36KLxAeccGvXR5awWsCmggPEBJEbLryVf8+azXMBpVOPBzx/b8iFqA/aPStHOKfBNYK
BNdLU5pmlwtsUpWaknHFdQ4H99JjUSouoB/DRQ8n/H7IQfKPpQI+NM0Kkskh7Anf86sHbupVSSob
zn55LNaIXR2/HO2XLNa35fqLxGvYz/Vfcp+Wbm2TDMUJjV/eH7aTwC30Qm48D6LRmMFIFKJadJRE
9NwJhjoMCpnjSPyNwC/dTkirb3iV1/DPvEjcX8Tk7udXjaG9oEIczeolDqzoheJ443ltQ1XRwHzF
PK7LER9kZMfDChblVdyfkbQgbw2cyqfQALybUWiCRbtK9deUVLrvwowRZn0ez5RTKdusetd4m5hF
vGX7NVSW/oA8n4b98DlzfcqzBIQISj6tnKUATQUwry8kGPcmmOTnmuukvcVnuPBsaMSHfffkE73S
/6wyMB/l0eNH0v0dSW1jOB+lwjjJ/L8yogyirz7ALloMIMCO4RNNehDMBk1F+JFbh5s4S9AZ8D9q
XwWGv9H8x1ifD7C6jmLNUG+LOy8jcgPhL6DSZ4zWSyqmZv1xwhC9uNNiNiT187/9IYnqmwptDkr9
Y3pVEdEde5ljSrTCtrj7W8Ou+wrvSoSaM0BTETShhMGMYowFiVF4FPX9GrVJBh6RBuLbx5rTHrlO
1HfaSuM5FFnIHfHdy756sjNKu0M9Yp3mXODDs9BFIHoIdruG2dvB4T8JjRUc4jLsSE7vad9xQpOz
+QBkDzaAzgck/pgYpPoPCR3EMLsYPJCwnWB9NcRaf7JMCCCNOgwc6l/L5kFpAEtlgj7N7AdJajeD
1cVQYGkzkMdoEoi7OGHDNuv6DhwV1CxOURx0PiIjtXNo1FOFbwMGs7w+54gNOI2v5V1UJT4bZnuj
VzKsMpXNAfPpbIDC4LHqlM7A4gd3wYZC3Zn3OzWfCOmD6Q3lHHaziSXnvsDckDG5nq5dEIgOXe3S
mR/UVKsoRfMYOXXn1uuurV/7dxnHmIu0nvS4ror5YVA3eVqSCkRX3U5hNAmtct+wttyhQVLz92NU
WH09gsyhncy/3B77uqtPy9Joi8vPuwwOSGyHRydHEjK+iLYKFgaITvfLT5mxODdeE9/IcqT1mbTy
JLNwWhBvAz/GsUGKpwXnr2RI89CKjHu2rJ/4Vasjumcjb0Zc8zpQi93ny6TqqHW2/F7hxKKlnJ82
kLQZW5zvCyvK16AKi/4qbkW5ZFZCthFRMTkt/PPeqMtpHRIKzAVY6TlbMeYXmi5uft4yt3qVThv9
1IXZzVDJEv+e3RdKB/gbt7hy7iNxSX1vhlKUqGjDFk7GBeeDntLPK+fng3tSlLGB5tJxj/7a6kwj
przGFQpOsfa4eryv7ZhQebrQg+EGF8G9Cie7i0RZCIuLElXVMYkXUCet5BfG+DJvdKA3D9zELC7y
7E1OENg2vX+ZdfOeJ1nD00QSPXi8LvBZtKdV6mB7wbFZ27jsFifvhIq14iidy3jeMx+2ZnQXAhyY
n1lA8J1NEttxsPQ67Y/XUKAQ+PtuvEk8FYADZsnIJIt4gW3wSMYycOHh4BEJrKySPL/O+Aaf0xEQ
Ny0jA0N2sX2YN/c9zbsipf4Qgl6asZap2pkhLy0HWkX+D4UYANIL2l7MB3NV1KQzIhHtiRNFT4Fo
g+Txwfurtp7+AM43noQA6hSqQLQLR27Uj8F9IrNYBVawcTUxKRKJpz9BLuIMiW7dQo1QJZjAcmx5
ONNNVWeBSJ5BD4TVtcVyKY+muIU/eCZr5uyB+CRgQrMCS9RqbZ36NNs0MPv6AkrS9Qr1+Q9J/NbZ
u6xwMRy1goXPF43Tjeah91vd1ZQGTtGELKCckqcWoK1+OIwhySw1ZeUgc4OdqinY3i7SM6R+xB0Q
m5EIGfdUE0NaglzWcSxPCt8HT9iJWTTSK0dNQwCGqeiqz/VqafngucZKpaZ4w243YTnvmNJDGRHu
UinyEsa+Z2NfyoaZxoXnWBN7VXwYox8cimoZgFf2PotZhGoEGSqhzY3zuv2rwSlPZObS0aC60FYi
vCOUPlSi1Gy6rhliT+BxnBb9hwgn3YEdy+HtaDEjlo5Y/YX7ZPkyUkQXVErUecsAvvmEw73W/Ww0
waCJyMG0OXXeGl0FC/0+ZqlFnzQe15m500ajFsBb8CnTGQhmth4S51Th8KCwn9pvYxRaNVrYpgYJ
SfNgGzgudP3OL5U9whM1YdElRS7ai9Uw+JzkcVL52OxlKFzfnXIQPIXFrSOVwjy30NNcaRFjgPy3
Oa9ow0SSdcgTHj01L0TMYJJ+x2Mg7f/w5WoQx39/n+wyZX0RvygCwmiJSG0QAR3GjBbSdTovzrzi
9cwxhP1mSviWPEqxpR6Yy9xDhJjCB4odWOyUF08MRsYBiU/QBwgKnPhkzTNnFGJAfSH3h1PEAIEo
EsCia3DSxtMxCkULT6l7tnDpbpvzI0T9sNGP+lnY5P1iVa2+N50xL3YTCLKsnYTR55zOl2+Ueavp
uwINf5fRlOzVocqWmoxiVGXF8OXczkYOZy4CpNrG6VKGG7boGQxVU1HMQYxcU7BUMQoOZKg9PIQK
kAW/xAGeajoOAYzo/3w9fjnuVbGc8u/CvOrgmfVsA7oTtIas5y9raLmrfVlo/Rz0/YK3UtVMsJx2
d+NVqLedXmuIuPDqXcqV+LLrmVMCa1f4FOZM40HZyvPDLjs5v2rafgDEaqRBdZIiC1fAVGkw6p9E
VH4nW+tsnN30gqIYm76wjpHCDU3VzGsd0nhcuRVnK8VUpzpvQ4890y0ZDwaSOgG1UgvjMKd9XcKF
2PGGiYdwIRz7LZl6ey1+VNTc/SU+RG8kzyXNXkM6pdvIVQz6pBLjkOaN8MmmikQNThqf/HYC0VCr
bnx8gts+howbffIOSC5H6wpYA2ZGyWG7bfXkifPt1pC2u9PkPrgVb893l+ZqPE/RID8EYv9EYjNm
hTnoJ6enjrSmhVfO8avsWJnIc+f8QS3j4oaQwLRyk32onFjC1moqFouF+pRnC2KQMZ4080WT12Tl
Vh+wuKp3BTWpSIgTTFWAppTZQcSjqnCdHfnQPLThtmxegQox6xE4zRx+I5o96CTwQLRE850yA3Fp
DXf3n+dUDMeRSmQSmgwgnbh4+ZSO1oW72PeQMg0HHbVOo4fzJq/EfPqhVC0HGoDPy1KbZCIpVi3M
B8XY+XMq726kgrFHZ0gtDK2QwHETQPe7CQUpXVJeyeTRpyU32Ah5PtS1WJpzaqRa1I1+/299g/7k
w1S2p+7YdMvVQ/h7NzwwiE7Hsqu8HGVkkJR5wkwFfh3RcXA+5YExWQI8lm0pzRnZILZQNj9HP/ab
xrpppt4YXQVCc1i2dQd5ZuLzexLVuK2rLndJr40lUmZlt5nNPd+OCGaUend1uNiZEiD7flhTH/8p
1l1xQGd1MJJNyEqHJp80gVOLfCiSKxW42kfbGoDMQg44sBZ2HDKQw/NoejribARurCw9gHoTftIx
GP47Onl8hhuDrvtG2gGOeD9uKXX0cgDoLTwTFQHBsvUb9ti7FboTxAi9p7WgIu9yOZNN4uBuGl/V
4NFki/3gc4uub49f0lvDQEnt99q0ooU0zgwmkAlRGf9Iwix4m+LrxQPUUaS/Cd44vB8Mw5YHYawI
wRbaxIZeRotVTwaCjkamAxtgZ60OyKtKDrIY7P5QM6sAYbj3d5u8tInIilzz2FCvoxXUY1bpCqo+
bUr6jfH9c9R1uW/VCNm0MAXX6lS9TNPrY3Rx4wpVb20KNM4W8Jk613J7nhQFM79lpSRMreuQiPMr
OsON2QPOLuDuJNfVIrWNajSxpm18Ow11xKJQAhM1zAu1TTBhFvRgcfMmAU300IUfPVdrb5ENzEZK
DkwT9lW69O0IpA34ycfrt//RbTw2//jICMLTNTgPJelc2axPBRC83EcfUCauwdiWO9MGz+4a+Nrx
xZBqKiaGsVuUQJ6vm6Oppy4WdvyOOmoCMDGm7pVen2jX4yVOxaH17NV8EIGrY8l6vKj/T1k5rVrH
NLeVkefXa7q13toOTZgXzZot8EEl6cOP7mry377cOOI9qvNSTzmE2alQuH14KQZ2BGmmQarAm/8e
dY+kxOlNbrJyFoJUXBHBNO6n/msk2R/2CpyodBsDbAh6nrwjl4GDQFfG/GQxDwDBv+xAVTh/9NUl
t0F9VxQla1j5slnDwhvABeLxDrLHcUGbBTRshylFhgA+a/0lDTSwHbYKj7+xcml2LgsL52ogMuyY
+1fQgLy/FRHlJPFOA24pYd7P/mh5sd9EM04dtG7HFvkamMDBPsud9gWgVU5egg0kyq1LjjVm1N+K
+hki/U0Ct5Az5NcbmK/71hhwAzqATD2ndQ9fVb6Yki32wGB2rTBY5opkEa9vIMEIPY9LUzCgwrMO
UfsaaqCtn6cVAg3UtxYMcrFj3r9dOEsHy9Icfkf1kjtBc2canVqM9labXLT4k98aSoJJI5loXoDI
jE/4up0X5rjCdFpJDtYJWt3ekMk4onw7vgs7qWGb4VprqGBrLvtnkAXu0ItrjQeJAC+KLIB7esq6
yiwUNp2GbSkLINhdv6pEEzX60f916eB8qfK6wgLiAz+tp5GktAdxSO0fSjSpwo51QlwRhutDt0EX
Yd0IeZCww2Pd/e03SZixOLPVy3JlTrCqo6omO6/RMIl2snku8UCLo0MgBGkbPk35pKHzWCMQSnL0
WuSgD5sjuZHiKajNRE3rKSatODGKTc00ZaxMT3ldWbT/jOqCCKL10WDos/qLxYHVhTRQQntXnbbz
X9/joDIpGHpi9vTVbGXDi+f0Hdd9Sg1S/sINfrPJjKAF1tzQGkb855gtv8Q+0FcycEcu+fnRlrAK
63StP9nb7QYIyCs8nFlomRYWjQhgqxC/sD5YW++qaLXJC3AMTve8lEfFXEQEWMLWPYoxvkzGm+PG
cZEWp/3LdjHIukgLm/BVXSeUAf4Rt+IgQ4tnCd2HHX55ZquDWm8sN0swsEhnbE8/dEUrWcR6hv0G
TE4I8+MJCs29W7ihm2SYY8SldzXW2f8IlDFa7E/lOpnhftmFRHztU2ufi4ZcAPg67HEu9m/A6Kqc
lCuTnjqmwfFFhRBDlxdViDK5asn4fT9XTPt0bE8sS9zYsaKRiWlrB5mIPSXrT5GGSyQISRtf8UTE
Z+2iuZJdmnqJ82PLubjEeio3wZ6Quh7hewpoTqHxMTB7Ytex8LifdXcAMMZciIKdjIEuG5Yr1kO0
Gk3gEJn0KvXuoHenH6fq4omCInwZY8uIaOIprY3R/5zMzMBa5AvjAasaXtAcdSXdcBH2X/52XkJy
kHQYu88Z6HCN6bKIZxO5gugcP0V7Q8uGsp2DcYAl1XtSDxe5DjLk3m+VuIScrgMvizRDSXCWyga/
EZ3Tv6G/r6kexwvw2nGKgigS0p0StCwqi3G9UFdxLD7zaGWbIaGWNpjGfEiNMELhguAOeV5iIo1Y
xqNTjxapx4AHf5VxrQr07Al4/ub45QUtZ0SZseUJkU2d4tadAldSHH8QCn9z8NyrlDJPvVIxiHb2
UXDxuJNek+SJspv17os45QCEQaqRoUVEPJ9AfzOefNWgjShTp5zjdA+vejgMoT/fRIMR5V0RhqXW
Y9ZTI2phjQzNzyFamoiXNcgtMhp6o9RZ3BWTwpCbG/FyZzg2JBUK4p1s3hRjlqRWNrALDjiaYd9A
0duJOYBo8D/ggD82GTe/VJxH1K0lfWA7n4dxVUUBBmqZH0YiXJjj90GqDDqlZlDqcg4I1+aJPhz5
/TS80AJSbqACD56YdNug4SKTT/pjntnfcKgy7zWKvTiQqb2r4WscpNXjnErZr4l0N7WPBvELJmbg
VntgJeZh3AiqwISnl3md/oboYk+qcncWq7PWcpwuOS6LPWygx7dYY7dEO80oVyfSlqzVhOf1vyxW
mgBV2oKXl81bIkpP3rES8NxYcdThEHEcv39s1KFB9ClnbrfCNSB/6YFzy1RYp569wbMVZAyN/QCb
MUidral7zOhCaSBYDmlH5p3ULubxKke1jRBzENSxisNZ7H6o/gp2pWT/VhLz1q8uaVyMQGnlVfzG
Mr4kbJPzC1qDg0JTHYHgU3ikPCR7E18WsUDptFCGQ3lqiQ79pqMZ4jFBkqiQMApvGSR86hfOkRJc
PKgfee2e8nIY6p/YVvHVCw6laBIAP0ILwJs4jqrZumuRiGvtnMGjwjNy82dVNfihR6cSXiaQuBVN
anoiTNrvCx1dbpAM3LIT2xOZSKaVnr8w1P4/5fiZmAMQMfF4ICYVkUg+fgI6L4Se6t7Blvgi+etH
XCD2l4cnEpC8pcn3Nr5/O+ZypMtsAaku4vD8GUb9wHudVKjbnSQDk8ku+AuicSlT2aV+k932HRWc
Nku4It8w5ozkCIkpKa+3jR4PXXGdMe/eJqu3c1k9nMFMsTSFis7CeF19We+CuuF84OuFoO9bPTgi
0NhgGyCg2zNEKzQsLH1xyxdtx7Ah5Rr1+3LC3yW69jtdtMu1s4Yt/2BOo4YZGBR0cpGieJVhtK8o
naGY9CW00tINbDdO6nw5yZMFtDjiwVCWQ1TMqla6DodwFLWBrqIKMMCZNyiuBzXdjFp39e2W+tDx
OzJyJaF51OOoSdLfPVFRYkoZLj3LeY+wh+5XKdEQyOWuVJX+bvga6Jy02WuYmCxVsVcLWkh7oB+H
2+gSVmHygf85h1vxvRZB4Q1a/k1mHeG/+HWWUOPR0UqnuqGXEHfkyK6hEl7Let0InOJkDLwQGG+n
aOoLfRh2/dszSv6pr6tiw4JpjcjZJA9PRG83HFkWm36/wQ1ryCfOVxqaQSc8MCqfViW3KiH/DjPU
fXmUMu2ci7jqLlF123NOwEZH9L3/14uae5xyAmP9Yk1Y4SaTPsV8sXodT4lZ1MhWOwSgklTsv5BS
6pHzwTJcJ9iJKEDeoYJ2AEAOxjRUdjn+cU6wCD29fhYabOULZcuk64MwN6nUV+Np8MIeyCrm2vQQ
zmeIaPf/gyK/GMBANEo9FbpKJG8HLcyoeuDx3MaZVRL5Mbc1Lv4/0cFCWctFruL9FlyyC84WAgWs
EqfPSi31RotKMIhB2q56DHoNTrQGBVuxig5hM+LmT9QPtKu1/4H6z9MwIuw0fDglbEF8Do/Ifp2J
GOGbdJzpVNqS5wE5LNHdU6OPc01ymYI+t4xpf+9+JQ17r2LjtElvKphVVtl9FnkZk93LEVQrJuM7
yD04JYvxWGb7qHVOPhetvvUcxZZX0xazPk9CaYX/SNOW1L6YnSO3HVQxMGbwPkF9UdY8H+cwCi2y
NSxMt0JFyxhrK45EipIG/fQjqBtP4ToFJYTHywXY4Ct10VvoxorCTUfTzDz29ni4opE7r3aO9jX9
DVmgJtihfqjyJW2QbbCHgYFNqcIUeQEY1fJZ3vIK7+NN7DZRWhLAM4nvEzTG6aQzt1AJCFJh2HLo
g/HgoF2GlzRwpqX8U4cx11zLihVKRV9skshd+7NkFA4Woh/EE9fvfxYoBrGCXTJy8VFHAetPADyO
duKS66I3sh/OqxIxToR2lCumhYhMJMXpE1QnKa2tuKFfjlv45YlFsRoXtAEVhFx2Rv+HVJU4vJTd
IdwtPzVGgvQsooPaQK8pWSfOzk7fhIr3q3D8J33jV9CZrewT3AI+a69N/doL+iYiE9ZBWxTynwnM
nDmEcJs+CU7j18NTRMquMDjoAijmmi1DfE2RPrKx8TkJAllKPJfiFPgAdZdEF9AfjbLA6LidKg7v
bCK18K7jzd9lOSSvucbVOTHj3wMhtLc/ID5D5EQuXNKzBhheeCp1pkWDnkB1P2FnDO8q9cBosqW5
2lT04ZcRPvIgqfAkVtYhlS8pdxiZjSGm5PnoaqflFEgP06ft3BWch+WvRIivihNHsxatzRgKyIan
LXb2GXTLoGZdjjt0p23K9W7DoXdRbe0kNVsF0I6L41ArPdQGSSeB6EA2kFlbOB+pE3cW+cAIcGm1
mh5wy/o2SNARX/dW3Xm4VxOqrRwTkf2bJVie9NO+lTyfjf2jh7aumLZLJhk+reFq1xHO60MUJhTW
5cZZhY0MxnNoN99f8SqIIaU6NS25agENUeZtwe3rpaNGKl32BHw9lfLc5qBFfvsN3wEjo/KRTxI9
euhHRhgkpzZfFljsNnoxWSO2UhN8hqEfbJwApMgg+9WEckOSuE7c1lO4owtqCBca1Pu8nGeoPY7S
AReSvJ0wF7ZqJwlbn673YjHZJpMefOIWymIcYKbQz/4fO8od7jgNPYNEZy1Y2DJZDezi/+evIKeE
VobNVvFNVprfWUXCgvHwqEaRntrzwaUe6Mc0xLMvacTJvmPIrTU/op4NQxb0p+XQ5UlfcWQJD/RB
e4Vr8BDEZLAYkseURSEQ2Q9J4amytey+EegkKd4f0ZLY45lY74Sa0gZXJ7sU/G4vs+WaJjiPxnLA
9VWeFykdPSVxLSRNUp7EE7Y1VfYB7O6pJaS28HNxrkIr0N104tQmpVOXqBMGpA8XJJfh+vsvPHag
nnbNJu9PdHstIFDdOOp9wnmj/GAp+BbDsJX+Iipa47Zzc4l2QcXIZKDbM6wk6CbkBNbSaTZEdB/S
BZ2dH9y0PmPMJ5E3QWDdxUmB8bhQwEAn3xNwbxU4Yp1eHkDrP57jbbq8JCJ3kN3LWRNJPdnYntdE
rAZAAVkvsFNCAwoMyggAWsxOYijVc4xGqbZ2o92tur1fjn7p65kC3MwhrcIO7RB55Pk9+Yjvu0iK
AbZzT0qq9sFA3LfKlMWr7kyFZNzEXv51NspOR594h/T3h15r9Hz+ui92bzzJtwcevuZUOvMi14XX
9RCLelX+LCM05et2Y4O/xHi2kDLRz/uM/zFYXMijCt5Gtz2pVvL6qVmJs25c/GQBfdh+GdVnhYOG
I3A2knVoMFwTudi7SKZM+qcxHzi85ivac+KmwxO6GHC9QjgWGmR0N7Wf1rGoccTR77fTe2E0XLZw
xTWB2k8VkIRJgqpw5GMTJvBSB4uuNqYv5uoB+M0jbnTcUR58RYEPSHnNA78XAKrvP0RxoRaRfVLb
Twi4b6rYfWyikB87DuTRG+q44ctiV+Sj1eX5uWCg6riZ7pf/aQBGzOjSws+RBvLXu2smjPiZjo4G
sorMd1D/tFMyx5fRC/98GRiYsn7yBus5wdrDHZhp5WF57j/QjU3W6CzV/Pc3aGC/IqhaabkDEx4u
6YHQreejfj6ElhQTZ73riFf75ymiHlBVCBcts8HracB99hPvv4BrBVxe3qZ/nwUXKqq7snQ+nrRK
akRHIRlabP+MYrXUdZQBS385DSx8mTc0UXLigteqC5Jyalyj2sgbSAwMutWrITv/gEKXXik1SFYo
thZuAU8iQrpJr0U41BIvrGW+vCOEUysjH5TKFaeuMiM8qLYd8yl1W+30bZDoQuaBVy0f09wajepQ
vcJCuvn9UWgWfNH1Ua7kNTALg+4ZnUTi4HDJgltWd4XUHaetZSXVCVtj8fQkUo5CugamH5ct1R+0
dv7/YXDERuIBjLM0R7zB+/4MK+VMGV/3mkxY/Or04ol9K/Ez0lzcpl5eGEIYWImDvfDMElq7DrUM
BYAAQpG9DcOYxS7B6mMkvs70YSj1ES3UziLWC66gFV+pYYgDfeQ630RBf8pcu2mV1kPR99S/8Mgu
X1nh7uNurcsvM/1b/+qAgJA4/2dMgg+rzSvALeKpY6A9CzZy4KWRy8qHyBGFLHBNs1EbcAvsjHdj
GgFpduHfFVTzKrqvAyoJqHyp7M280HhJTHRH7XMsdjxs44IIjj7ixhhlPQVyyHGnt8Mq0H1/PT20
u+NHtLBmopHSN0NKPEDe59jxsl24VPqUcVPWhBW9RzK5opKB8VjlsxeMoWQdlN9lJAE3yX2MxHyO
GbsLjrhaDHhxS35KF1wXQtT/g36yt+YImBZDOP0Uo0KQDQZM+BaDABLmgbOCPRxHU7U3fBsDLb8C
0jneaEtBDS8wfmCvBc09EMHkeBrKuN/6KnoiwgYhlQuBnpKP+r16fb1F+NBqkbcwF+JHeh4XsFue
vu5yqZrn9Ymbm74FMxViqWlZ638RTM2aFEivymODizyWfxMuYDTKan1s18xg0F6wgLotYXD5EcIM
lqkymxAaThC4n1UlDWFu+YyZCbsUFE4p8YehWN2nxOhhH1EZzp/4qjaBr0DFs2Jo1STv5P41wOSm
x4vLMbvaTIdWSKtZPIBX4981vQ7QRvqDQpWqXRLFHhrL3SaCDIqaBh5uSoamE7m4DZSJSgTE4csc
K19sgV0dEZo69QobBEtktFtLyZ2Q6WbTVyyXmnnX8wkF9BRLqJWTSNlpvktO5ZJTC6EuobxKZi8W
iLPcI4O+1Yf4ADkwLNvgGOrZzJNY5UnJcpZFvKQDLTkMvqFhTYvf+oWZizOswrUZ3cB1WT2kLyXk
6+kHSeXXr3AfpssTT177fqYqSWEqFdnNN1JZ5toR6C/YArsg6LyKBg9sv3lqWidvukNUV3RXrPwd
g0BP85MjjY46HYBB8cGWskn5pWwoRqIutgZ3KIlg0/9E8WjnbKhqcqgUpmltYtqZ0+TJ0qKS9xnB
GkwVRlFjn9DsKgj85TkiuBiFgs00wchMJOvY343JUyqDnCj0w+M+IE2wBUTOhT1fxOlkthSbL3e8
yU6OyGV4kAF+Kf3+VYzPaqZe3O+gpTmkC08ZMJxEpiWewkb9zMV6zPHEs30e7tjvimzqMY2ISNsU
wYG9mLDgyxm+73KMAoTYnArHhaWDMXUnQVJ2dufB5E3AMknrceHUVNUzJynPDhnxM7/cdUPVJj2O
5OXVvYFo4gcpaVPvnvYnxWJbKz98OtaiKUYRgDSmpAjBLhTAAwWp/PpmmhbT9R2kdK+C6wrcBk80
yF1otIejJz7160R480Bl2auIRYP2pcCtJKJOgEsP6QXGnmo+HTC+pKa2KA3eHiIojPGd5/K7cOjg
T6NZvPxfCKKKltixutKDmgM/U3T4rpm0gWZ1SJtyiMSD4Fsw7UILfhRtCIGHOS9kkQBLC0BEPUck
5k7R7P6GCferpfM5Xs5xg4xA0dGafImqWoJZz1OcqE8xCntPbKCVMtGO36R3iF3za8iORl8JJM/a
UdkR9kg2R+RFMp1zQjo5qdzmBJ/Nm3swPk+85qU2LIpA9+QuSdNdtZFcU64EUeAekVeJJ5ji3OG3
lVur3iqFWsJYMa3YAtBUpFu4sG3QMvWltu1qtCvwLMIm/pqIrDvPNm+KmZyg9frrXo/hOSSg/YOZ
f+E318zUFLZPrjYfBLXpZD9jdUAdI7YzuTA3/tjDHYVyFvvBD5TRaI3+TvtF+J1dcXUA6Yaj2Mgw
4pNBgoDs+1xiKEzvLZ/vAGqHR9huf8dUyKN9WDzxQZKeeKbTxJLCZnxtLYL4NxqoItEy756BmS1y
vtCtiE2j/V9DXab0hL/I2Yp3+S9Ip/egqAsk58xljoU2snhh7UI1ChHGcz9cATubX63rtIWktCwd
g1yl/SI0XU4MEMb4BRmphiOyuBHGusGR4XIVGrTQ2BzFTC37TLHpOmvcfXgyT7g+IsUnf/zZVks/
NQeJNpXm+mO5w/xXtHA4GpbCPvpZvvobWFrUMo/mjhEOPmiqi83JekRmh5jqqtyR1wrXqx2SRF9c
SENYijK2WROnoTYs0e7TJRvc0T5UsWSkPM7BAd+W4i6TFqwUArmxAqJYPO0mt6bUqscgdg+ojfbh
T7mQzLRlm5k0TMmmdQRjxB74gu9H8xtXjmffu0egX+hyVdiZejnLkvvDvZqI51qT6Se0HGJ4hzeO
qNNBn76uvLsJj/Pv4uSMY3QCSWEmy7u+6WLMw+SphVEwL2zeGxlQFmosEXAKFsDMHJ3w+5KHEuuN
Lg3E6PruhIV/QAUsFkAew2cvhhJEFCaLBkBZ+Nzux/zpAX+jYizJNnZVL+FgXM4xG8lzA0yk5sBt
NOjYwiXcqKw9BJEoDzk846jt2aliAAAih0U0dmlz2mzY1rh95ysumgJmxsNYOYBogtkee5CKeidh
ijTfDsZ2mkzymbrt5RQxs9Vc8MWAhqEolet7xMOPMwlsp0T4S/7lOwxllbe027NrvUH3tvrfqVrU
X6WGvNMXaHMoBE5OSHUC1+7NmqojaLx1T+OiZdTirmxSwDbvYJi7VWeszLk1rn6KZmg1zV2y84HD
n+2gF2Wcfw0pzEj5qqCjlmSwJCvucxDDqreTcYBRIKCJUDFdmZ4PxaypTUs02Jwj9eJIH0uQ/jvZ
mdApWusLTTcL+anHcXNI2tydBUkIrKAF0YDkhwuPbYV2hKYonBQUQnuuy3/KE5Z+zsBHVjoZzvEA
1+z+ilKcTzdST5NEOKkgs6oA9hRJR2t1PhtIxAdKatlIj5Q7J7mrsmPX2dduDZZ4iz+qUVM9wt0M
4/1vWkxEz6N87JETN9NTRaYGdSlA9hfc8Om2dU/aAWVn3vo5KY4bK+HqbwJa0IGBumdTI0lhb2Ss
Jm/GeTaKA2q5GG1Z/bdkWybuu2/xf09QPaqKDp/W2ndemeWRGq08RQmp7bCzFI6hsXJKlZOPBx2m
6BI3Or7jUiaZmJ6iDndlRuV8Zqq93yxfQ4GZzRCcuXEIj6mR95RsGG8UTwZIxGD6/N9CviApKjUq
Uv/84WAkds7dr4C2AeWLMLLjvsIllW9+RzJVyE1diWBFMGB5KXPHWK8rne+xcZTT4XzJCGZyNMrJ
ndsH1E6K4uC/u2tIByJ2On7D7+UzgGrjucrQZ1Eanx55yt9gyE83qP336aUI9nDOdjiQDRk6Zuk6
3Sbg4VagIu4452kTsBQLHvjlkFjP4R5CHgYU/TJysNOuURlhB1Dnu3mbGmegd1b9aUdXL+oM1RjQ
T6fwSTBV2X5DAUiFHaui7149WHZmXxGrEO3QRtXB55VKpfJBrH4WGOlKGveVyQxqrwvyahRZXGXx
FBo0rKfWTuJpICL+I+neTnU8If1ODfwU6t2SQOmnkEfKvJCVSWsqNmcEZtjY9oUEp88RnBb6zsTG
ZCvHGdgO/yr2rVRRi0Epyam+cFa4Wy0nNnCCfg94X4q7/0VrzAvztdXV11Aj9eE/UmYutexqQKGu
59yBJ251pDelnJdV95pAjDj93IUCc7zANKMQzg0KHKn74UF7whl9pg2Ri9WxFRpgZG4R0yg020fg
rJH/mrjlxIjnfRmDxgj/djwaLR+iUVPokNtjsbZ742OM0aR2vuqRmwhwup4NgvgIWFdd6Cxx8gsr
kaiQsW3A8TI8M2yNhy2wlZmgM0IAXf+pHReJzCDZ9QjwbKCfohQMOGsD51UpH0IA3OZOiCBoN5IS
UN5fBvIAtM0Oj2yEsjPuupK+tAbW+Bf2CgtPhWvq0msZ+jxlMrqul7eqOVR+4Kg4YNFMwCgT78nu
NM9+L8DQ19/EY6Z3cxpQbQVMsILsokqjN2RWgxsUKkNJL+4KywDCw1GByv0gdXAbx/JsgBvIEcEK
2qg27+mM2gT9FMH4GKBj+OJwGRJMnlHnIdc51OK2nWvLEoJQ0Oq14YhygBttI4n6RxDxEfw316xh
0HF17uTnJR0mUCtTpAuFxQsMNedMHeV1h5bp/GtMNfS3pKu23TcynQ6R+RDV7/sj/5RHFq4PMdJI
gNzspGudEo9XrHaLlPI0/YJCMrV6iuoFVB4AenZfF/+vKDnlINR2FGgszjB7FIi2uPJBJVUm/a1X
raNjG7uqDROb3Knhf2Cvv1zqi+0Q3X9TdWSB1dHiEpjtoy/oRoWMv1BUmy6xg3ED2QUpaxE5ZFA8
C+BC8VlmukeTCMXC/Uc/3Pr5MLA6XtGHv8zmfPDMILI87GHQTwzzp5F2yRxgXrwnjOsJNXfWm8pz
Jn0i8uJNyNRV5s2xKQkjvEeXXGzHuuV6VGIDCFAWOd8SP2dzM+e5n0Km1WPeRv96wt3y2hAJYfKG
0l1R4xoLMj0N4dtDG40bpYXI4dh96iddBGOZuFkxmjkpN5RFcmnffNpMMSrRAZKJSWvCgqnDNGvk
90izogXRlKFrU2gACa+aBuLQzXYcyowIujaZrLJ09ELv9gPrHSkzPSU7I+QpHACqVtEs3RWMgona
twsA7QGTn+BAysg6Ftyj2y7oYsc4J4H8UmNWlMyO+Z37sa31cY+OTyUiIjq54BMORjlO2cgWvVNB
f8i9mRjGu2OjZDzwkQA7jj3GP76GMi0fPqrPjrm4DidFX39hOBP97cEVaw5BRqQzMENdo5vRlZ0r
JpvP9W+wvWZhw/FoeH2CYZZUO1/dpEyeBBeaS4JCpFj2m+/JxcqGZYyJ9BWE+q7G+osfZuAukaa0
KurqpSoihj4sMLq6FHwx7brGBp/Z+xEtqcjszblUaGH40zzTGRdP+s2kBT0c1S0pG+IXttVAaOPc
SkW5u7hc7K65B3/nUNOo5167xJWYtp2BBd8B4sdcu2zuT1YWbrAep2ntFRD+uHIPS/dHV8QcCeY6
N1WufQizybN3hbJlZix1R2tsNlEt21UUS+aM4hn0DxZ74VP34yLjLJh/0YodNHacuG+wRVsC1Q+9
X0pfCSDazYkCe2UGPcEpZg06yA5Z/0rN3fYGWf3cyEmMXKi4/HED08ddGBNQW4UUDws3xykEhXUY
hNDfys2WSVYjhksn+5w5CUYKZxsDmx1dezZsFGnDEFQCWmNBrf9FNb8TDHRtGi0As+oarb2aaEvI
meAy3wLx31ezscSSREoRwEPFeTlFrC6Q9vMOGCbHgwfBDCXeK0bO35oX09hyXH9WWJahYa5QtazD
NoW5YVLvVRLdeKabz19bhxY2qrjOJzQPSZKjYjk8aO9mZjRH7Vxh5qh1AIoi7SLihAh85Gukdp5c
9T2L4CnxzQvG7RXfeQwC3JGJKbDDguCRtGQbNfj9LSuOoTxO2PDIAHXzVn/w/4nPj5VtLv+rs3mj
AYy9x+T3ciSsixhhRdmxKrvCZDq6Uifnkt3OhlWMuXyvpTnJ/jf3I0qpevHiDSxHqyhQVtGf/YhA
j9y9CJO+1HWX+dGmDlVROuq0RV/R9+5U6SpHU0tXKXZzEpDIgjQgJ8H65rqkZ6duzq8oOIsWfSVP
QOK/QstMcOthV19IDblJW4MmeK8MILloBViMk447EIyf68tLbNBQKvZ1gblYMYXoVFrq87KxrEEZ
rBUlUzLY+g2gQaEyrbkV7viHAqrkpNkWcnI1OJXFtvnJ99/l1R35wpnGusz5gjGvCJO8cjdcBjA5
FvlMjKxssd0wDB+tL4eNy+nR4cOosXsKPuO5kXPEDr6JfNLPygrYvJHirvZwWNErVyziNZnebz1u
b6fkDBH8WgIZnxjl3ZHCma/n3E2TCehYkiK3CPs6uLfBKzTb1ptSpN+zzECi4lG+yu6stTp+jWT/
PWfJXjwMJvRt1xDXCJazKql/397MybquKkVS1lklsjN8GWM/UcJy/Ihuiy2YIptosjYQq3GY8q4C
FulTLpOclBfEYM2fLRFUw3FdJAwcMVpDkiT7BZg8sMNLtJPPYOPUSDVCHkrRnFzVDGUFfguBX3hV
wzFgVTnvgKQq0nYcILx+he70fISAzd04tm+KwKIHZd/7QzQjZ3mMltsNVI7GDfSbktRU6CsstjeF
TIPPWFZbQcX0UBQcSkWxL/lfOwbSU9gnwvWcrX9SOMs4uHOxaBmfpFNoipgpJQLY1KMJrwFIZKrp
a4MvKtOVrPq1SyznxlklJjf5bx7+kPVm1+XU7gRmNWcnTej0OnmPuaSsePd6nX34hstunjnxLdYE
XtRXWk/WMFQWG8Q1AJGOcTR2bDoVpv1Dsbfl7Dw0BLQCpl9ut8h8e+g1GcxaRihoCg3LTvi3G+HU
cUb1os4FfxbUtIbR9WyRiv+zQNrXebKLqtXap5G/xlrCDp9ZV3MjrpZ1i477didUXXAB7ij/Ay2B
wrxSDwtr1N46zsC3+Vg4a/Ypk59pbMQTD7J/6PLx/y+9zpxElxCF+qm3tIbsqV3vQJlx5ekCXSfZ
LETh+A/FV294hFqUEafxDlK2NNKMCgLDL6fL6NXH4u5642w19XoifvcZy2y4jXl35kSbjeuuU+pY
RWnlVesS8ROSz0/u1W0+YedDjqB0KML4FNCyw3dtv63I/kYRAx1I7etNg2ZFWAVvgzn+k/zreea1
BrwVKk3g4Mz/1zxgGQzltFK1kqpV83ozMUPWXGwqYcWd/tE4zga1RhLKDd1ikEVV1uhItUuudsM+
zb/RIpHDHtgT5LxKyfRIcL1yP/GMKmH7s8EtjUWPpwFZAgmX+mUVgR7j/JMh5JOShH5orEfh7rUy
/imS1bl9EEj7+Uuk9LYrGF8hy7YxAC0+PGy6+ZIAAvaKyMX71KjwL8qIOEi/NdqBWI+yMN03emYL
Ka30xz6AMp5CjJSs7QgKTk2dvlLjGOsZ/nobewtduVfP0bsHmp1Rq3CsMrC7Vl5eKXvWoRYWJsni
tN5XXp6uzVNk9QzVSF5Hh1b7mbdTDPjYrVnHjJaPppqZAe6Z51vHNwVKlNbenZ8o/A5P02HsujCb
aTHS9roy+2BA1HBlx4SeF9vhCUxC6DiFgX5Kf6CR2YJDgN/pXsZ5yvFI+MH8m8LsZ+4rCW2mSiVe
LCPO/DPSgwKx4CSDJXWzQCRouykBLtx5D10G0saxq/mu9E6Y/WB2y6iydEWCqsCj2yhG3tlmR604
iMiu2mOJUFHmjAaIjC3ZoBQeMbQSIb/UGfoJkgCwubGDIy8gG/Y6BmmcNWqEeGWK0jpmKzJpyOmq
va9b/eXVJYMkzk9SI+73d2al/X7H5JXFthoAXSPff/+sQ8yyGPuH/jDpPd68XHWxlAN1EB0rcs1S
wZrzSwW9xGSTodDbeK7tD9AySL7/y4QIQurb/gtUJsa2DSf+5FMl6FLEhtF0rqYnwrLB/2trozmN
8o5RN88tu3Y5mUC1rHjzeweIzZUb5iit2dlkVSOmf9flk2skB7a24iuUWF16ttDzPbHE/deZpUW8
1dELmSU7gbkQnXVt0Z8JOEntLMiqKw62Qehh84y3AW98XnQokODPSYkaCd5TteDbi1wHIumnX8kl
qgcD4IOoOiNmRG1IpJ8WQlTO9FjlsV0oPTOw3C1VDm2UOEOZsFO74m/woHKGUeP4qzfrE66d8EAk
Qp79R3JZHb/strzopw/BajoEsCfhcB0gu8Ewu82vfKMCZD+HxzOKOfziHzJ8+ZXB/a7QGGUIWbGe
jzURpyE0wh140mn54yzGoqlV0ySN89mltMX7eaWPZ51lPzt2GQ+yJvcBM3Ntr/3MWAjCdmyLFz1P
Kp1Tr5epNEgDx6wwZSGwHI7vlLcepSMGnVbsaJA03hPPlYXedgJ4+YiMnl/coMMGhhaUJHRDghsn
RvgLUbuv9tVbO7UKdo9A1wCfcG/ajPVlG7ep67U6L2EPgOY4vl0aF+wbA9zEgQM9CPKbodqNVdLA
8t7gtYuRZ52Hpyq7Au8S4SZGknp6ZJ5M0EM6NjISTogzqmreGmBARcjNGBb9zWFm+ONt/B6WULqM
FZ2aWuBnIJ9HPsy3DuUzF4VmliASmPrNY7/NtPRQivXs1URcU6UBsz1CYgle5BweKaqFbDk1J+AT
rZIBTk37IPxdjrCuCvcrN3kNSP//iYAA95RU091TgSQu6Fn4ENhr8uAHF3YyP7l3Q4Hb9+fn+yYx
k4PeZTc3fwp4XuIYR0Bv2wrWGIe83GynhtQl45e49BEYWFuR/GfhuW/6g/C4fg7qd7fQX1m6cKGv
xAsL2mwNhKXg+tSzGVtkBXCO+43eGiU4WUo9IhAkSg8FZiRX6jThT8qTd5oA4yTDtQqe+1IejcsS
Fff/LbltMLudHJ3Gb6T9N5GgYrGvbGbYY6edTaSGn3HS3exl9KRi21GfqA6bjjGRvif24GTy9+5Y
htaGeUzje9Kgpql6lcmFh9+RsVGgtr4ga/KCKg80bkDhs9FkcEtkz4VdABa0go0QnMj7MNTlK856
f+xzE8wK3XOjF7MN+yAoZKPNtehv1Jb4zp1wXJOQZ1VzWNfOo9CuFSzpgpDEaP35fX2CB6as8mOS
AdjAzz8v0xClLa+ADYctffaSUDz4DdqMY4whQ1ZsJHCgqMIZOugeh5FvD+cj1sthbhNXgKDKoNHY
F8jKOFbcRqKiyZRvj0xUyKPH1Le7M8/ewVdPACKzGWLlgbo6TJ3Uujih+ZrrjhrxJuwfd+4MWcEP
Ci65ACuOrWJOwwxyjr7ImFTneDaqThE2eW4By71mS1B6j6EDO6IlMtZn/LuMwBQYLirPWlisHZXA
EueA2eIHkissMs0w/FGe36LU6o4J1cpbFaURCXc7BoJIDy5ssAcVrBMTrcBiZdg5S/WVI4++xAE3
BADRZCRp/cMSFz+3z3FBotiXN2OHXD/KrUaNQo+i3L/m/gTjubRfgKU7yYn6jX9Y+gQ+24d5xSgF
0C3+il2d7sakddcBoX2PtOHc1hwyYyLqrIZDZd85X1mL4Jh2wq6xdQ2pel21A3g+ym8GB34T/TnP
h6RpRK2KlCbd1/RVZD4QcfLLnAFxsgpTKF/OSaTWxrf9XIQGibCMS2449vKQVj1R1WutfcuY5jCD
Q7nqroHxNAh7XHjOZ134dQn8FbFGjC2t3R8TKS2QUna9VK64fBvKvgSXMxocLXUnsP2VOoZkHZ3l
WAP07V7R1/rDh+A27EDhLKK5guDLSMbFgZcLSHj1EqPle77nr+5Ygg4/shVItb9Gcx2h+Je325Rk
3qFqLENN/Md9KVUGsqLTGuh9wDEpb0bGzh1PnyhsKDUuZ0ts2Paa9LLp0/VuhJJQNZfVTKrkUJ9m
HHh4YhfGkC1IvDo0AoPQIGL0KWfbe5d6zOg6wuEBToM969qgYBZP5mK3tqoDnkN2x7Lnv0smQP90
OHHlf9+hWlxgMx2beFmMbyvNCzs00q4qyWYM3AU/3tciLwF332NscyiqGk+aHkEfat8YRpxSsPC9
uDLrrvn0E4maeiGIAZee1HZjQOLEuPL846IaiQ5BEg+j1Xm9pfF3PdYcgCI4mtx/YauaXVNjY407
TpbuH0LSY/I2oLnOIOVcMdpVC4kR3rCiaujZjY1liJ4noHW6uVxssFD45sBi1mzKp866ksI43KMe
cAeLKBLalU/JDFp+LFzIOWLIuOOrlqcsCOtT7DHEVYuWJteBQ0tcCM3ZnosEAprvhQSmJ4H122+M
E/2hsYhg4kBokav5qPhpljr9Dv/FEOTQ+s41Gf/onr/W6n54ayXmJobwwb9ZnZ2K38dOBMpCcOXx
ZAlA78dMffh3kXgdxxLTYK0p2kNFS7UxTMhM2Lxy4UtVkus34QPPuW0Rj1Lqv7Lmj1Wo1wPgopYV
PHczrHEDozm2E9PYUaxPVvOis6R0kYPNB1/QhJjKezk2WwiCyMK1Uk/qpIReoDZSML6a+Yihko3x
BmuEOpvpSQoGctD5o2ZJ4WmxVML2ZhOkZUxEWD1zSXwECGqAgXhF+dY6PilcYxhUoK1WS6J7JJ43
ghtCCtD0v6LGxAt9uN6+1339AC/TIfEs6BB09HCopW3/Ss7qaAxnDycGIteHqyKGRNCKe3EDEtQ2
04OzttTZvxqvzOqJNmHGz9tKchwmSN2Ior8L1STaxmTVnrEnVznRUGXtYlC3eTBC6Dd5BuMoknHr
gdXh4MUQiu7y5ee+3Ra2veZSxAOE1ram8mXJMjjJvsYs/fq54nFscLh58fd/7bZyUHUgSFNO6CYp
Ru0jm0RbsmRiljFEtaeK4HthDUXK1R7/FYUmr9WGuMPaC3YkHlXbiQJsbuivGbTDbSlNnV0hDzdC
nzGYXBvD5enEB9LnQzFZz9YuqD26FAnWh3wqF2aDi3gLFC5v790HjeYFx62XYKkJBsJWgzf+luzk
FTh2Mme6My5ty8wzPARwyUP08PrLagbzRcdrwqVS+IxiUOs7tWZNN1GSVFoDKzlPELtslXHdeXTR
Sm6f/sC7pummM3LdaK5JnvBgljEVMRtDxhBZp5PfqmH8dOmVsjK43TctDcObA+6ZL1zLILk3ejre
JKa3yFvgglmUV6hjSScFA/+hgAItZG7tQVOi5DgKQpJdn0MnHD5zLqYr8SaJzmpLKDC6d2Yg0iE4
KylCp7Mg7xUwdIZxVac/E6NBdixQQI6L0qY0PijUfTMGF3gtWaLUFa+9hXS8Z4lGw7SwM86iqVi7
V3A2JA+9jU0XGsbSHuMZtbux88dQu3Ym+YOEaL31cudp3oBxEOHORiEVw9cWYQ7qNbF4VBxGBYkm
2iPyGaVALoUcKLlxjZVnDML8IaAWe8GnArtiP0ePUbKklc+OBGdKr9v6awTsik5ZNE26R+BDmEGs
LymryqfLMLeT/QuF+P4Bz7OS56Jvg1iIjQp4YlBvQA7z6nAc8AECx+jBt6/VJ6ZrQu1irqeLOEBc
h1eIv9Zim1iTJKqVYoODjQ8MFUPRWPHVdS8MCtPdrf0cqfeF1GUI9Hw3fu5ccWEhF/9pcUgRwZTZ
yA6qCJDue+9PmXZZoLfMVl0TS3uZQ1Zy0xnOVAUrQl+fww3TxOVSF8AcmBOpfmOhzxBdoUMqBmvf
XIJSLUIzzH+7mRMHaLUv/LW6NgAkCHYDxXV80tOFxpa9WtYwYyMAcVNsUIWzyAVapMOXhIou9Hcg
HfIHCTUhXDwS33tMyO6pjk2yDrb2qOAYzn0cKZ3MZVz6FtP0Z/OlqG4NVwrC/juGOfrsp/HCXft/
tTt+e/KIh8lq8e6+yWcbJ/xzkZHvpwO+gDBZ+HuXOklFjZT3egSyPemPc8Q5AWzYqSs6LfiCZ4LG
lflLCB8qAdnQ3BPPVDZGcnH3R7c4JuQ5ZAqQwG53kTzcGTInDwssj27yVZXNdF6pli2UGBOtzSp9
bTQNNcacUz+xl1QNtKVq7ZXgdyZ7QBT6m9kQnJh7ODegWDjZend6RaFaOLpLERsaDjWhKr/3jSpF
GaaObCc4emaV5QyiPuGUVaGU0WoR1efy2G61U4TaTjsyn+dAe3bKHiojKxywszjAD1zwKPdBHHRl
C1r6hwfMy9sGhC6f+IqDBwLG4iUD90Zu4XMQXvu8HPYdgUkPufo05NutAxGJJHE1gRb0L3M2S0oC
RZ/RWMIvSZLo3uINO/1aYBNq2AUxJuI7Io5zJpO5OVtsYYKem0Pl5l2u+6mMBA2vuDWpFu2UqY4Z
SSb23+l4oODPCW9T/HfpaRFinSdpXkMHE1xsm92tW0I72KtZ42VggSZMGxG9eg3YThIfAbFK+2Pv
086hTrx4d1Dhd9t+nDrDwmBpgZtRWsY3rciP2CGnN22OdfKP8TWotzGj9+CFlx7+jeSiQ2QTzXbA
UA+xPxKvS+aWjQkfLa0tPqLw2ppqVa+IzvaszKvnOcPsXWNcAVQM+cd9T2ku3mf8udG+HnwRyoDW
CNzZrL2R28nXfUZ0Oh83DUQ2a9sbaqQ+8s03Q/9ptiVCjFW2WzeqXKUHvyGHQJzRS+3Ah653aIN8
U/c0xFq6szMaVah9ErD4LknQedO7xpMu7ZhCEUwB9bAAdd7g+5kY2BJwE8P6ueAHlZHE7VRwbmR3
i4DCl6Gj6+fB41xDEVxtEis1VAC2CqIEOEOhId82A948PkiPiMagmYy7cpdJQuTdY6Hvy4v4OBdZ
W2tr8Zfe87RrwmfCPDksxRZpiH2YrnhxBoRkI2Udv2e2TRLPWTZJtZIsg9ILDzWun5LLhU85pEVa
+8gOiosLkmZrTsH3ztYscG95ec4VFQ1G/hUWrT8z3996gZt5/zXQAXXdIWMc1wG1IGwq6TnZ3z/o
AICLh7V0fmswv+Ch1MjpDgvCLZtBGBwWuV+fgcZpmt1tcVxkx+id+e7ZsyYWrH2UK1Nq1zrchQ5k
/LriNwjoHtmg1dro+7O/veYT0FAmcrayzPGGmBWhoLYuBFYKOOxKHtze1T2rmemdfTiff3/Mf+Xi
uBcIKFujwrjue10sKv33n4zZlLoeUvleHLzI7Q2l6CxGPolgcxqnAWGiM7f5jxnd8AfmikohUPQQ
JVZRCr1TVa+ok7r14rWGpAH8Qx8S2CIe/jzXPg1lTM7Z/Ip/wj7FT46b3iJuPJIWlUqAbC6ObQOZ
/h/XCEjPvIBa2gVjHtXU3wG6xDoSiZjQZ2pNfX0W7uVsE7oetpdVlagrY75Qa0nhLhzly5Ykqj6c
QE6lSctZsVYgiluQgpSnyRMbPnqekR7W8j/R250XIWI0wk9m9a5zFqOJbmvBrB31kzb8NHX6kZJK
ofDcfHaG4lRhtPvcwKTM2CfXFvIph14CrlmY11Nguv+4HOsfW1Ob+1jN3eYioK0Q1RgJngMZhVcR
WjRA36CYLvFBrzH1m908l1kn8Vj18gg662NnBU2UMAdHLbeJK0ewtG0hxR6KMe7eezSv9FAV1iZZ
OmJxF7jvMN4bniAjBRXOpu8wITmsg5KAngdeB3JeooegwfcuLe6hZuCYMyWUtRe3qlE5V2V+vxw4
i5xc11esM+QdmIZQF3iZPsLz0pyF8mvrOK0zUfRs/ptng3aoSQd5UK3O/2x12o484TL727WwgZr5
Z0Tu/uBVjud30R2xgVXskrNCj5wl2KrrGXjgb/zOdJMqXIfeLsGBimGdjJbvWTYQSsEBN7UtSm7T
ZLMKoU+89CYm2GI8DsDYoyfwk15QChFJTzo8Dv4O943DNLUxKrvp5iLL35GEoiYvCWHAWxQcMwJf
gaD2wbudDOkUIWCwpCLmEmm+2lKNqXicPeTT7yJAR2jd5/GMnh7MSuxJJKVN+opkUg4Dk0UUpvXn
T7W3nK0mIgCKWIKnfwogITVmct546MtTwdqMmXRsgffeFRowTu+ibwMLQY9liv8gOhQrq1/J0ETr
ZJamvPKKBmwrbj31R5RpkijsFaI+7cYO1smk3FNOyDYWjg5ZHg89wgJe30g6NY7hBF95AWoy/7cW
3OYZV2MpW33gW6RLZYP3YbHG6KOWziXGp54P5IBRiKRRmAfUbnACiuUuVuXtVLusUACmC8wc7DOl
2bOlyqJaEEROFfMrGgHo2UzwTvDGk1Qgjixl7ZZmYkNMe+s9XiKNXQ3TiXA/ltObpyya7ncOVCRp
mav3Nm3LWRJcE3VLqryG1dJ8M550L1txo0m1cHgHyiQH0uhiWMzGoOOnBAM3oqwiEUxllXpHFEiK
9ZG0Z8XdTEIE7OiFUQSrf4Lzs0dSGVc/SvduqyO1MgJ8ImqyzI4W5BVK3Wg/rMMMjn/f2smiSlgN
/sRy/4mkEiBXMgL7sGHD98RHJEpZa2izCsV/oag5n813nTm4ws2MDbGezPFncc98DHj0CCFq0Zks
xKDypJASE2gpycNEJ8Hnfb3F+T9JBCgq4Dcm7hyHi1tT4hRY6Ws9ZpeUn/WCQF+zPmORCPcP9dQb
g0OnGF0yMaVfiqeyyX4CXR3bmYBLs/COD0zMriAU4RiJyeoRhHgqbcV6byq5VePSkJJVRQR1dtw+
632BCFbcMRG6/fOqImCGRF/xzeSEwSMt77i0pIAPKH1wml50WTcJEaK3oIzNxqF1onrlIQJIU0ok
BQFHSLbCNR6u+LEyBBCLD19y4cEQYtfGtarIxlArqOcd6vy6l90Y81KI1UHXNI8hRXBWz4OBRTvV
fc2YK4Q9Uxp2Z4nron5BdzONYnbMzRStnGHUCjM3N/GBWZtWaaIcmkcTDAh6Ts9NjOXJe191Urw8
Rqkhw9jDe0ljQK+ZqD3H54p2pn9EvdMgVJVjYq05RSAWnYiaZxRjAukqkADTgT7zHhhGjpv1RFvZ
SNrY0IUdGMQaDbnVcqrrECwrT5wXVue0ubz9jARxmst2wjW7JeZeX08Mo9+c/kk9DWprwUrNbB8z
7yFEMDt3jlYTBzZ4YrLuEhroaYGfvK5bNc0/7LSh3Ktk0rP7hj93tmRUTLIL32+0gaU0F0e9DnTH
7+14eUn+FxuNIQLLwMR5raVFJq5+uVH+czebgp2lourIrJpGnFGXQMZv0bwnniLRg0CsXO9BA9i2
5TXAKJsNDwJYz6DcJLsuLqrVm9jdO/dmSoZdO13zruGhG9qSFJiREIBhd2MfyIOLwXDuPG9HZPq3
dGo1ZouKnHpdUfs2WeZlkJFQTlb97EyksO9vGxJUbTG72Kbmu/+BXAS2O+hXBxYgaYhixUGaPHpK
qA0CbOsn06wBykJnGBdfRcjy3ktc6/MtfBfS//+JJkXmXrR2iYL+uFYkqWio4TsoVWff5OWQl49b
lpZJB6siFOMFrgbPPsNSeG9sQw4AuSkHLgPLA50ZeELJH6+8WS9/zvI7eqDW2ry0XVDJTy+KUQCP
Zz3RscI0FF6czZrV7NCo7QEanLvNtfngbvsyjhCVqSBcZbzvRtvg2iXnjlTWMGStSk7UH861wkWu
yxE7JUchnd0055K1jgXNQCFxEwORnerIcAWzRV+sVZDR3CHINLNaCf46J+RWpIoc54PCar9WorwX
vMkI6A3qlxGQK1H+L5XVhh7Sb/cfyotPpk0sCl43TKeL/QoGrnaPeVwc3r0CkPAUGPcmtCJX+Adq
OaT+OV6J7Twpvn78TvwWmIzzpO7gc4wbyHlq1kuzEN43QKzb9YNkI+VKOfSG0O8UX/rt0sHvklRD
MCXcgOImxOxG1O/pIO25FLVIzUmYZpWzSdAziY0ovojcMdB6BghqMs34froRNtz0QQM4cnCfIqkd
ZhLZtnzCxj/Y/YiOIFzj0RySMvfOp8dw+0Yy20Ap5ZdVKWMmJnpZzyz7yV17lstW6h60lj2b9fkw
QwUEsHjR/3O78OWokMbKW82ut3BRIHtY+ooLOYBISNkhrx3ugq0iGvUUe1R672AYpSgtaT7efaLh
6Rvw8JKevYmkfCZNokpNSHiE+ZTUrKV7aY8n+9XG+nVuCZQ0OoFp1a/URyLmzBKN48cLoJxKba8A
5GTPLxXH18gyZrbeDaQeMZvDDh1F1BAbGFPFpju/lfpKI+52hYcSQNKXc7teKm3a3FMFKEDwBx4W
WFx1vuTDR2jCmYI3gWnH1NmnwRbanY6TbGHZwWNkWZ1ouyMoe4R6qTzyueRZhbHrLbbzrg+/GyDt
ZgzQ8hTTkavXRvfDKmxIugFyLnGeGSesbtPPllAKRh1/L5syueoYnZssKVOlq3GymqfaySf1DvM6
OtBcnaYccst6sGQKdVjpbBFItu6ZuDmZ7TxglGTIXn3D/WU7Y7J0rmsajSLwICO9ryprv83UTphW
cnNsQKy0wpUUjTwoCmlz632jMXdsvhlruw0Whi3BW/evcr1cx+MPfxNcWSIE687gZtnuzs0SD1hB
BM/Tvnbv1QWgnJEr4boAZfSmXmBfQkLQUKi5MNyN5wZI3u/9JW8ymYuwwvyuwRkcEEJBFm5rD050
7bqq7SmCmd4a90E2cab1BHPofqPRRtkLtfLnXGK+x90rtoGneY5xt3wO6sOUyi6LuUGsmjiqKu58
0OBYs6325BbgAHI/NsEuifpVxF6WEGaHsIhcnt+06cZGuecAGZYZToqhFfbkod2f2PvvadPxlyce
9BJC/0lZlZzZKpg6QCl1DD+cwymPfHlIXqCZHBAduO1hySL1QGSKpoX+GCtCHu2OJQMDjyJL/j/T
JI2TE2YLiBwgzrAMMeSF3tfShTVGCz77FIklneY0whxB08zUpRUcXtZzfwsj5qMAOMSHj17BfXjF
KqFuBiyg+2OtD6WjRLZHSvn8zLXy11lrq1oRmNQ2KC5IFjCNH6gYFJwLAFOVa3FUx+C/9itnPlun
bnSoqQ7mZC2jocW0FOfvqtiCsuw5MGmlVQPb3EETbiS8D9wxYerkmDJyCb/TEE17jk/2Z8XUzwgD
+2TF42zO4IObyKbRY+b8VktJz29ziDyxM4VxWTlOPIo9No0jB6ojB7l7mW8KVYbKbfNsRDUZzA9C
jAZei7ccM0y4kEMEWIoYw2EtIiQ+61zK+mgFsf5p6sK3gjHhpd+Ud4WV8TyQJn9VAtcPfGbrCztZ
rkCVZWkPDiJoEFU2x8Wkou9JPab4SuzeL9GGTiA4Yf2XfKOyokEYpKa1F2jpE5j5sigNgxf/wuZT
ubYXAicHN4crqN2YRDrOSMQWvYYfGy4DLQnZzePcskOWfa7EZfoybq94K1qzxoUdcwDMsGX1S5uS
GqKxBUfB3oblPdLgYmS/vPBnqhuWx/jO+f0gowHLVEKfkU1ZLOvBJWfbg03YH1Jir6oJxl9bODlI
7w7CIt9ocnFZe5fZqLzb8Gh0QpodV3clB6pHD4TSAFdqaU0lJ2MRW6eicNWhw6+MS82w8gSpDEhT
r+tzshE5xyEssWBTN37SJQsYQUfvHrxYR7E2cNaBdDe3IABuV7POkE5ggW6JvM8MNL1gp7JqUPF4
STHxirll+A2Dwbp2vtOO1OSotR0CgnY6cEz166tG7dasj1Z/0CmQrTFutzQwGWmQGuOYHoyFh0nJ
ctQMTg0YupeVo17b7Uce+dJ0r+Vv8eJOFogWdsh0W/FWj17rqSrJsTsVQE9sg96m6J0e6YjysPLg
k/u8+08JxXH74H/vSiAL8bCezzNgy5l0s+n/zErPpC2pM0q5amL9DHateFMhfyTlLxdc1CJpl2aY
BrZsNVtNaa7e0MJYqPrSbdVSjJMvji/E5bUkgFUq6AXinjBpRTBTWgVsoBcfaaqaFtpFrtX8B/XJ
vulOZm2nD5FlTVx6cdK8pVqmQJ/NAlDOVx4FpbIDdvjjKMIGcn2L21xZDg1qBsf4qeEzqPC9098s
cJlSe0yNh6ojmWRxzc1AaZQl2MchnFgnN8n2RfVvgS/gpXuyRRwQXhRPhwwIXKsXVU4keDgWE2D7
TPzZsHpWl1CxKCLWA5dcQ6CZedxWnTigxNxJmcS7+7eSOBp/5kdnoInuyWTJkotReXwi6uYoX/KS
kwuU6ot+1XiqcuXG3W2xswH4tFe74tsjDSFw3zVzbOAdusSdkZ1WbRACcpgz39WE6uyi6bodCRM9
PyMcGZDN2vYAOl9tY16GoNWOQHT/lG1mcGb1RDvfT4ipF14Eoo2cKsgo740Vyefpe6w/Xo9VZyMy
voKTz55q/bqIvbLPyDTJuy1F7RH/65RVK0Cm70yoztM8WMgR3QqLCQ4dM3/kNa3Ef0zUWweEoc6W
RD4ai3BBe1TvuBGjIFQ/eI+OAKAF9dh/mDErUN27jFrI5v3OzuV4HAUkBvWL8C4zFy5uGJS5xPRj
6KVCxlQ7bCpYC25kZWS7E7vJIPB7r1uAF3ozy1dUigEID57yAHy60luYRrhJB+adI0wFte9nuDRM
h8kvunq871yIcJx5eqAIu9SC/6GPCEGr4QxEzgicYEuKYqUjhkVBPVf3rfqv5YY0wMAdpgRsdvL9
fBojhe9mFjGU4QiQWqU8jTmzSlf24+YP9x71NZ61+1OM8CzHd6U3K6Tc3gZR8nvvEbvsixYtRSvn
jl+W6w2o1GL3AcfF5Tw4qXPgCjJP3xQg7/Hhe4ui3GX/ugtoEwGSKljch5JTmWNZIlwYQkxXQeyf
XmxHcq0o1Db/Xt1CgWfycyQWuWMMoRwnX9KCXB1OdDcA0h6+OsPeh3RSLOwB9/c6pLY3+elIGHhl
neaMbGD3i+3BjrtISnutlFuCXSyrMxt93HRxN3iIKndYMJrzEl46FwhyPDHAmMMvx3ZnnVsRJW4Y
HUnzW/umHonfUd6PYx5za8sDQWk4++UO/TUnyV5bYyJOYsJAYFv8hY1s7pIz1TZQ08F3RWu6FP8M
hshd1wEWIzy40NoJ3rtS1NARB0srTXrWsCJ+msTxYHioL+GfJw894N0RrENw9H3YjAcqSgfsJ38Y
8kRBlvoMxjbcqZk8mn8J3u+rlDPv3KWtgpHTW/5VeN7PM469rhOl7QLDPoMt2gjkqLhwzZceZmas
o9uVrkphIM58L0p9Orsh2VXvSHJwGX6jCSLNmeEPWZwuzPsy8+/Cx3XmlzugdIb9lfzzSVDlyx4U
Z/MEwQ5fW1u0NSZtupllla8lZxuKWrOJQnBBJXtCRlLJeaClCvFwZdMSP6UvvFcGqIgpCv3KFLKO
p/AXDFB/YCUk9ofHQVhaLoWHCRpYrRqcs8tICYc7bGvE0XpwPfbHpcEMRCX4sOgfx7coHwHROlR7
okjjx6eLzjZu5uez5p+UC65xhOqjhgyXOezLUWsnpyW16Dxu431wEaKQNR/viqig7DHLdbJsK9dz
n6MtwjExOL9uPdJjp+XaDdF3+FhSbzNW13HbgaQf/LcAXPcnqgi7IM8xsTBj6d1ivnIxfFdz6BHg
4cn0Fw0PU0ooLmB1Sp4zpnV/msGqv3WJC6PWdG0nQ/BjPhL+THxUVqUhUmLxdgpdMMIj72ZPrYv5
bC+muSS/Pd3A0nTPYOes9JbSM3nqkZR9kshGx331GOEsf+ZBcXpv8Nh2Xz6QxA1oBXyKY6xHis/s
lRH+qjVCOl2ACya9ewJ7OgyozqbGm0o+C6Pk27aZ0dlsFLRm6FJKIn6JUX0XtF3XOvZQ7OT03Yh6
w1jN1vfHEsznydKYPy6TRO28oZVTESJyta+EbPLu/ySiM17LTFZZtd6wEbJL6nTYzL/hwEcDzrts
+OYt0EPb/WhtBzazDxQ7Peiy4E7aJ+EAXHo/aPpSQMEa4u9VA6dbY1jHA+GmbwK4XzouQ14G5nrK
GDV0jibh+yMTkItfeyRpZuGdNEDAfvG6JDKSbQxZXC+MVZgvezHzHlMvU0YEbivfy1CxTG4lgW0h
Z1Cp5jsyjVd8yi2mI1vmK4f4wsWPt9En4NgwuxTyLMf64GtzBbVgGjDFR8P/fH+iRzoI8u2K7Zcy
F7C2jClW6OoqeRMrmWa9EmosOBaJTf8N54RZz4XpQa+zUJu8Ecj/8bGB8LrmlARazGbcbTZRhVHd
resQf5BYfCuSKaKy+z3FeoB8WuIyho/t1jvtZMs5uAoux8BHpGqBhAaicKAiU4s6/sBkTIvKAa1t
/+buuGX2Djl39OdVVkmk6aH4TnV3Bu+h6nz1U1SsaCI9K590piWmGBrWwNVf19Awe5cP21Zpz9VK
AKSbo34R/1jF0WLbG+mjcOZjFEIXmp4EH28BF3U83GxQZqmkhKpvhLsxLZchlrGDiaBt1ftzwnHG
VUqyjQpeKfrakVQymVOCNYorVA831l7Rk6Y0n+0ZFx5y74Yx+Lg8+mpyUg1CKc2au/fqVay0sTlB
lNdU5d7Nf2ehKcw9x4tWjVkDEh/OCz9prq9HcNl97kOB+YD8aksBVwVD1XedUV2W7nUhNjCO015N
hzOLihIZdjwkkTBcMgky549nYVmZFmhxgLnPxeiOC460BeDWIdht1uXEbHDLn+0bL0ODJjfodNOO
Zs4cRdnwK7VySFCvJJykISLDYlBKAa9DTPLBqiDz3qswgpEL4Ca0waeLmfgDJy/GnyVlrkjOLHjA
ntCifkNts0fpkMMLGG8YjKKRILYmE3BIUNAApWuMQ6CEkroRbvDAgSjNwbXCQV/IAhe3gHiS3sUu
nASoMhe+m8pu5FDaWHvakhbe8MOCzGz8yk+XO9IjvFHMhRfGk9KKLFVr1ewPYdwTAAOVShwgzKwf
nVClAUcjzAO2284jH9324I2TwBoDBSUS/GTIGGccvTAM4h26qwfKHmfKMXly5FGw4KnmYcfI6FbS
AitnwYAyaUk4lZSErTDr27S9M6UrNEc8xAw1NE3uo6ey+aat2FODV/3uHHUF7Gn4dBHGuvIHvSm1
bb/bm7PDmic7Ko30BGDjptPKZ6qgv2q4PJKc1k3I22KxQQNDVp4fd0Vwq0zRCwyfcwgR0eLeNYuF
NAqfgukmFGp/5K1dwNemOw3uahmf351fQ4yZa5D1PjZQqcdlY6TxY0DfUu6UESlaPbejmPzj+Gcq
FCu5DG01nC3c9jHWF7f8T3kgdoYCFdn/vKY1sPLFWrkaXaBHqv0QdC84ZtVQYOagvDGTjJyjdnnw
4DZuTtIpz/H4cTOO53192VyjdTHpeYp8nlZPtOvCxBlrd+GUqRatf8MsGejt/i7SFfoU5lmak9cT
2Ado9FnWaHYKNz0z8XUj7iRVlIHFM667Eq0pHNrYyprPShR3CHJIEoAm05jkAXZ+B/D0AU0ti3+A
9BpVRc4V+wUJosRk8MD/a9gG+u9bk8i7CEf7mFe+K2HUkx2OnGNFE3xxDETWkARfeDZqH/fGcAFI
ZAQIE5VeB16r2a6tS6zhNZrzlK7yB34lEyaRIT6GbuLFNQouL98b4xQpjAZVeaMjuGvZAhmcS616
MWEZWQFqQo+ySrCqhXe55expyFf+ltk61i/jnudzxRi4Wh4Digewhdj7+5k4Z+ZBB/TMEckDLnDQ
mHD7vV9ndUhzAuyCEs0l3dJq7GyllS08xXS1aVp7PGFjGlGmZwkNyhYB8EVQf7vZmB5T2axZTlWW
iCARb4DAi28EU3PexUAQZbJ3nHFSX1ACpnYE113fu3otY+WU8WDU1FbAE++Chnk0S9v2fr/gfLSE
teCNzbAl75AomMbXosr/mieZCnTQgViGlrKV4DfOzrDI+HIW96MevuAzgJrl5Lf/ATmDnE856P8b
krBA270ETnaBz/5b8Y6ikATaqjoCJsgdm4uYGkZ9Znp5IPshf13EL95WOIXG2kAjpievC7A0MY6v
u+TaQbNMoXpp/Pw8RyuoPQ69WNl1ezw7XhjVjVHkkiISYC4uND7v4wKHjgMNWdzLir1zAsdbqbyN
e9MedPL4Cizje/t2MbaDyU5hHJTbphJpTaCncH6LKt1hGuKQDt4NGdPAWINC8NSAr7PZq6xUMg7A
119ubV8St2VtL1q+auVDUJN9m8QrsfjjL5Sg3vLrbz6BISNrzdKpA/QxeQ9bXNfKuQ+gx4uvu3qO
qocG/+vVoFjMAoJWUEpHQuHA4bnceF7ItRJOaPPKXRK9l4Ew1xj/IvzZ2Rw+7kDH+9f8U2/R0xCg
z1SSE3j4RFl8khZ4G5vZF7kde/mUsjcdZMapFXFevtLp5NuNr0u/EKfie0bhcxkYkd+bDom5L8Yu
wUk0hC2DNltEo8D39j6H8u3dGo6ohiv7kK6JOy0RnHE1NvesyVKQ3S2gEp/xElCC15OL2Lx/eQC+
A1/5F2ChO+iLn9MHIXaUfFU9cZK6k13jSbl3o56T/eE/6CbVa2Sq54zP8NuZ76cX5svSsv3qroLJ
fFdo2D8nkQyq/JrA61tTR+TyubLHcrJa6v3NDogGV8+J/DdAxacfa4qP+Eca11Jnl0b3kX3WTkHh
pTTrxj/HoEnUHikROfebbfWoY3WvpDIImhZD1v0erldqYSXpXODciMjVMBHqJ49PvmU8vWfayJ6P
V6yCH8DyH0X2tsbF0J+ROQR+K8kHg6LWAtdZMpdlIi5UCPf+NIdvCpLYQPAomAI24Kl2SpUZhPxS
6iEvysmg6PhTGyMJoqtx5nwNpmqSyu6rOfh/KucDyOXTusSVVROBrlohPcpQ4KmepPWhqwTecE0L
cFitFxlxp3kTLNfMuKOf2SGUSju9an7FJDRpIMX0zZCjOmDX/pSd0zqG2dpIDiYl4QiMpHZ89/wP
ceio7yDd2uWk8L3zwOgo041Fh8kWQ6Q8KMGplEfaJfLlPclhqU3DYGbBWbeWce0gApgY1SLZJNYL
viitYvlViiqF9aO201uvXpUcGCoTVp/43SVJJpTCyZd8bp47Knf79ZGbuH6ItKzQxmfy30qQJwqG
t/8LiGB6NJWgFZ2QhQ4SXh+D2PRzmlXNC76425cs9+LxRqK93spD710DsH0LfmWZ6tIY3THmdJ5k
TTTa7S0jOM4jw5KQr5IRcH95+W9ActNqcfV5BndVQeEQxHcgxS+Py2CM55oDdFFrA0ONDpAhTlJI
6YbHfwyjJUD6mghoJvevpVF0VoXr9YugrlskLlCT+iuhFZeyBoy9THBNt+7KFQmYfoKFeb8WlBCQ
2mThlio61/I/M1TjtZjiIBJUCm5sIoEjjjEH265a/fvTY9MXX15NOiWF+ySNkZ8rpW7POwsVcXjK
Jr65nsvehs+XOVnMlcVXW7mI+4zyYpJI5FW/o3OWc23/dd8weGnXeX/WUMIZdrTbP23WKl7sTw11
ZeFwpaAJTuTcdak7BYDX1wj5j4nwTvinKYP51/UTM/ubZIlrxLW6Z/zXxRCXUPJ10bYOO30qRLJF
dXJ9DKbTOLgVTXL1J0fiQqe7yaSHVGqxfsCb1HbLqc5ZfOjaeZuOF/LctBhAZmt6CbstOik4EFfO
HjszFQpVguj7pyWnTnpwN+1OfzoY77Rh3BZOxwkNv4c9oQE6tVWapbLKriL8AxeW+TgXRe2GrSR3
ub6ehk2ikE7D2VDLnAjIB8TsROSDQr/0vxitNanCC0iiDNg/xiXd4RTsKX6aNLDL0NX8Bf36cyM+
+WJ2p2h6FvMZilpxkoPvm97luRrqI0ktSFEu880QRDWoBTSpt0skyCx5GIECUgb2xJ+Q1YbqvqJ9
1MlguJsAK6o4B9f9duAapYGHUilEXQcKEfM704QONkmhctcttB8jJQsfHtXBNzwRIVkDj6pCiI1h
7GlEUM8WbVdD3mWt2A1atEp0hdhlsD99kwKW2uR5KWWJdJr/PXd7Sv8B7Il6PzTxv8BHDMG198x6
Yekzartng2gqm0MeTHY2/kGCA/bI7mWUImaHpow9h1EYbQCDHK+ESpY+Saskc4bp1FtsHkSRH+72
VqIIQLhNFxsybUI1X9CcnbmOB2jxUuaJXz/UzomvzasZuocnYMqeTk9PJWwt6vJl3YqisIfMYA1x
mcfq2nTF/CKHQ/oxKcR1y0HS+11dDMOKYOLVZOfYnSrQ4tA6klbUfOu8JnNcECb5N/eLzNlV7rVh
OzuD1nEnnvzCq3bczZjsMD5rX13VGaRW22jqcGaGWfSk1iu8SANMj11ckg5cAV8SqZhyVMzExADM
c4SHDEktNWx2FDlaBBBPJjU1Y1cfPsck+KP1+8xvdcXlqdDnlsm0JTSjSOjTQ1Cui3iJu2MxaDJN
Y4GZkKxI0QkQ6EyHnhIblwhw9xnaqxYDpywiVVXYPvy69kw9z6cKL3cPeHluLVdce61vR7kb5urS
n9oVuE37DVh0F9x8HVBfOWIPUjqC1uctETwCRozJaOtk3UEhGJheOp3j0TT0ASElrYcjr7h7KBOs
bmLww4IDqoe91g5y2s8g3wNsbiDhaZKA6J0EwI1x/PlXYTDXZXGu/4fkNTTfMpAYtVjLBhW0gEOz
SYIz8HfPmJUXDMXHMIJaKhxo5RK2vdieTWBB8k/FLPS33vSP/EXxO1daHfyX+Hdj3Jmj39vDSRtn
Orz1SS7p5s4ZxqWmntvQOn9gcWOfRZpsqjc/FcboV+NisGyhDOAyOk8LTEkH2TO5wBqEa0duH7le
qDkbRBQPOXEOobZBLVQ9B/25Bb5VIt9ClHJSw9RcfPcc6HccCkoJGWhFOhlWGcKPamGjDOqs2880
GXnl1Ugx7hPMdRRfHcqs2mTaZCyzBnXsp/bcedaVlXAl0a01KWofO7x1tsmuW3DFtowj+AvRiSzb
v5LZFCR/1hD2bHgjPyw60l4rRGhaz4vs1l88C41mGaLv8M+nhBXrxExNgKPdZWK3+MYalZH6b2pT
ii40odWYDo3ZcNF/iTBZUWzj0ykrgD78UfrI2oLWztjFjHvgOyGh2KH4o+nQ7tR9+bhgOq2eHa8Y
h1SNghSQULB6QRpBkIdIXC9+R3M83hNLFFs2sgj/M2TdbQdy2l4ML2VFS3wbcwWFxNYvaep4nZvq
iJV3039ksV1ZCRnunVm3W2AaDOJ0E/TGbTCLYkCzNlalB2EWyK2LC/4Xx1OKGLM0Rn9BEm1kwuc+
1ZeLwlRC1x4RO7fcQ8ub/YvHzd6CQYPe5/oDpHQPA2gT8ljZahR+DJSmYaIOfMFoq9UhBmFP2qh+
HCtTlmAk75mYS7yvi5zF+qn3A+AC8xd4br3KdR4ZUKQ7WAz5AjF9yp/TKKM4sCpjgi4SGYi8sKqB
4nA649yKuG2LLBWdoSC4FVaudo6pY2m6QRkzrRqGQyq0SmVtYbsfF6x89IsesqCa05ShsmJ4aZAp
v3IhAVmcw5Zk3XsdEme00Ji9pwESm7dZE8P7koiIDDISy5ylD/KBjQBXfmbC+I1ZLwF0jWs6sXW9
G48F+bsvgnCHUH903N5X8WReNBrL1n9EsA18nibXjU/sn9Q6bAkCWegAsCX1yLde5+SE6LBJ6xEx
b6G//30zUQsm1dgv2GBiJLeFWx7XS1gjWjMa3gO2sO1KRO7LoiwoVazkrLQfSGTE58WJqhy+c9NI
hKJs4KoU8H/wWUcQYixleSLcNDSoCBTpJFZ+kgQZjRU1BTyLeX+pztT1j1gL92mZ3uFR66sFfjUF
uTlJtH035L8C1dEgbkCH/xxEdHXODXv8NG++5kM1dtNwfwmX0SbSdz950rnAtX/tTdctxx2y53D2
eeyJASAMN8SBZxo/bE74IGkbObTs5cBFAK+v8rBSfX9go2yVuZWWVCpCSy7573LHzW24e+s1Pr94
3yNPIm8uEs2i7uE9kZNVJ1yQ8pkC+tRtxK5KbeoxBBrE10ljrKahXQarsPs50Xu4GnPyv8VfTR1p
kdmJLYM2D/3A61HyQW46J91rU533xFtrbKTR4SsLCV8Ay92wySk4t1kogZtEo5usT6d/D0O9Qu2V
+e7mQBeKSHaPuFH2LJwAjhcQxf4AqtdrJ3ZhgsAQKmF3+OdM3CmJ/S44yCp3ZJdvspWORStR4d/1
PU/7C4uWwyfQh9lINOwP7dqtY8iMdkocmoF51sSwgFIYSExi4t9VTzf3cBtX/5lTx/ORQ6vw1gNs
59Q8khkGjzz5npg/lXcNr4xLOriD7KF0TLDbWFbZmpchqSN/GP/n1e1C58nIJTQ0d8AFxozagvJ8
zrzkw+2TGzy65kD9QL/VflnILVE6UV/Xv7nMfwZ7ordEVEbuD6Y9Q5uCFBYEjRwFgNSTZJBLjyqE
aL/V92CIKf2nQvARBXAAEZoh55XQvzUA6o0o0DiYDXWQG4G37knZAGflVr0jbsK5ik9+wvh4ZVr9
C1WgP5tEz7dYkKuPEFz+jWAY1auvFDVZGOECvvQEY7TXeLVrscbZTUcYtvKNReg8ETlNCyq3Jfyn
H8HbX0gCvkX3/53wsB1bkHyw6sRPnL1siMDU5ZnkDUNA7egpDeZzi1AzzKNpMS6pVQ4GIZJB1NDl
GunsoFQLQ1o58Flhde6YZQKVbVxMBCPzt8/nG9rb8d5EMDnL4Ib+TRHJK85VTU6UJphDhtC4XeaH
s5LcK2UbJxHKmSFxflWG/+Eot4Fwf10E6xHQGDkE4wXWFbAhtluJkPaL7KloArnlcz0u2++KYQLX
MDEQXTRhYYq8xDkRCHrIJzmxIAddHpKkeXajt2UHxls5o2XTQ3rafvC3UC1Ygn6K/suwSOxsF7dn
dYxcjlN8aUSn9Hd4yZRkYq6xqAGlzqHnqNn5uYq1kQz6JzRCvOq4HqZdN1i/t//2e95VCTyAWeWR
+qTkILSdR7WNP7elZmRavqjOFsKf02s7ilrUcbs5YcrCV88xW2jFlMjEeeSpVRGXLTDt56JPvxPH
fWJawYYFMQ7iKTC0tcdOFtUe3pqJOuIPzJidIxTYZ3cKdYlmDEdDilLA9sWqpQ2TNkze1zaDJX/E
DlBoG9p0ErFwDBi4ftA3vBlx5HK1b1uprpZ5LHZ1B/qfI3YHz79b+mnoTSbm0oHWcdNphwtDjo4T
36ITE7w36np+lPSzlNVdtZQFdGxjdWOJwi+jyZrQ9sqxqhtIvQhVoyZRBklyeEMTt7eXLRwzFcEa
tEH1E4Gi4wny5rIE8beS/THXmSZgeTaOJ8CIbQb6USZ8BfOqo5CDClczGq195BeJ784AqEKW6fOJ
IiHZX6fk8NWrk3rkjb0F8B5LdgyhG8BRmTya2w2+e6fuydG8IGPpAyZ0MC4p0JQ0NOn2W78VCkJe
opq6FsB1S0DEQAPcCy/RghxtkBlsD190JFHW5s93kw3ok5D3rGS0b7CubEAnDLLI003+7YpeEVs8
cyhjGY1ptYVtOP5hexr2p1DBBEqTuUTeebODHur+KirxNtj/JLbwbDZD7PmYSSmTVFe+PUNpAP3D
V9tqRTEAXy8k+LS5XyrUDVYn1GTNn1lANcHBQf9N+TRi6Vlbb6VAYqQ6fmZR2foJTeBECMPmiqYO
urzhUZqv6yGnZ0g/Zn8UUWfdzVAOgrKZJPVXL6xf1Owf6ipvSfdSd3xtI5b3V2vCYVcpvOJ0IHLm
tgJqI6LDABhO6XP07qjvQJ5fObLf0tPNx0RHz5S4R7kQk1Cvx2mik24wpe0Vvs6wQ3IvDNj9LjqN
x3eEgJ9kuzk7otPgCALP2lSpnbpPmSe7GzyUmz8jld+Y49Y02vKrkF4raYV/qUkvJhyYmGIJFl7Z
QoFLv/EN8cNwGnVIfWE0C25ZCPuPBmc9nDYwX4qoJPPv2q2fFSzusIn+x5XQfec2kjKko3KQeB+Q
FIO2LYPw500gUDTB37t8iyPUcquHmVppdHBrjSwlZ7NwZQXjR3dfNAHrlojdGEszrceaWwpJvL35
HdR3RiksW47yEtNVoMa9AmZ0lApf8CctqhyCgqk74BQS/69/ZiVex4XoDTeQwR34uK0ceVcQkRbd
gtVD/tFCti4bFpoDzXwyXiypjz+5AZoiQdp8ohXvaleIUlxkV9ueWVOp9/9XzkGWJUoLczZeokEs
sQGTxLoXYFXA9mXbRPDFgyQdXYqH827R/o2/JzcKEuJfN9pqkg0n4TmtK6r2qyACz8tLHEiVrI+h
+YXzwIEomlvYGhwkaCy/xrYmYoveLclM0sp9bGO4SZy9c2SD1KS26qBv4eTP1s8QOZuX688BeR6H
c4TDT8WnS3vQ4tnv9G9eXjZkr3rkgmIjsd5KPMorH2NCkd1XSvQ4LHnqpcpiXzv3CT+c/df1KoSD
fnneb+rDw/2ZRrpNhVmGeJvXPimcl+kJeLhiRaPP8DcCJdLqG5AKDoX5AIqdrzQmOeQCJFqmB7uI
RtHsqy1ZmoXsa2NJsUBvJGz5l9WwdqysG4E5qvoLKNexICaZ9OP/NR4R/lp08XdNH6qtTufK6pln
excgGKpHCZxVX/p+GpIxxX/+ga1FAXU/9eGmSafgcXdEBincFGMoC5m3IzBfikchWfuLjYjmPjFY
UYj3rg75GRGf1D5twdNgeR8j0OydVTqrVVbfccL5mh9I6MGvZh2up9NyL3i9JpEvk8uUNx6a+I0T
u6c5ur5lnt0S4bP4GVi4j/WWnEoabO1ArM4CVwtnwnau7gH3etR0uieGD5xLP03JDIzzhHqY56CA
v6dk//5XPSWGTFedibNKIfpE0DoXp3yzpjjoNUFLdQZQmLT83vrtxbPEn/auJxg5p/h57vm89oxC
SCA0kkXABH0+hWCVoHhLiS/DTvIHhTBiOb2M8ids6pnPFJE0UW2g+t/Cb5iOkZZQQkLkvCKeAI7+
VetomvJ6kITGhuEEuVHl3GjRnH8OeyGrtUPsIrmEDYIrKWdYEEKQJ6TKI2sSQ6fRvHTQ92WWad+n
Dvbsi0H1fO8rS5Hjml/qImJDMbWytARdUb5u4nPIvV3eBKoTBwV8tN23iQa4bHhUDgBN3FRVYoUt
e992nJPHeQrOb2aFI6TxccZ7bHk4Vut0C9MnrimANJ9T01WbhvA4RkwZotX+0HeZBaaX0dBO3BOr
606rgtA/T3JoachXPKvDOqEikBknNe2U7ITo9LtjXdcipQTABPytqGKq+CfRS5w22Ej69CaKwYPi
P8VtC0ufqioEhSCAXoqZ7dCUGFAfTj7Sxfi58eSaBf9njNYe8ju6Cm+cWCezHAFGh4hd3ad1dZ9m
DE5/GlPOfnpQS0MbMzM98L2FRuj2bwHGrO8vgKNJEZXBPUgGCK2fq2cSkaNjpKi1hEtgC30DFClB
2jNdMH0sz8mUIn20nGsNkfec1kC5XGnhRoL58xr1g3xvtxURGdd2RbeXAkqw0v1JKIxSdukioDXX
joBPlO35EDBzJn/kLRtVt9bk4qzrl2H+ZfiIzvN2IaSXin8oXMKFiQNCmjy1H//2DYrgBCFJDrXH
B1Sg7P0rQJZqLajyNC4fh/cilwew0MBfte79fjV3A4I2Q/tqhDgLUZ0l0rZoT9egPUUwlBgSUuqu
95vu+dItKwnTTsJ3k0P9jNchnXpCU9RJot9MWRVWm8lG7ABMgaCHcSpf/L9piuUZZQzmC1PNz0ei
P7iSwIPKt0j1CVmOhbnsf53UCnDD5v1Fl4ZWDYYS16cnJhNczy2it0mrWeYdFqVSLkXJd7CGdKaK
j+gJoNYmD8qLhP7Vo7hBvh3ZrQowNPhjsHhi0iwBCijHl4i9ku/L2UtlU8k1Z/501kAOAbjKW7qa
y8M5O2NRO2l6HISLjosN9eebyFXB+zgCgzPxUJRHJ0EsIgQBA6rxdGP1WEIkBkdgfmZzJsqdQJjk
I0KickQmDVufgktkr+cI8ijWwog2hdm7Vqr6ewIC0sC/cx1fubLprLCMTVd8tPv0tUtchpMcMqQf
zxreENM1JITnx1kQvj8GY8QuWmur9uASlRcH/jQ2DzzWUZrCN9XBK0EqhJS4O3+RwnbAsUQ2Oa8R
s1mNmVgSsu7std/twv7nA2BoDpzrkgTOA/4WjeEkfw7NNW+ufdRbNmbjKhtzNO7uFtDOmQ0XTJn9
Q2SRE41SEFVFFRp9RMhKWBT181oSdDVGR+IgIK7P56NlP7xNO38FcE+kEut1MqYCgizHECEPsSxR
axH2KDRupW1Z+zkm6s9fMsmjtoooi0rQw3roMU0Ro5iD7O35B1zzlo5/3QCNmboszm7sQNmrr9Ch
jKzqZ4mFBiD4vV1CNKjHMAN6UCy3/l27JfIv4br8bu8CxDlAJTeTdiXq30wJOrYxO90lrD7L4xuJ
EipxJxU1q5SKmUcWvrig+rK1CvgGNBnjR1pf9r6/hokukQZ3/4RXRFXwaJVRHaRqyyiOkIE1UFiG
qjvheXomLN3HA+GM8kRIAzMbeLWkdISViAfMsvsoz+LIGVPXOwwY+cyFf+EXnUtIFZ5KlXZvneZA
Gi5JLdIaee+XGNfzuwTST+Be16to0F8A8USlVDxtUwGAo7oDnlxIGz7teRdbcWBT8P+JStjZ7bFd
1eafhH0LOOhe7EaPhsBoYuZwLl/fcreOJz9hPCjcxM/5DTG98XBjTAQW4xgVsZUJ3ITxNU9z7+SP
cb8OJqrhdGICBA5usPjoFw3KJijSjx8ujgxjEUO2K2jlQ+ZgoHB94989htbg0ginWmH3vY8Et48I
o2O1NH5iyeUFogG+jluK3c8DupFCGhE5ExKDzLtcVSwJ5+neKF0lqG7rj0LzxBdHRGr9vtlB4dhd
zZezr0YaojGfLIWlSOeKFqpMR16oL2kDEy+UQLH5xR/HXO/EC0sLy5onc2lBe7lbKTCgEiGpCRzT
wmiU5XxOgNeixzigDedl7TxZTZs50oQUv54/5zuhPjY55fdfOarVHvYrZcAmT0yrOQcYOGKWv9vY
Ryl61FdckSM8LEdyNMqhwM2nfDI6FfuokyUNBil9yzUCcPqdbZjSgA/dtQ7jXJ+38tqfg2dOrLeY
dtq0BAeVzxMjCoe6KQ6D0MTqv5+JvnsUGRpU4zt9W7UEzx4OF55fYROGjL1p1/C/n886VeWBt5tc
pQkYK0nxgORHapUei2aJkFfaDO1/ZuhYztYLkoNuBpvHqo6V0aZpHsaEU8YHr+waeTANaldyoBMk
6MljuuQXzxVrCrKxUSjvUOPR/DbCAkwldce1w71HU7jPxeH9PqoiAB5fEEfLn6UyQj+vr0qy/Z0g
3Fkt1LCjk8kptdC6a8DBPdP/jPntJouQagTBnPFxXQOKz4d0Rlt2Z69w1Ph6TyLmI1BdQNOeD1kS
ecv+mr5jtvtWWyws539ontFqPiFnl0oRbj5fievIGJulzKIc+a5sxf4SyVeTIevQuOK2M014SUEX
phSO3Ls7cHmWRAqiqabVpH/dCsz77LoGzX2tUsKa+lInP7r/XbRSRHN02BwGMDobQASbYRvfZLtS
zgVaQ48rfo8izy4kP4+3Egi+KJafA9vbSnGMf6su9qXJchGXZz0fhYaDiqYwyjGGEYR7qa0NYHCJ
fGmNhZ5bDTRIvZJEwcqMtKAabVPO9YeoVG+ZEsn1kugrZutEQFNdWYpqoOHsoDanmkmVSCw/KlDd
YD6tNDGXyDLTVdN1yUgb/rB5hKN+PWuKYI/a4mfVbGUF0QyXEyoDxz+b1v/Z+S9ItnIryVoNZVe7
8eeBDxiInhxIe+DVtwOTYCaeOdHZkgYbrvYmy+bGaXTAjt8CR/LNtaa1PsxX7giUoBlaRKLT9dI8
rg9MHyj19gI67iQwLYhjGX6v12jZcH/nQIzEqUY5Moo/kA39iY1z6m3NTCh1qvbbvWcwLFk467W1
rMOC5LxkgEyKJQbEQZgN5NC6Yw3yuINlM9Nit2O7OHZPbq2RVkY13+nD91ypmCSWjzvxPP7aSGE5
JbvFw8a5ZTVA/FZlKe4b5JEsVYA5ThmdiYFS7vuccPqvf0+7eUbhCwxoMPHs8qd3kr9ePQzLk1A8
TxD6ShLUDP4fTn2aImzg+eWYBxK3huxRyNQDz9xENYQDHNPV9j7eCX4fFpVYZujUYVcliXFkslKp
EE86rI3K7LxVhLkj4skPJGfeHaIXeSRcDkMuOJuZI61o9o0MVja2Ayhzt4GPzxfv06+6G3c3pOAB
Go+I0/rS+it5KQDDUS4Wu8IT8S2Bikk+x7l70lAkDA/D4AGL9ImPceK4QiHUmWEZYpeLtdSUIQip
avkOAB279zkkr2BT8WYWu3utKvhViZGyUh9WlKW7+LAE1OAW8GiKEEU30mM7QX/2DAhoftIpX7er
Sq6OU3tyVzTt3ebtns7B1m7wp+7IoOtKnoateWi2+hj6OJKoPRCWWBay/S0b/WJZIqh4hcZrD/l9
m8sVtYZzBVdMit4e7v1wnjyPdLrldLGHYf4wb5m3L+4wmgC/2rtxSJb4QRncmt6NFOdio41lPJTs
4Pm/gDHs871vTGxdiWOH69OGwiOGMaIJLQNKvvmEsz/odc5s7LUxOjn6ANKHQWWTPIqnXfrjn27w
7nYbfJyEWibV1mOpfhFBrRQDW4/AKuFORh85N8h5BZ3NO5uOdNZVZMf7yYEI8IAnX3qC74+v91VS
Tyv8c6r0UpQx1RdqdlpmIgJLyF5xeEhUWjCV8ZsJzg6kxU7YACeCn2nqNXB2p8iJl57pSyqsJA/5
fal1vifj9x8Ti+IjkG7Y+adwGVpAX4BfZ3wGhAOkk4JNy1MaBRM1I17gOwbEt5zdr7GsxEBp1H0N
ewi19Af59SDpYaScWOIlTA12y8TxWRvqjD52CCL/O3ThLNQyO96RtnNLZdCnxB2L/dNEFgvo9iuG
Lij4qOUwACbnj+1/EvWro2afJJ30w2N+k6uicfN/+W0B5FehuNdPxqokrogtGxxbSyuEsGoMYGgW
FHsBpMtny/ra1/+aP+S/w29MCWYwTQY6MCT0Te9bWVrj/a8LDJLI8t9hOK1opB9wZLrFSm3JdPbc
sZ9mUQRP/Gkz6tv/D3JyEZnIqKCLJoJJL8AwbiVCHIY2ePIGWgXcg6ygeJ10j1c6qY0teBsLe9jY
W58LVe8r1PkY8pzBwapw8H6V71ELoydXTvJPJfXwBz8WQyRrI+l9GEiO3G70vmkF4huhwWfLJOle
GZyeyV0NA6mFa6FPrplIhty5KKyP2ruNmzC/71sV12LjMCWjPF8gDEG69QH6D3DsoPXs6bYo9z1G
Un5LNwmNKYM0RXkSNFXH2gW3015n0HtYp9avPAh00qSwqofpFfRoc9Z9FM6MltKr/J4OcQcq5qJx
Nihr7mWEWe3YtquFeXKTrzoSSnf3Oaie5bd35jISeDEUrNqBdGbi8NuJtYND7SHwmMtQ2MIBV5A5
4U/af7R/Tc9AdQbCp63rwIVonmRXYaavlEeF9PrW3R5qqmLI0twbeJoq+IUST3BpIGoue/di/l//
0pfXPqx7dHYXGTZn3yyrYlzc3rRhnMaBQ+2W/rKhsXLWDiFuFUJ9tvJneHIesFwHnSFfKooI1mvp
t3vcehPKR2rzQerZWmilnM19WZyKDWlgRM/i8fjW6SBW8NxXK6LtL5uJqbzHavRXwBvquMWhR04M
2omneNv5pCCwQTtNHSZnlgG30bS7TuC/yqLwKcYQ2X/05boL/ypu2y2yJ4GxTGkvKL0gZb5ZXXxs
Nmt/8qJUUTyypKN/XC5t12QOrtdEBXAM+xSydGkjABXN5ahuWs5yJBc/sHuRJxkSYgmXqjp5vUun
MGrWOF609U9DOBUij+s0zcX1FD17Ol32ToGX8i97xQOvMXOPog7F/k93yOZzFEocCFFcjg9A9+hg
06lcCCwNvrAOcyOtyZjmR1e0Qf+MI5eP3zu8IQOFbJDcrHLWwp1hXjQiovsXhgaydHaglBooylXu
8t+yO9UKdnie/2+wMFCrKeVy+uBaMnpkdTAma2uwWXWQ7ZS1ZAYcOU4Nk5aubf9DpX35sa0wP45q
ZCdN8hHkjdKAhVOLzHZo/GT//0F2l0ASxmvqJgvCUtpI7kHry5HpJQZ0JFjwQjS6x7ZMWP+EFSf/
GkLizhGIFQkNT8mVAFnqdt5LJOkEGqRGKa7zVU52TVRm9YMT/hwZl437sUZ7C/XNKYWHUjdYsnQg
hmU0m0irxoIR6iQmYtn4tGgQKOpsna6yOtX9Wv0GB8lenjJYkYV7gFhsUf3fqaYbyU3AbjhDpYG+
RLxMUUNItJQwDICKkJCLe1qDFHhsHaTjd4vYZ6oegEJXpdu7weGXVv96KosI9N0gKQj0rx5+NUk2
PoMUaFiCy1OkC5OyFW+EB8TSYJJm5I0gRXf525ZS1fx9/jSOC2BxZLYBoaGUcacglfBWX/IA+/j+
v3/jVDFbfPQF8tnLkSU64TK4tFQY2hgBJd50V4kFnStEpdHD6S+T3/usXSGRRy6+qupNx6Gy7lQB
2BkjZKV/+LKOgYYJ4EnfhF/X99iu7FqCSdSiw+YBYh6bcqnSp/Kwo/YXbd4ulh7elWfkbX7c4y07
pPGHmHxTFFAxdHPR03iIhsthe4xhH9KhsfJaeQjdFhtPs3E9WQ8Lb+Y+idtvnrVZpJSF+kFrz8Df
a8F7jdFMCXtlYuIRfyNr6FWaD+z1SOJzdDcy1rUQ72XRqvv9Z68K9YE760KkwvDgt8iJRaiOGRbI
HPqhwi09x7xeZld5iOZNrU2hz4C+FqSjzPJrEyOeIZDXztfnExtqvegIk/qwElxpEL3QwE1K5ITz
TWti+/JYFtoFxcYakh9/czySWzdI3p9c+VG2rKzMUHbYL12VhrlAwLZqCv8HLdsTI+pR3OdLpqHz
5+Nfd3TLO907ce6376m2FDR50Pl0GD+4fcfeU9d3wARsmjQejCxOKUFaX8vbqFGykPZ88UmJrNH9
UnBDeSVMcua4CyJRCZWzuPjuict4MHadbD6jiFHAKGiVHu38x/W+TrezAPBWXGio3JQVWsx0EoYG
8IK+40fdVb9HbY5dRLQ57v0OXUENbBYqV6yy4YPuJ86E/g8CP2qFLCe61bThcNEf3ufAB9Bd5CBb
fPGFtvXGkDPiaOSa2Oif+V8zUBtaYPSNBuWZarg+pZZuHlGm02S5XdGt0RlSDBtFgsuOUpFxAnvd
jKxE80BFLIR+oH2KTQ4A3VHx8yJ5caf4t7SdoWp1V+9/qHcNthpspHrNouY4ljSqbKLmCJ6kKcEi
BNldqUw0HCxB/bQrsvzW1omgnhmfgrBiqH/6QP6lDEnmt6ZbKrpzNeHPTLqeZOMsTDzViGRMm56h
+kEVeNNda9qjoh6XpTAAcfTFmCc+gcj66zM1AtvpBy6iabDebEHvdIoOXv6+kfEwMq3iraI8J619
EnPKZg3zDX6KDrQmxN9ALF0OVomMpFD+04Aj/oJfj5RLC4ihiXlaUTsDbNpkJ9pZY4ghOWQzoai9
s/bh4MWEeHHUBgPT71aod5a3Jn7PbKyqm9Ge4j6vxGbH95EPGS7aASBZr8n9/lYine6mx5BhvEGf
43AW3p9f31oIdZw3TY14sR+BtMGsB4Vd9Ql1KQYkRWpU7rgy3dlBtml+xW7wCm3i1Zb9u6bDjvbD
obW+j8nOCL4iIgvE9TavG/+UlVfcATOy0Yb/yMDeIwaz+SyFFZw7PxUMaByA/uI+hJdHj2RjlGIW
ozIuLc9hOpU7c+iXEiFfTqqUnq/rjG5PQYfrVN/U6o7L2184RW0aGZdDieD6++cIjIej3XofI37c
1rALCfnAe3Wvbmrly12BjCL6ZerGYHDFAKDe56YIf4Sa0t4fsm75fkLchAGVmrSJkc7l44y20nP4
NvKeBf9CPuCfyyw0bmXbGOxzRauSGCBPuAWyrSAKMqOdeZJXwTIOf9LMjjqqug5ZEXVh1LUPP2UW
/ByeltcZo28WtK6KmhZHFWJtGRAY98aMqvRx3PIKzp4OG70ct4b3bni5+Pfez/3LE/74Ik9UKDjH
Vn9HSYM9m/qwxR24wt4+fX/403BhK4WSU5Wyo8XhwAfE/L1AdlFDf3ViXBUWdsHdYjvicJ5e1yB4
OJuo4lxk+5w24RJ4OgHrlcdh+QO1OXgsT8cHux2ogh2diV1ypiO8CFj1qnEtV/53n5U3+ajn62nL
OfHPFla4Vg4XDwQO4xF1C8ASiWTnrbmcuWiZ+/4RhMWj67CwolkWh3NAKlwer7Zv0kTaN9nBYc9g
8e2dRYKhJ5/7WD3UgNaAPpI/Iy6JqOsZojwQkAk1zQVAkCNljbNAOkxY9DeU5B6LSGQ7+Igwo53R
uf0FAqt5uKzGHLRDHseY+AH++VfQccJRHT2bgJVSiemIcG968SQ7/xoLjkb/RXtkQOFcAmiKhk/t
hZlG8I3546BClTB3UMxzSlqB69aPGvnPHU3027u0lCzI4VULJiJgeIFcaVoS+4eyN+hD+3ht6pB7
JPszEAC+vhFpcK6Kuk7Twf0IAIQyD0cBSGJedWHupoF4zBD3AEs7kdw9fK5RNS/UV7aLtlvfS2+k
8U7Lamf+pOCdC3GsshZ+aWuFjuDq0aisrcGkhHauoslyKnUIRIz8NA8JhnCYNkokr+ebzM/L48jQ
VSiPI4Vp9xh1W+FQvPBiyGgPhaZTpkcDiG8KVe3Gjijh95fIxvz6R/yJnz1jn3fZDEGEdIOnxvnz
aXZzzy9ynLhJBIazOjlNWsB5/2SO9PHjHfjG1iawJFA2gD5Hw0OmysTn2dotR4Mt8atokq7eD9A+
atxArNh62DOFGHvmlmon7NVu9XQFwjZmGD6t5h8z7bcFdUbyXN7gu1xtF4l4DXeJnJu8XWeq39gC
e975hcxvGjAE0eiAzqJeg5O/UXHPl5+tQ828i9kIhxabm7PHhyuLxsV9mCaCQgH7e92iz1WkBDni
SMM3znopfbAHshD5+blaoQ3rJoaNzbzZqTsvx2HILr208PE5NvHaYVBtpqDdC97GU0ZyG2z//UX+
6aCz9SpwqjLuFKMqH8J9Z1NW+vYn8blkxH8kOsB+KQLHB4PryIm42mdQnBGh9ZFvMwsgpbNsvmgY
iENeMQlBmbfCXne0mek0MeoI2RP2i76J17FJ4ZenOhxIAh1o/WguL8w+YUtBxXjH4tWz6LiQ0ssN
m8m4zmvxiVmibkQ+czwdMpZb07peXRuQgJMdo6CXdumXR3Q/Xwt2nMORJHKOya5ddHPzYA11FAZq
z2xdBur7MM/YZZF2aI21V3JJpOXkLR+0l+0ZdNaQyXeHpziHx1AYRjdR/DZxM5lfxEnEqjKSqtJj
5PgN7yt8bTS4s+N2o4RV/f5VqKdTF2hdBVDwN+XypuXzbPtTbDASqC8PrrCY1KozxoCiFFiotKz2
nRixmEOqZwfqhol5ajEt9yd4Z4kOqEUVloO3lzqwpC8DGEmoNinGew4ycId42nilE6VSlcceTXWh
q2YCJStmJ47p4DmqgUQGQt9D0/hoc1zRS0OZlUbExwf1Qi3ny5UKqZMY+cguJlRELV8We0L/OYi6
ykXsea+ussKWEdLBAjknSCks4BRdycr12kxogES+QJbTJti7384VZkW8/PWtEFjP/oBi7Vk+JzS4
Ma10WPFTwh/seCX8vqus3rxb6CvMb/2ryjJXd+JZt7aZaxXVzih0uqef5BQW5xR75y7aMbgzgP4B
sGdNiTg5c9wU069qhiwuc5m4wi4PkYRmuQZge8PX36kdqZzI4yAibtsm1YDwbNE9LrNs+7Xbwk2W
VWNvn8tOXBxk6csbIjBX2W6ncuBlUega5qkfwJ+r+J4bwTf9T/UdV8bWs+E9J4SYqS4NrPo7c7pd
VJZSn3FRVhlqaqR1ExdK3j/515pK8BWL3b3Ay5jm1fy84nCGTmGv+xCcNA78COOjxKls4eQCuXQj
C0lHTngYbmzuV/QBCMRbTWmEisawjmYI7rOihUQNunbSAHISaTrvfkidgqGu8QZSnfiecA66U0S7
P9RqWymWojpMKtBxQ3rgH0JewIsHcQHcpcsk9Jem/HTKU9W5qKYJl5oxYESZURm2ZumPNaXSF1Lw
Rs2k8zZQg2iZtCqdr97A821GKT+pym10GOE5cUeC3rhGkAlPriFjHkf1p6+oyzH9W1GTSOuhqW9u
1D3b6vgX8E9rm9BwFSkGUnWQL0NjJ6zK/f4+2WEyMksLj7KdJ/18xUT73cjszwfZDyyBXot+gIGg
Awm+StajW/rVSAtP94DLeG41h7K/SjcjH1ELRGfPyQqh09v61ReK45/YTlPGLsQ3ZEaC8nVgP/r8
QNT3aKb+9Ky6Cq5Spz9mmg0t+jP9QmbUsG3XxBIoQVMwy6oa6muXfvG4gkOfYCzhgZRWgvA9ePvO
lC/kGYRZZq1Vg50Oqdw1meNB9jOsvSCQxGAx7s0Tg0jM/13iC9Ap50CIym1a9PB5KRlPIdyVy5na
X/Eh99nx4iPgdNgNzuXlEEX50LGKOCpdoA5Ef5vVnNuNMoJpovMg39VwJPzkgJ0k8q++Awf16AR9
bnPJDVfN2vTGwUiPxA4K+vMI8gHwdlyWps/HCFn8sebov03YNqbQfOfrxi6DIPRVk+4Ax0ha+5Ax
gu7zvY/ZkbB7CgIj+MeqS6OHUYgme/1Sq0RmxVIHnYmeAqn1hovBC9NkjeZa0/EVCxfH0W16shbu
Kr4arMDOSxzwUBTsNF6IBak4jS4OwCA1JknG+KTXQWrKCv8dTNM1+d7qJH9/fUSTX4aaPRh8s/LQ
n5gL9KYLmC6DW1QxXSykFLiHWgfjM9AoIGWUxAd2TA/Yw4cmF3pE/ROQh8Jg9KyIu+mFMbTg6oW1
qLzqrqmfUoIngHJlSKadDQE/c0vVrH0dbUitCyW5+RiZ/X1OEBuelCCEbCnte9fK+t+4JtAhqs6t
/97o/F0V4yhT49NW9Mq86SQmP6ttEOsIqUx1CDbnlNlTgfxNZ0n60XTYWlFHdyU451/0HSrOAanV
GVGMKxSuiWyGJST+kUGfOcwGSHpDu4BwFp39gL+vKMeZYFEm4jOsbOiI0z99vxCmL/ZHUVuC3yAH
V8wJrsbwj5y+HZDg1lhDLDKy1wwnCLZ9mSko8n+HAi7I8Wok8XLiZuyhmtc4LllG/C88rNXOqyr/
+RIm5Vi8TaRi16PMm9N5qLDGoGb7ykSBFmnXxEcdhC8Fc91xdqQcXRQwjOBJFBihdTOVcGytwIac
2Wbem1uVNTUeoWnOhTCZBUPymJ51UiwfLjCDs+ElT7IDRymwodfGoqOvX3CPEzLccNFPw2/08wTO
kJtCMxNFTklADY0MrZQ3EqHBnmo/weynXepd1Qz5Obhm4bRd53Nm6Tu6Ok4660Ol7d2cenZwg7Ps
GHu7tOeAJOJzzLCMoFF16sltIgVxgZ+X7AfXyNRiCfaVzWVjNY3zCJnqCCvZbp87+IK46TGcDGB4
uBXhtHfE9orhLcaL+rnN+dAi+mHQx24qSU7TEYhfCW+3Hoxt4AKgnh2eRCZe/sCgoi4oPghCsMQR
Lh7PzafIe6XNCmR7+5MvAOLaJPFfkNAwWQsUALexQgtTja6B5zgV+4SkQrmuHvEyfpFlRV0JYu1o
QZ7f/0vu0q7HJICuJQKTBJ1+VI++H8IN7TjJgRvmen44FCNLPuzK6Q1tUOOrLiB5UR41yam15N5J
cl92w/rKClU6tTnjRNPrMYCNL06SFhptIXKMXPPV8ze1Tcpz1EjtshzvTtwyZAMY7boLiK42SJoi
lKb5V+B5VYc/xycuzoOn2nxr70CsliOdGcBIfGguy4PZL4+CLiVwm3fmSTKpy6yIpAsPZn+LHha0
XON6HqU/ZIjScpuLVVJ1563IOn3i/NWFcQAAjlOMZj/m4EISayzY/taQWyOQvhsXJC2G8LraLmR6
YUdSYbKLnjKx46fNX1Q2hw9VG1PU5eI6+c/ee/cJwwh15T77QQd41u3pc1geEFS+jK4vY31KKrPR
YQAPH65AKOC7ITCmG5ftt6H3QADkwiOrtoDxtpahib85uqrALpoF0f5gH6EkcDpozJ2TH35eJI0l
+9oDOqyvR9q1v9guMNDUOitsTcRgH2OZicmt17G8jDanjeIpaMsaDx24la+fRiSajIcLUal/ofs1
Xi+RnwYwrjbojU+fd9U4r1XWSCsoIzlYisAExeV8fnjXKn+PlyICYM3Oo76avpRqKvjnABur2uLm
wEbZbmGObk9c2aP5C6wfVC5HeM8waRvRhTM71Pn4b3gP8pj2VAgdjyvJbq+BM34iisPK4Jz69XQX
LdQ/dPrX1ExHS9Uqhy7QJ/b2J+P4s2umwepKHT9Xw5C+A2dGjbKSyyqDCY0CKMGS2UZglqJQhQzO
2OtASfONpAaM32vzgWh5NXd1o3LklhxeS6TTXfLM8x7vJOSvc/xULmvwIyO7Tb7kqtlu7qIa0H9i
sKGDyu7Xndw6mghPNhklyP2gOZ6bKnM0xBQiy6ZDUpbGKDh8MjhVQXVCz7kp4cvHrU6KgQ2tAfcf
YAP++zxgIpDeF8nOKdhjUR3dgJqnpdL7MG+cdy0AHMJvMrgQgQH1/tF/wxNi6zd1kvV3KWwuVRzV
7cwAF0MD/ITFe/NQ13hpW8PPd7JHTwkOzkzA1PmuUpDCvjsO/P5Gzc/o7lSu/fi60z3DZr1QlrgO
R6W0er4uyVD3yZqxsIZr99RC2trbMyqVc4LDovDouPflTw2RAgevFouuB2gYapRfQr50VdlrnyCC
SJEstIXLeVUJcPloKSo5b3Ziqxy7f4mKsm9gXoOXdgUlEFLA3H0EKhw/TEGSL25KDLOvQFbwOTDs
OsJvPsK7NTvZPI1DIrFTK0LFTodeTfduD16V/WRgW/utSBumZGskCUtujgvjnudJL//nkwT1BuDX
fvl0nZhKygz6llgA1QlM1uRXCfsnj0g/FQOWHjz59VamRYnTE7z+F4ddmjOTna5fFodNW0Cg5G8q
rZwlb8C28d9QLQnjeKuKOENfv8Q0HOuK/zUVVc7f+KyFi87Jg8nBd7Ux42kshiBy4rpr/4HqZfr3
CmLxBZOKnJYKqRVW0EqrUBdZd5QVDBanJkhbZqIFBmBxzV3aYfsNYTFSKfPqsviiL7LiLNiUUBVA
1SCN5BhxzHFj1FQg1QFr5oANd/R/s+6ivWwMegGGOUpnPHejbj2QW1E6sop8G7oMo6ao/138o4cK
qXsudZKIl/tmKTYqfmxRtqAXYQy5oAcdr5pFzScb0+s8XaT7iXtTWeLmsTVNyJzW/yI+iZKZSRvy
ldEZLWuh9CiflNW3bRYeI1jFAlTbg68op5SLvEziwdCCrRvtA1P3WMj+HYN4P2LgHy/S38q9Y/cS
8gw82IJPllUZF8x/7AOHSre0tVC4cWUwpl+4hPV4Y9P/jdXIAlhLAtjrlYfgA9edkhxvECpY3Pes
1RZh80upMAtWJeHQsOyfRVlQFFCBu4dlueLEeAxBNDhmMYxUXt63M9L+U8hWSLys5K8lu5gpvYu8
1WPSho0FQWhdgPHp1SHKNTj8lyf2Naz7cgpbktYhIJ/vCBEW3hvfP+eU3Pae3GmJ8Mc8FPOiOrJt
8QW1uLWU1xf0+OieuIMqP8arCetIkgAWEl1448PLmVR/86IPOvyHXwOOaPTQwIemqNEtL2bYuKy+
W2fg834wdDDLHgA7VHgWUDPd7qlKPO7ZVxgqZFChmpPx0uXsAFOcd6jxrkIJQemee5ByWyU9tQsx
dvuNE/nOlWXTwEt73V3ecAbWVBDfstTesSOu4VR79AXT0W7TA1EKUXozIm2A0EI1+Yg96cSP0isD
z/Kodr6OScfzyg4Wve1YJr/8taVKzAeSXek+2MUhOLtDHzj3P7Vu2sPU7AoMG7by+uwk8ZZi+p/u
DdPwz9gpY6LBsyXgS3tuNzZ/rbfXeqzTHMTJrRstQm9b8nqvB838bPXU87qJjphLnSGDOxgqT2vS
suXnTnuy8BGG9h/xo9FIBLAHwZ3dDX0efOG08nVRWPgg883HJo9Lh74LQlqmR/98BeDhi/wsShx6
m/g/eHqQuUiWKhOurnDXpFQil6Zajn1GTxGNmDjtlZWy0DZINq0eCGROQlF3iubuupn949FF98iS
cACrR/Ls0kSEIjSxfA/SpB0bNG5m0Ghfy8GiNJKE+fePyBpEE1XNGaQ0JeghP+NvAlpXK/0un72/
xWaOSTKgTkH7e+HzntMh9cn14pHxSISjNd8X5jCTKSlwzCI1/P7GxSFcwqE118l7G/Mj4mIWNafG
F5iejQWZAmRBTqeIVOHtgFESZB0A5w8lWa1qaBoUsQ6iwo+vwl+Ql/EV+MKSfa6Ih0va7ht70wwI
Fx1qhyYS5FJtRwtCdcwh4rCxXV2N3BSJR0jmu59TyTGNRGUaa+SRVtUH1r7AfSJW4yZDTwjQt21a
DVCOoSbmXxYyENSZ26QQNX+WEha35fZWMu0wWM9ctZhTson+bAuWMUZI1NW6kP7ieJg2CBvPCi5c
XgDheGnDYxQf6wWum4mrdFCJe4EpeCq4eOYUwOWzihPd4ANRtsYdcZHfHq3F/jI7Bxo9ot3Dnebi
UCxyFpIgyYEEUj5xvTFm8mgmpSUNYCxBknBPUPKoIb0iELbOB+DTXHqRtgBUdkGFweMR0cpQXFvv
h5sRFmyIvQ9WrntJ4nYCgkAFsFKh1xYnLKGOZUHEdovM676sFTNMmy7nBsZBcYOeUm2sDEEI+RUc
NxhW1XZWig96ZvAT5BedL7cZeYokAkq5HsFZPpwxj1HaAzzgmgHERvqWS0BM7IeYydv7vZh+NUBd
R9zQ9GcxcsSHALrYR4MoXhiN+AEoZJGoAD2m33q0sxdDkQ6JohOq4GXqlrauudogpRoCEDtLtaIr
7+/60OOHEXWtGQmSpMAPD5fbEV55HZtkx+hx1t++Yt6aoqo6ubQrLo7IqyFZD/DElNX4Y/qsRgm5
/3R53lDswKW8z25yYSIAIPlHZ432Z95EQSX0j5MDSIc3GUa4Z29DfOdeyPKuNvMiY0EkQpcNd6mW
OpEy7qhvoInoZm/+AikH37PUhJo/eBbABtcvknkv7Bpt7AeBsmb4yBfmu9hDqDCARCjCcCVaEQBw
OQepq31kuqZkPF4+amHPkZcdp+1mv0ckO4EvRN9Kr91uCGI9aaw/GjrF9sNpRjmHzpmIvdfWUG2H
wGwe1fChHBzukPpiW+g9DWdcrRrbexFX/iaGsG5gTsUg06P77/Uvm3CKLac4IIhQlAzY5XgtKSvk
2jr/+TdqiFN4TbDw+WfRQhtQwm12qwyeMCUwNPKSo2LXyZx2kE1C2VepSHCH3XlYHUjvyTQFE5iM
FC8dM7qJ8Gdz/GV7Y/fUVNPg9oeUfyuxyw+lWzZyeEYNAELfCDOWkIwW+1rrTOhhcCZRN30vfkIz
erZnwWspziQH6/deP3Mg3mLkpxnMPRaDiICc1n+LRAwBR5Fmq9z+8sQSc3m0+7ekXndCc8Zse/ng
/we/F5Efb75LKshwlMlg0q7U4Sx8kw4tMHfn2S4gIZzreSspXlInM424X508p8iPpbGSQnLzkRnO
I645ECB6V5eC6ikenpYEpmD5gdcyC7OIzVpH+AjbWrJa5Xs0NPfMo3RppeLhCAmwugnMOFVR2bRv
UW/MWZDwRDLCTIwxTFgFdOGV4oJgT69ctJs6VZGKSX0w9VZhUEid/loPfCrBILIdb/zDDFwEBLnZ
Xz2sEZrf1HMA1rscrp47GVrHHu1ixPLtU5VhoQoVjACCC4e/7pFjSrnrqhdpQYgtTTfr+h8BPt9T
p9KMXDBX4PlXPL5izYGVHQrfMtbUQodfUW4E3oY3uUW6NBg2SC/qQFv4JcDeY3swo9jiKcZdUB7f
+8h9hjSU1suMXCTxDTrIjbOkm/lTiEXd75lh6ybhByhKVSSME4QrHe/n38Eyfka8Y6IU1mnlSocV
9Cu5nG77UR6RPNFW+jG7wSYhQS/l8yaocy4bOYyXNZ+wnYbWWuvjFqgpmJkY6GbHtwOhM1q/jtjz
1w1HisVGNllhkSCf5QKWhSK3c4DWygV1hsEEtL1IijTIQdGWYksStknP6fxEGnTMIHs9pYMfbDCo
HiL8xVX+3Gw7PzfbP9Zh+R8GYxMXZoJtt1RChjhXHcjB2uFLHb1jhAkLBLtdDaVm0+bRKVanqF+O
r0ByHmPqJDn4Gaw99YKIhbxbOqnUclK7MpKvn7VO7Bg0ELT73FD9dzY+CBJQqgdBzEGf+vJxRK2H
cyMPk3rR7IrN1b9kQsXtxnMsUKmB3bB3Q+DD5+pyXDv3VDSFhI06gzGh2KPYdMV2pT6xtOnPWieR
jgpVFWqTZPB2f70jK2d9PVznon/hUK1CWB+aB22Xh0LhSejRqOFiL+kQ27/4a+B6UoL6qg0UF6Sa
u/4R8iSOY7fpdqHPmgbPLFTkNsm/5leAJW6GxmrY8yrDol0M/ZotMGdVgOkhZFt791qMPHb+Ddhk
yYWJW2CIG3aCQBWNXcFpvbSAwLNKtht1Vb4WEV+W699h27z4quqsZMfWM6lreR/JYU6It9GXRBhu
UQYm0gqkH164pW0d8CkAmK22094KxFzfmkSpEeYcyXH+PXXCWnLdR6bysul/5Wz/RxqXbMYeYmty
Ykgr2yGVrYluOiRhtDPo9zdwx4dXVCwQRuoVa8kvIW1nwfUK2CEtV2Ya8eDn2Kf/Szpy//q0ZgaU
0scZGkKT7woU96vbJgm8XSMIXEU+jHTtVOsd1dAmwRo3pnxmVSU21FQZSj31kbsY2gA+hSFGFqJX
M6kTj+YdI2P/kih9XofsBLJN1CtzAc5CuObFGkl7UOaFFhPcwxf0GyTx4yd99lIXfFFrWEMbGAS7
D6tAAtpbtLkiJHGmFpjEw1q2mmIHkDsv3W6iju87wWET214f8ZA2pEoEUPiw0bePVVid8oZpoy+U
12wdb5OhXhqu6uaC1BZQGyjZNsdzcuh7c9Nnw6B6tCB8AJmX8Sc60Y7oA2U2DCCU6HeYk++0EcS2
NQ3Rr8rob179OuL7b2bPFGA2caVWikYd7tkMvgNgNa1Fi4Q+54nXsFQkHDa/mIO31tnVE92Oj0Zr
mfESKJtkZuAxU1UOOdvFmn5/wpU1nV1S2w9yygF6ehsCAow0AuwVahpWWKnntZuTzmVVYNzZ2KU4
LHc5f8NdpmpWFS1+LpIgK+QJVDrczvcRNquAywaJoNEfn9YcC07ETnNlsSMujda72n3U+3EEWkU7
yqRgv7iP/2dEJVTk9L2pYm4DGLUABaTIIeqVL9EXz+bBF8b4GzHKqTdXjdqS8v83Go43rO8LfJtO
ZncyOYapjsihPGqzIHfMEgHhP3LT1JSldzlY/chPQhkZomvACNwq19LMRWTCUZmSdpgK9B42ySzz
nY7LcLLNhhCguKcOE5ZW3I7RKcOjCVciEYb+MAgRylZwah0qbcT8oV94LA/D6gjYGkGXnjQfipX4
qauiYVlnbTeflMNzfvn9beW/6jv/63O4/0GE9B0kudEudXDFjDqAbHgZKG/I/GAh3KuSvxm9uSB2
vuh/IExarVM3ejXLBaKa/OEq/DEk9p68a6bWVMng9C6B7fgHLsvOAFehmneKOcKUkVKjHVro4HLF
MG1DR2eoEMRXO7GIsIxdmcVPZndW+ch+VzGrhSUqb4ZvrZSx1hP4DOft0kw2BVeBdNX1UYxS8x0X
5bI6kwFqn2w/7rDPKuv0OkXgc4vGjUBFuiTJtYD1PlAZGDAszUgJJ9HYrqHNLWws+76oyGUAkWh1
hNhEe1458wm5KTsjHBWJ0xSZeJ2AoyXYfIo4TM2y0NXjElS99oieBu3InQg0PhnCNzZWnXVJNfTZ
MSevEOe4lwQK3krwPENu9QsEtdMK0Dnx/U56P1mpbqX4Gv06kTxfyWNo6AQvodlIeQr01qaNb+NY
LHxFFfr++vNKFrwQ9QpPERfVPeZF/qGGO93GiMq9OaCBIsgAttDjlqTa+XXdiNqxpNjawR1N2Cf+
33IiKe8xc30CCAiNCkYTpeeT1dIHqMuNANo5FymXj5fj8uEjNvmVSerJR9d/WgbZPwq7qVjoTO1Y
a42DHx4Nn+j6c4E409zEj5ctMG4mjkAtL8SMDpb18PBF4i4scyW2c2mAlAXONq3vOKrJPDk5r4P8
CFiKLyQwbZxe45ioCgGWv7ZR4XjXrAzGIBhbtsnUa++DLXUQqg1CA+Iimb3CpUp0CoVRLyFxFaN8
KRPcYf/Kbiy4jv0eeN1SlPTN60vEG/1rjxA/gx6B4nXuu2woo+HqPUOAWS5XnCM+gT7K3C6zaTpD
AOaG6hcL7ktWhEPo6r34JDf3fxh4tZinJ8UwwhVhJZJdaYvQjBmApjQuACS7+d4xoRPE7sYee6we
GQrtbevqXhsTH5BCVLzDNv+QIs01GOG3EHopwLuYbyNcN1UMJ62G1Yx25U+jM2hi1B1NGSofy44l
aQIVL3LCxaVCMQzPAm7COe9S8xCdNgK9rWasQ1X/8OIoCZwI/vCEv0L/YRFlLfUTiw1H3BGvmM/y
HGgwo54ox21i8+qO/FDwTlAFCqnnbuyPaM10F1RLBu8oE8CRghLb/cBBgJ6KWx8PSk8galr9H72B
A85pM14rfMrTL2e4BTEmLfTXOSOtgDAdU0bVH68WbYuAFxgVZHrwvzZecQU7zVL/IN0Ice+22OlP
SvJDgF/WADShJsAKPZ8E303mLCfd8he+ChZvtMVRQ+hdOagchHkv7488yoc1rpstQ2bHc264Lxfm
JCN8yUFhYunIAieq7lPlilAfrDjUE3ithgDThRbEaL5ZsqWaJrm/xIqVFdXJSIEcVy/lUcF6uCTS
Zm4O8cXD8JN3dEkkqCOOfRW7xNFhs9zTEetxoymvqlgkqgev0x/QU9TqjyeVY9NRQcEuMs740XvE
7U4cOAbhtEGIXKmENKwZ3PuJu6axvIs76IKFGlK6B/KRm6FRZJGgmNhEV1faBAVgTVzfHumWjNh9
QrF+uGvPC7u+UTPs7lfVxPLohD2bGXSg18XuKvxSUyZPlB2PWqQVuBINV5AdsgzFk7qSo89VGby3
8IJwYczW1xZDzAaNg4DBMQxDQ9kTQ+HNgpy13zps58YsQWfMni/m/XnEy84OKtIjB5pL7q5ReuxY
0XUaCBusu0O+ZoPwPJiVMkE2IGPrvDa98sq59tzWV5i1f0kFsKMAlIBCUWvZiNsvcNCdSzkFIogw
HxQPrbhjrbEygjvoO13BugcinSI4ZHtam9RIuIkVk2J0tHIawdGDccNKjeu2pOBVrCGkohaXqpJq
aBW7Wo07vnli9BgQQ2W1+UIAa9qcPefBDjbzyx0wpDFS1N8iG7tFi/ue6y4YNRec08kZxkziPrgA
p6U+mgPN3PVhm7fqVz/yWNz8gK5kNUQkXw7ZbEy0NDZOuSLw9/GEpXuvlKWo3EaGB71CbJ7mJ9Tw
xr5bxcX1mtzyDY2O6eSg/V1Dh6rBGIW6MdxpxhosvwyLKjFrXYh2ZrD2lYp4v9XXbaimKCRwlSDP
O74uSLIpgDqQZC+k/ZP1DIIzHyvYqu763kN8PxXHWw+b0Z3GJl4iOfwgtrGD4hX2PWd3OiXCxqv+
iWogBqJAL35k0+xOQrf07FMR2KgG5d8CIuGfd++xhvm/9PFFBqZOgWU6RcydpLXB/sGNJvfzKNea
n2Tv0k8+gFZXzXHJNTe90+/SuPiHgFBbBBNa2pz3VlUkzj7ElDWELfNdTMHgtuIfXrT6uMrtOOrK
dFAbiswW9aMd17lTn1U6y92UqVFzxQFjXUvFZGIu/ymzVjlMKUruCBo9IdxQMDU8aIp4LghXqKV/
Vv6LjirryRrrSTkotYcqgKIlU5+dnLRhddoVY28KzH7Pq2+RkijV9Pixq1sBpcOg+1Vq6urSdr23
hgRgpa3jjBSH7Mwb1fTepEWcLFNW1hQ78WKcZKEK8eN5VT7o0B3XmDW4NiBMg/03G/89Tgnls+bL
KD6QvGpefhN+OmWZE1hM2gmO87SRZ7W02n5iHZrzXX5ZkikSls0RBbcihkWBXv2HevVwehFUebfq
ZYAADYs9qBUTlSQI3VjQI8eXotjw991c7ZQNqrbkKz871yyMcXbYJUl8t2DM6trVYoR+Eit/ScqV
0JwX4XH/ZmuHuWfbFYgAPCo0z1wREnsgsKBxQuRLUdsal13sXdRBDMoNE2Q9BT0XrYc994QPNh9K
jDWMR83g6zYLpME5jZTx9z5EZFlnE20BfjK3vAyUO8o/38Rf3GMJTYr3PNIU9KUNZyCvzcditVQU
SOm4u5WwKEhPVa7Krpa+L7kcTyFCp0lddyvtwKkumYyGFWyIsLW7esBaRD0Ww5gv/oXyBzi2Dy6H
gMyc9+o/8fUkWHi4IFXVNcUwzhlOPQ1uHQG16uvCWR4ELLgnt+UIpwFpD0QY6wqfUEmNn0X0VCyq
BSzh3CUcZ+VLHd3X99G8SU6nvee1fgNctvC/UKKo/T5MtgRTZ2lILv1kXBnT9OpH6d+GsQjhQ8QC
Y3xXg5n7/nk7pAeYaLN2LL2iEJqMGTAf20uMRU0QbtSbX3AcT5K8FS3M5WAL5ok/3MR+ojtR6YgE
UCjMnnoOJKnB5wtYH2zMYV1eDQdmAaMK/HySEuXWdWkM+SaoPWTdsPQWrUhyLVW/CLm6YkTWeb+N
YbckHyRtREeu3aTxvyZb3Y2gP+IB+i2ZF2uSGXPT4lZ3pR/mMebeiDjaq5LQT41kaDoyBAec75Yr
snLea1kSLqkasKkQ23FsbB6UsOhnQtZ7kCVX8lzItbT/8rxLjVJvlvkkK9wODGmQJITY0NQL9USu
cLTjpWcY8BWD71EJF15haH3kHHkxYEnWzemGYGSvyAwLgrtPlV5Gk5rh5RzSxTKyGjxTk4YCnrZl
sZwkA/i2By8h7rZ/LCzdFHjiYyDUHORDBvFBECo3UjJ4hIcPw640/ilV4R4tUTmFq8xTwTpEygX7
vwRyyFqHk/w0tjPTxqFwMxz0DMTGGk4j6s6ceDPx2Nf35nAxtMBYf25ifvVrkLUuLoREVqQpAE9F
fNENscFypsOJ5GBI3Y2uE+7OcO9eY55TF31wMconHxE1LX8xmEVoyTeo/hJbdOZSxqldukk86OME
DhXPP9Bc6OorVCiBLtR/PaH0UIfzHwSdKE+SsIT0/TTi7W89xPeQALiSi5Ximceb6jX+w5IALIEO
H6maT/GJi7pJ27s1UGnmNp+2D6aW1oDsdhpVy5uAU4nxKJuNP/3QH+GZuwiXbTZrv0TwRGwDrXfM
0YEn4PBIP7lmdCAQk9mMsArW6XFtpgbGWT+SRVVWojQsMU7Rkf10b6iWw9fI5XWgFl5mXReeTHjW
gQ8KUelrHqyId6HQsqcrJGrX2foVweB6VbucV6GkkuMFnOJUAWMSQePik8avECn8Tsm9yTg4nddL
eonsJJbjX+foAWzFEjSbY2TTVBYY01dMfHZRVE/uuWSZF/MZ65z5bK1BA6du6DMsqltqkWxK/mmw
yNSa5yVCfpIqou5ZPTM6lpU+eOR+nmV4E8B7z+H0W1HzV7nbiRJqB4ntj9lDc8YaxNO0IMIlHTir
P2H1A74BjL8XRWsaGBd6YjGZUsZklpr71eYGfDplDTWxE0CKzyvwQhPZ065Ka4vlrw2izWOF4dRc
9z9LLDHGdHY7b9YqaVK/+OGaDp+70N3sUu/bTiVOToSooBldJjReJ1R7ajZcj63qKWcBHkjck4Vc
0YrrGnu+Fr4v6fxte2snh0q2VzqSk4vTtadtJED9oS8vCi91LRxEAHhtQfWHTIXSSBIXHhb3eB1C
48VDBtzdYSS+hCLMcZ2Dy20Pd1rb8cBFG1sweKDk+xH4FNi4yMSC6fPv73tLBlG0tVggDcyBhqHl
/9OvY8tWj7rps188jTxLYqkK8CPTUXBhSdRpgWycIA5WjL0GbhbLCBfE7hLKCwDEZIv8NQ9N2/DZ
dqg7ttw0VRpCoPTjHexNVuyj9R+0qcLQoW+JYYSQcnYCPaSLp08H6roNbFXikpAZ7rIKRnNKryyI
VAEg0fhkk9eoXLzYIhSC0qf9O7yl22EAc4zIQkUMvH46vp2/D2IfIa0/DUErCMC1PUFBWaD5hxPt
CHnlMF6SLXwMKqDP6xGrt1kjySh3hWu4ggJpket+PHcwIfarLMwkKi+7UfZx3pUqmuwyiswJ3DCX
TsF/QKMqAQuQcivvjul/9g0us5/MuCj61tuIhTTGHqvsO0+8v3Y/1cfNQvCrg19g6xNpKCB9ZV0x
czmpcMn50+0Px/r1dUhLfXWkzrZwIlyvGp4RWECG3/XupS/TKtXFtVInIS6tsNlo6/0l9vy2woTl
ApDlnjCD21NZZh9w8m1iyEXgGMwSTbqx2J6QA2semav9Ogav8F77HfkzhaxoJhlHIXqaGhqC0lbW
WcSB/bCQXt5MIWiAwk49gaqOdNrINKp6/LyLSsMiYlIOfl/LvJm+I1WATnnlu0/1H3sQoYnQAUgE
5mgYfSe3++IED0ETpvphj4fZogwdQtw/GVUK6geRwhZe/CWk653S9ona0P9u6X9flGPw9qCqk77j
98gJtZm4bT0uWTje+tNdsq/J/SlUEWEivZzNlFHDK2zb+myst/g5YBRHsllp86f4x1M/oUE5cmnv
oqNXj4VGdz0DaNOcF8LQFXHynPKxcHPU+KZVQBTeK1E8RbEJD/ZIjjtn7Z/mn2oA+AMxBk8spc7V
JEsJssi45JGFILa21Zzq9WzqFLNjRAmYKVNr40QGFGlLJfvkNNTr9Ln3FWW2do5QVwxGrg4SpQUZ
mvvp6VhEusNAcO6iUX/mXQW6otPiFUFRe8Bt2f8dXBx+ggUxMj7wsPFTo+axlj1LVyr6tUMCvD2g
pWnNMtZ1SCoTptdGFvIGCx1dJ5C7wY0LBZgJyTZwkUzVUxhSZhyoqDs5v+dUZF7EE6drfsZDDReZ
tz4AwOeZavb/neNTIO0Xuor6rHqhsbjl0pDXkycUaCVlGF/+tzRoi0EIz6Aztu/PDoQ1jNj2ZBCY
l8j3CPm+djXKc2g8kRpIBJCMVuMu2KVw1CRpDpVyRjoS7OIq1T42CY1Piq8qAfFycODlvuTsYLI7
+l+WfXRBUjaVzUs8pympcuM8kogDRgT4PIu8ObGMyoM9c6rZ2heomztDi3P19AwDtqX3TEnvV3wf
oo7+1yXhzS+6pdCqhSC5CIGd0nyx5ApQEAWLc9rKy8egtDxQOTS/4cXJEAv5cq7nxd4BsnFTCYDJ
cHeOVkUGb2algy14j7X5gG6b1iGLLKxdqJs3xWWYCYOoEzKFpArN/IDbUP/HEEwSGvGZZJrl2+3W
sNphezOE3IS5/yfchPhwQO8t4hbkC7gt7qYeqhQUL+NL8FL5E+R18IOeBvU6DofE/ofCTgwjWgKR
PueP6VsRu5y3lVvmTtOi9hjgN028ZHjyeoG4yr88uSNo/GGQolOp7RVt2AjQZP5B/xHQVc23+Xas
JM6m9XTylqvPsUWOPpx6OHdEzH0Mnt2liBdr9VrrEaW+ZXJey9nX/vR+PN6EjKrnmX+X2sXz7UC+
BtRnQCSxruJrmK6IT8SEFFPNlAX25QcT/B93Mu1rBNSXzLF0Yy3dnNh0cXkjSwH3iIh326vGBBhr
B9njPRB3vm//KO30ZfuI78v1u6L/T+nOhHiRloDdNFF6NH+/jTD9CXnKyoFKX0joUUDsLS3C786s
1tkGlL2Vn9llvD571spI78FC+MUb9ZQt5C2cHsDTWC/K6oD7vpZITLeDj7U764xoWWN8e9D6mnsl
cJjVP2Clj2WcwCRPBLGhhM5nFVQwZizBonj5qplZbAWIo/a+4XEipR1ulgjtDcUsyWBurbQl//29
AkCDKfFPL0W9QcJJjGVxzScrq9ZMPNi0tNiXSoBy06QtHj/J0AwE3hqgeDMVaJMpnUKMQXH4Lluc
XoENLe5ei6dzdNGvssQZ19uhXDPTean2F5YNIkkfL5JGztZweQKwMcAbw/93v2vW66pKGKIWSvwK
uI4YNW/Sup0ABPBa/GmQJQN0tQFWGnoBqVtOgICnd6xSL1XB9izffyH2fuI4wYUOVi0uJpxkohFz
giPa6B6efDdMB8b34/4I+ELu208OVB9WfGr9n4lH4DSo3rf8I0U9uTiCE3d/IKEuCXyl8nm8tTHz
YfJgTewCi14l+LII856ufY6nJ9Vtu46lGTqouQK4bcuV/a04KzOQo+h3Ko+vSffIW0K8AL9RPtMK
52lMX2gzr6jG7srqrZ7diLueu14NPuAkxOphugpZVZyL6y/8IlBY8CC5MZwD3zEK3Vjl0I7lvnJ+
pUu1QzxtmjmwkPYuO2scphzqYuE6tMOqExukMs4M5Tux4cVIUmi58Va23q/iEwdc7rB/9tZ+3ozB
e9XiUE0xSHK1E7T2upHQg104Pd6Fq70D3O3B1lGdKGMWtD7wrZneMz5gLidlngBIlZqX+VmXUXeO
af80WTOUEsaDusIgtalXQPmtJTPrALy3ysx2w4CXOp/ut1EfqYoSbDTQ1xthHy9zC1NLimY+b97z
DDbmN+6u/wHGCPP9i3oowrp+Sw4hyz7Y+WwhSloYK8b0e7RHdp2ZvRuTK49Crs3OmBYfRE5q8Yxe
OLifwEPHnETuVRrIHlho1XWXJY+sSZtWpI3IOfqXZDTZhvGC1vbZ4ztuNcLCJnbXQFXVehf0kQy8
muOoVUSyEi3DIYAP9ecBFtwgE/t/XyzNN5gHvsxbDM+1pcKPduu92DUhgPzyLrpda5U3vOxki3/x
km762cDM5Pbl6tGb6RtWdZESj9dApuXLCMULeMnqNS4uQRgwDHcGTPYFxQnW69xY29kmHEvQf3sd
YuerF5dDZR08yt41PzavIWQu5vJ+v8BlHtDUoi8jW/cfXtOkkcSdULf+MaHOgL7oRgmcIuu+09w1
RvOR5GF2SiJbvBFqvuzUVGnJKQYp8IqmLFUxA8GmKG6YAGO9EkIVgYdULhvIMvF5qVrIDXzTd9fQ
06dfFt90j9+yhAGcJoBaF4QjG87qpwxRfqAB5lU+JobwV6Zkg791cfjfvlSZAv5qbhsEP0S713PM
4K6II2pGGIMwefHdLKfSfZtPfn6yGrIZfoo7TfLaEm6EiWAO3yAKfKvAz63ZZS/57oQeIjCFZCg9
zElDsamsdjBM1q06o3J04NkNjPsbjA0/1gMw/o4OUJwzi/NV81txNhDj5Ibu1ZO5XdhxMf5sBwa5
2Fifmib/a2xOa5AWn+mhBGbQu7O7XGNYf1Ui+YR8CiEvLPD8TpESCJUov/FswqLI17rNUzs+BbHx
roGlHH43poUHZvaNnoSwV4UXkb9gXotvg8+dLQ7zA803u1vs2QD63Sg0GdyCz7kvtbvv6132JLxY
L1QsE4FAltz2qkDLdQ82KU4+9dFfdsPcMq9lVpHRs8AbwWSVfO/jOdtd7q5eRYJDrCwLEt5QT9o2
JhH/w5KRV7GvFe14RVtTmuYVAEoow/y+nCKaBLXGKlQMrPyfhOXZY7d3UPhFaNm7yuYeiccETSX5
uW6etBKsmZVVSEfJ/Y+utMM2FsffRONcdImawddM2qIr1K88E1RtR+n+Q0IA+vcgj8odp1U7HuHv
5eR+hU5YA+I66z4widtRc/nboetoyHUnlG5/DHROAGeaHGIeznkVu4BIxBSSQ2DAeI/Zyl9IYjEs
GEB+zdJtGVgdi1zf3VNcxtB2/CjGm2i+sryWJVw4Geh2FhSYUGqLrIXlYNctcHvsU/sR+4wjk430
8lM2B1xVaWhUCqwTYZSas1wH8dvy9IjosabRqlZW2/6kwA9kZF99lqpTj59IlYXD9wKpj3aDlJoR
vOP66Cd6Nkmnn7PyZmS85wwkp+2ThGatn7uJ9bk4CDNYetpBLOFXwCqPHhMbuonzDbi58JPNRtys
M9+XqfDXRXBG9cmjMwZYj5MVgWOLXAr+tP3OvFWebdBy1d5zSjEIbkjNSlwVtHKsoKGFqvHKmOqo
On48upYgr1nuJt1uzpcESPeSws3b5eat+UnyXPGI37tZreNnYvKPQMBBG4WtYYa4T3fa+ij00DGT
nTDZBawytvOW/S8cL+Q6YrYFEGwZC9HSMy77/uCsBItr6sqtdMT6TXNZMlMKP3pJnhg0G3jON3Zi
MmjQH9ClWyZNSbpVEv/8mejC13c4ifK4FNFSL25nzdGytdza8CkjuYbQO0mjBLy/gdDteafL2u1u
fthLz4AaJidC3dcxork2zhKk47qr2YgvSpRDboxhMEoePmKCERxo9r1mv8hQGQ1E3dxJxWjXdMHJ
8VX15ZhnbQwc2Hwx8IgLoRp6Vis5HDF1RCmnmH/HcKDlySsArDHAAM88zGGLopbjEVDbuHo19P/6
eLsdZkrEZlSV8e1RNrwh8nU+ZymQtVJdgmKc7n6VCxO3bHpqTlEnJEd0eH2/ODVwUP/ys8ILOgTF
neQvmmOxwFdCS5rlXaZa5VTddSe5axnmnPS+hS+XRf9dO2rGL/o/f5TzxJHn1S+jNR6okAAEtLyy
ZGLULICB2R/y12M/SH4hxIXjoXMa1GKZFXIEBViHrkJZjiZOKAT8iKs+SnALhKzBsuETLyFaj8qd
9ur571V33OZdBfHnHzQygYMkVimh8M2ZWesVA5/ChbzNZPVcGzIyRia7+ATOhDvl9CrR+cHFFmAP
CcTf4pofb6irE/gAV+Wgxfd6dBnb2R20+6GItx80aNf7q7gAzuxKUN+idbHK+hC75JcxhmwjSIMr
pSB5yZCvdccCG4Wo8h/Cn6WMeMpxmktICrcdnENmrFYMT9Ve0LVmqTzDaQoVHIwDV+f8iHMY0wCy
JKR/Qf64qYL+W97azY5xMoZfipi+zT+Y6xL+pKs6WW7FNidHmtK5pEseebDL5XZjZUtNibmWeZUM
cm6uG5EVxM/7UCgFsw7tO4cfiJl4RsAJfYtWXdo3OXbKxBjNOhNH9byF0hBMPB1b8kQ1yDzlk3We
boYcrzCrc7ERXc4If9eVlEtGHamkxJUmrq63LTEbbgfgr4TvwMA+B5+t+lKthOsqEorRYaPyNHCd
AaxipCjXIidbjc9FPTX//sSvERspAGYiC046WuulyrEaK5S+hoxQEFGcDZKqkiJBMtZoM0xq5kYN
dYZ9z4whctJoSTMyg16AaIcc4I2JIt44uGqrncMBJsdzYaqkEmur7nRNE8s3urm3Q7gguHRlvZhM
hPmDHfB7lvCXo49f+t9XLmqRxh5aC7NzpOueygBzicFHImerwJwEb/j2l9kyqhktlPCVUX0ExKvq
wqmukE9O7wE0IuMsnKaGKbintrqIIJ0u8la813pR1cX3+1JwDAKJbrl3+WamqMNjoKvfKWQ60OUD
TpowqqTkTKD2vUUL/HmxEnqGLfe/Vugg2CC/ye1g31zXKgy4RavXwyXSIfS2YRGhvYIsfI4kPIOu
SiT5O7JRnc7TeLdxcXWdIbmzA8PuILysaRP2CB3B3bno8VdUXyfFv/CTCmEoDPaosB4CCs3yTKsl
4ovNjWid996gv+x+iTb0n1CB1Ou2M0wuJToCbG9jUDgm7jhacELDeHIZwtDYXJvHwahGaary9p5I
NdaQJ1msSoHes1HAQ5bS+Ty/g5LbSyyUNBdohr6/GZudggp0KsQv8hmU1L9DKg54MtmfndWlM0aw
GjdOYztOezqNnYrd6F2EJbMLZzvDtbPbuGakREdYQflIb8kLwmTC4t9ftJYBK5DZAZAykbP3jPgO
C4ds9l4E5LoMCWu8EJ7xXiV5JJ/SGFYB/qvBI+1kSNI7V1E5Sa9vn6BbY7jrNusKc91q9GRb+DVK
kxBLtjuwzCGx2cwmxjat04R6D7kxQe8Da73E1nQ4+R6p1luq8PIKrA+7i2MEmTDJoDyu1E3AX2Qd
yyfg/1cirgm7csGewJhWr/szhYC+A+qfY1REAhPFN6y72lPbTuj9q+4NWcQHfCSzTggVMhKp3AYa
8CkowHi5yAizvXwumMbSjd2HT+OiGA2EG/Bj0McboBgzxaUF9f23nm7iBhvyLeT6CVHriSnOuXoo
8eiqiJoD0rM19YlrGchek7ovQJzvFYKoE98/wEYrbsmQTgvYGmYMRnmX2UcN4ClyT4wW+Xq3qsTM
OdLifbnYL1rMaEgOumYAfKJs+aAZJYmmBxfA2gvUmCSUNeo/RUikYeNkX31dwxxrSTYeS+z8uey8
7XrbvijWIcTfNX3VHNLodfnyl8xfK+WmUJ3wOvGqbjAbY0cq7Auy4643qSawwhWoZh99Cq78mNHa
mC7KZj4l82/jx4z60iVOrY/HptPwvrEiQbXFYDN2dICeBchH08tZ0XTUalAbfyXMUasTWDx2IaJv
UYp+6gzUG4XUXRxnDyMDU/VnOXSKdkgwWf4j25J047acpI0jd2gAcdHPyqNV5QQxHw6X/Bj5DeKL
9iLVywkYd9gsX3DDM9T+pPRSOHi9Dl05HA0mzPS4lEpNFcmQh63tQPydXAe+rghCDFbD48BZMhrn
fQpqvk/150bjZWEwDI3toE+63QU+0tPBz+u+GV8tY49SqNuhdCxHG0ENdxcU3hff3QRoBTN+72hT
ar0yMfAnsozB2R4irzfle9Xt7JquVN5F7lBda2XPsXeGqrUXpHScwilef1BRAysX3Tz4NYDHMQxF
LdKU2ps8XNECq0Xib7FcbSxyAhOO5EL0jXHOWHh+OR+OPoKskHLrtOj1gzwi+NYPBzpJoNa9QOg7
gABRbYztG6xC1gu1oSCDHkyt+0kJ+MYbU7CKzRrF5vvqYqdzL7YimdksaMHBW+Nf/0vV7jVAbOKh
fozOg0+6HJJAU0wNBIjT7S26J4BL15o6Zsmpc+6m/S+tsDcZNlTrhohowmSHaT1GwFfOABwp1glg
JDyko4WdwkZNKWK6jeT0l6o0Fkpv7wZBK3sa5xVTYWFPiI6gMGj27tjnmHqfsWBl5EPhl7HNPMBs
esYANeYNF0pgN6SLKW4K6za1Ydjwm0j6bbixnlOW6yaX0CNinQEyiSLWZe6gP6koxb5W+czDHSm9
qc+kYkiIFR0ax7Sq4pnIqOqtHcpV0HlKCuh503vjmZp5H3I3B1LJeD/ApC1suX1IKR4yvmpbzsCl
Ny+BPCHpnWxhGW8ZqbRvG5ZwojdwqFkraYIcf+o4NTxrW/w9TFRFRfJD6zORisyox9uVgxFWUHzz
cnRVBkIpjh79kKEj1rJ236Vo6TEvIEuu71Yba/vcBtU8BwZ71EVZ4pHboqUasyty0qTx/7RSCA4I
N1CWNKWJOzUw7i0w0HULdDe1h43hEJkVGmumfhMBkk36pK6te/92EmqfKNnArm/jrUXcJQUpjMpc
TzXRY50mdpiJlY0fanspGc44xPOfBs7rtSfGl8d7WwXvPWzvhC9EujWykyuYVpvlsCSQSZZZ8EOl
8hkhvFrrEHP4X3xWG3rLKNNeN14ELX+I8DUy1iWnDa9qikyTcIY+/WRYkI8VWPfYMx2jS3ZVzXZu
rbnFJZtrKF+aXALjZcIUrLHDQvM6DuEVnvLa5BVJZ3T+C/2h9iqSYRcuXHxTQbq2CPTsv+j7xO6w
mn9v870wn5EqbCGtkxKGPKoPyj5TG9ZnmmqO1YObV4nM9cXlmNNS1prKXKdjZ5FaDb2Y+k+u6+Dx
EmEsD4C73kqkneoJGRaWSHBFOGgrioviFo6GaEPq+PS6qtewWkd/1VZf0AWRT4CKD4en/hP/6Iq5
s3e2/LrevJbcy8exLLxJCr/XLlWiGCigxX7DSAChkRZ9Yxa4c1CmON4JOHtrmKWUxZ7RS52lI2uy
PalBvn/qymDG+/mncHYymOLQthj/YDVmEpmQ5EGKoAeuP3QtUerNsEB4TtgpN3RrEfYitdiquvul
AYEdoqO80UCnn6q+Ioea5KvyLNijPn87mSjVBeq5ufVQNPaj8RFvbJzRddkic0BbnKVhGVexS59z
HCegRyw1kRHTRt7XlcexJPeZ/ZrMaj6xj5PKgxdQMK7QMPwLLD7xsGEeOg3t9u/xJYwc983R6Sgr
whRUZ6CI1ia5PGUsoF2vYIVlsK1BKJ/fxC0wqRkuZ1LmupgdFUBeeNuXvFjVoWESWz3Jyrw3AfLH
refo1KymtpJJmj+JthTPaK/fnqCI98IGw6PBWxTrfdYNrtP/9D5ADXrgM/H3rpg9aOAdFM7ndDMc
+hgNDqVxm8RTmdGxKCBQxjpkG9hDwMSuJbHPGR88mNVCNanH5DzkIY5hzUzYWU/+O6VmXb5huyrw
YeYm0VloD3B0ZiBhqaGsm5omxxvaYW/XOY7180NXChIxbelmVUWHBqk3CvyZdso6cq298qFYCyPP
i0RZp72P/nl170FfGRXkbg5a0Hfo1Kgqa2AzkttQMYqNBXx0z3pjkICJg5lptZuw9FmVqGIREmYM
Oio0+fLuto5DguGXHk3bKUR2rEO9QLwoHSQK39bdXcxb5zWGEup3OkJ3KO+AgeOvQ1H0IyOTp7w3
YR+yzzmYmQyWu48QVuyeVbPx/Vl3+FWCubhFXsy26oGeI6TSa355iPqGH0ddv4HwX4wtfQ3eSM0J
VWEa2MrLrEfKZ2MveLTbbvF7DOaH+qm3kst9fkbOdaVRpUb6Jg8KQYEkgNlId7E14iMQout/qpOy
3SPUTx2tnxAfecrBr5oGX/p841yJjYw/SW3aRvmql3CeyTBjIqxvY/JPLobfUa1ZsZ6Px4T7RZ7i
D3Y300DZUKuE5uIskmWULI7rAduWkgvz/nsLA/E8BxJKRPRUI0xXmz1SQSoUVnV0d2d0wFPid7Zj
Shw49HiH2toIG1vEWyArNDA2k80drMCd4+WNlHCQ7vqdBqxYPZL/ClOZlpcMSSYmq0d8jRpGKjMu
J1PtLgu+Zv23JkxDFVxAzBNbHe0UY3WQ+DLuAFv39BFb8DQrcNSN0p0ar3JGPYbTZaGgd1FFhPlP
y1yKv+9zUmoqAFbpbddctiLin+Up0NRpJEA5JBFll9bh0RU2bN2eX9UxDSl7CEsEKZpTlpe1hcIK
31CZjNsxkdTOnTOsKW182aRLNzoUUixG7h1OYLLK3qlj8aGnLSwTbIh4BQTcTz7ZkDFu+31zRzgu
JiQxf+WjzdpFZz5zNFbYPwVdQ6iK4fXly15C2Oug3cjSi57jzO4AmrR/fMYb7rYlirczAArVJZUC
8dxODRVZVFCfQslKkJqPxcYcHba38/2SA0Ooq+4AMUwhbCR+eFbdh/UWKEPO32IXzAbQ7zFnIXqu
+QM69hUQX2e9u9kf++EeQVveVkgTi90kWo2afREX/Jy/f7lBa+PILyrsiej5nACbOwtcRRKaz2xq
CeztA8ExSpwnYGms0UnxG8a1wevdbKYfyG3HmOvvYsP+5JfYAxBz3SPi0C6vk3EEzycbXOrx+icr
WJIHErKliTOz7P+Ldv175Ect5qNRlDVLg8dg2CoOXyMC0kQVmzCjAtKxPUPDYdsZJxri5lOsKWUA
pmfVZpBm37+CBGwVAypHrc1Jm+R5C1F08xkTDkO3Pt8MVNGW1kVvANZLr5jYu9ZCqF/9ghmv6ewL
jer7XJ4hg0ja3Pt/z2/jr4UnioFiRHomY+B18e6KRY3dXW5jYP79HqRxdeyfWVX3SJBXo6fOEo9F
8Qh96ugzEIVwztCRoHGq03zIxN8cSA23hiE/Nh59COLZQ/U6PLSR3ixDlPV7s3Nh8WQXuBmObUP3
3fPUZVqZYuHTf7W2RIl5NlYaQdlR2U1361GfLW2ShRv6cyTT12FmtQpzi9/671CDtq8nw15ruSjL
pT9k4bhkgKkhzt8r6x4uMi41QUPit36KkVNJQskDKGjIKgH+EIHIhgY0K9/debDJl7KnRh03qlN0
sbjArtuhZqfgCET2vXVdzkSMQGs6vxYkB7gI0YDJZMJ4xkypdUXQas2q5tP3zLqvPIZuGIeFbLzs
1/0YmIyVLH5vJ4Vr8FJjMrTb9opz++oc9sYm0FEVbQGybm6j0HCpfjgvyaXtN8j8p9/0dj/l7i1P
geQNTGZy0D0dgF+C46Jz1bxhS7sbfiimnlhlz7E43K1rkL2KN9dp0YppmnZqICfOPVsZ9EdC8i17
M4kE+xodonRhpObXdbRtf4r9mUr65BhoVM0OpIq1KJesoWHX+KPaIrs1TjbamMgnDQdgemmSfKDO
I8eQvDhRhilhOT9UkzYfh6FtMTNwg2icmfnSmkpVB57Xy6wLYmOZVcWIm9O1D/2bubJt+hbjwpeF
N5JRrWzd6k1i3u3LkxONMgMIc26NEFIxC2qy8J2LuUfhSDk7lwgR8jwM9AxBwgq2qRsdiaNtm6wz
k3yck5VoeJTrEqfjcjx/R2GBNOiHjUZ3GGauwTcIyjsSv+ti2ILANmoiY+k6IBqfjM27oEDf+7Nq
Os1wNRlVaYClCOPxowlWxodEMd7pNDWRf1gtvyiC30wIPTuA8rZ/fu+UrqF++X3olbpcTNrbPz80
9g8xO1bB8E8s6koTSi2G0T5NK5qNsJBncq9OIRFyjU7gdH8NcHBGHTstTMSsAa5bLOn1YmWvsaWX
uh4VIHcHmvHdUEe9md3EN/NZx4Ywv/EdpQZdJ6PkkekQizS5wAIWTKABNfN9eJGlMz6QaBRvGDDB
xRbkO/0uOsJAayI0lERvGj9qp7sQKfKbHnJlfRKWfh1cDhMR/1npoBtB7uRX/90rhUs7ePeuoSBF
pugZPrrfZnAQdvapYoTctA9QoJiOZFVp/JVf1nXtRsKv5irV0+IqmYR/8qqBMGsoYeoaWKsdchmd
digJtVnU/Okj1b7TipA3ujduRbpVRdBg624QyvpZBeIk45wjZ812r3dL2U3PoUpgxJ1Y0JH+UbB9
A1W7mnlaBuab9DluvdngmpAhz9VNdoeeguQhCmqp6Rx5uD5L+fq1kfGln4iQWEcrNMYYV5Lrtxqo
KqvhHRJ8i+4Ws40s0jgkvndOT0jQ2yfkRNy0nvHCe8HShiz8+XU8zNuspMSewYdS64jRZSTZIFK5
+tpzJlN/u8uPn2AtoWWFUcYE3c+IVPrUuFVpIPdZsi2iY+XBcjn+4JWqp+aC0OKu+asCPdmip52r
5jKsRpUmPudqqOorUl09LCBlUijo2vC0a2GIUo4YsxpXGWh1QPWLCrFmVtfa+Rz0yL4cSHHT5JC4
/QHq/XyHvB25sNF2B5Axrk+5jHvWkztOaW8Db+S5jqgNL0xghXv9vF/FWRTe1JmzC0gu20PyUSgK
AOFh5KqhuLB69wlteqRK9yvndAMltJ6Wk7g6cy0pMrpb1tGpbuFKiIufCG84uIy3lmM3lMwJXQmx
2ILlX8ueSctJUah/Le3Txzu2YOpgdrbnV8GK1VQUmY8TKZI7rq3d8OsB9C+xMtN6/4D7sAuniTTF
IeBZ2W9tpvbVaQlAWxn7XM7m/7JoG+EyETN7+Y2FliQraHw4DNCH2g/Es2KfV5yI2RZN7md8Zf2H
5a8lOAdj91fA33Zxaa45YHCAkuXe3P1pDHgQzxKY0Piik8HYgj+BJb95Gw3EI/98VSiJ7d2WEHYW
3+69L4t2hx2vtzSq0KEUI0syWts6jpNX0hQ/EYFZmk4EUkANXfL6HcRKOD1O6ofHAzjgy/9H81Bz
I5lyaspUaMQkd9TywL07QPZurKwasDmKbmmiE+8KrLZyHZKT1Gu8KxTilCG7D1x/fW8gyHOURR19
VslWNCLgCgnDgDUd2jxMx07EX/MjbLW+nuYbwVX1uHCudJBfXJWMdelwrVtziGfJpHwdncezd2xD
sABP714q7S15sxqW+rV8m6Rl0ltAevLCO+FR3dSXDLZAH7HUS3/maMZlWsivXGyXivIcnpwWsyKt
6K5z8e3kCPt5LOZWP8ZfAupXEBm2D2E/uyHDpvxzTPhq28en17tIOSVIJfvrbPSoOmhb1J2aaCFX
7INN/z3+R691hz/rh98LPQvXPDlFRKVU2eXdf6gm6mIkmgkmqHPbHw/SYcPWREcSPUh5dLPsBdLi
tfTQG91bMkWjhZ9Q/KeAaFMm74X7IOXNf1fikQF+RwTX2yTmG2zyncN+BGDkEVXBmZCRw2DbEXMH
rC2jv08A/v8jlwNGX8KRzxREYJXa4CLwtsN70a2ak2bNzWq3TiF8dAXnaWd/ldX16k6Ze0Nqist/
VozNRqx4mMWUvlKc4UJRtIEP99ISj1Z10TV8mbBZ60qc2IwysKYk1+kiGsnBdwPl86Sq0DxHj1Vd
Vm8abTL/RZ78pEBvwVN0JKjyKOx7ZnAlPaaTpuiux6TZwrAmSfnZhI6bwlW9qnwg63SoDmGyOiXl
OjKL1MDlo2uSZjUNKQJjHMOtTbMGqigC2h5e30r7r+p7qIkX3sc6YnueRWPM/ND78+sPeOQZmqCH
3P/1256pUkSc5PZbUgcNUnfWeBxAxYQVN+r6GPOYikMhOYvOs0bIjgnNdgU2rNJrCarEPntL3SUC
k1B3Ee7YT0GtcCT6mIXuCoRFL/ng3LxhuGM+HXRiV4oUeZhtXPGSqEC6SIRVe1KObEv9kO4xBg9E
VvOC+VJd7FkC0INUMuUcELFvUfBiYAabScKz8sxOcqCFAT2tKCBKZ0uFux/hEHyVUWlGQhnepsNg
zkzEwo0ERagfrfybKxiKwIUPUjzwUWGKswByqCaFElEWhiIXjav2EqSMBRLp3xBiax4zj7r0dBz3
TMDwWMICwdC+Om3Lk95y/yVBKC71hyT5/FawLFBTxnE1CgKhS2WgBmSqSemcz8h7wHWBN7oWj/B+
1TefuPsVSqPaIx6AZXc4W/611xvxGzpGR9Iq3do8hXhP6opYkE6u7yEubz8vjfHZ339ZDg0o9mIP
AMwuRb0QWdED/y+O9Rj5n/Th+OXUhI8GnkM5Ms7qI3GxfplvLE2d1mb+slDKB+q/hx+xecUF7sM8
qhJK7wtgHmZcY0rE1HtDv8CLnXaewjeXpioiv3V2MPkwAVcVi/7B+AVWI3nx9U9Oqh0TWtWR92p9
DKgtxO68unEjmvfHCQwytocyfdZEj6VG/7ZHwvvvMogO6F3WHAEQlupOIRpRILk6wkn2qG3A2d+l
MPvoMBlQ7ATuA74ofbvjGuC7a08D1yrJTdK6eJgpGSuBNQYqHGFhXIPWMl1VueKdd6TlCevY/7PG
ZZ/3xpk2J4QTPR5owT4+qToUHF5zjm3MQzL2k8YoCUiQs9URxLAR5LUVGpi6cf2FV+cciS53r5dx
1OQ3uqIUevZcIde8UbdKETpgnVXFmLYavi69vhWdjMtbVAJvGqQZLDBfQVn6TmqO1ZahhhPGpuF9
lFNw4Kmabsh3b0KGKHSKaj+tOsKBMTYuchkVmZn7kaViCXu4eDT2bUVrzS3y3BthDtWJE/9YlNyS
PyOPZonzAyNQr4pI+JbuO6ZBMZfHEqTJ8R+WqjTO9If+pWMCGi+jUrdyHyHkW2/c2X2x+Z2MoH+h
MWJ3oqNKZM7ZB8OCXSHFSnJ1WTTrDWBQbBR3pGnGA+ZFpdaa3pbaEeUedQgxjlWTItuLuMfMTtnb
g1jQpXoN+SX0XWq2SoTNju8pjEelNqSt1zX+3Q6IWyYXPrZMMABEAzJ1nO1ZVwiclX1MStwIZEGF
Yb0D0S2G55Lblhq4x6ur4/XgiEywl7H+bWH33aI8kD8k4kmSyM5vaqWZn7+02SBi8IQBZ0YNRSW5
SW+KjVJ3br8bO972H0GTNNimS7arMqdBH+5jw6JXq2pRJKVYuvHapfbw2MY7BRiUyeCxuLJhV0He
TP4ckd1peiX2op3GIAhxp7OvixK5E/A8wD6o44TLosA1fgVrUcncWgGnfhjFDymXAA26g4CfjXK7
fVg5LXD3+zevW0ye5KEdNliXRa3UGy3F6y4zHb+jmmF+vjZPwiR4P1nD5oPdBd5npc6BTwZB8JDG
UjH9sT6t9sQ/47Bz0QL3A+XEhlFhEQlLFE7rZIaFdz2izGr6208Zl2VBwDUCuGdfO3oQa7C/5JDT
/jaqXhmhGLxpy/qfu3rEdJMNvMbUyqz0S/AUmhlBoC/9gjGgS/fjwbnMGazZtd/0Ju6eT6OZGU6L
Mwu9k86olWyOzDhDsbowwx7AhQto0rQTPdZ5uTV3SqwYehqiJeJQjuZqIYueQ+k4HEjFT/+8YICX
vhYytdHqVioLZUkgQiYzXIzzKThpf4HWIHat7fcdldOhSpx2jIl7QL8Tevf99TK48bu0djQQ069R
6pjAvnMVZWktEenVfOAnqU/rFMXQs03p9wZxfh2IM5QbOo+sf27WpwHwfCozHA9Q0HG5cmJp/u3o
m8KpoIApYkbqYrdRJk2YBXI/djuDkEWK0SKLP+/gMfXZaj0m6El67hBTkxnSfMlKXs/KgBIZNM6t
trQUWaYHy//Wm/WneFf+cV3biwK++SM3tn07aqQWd6ln/zUbpveTEWlOGlV/0srCkcNtJ8sCc9FK
3tHxzqPjBvF+WrtdQL7bESnAABzZdeQ2i9KKlJY8sw02FhnRz3zGyPQRSRSDIJf7ZYJ0IBjopTKY
p7/NgiJAlV7IK5zCfqBoBokBQK1Z0g1oqOd31vBvNiL6pUdOSyiVmfKtxsiIfF1gnQ37laOqBfNO
PYJejzh3cuh5fNisV1MzeWNwQpHozk4qAcck9G35UgdBRK2bebtDzJul3vfUwwARvMM3sMI/MPjX
KdMEkyoeuyloqfKMwZmDxfMjL96QZuU4MUsOZCZJnfvNXK71qpfY9AoUhaLKaiN1RQoJftv6e3or
Mx17vA/aa5tXxoTl2d+bpdJ9ZMVOS8MoCcg5NYbNe/Velhyw5lnbkmQfbujbPnZXoMaFG31JH77C
I3/+zfwfENWp/lmXG8mKnhbxskOdFD49fNEfwjlAxFEVoiyOHHF784WkR8iXN3lJWVCIIsl0RXGV
p7XOqqaA/g6vy8hYB/AIcuEs2jVTaSwbtgHXkn6JGDf9/CBVaV+EtYuG6Yp/ZbGPkch1Shj0lWzv
Uxt4R9xbHVFXOKXfwOJAQJSvZGPj77/xcNTJq2044bo83E6Y0zXTY9OaD9NEDFSjdUSA5hdAbsys
UJI2Zf6mSbMReTMm+4j4twb4gf8yOGfSAleBz3z90cO27tyLWgaiaeFtNnD2yEzmurQHgsS4+e3X
a2CDx3vJAUW9MTVCt2M1Tw0hg7hel8elU4OWL2aSVvG4q9MuuVNlJ5tIKccZaJke4JDJ5uNeIbBr
AeVxHBGQitljEJ7gsMHHUo+Vi7HuQTe8o+wPsXQydCatkBalu6M3ur/k51iAk1mc/tA0Wsba+YJq
gUdQrfWTkdwwo5aAi9lk0MkKnRA6zna7BOrZcwvBmP3Glfd9/nO5CikuW3y8ISaPvrn8qB87L+xm
roAKbNmuqUPFsYZyvcfnMlvLEX+uyLPppYnadG1sKxhs5AgrbhHsuPRTaClp75HNIBvh86V2cACb
8WVJP9afnqGKwEjb/GU3Kc5Vu3XPRR3eQ46J/0dLI9TbB8w6AVVsOyqz+Ra8nO7E9oZ1csPp3P5S
yAouwwa462Er+IsLg76Do38uRezBMLKYb/e0BBFiaXhulY1kmp9iRxcvJuAu5UWZoIlNyXkABiJ8
DXdmt+EnZxRSDTXOOmhG8F8TrWl3GFjhEAnQgErAuUy7NL9votaY1WQzAxtFfLxhyyzjd0iQT4yl
JuZ2fiROCL+TJGOJkeN2RZaMEvqgbl6DossAQxuOZ7mih7qW2c9pwK36xftjM6QR2BU6uQDbOQHK
CT4llQi9rQmzMKpS0LmrIAQT7kCld1h7rIDQEU2dFQcsuUhJ47DOy9TrvgpJkyNSnUToC9uJsp+B
6ynYl2jLGWcYYScoQcpFeWtAKfYA0ILyIbYwNHRhdK8pXtd/tQ9NfBBieBpsXZrStWlJHjWgGzgJ
YiXuHm2na0A4P1vQjk04vabrpFsL8mRlpiitq/8feHpp0THUHGZuHzW7P43CRGJQslBqhteC/BN8
+BXOaLDcRSqcIDtA3rjKGRkpAqaCsQWKhHRXUMm+iYWWoVr1+MXyQm32bmsI1bOjqxY77XEGKIQI
FQxqnfEQ4Xp/Nzl2dLjzhv+I8qTtI28zSHvtQ+FNNbm4akM1lNdmyyljqdDYTJYobRdMSgMnvUlE
zNXsuPCv7ElThlj0U4hIPdU2tmt5SKPFPMkY3f+8NwSkwrmlbRbJnAMBuT4Z6SC4TbgpmdvmD8yn
YcIx1n7JsS4YC9FhGthijAYywzqFFrk6BM1Ox1DLxnqD1lk5ztJRLTCueyB6UQALLvwsGT/uawyn
VVU3oXNyH5VcFyh/BWHXuilwSJRkRkzQlgnHOsA8sdFiy8J2LHKjmEI2MOpqeJNJGrd+I7zMuSot
w4UDZEPOp6CKBQ5hqunhnjwpRxmKEEOi5rjkHvhPasdtnO6UEpkKyj9f89FFZ7JVr6enwNO6IqMl
3DodThDKWy4TXuTCKKLGHbezxm6Zd++4AeT29WCKDri3dNiNQTmSVQAPPHFDLzvrAqsq1swQ8eh6
sD6Fz5y2vN54r/r/QAaZzbwGrP6DMlZPTKdyBBpeqKUSWzaY63JStANPPxqoa6e+DRUGdQ63UIrg
pufGNsx1G0rxgew0tI9FjQ19fXmZwv3TvsDA6fW2e6sQq/yyh3q6wm+jEz2nOs8ZkJoDnHt0Cicj
1AWGY5TjV/frfv0rN4BGugq5scWMleBye+/p1zMWSvHHIQbqbZV4XBywOOkZLXoq015q9PCQw9fq
xheF9XKhEf59j+sgqxKJCkspBbr02NP17ahKOz5cmCdNOi676+5SoCBwNNxIcDFQLYDwqIoJLmTe
Tb9P9UWGCgohQVv1wfhduumohYyuS3dFyoWE5ZDFeSFzNkii/eiLLNCVj8gFOSzxN/qNU3Wuoc0Q
R1qMPQ2y3PX6CCz5n3YJCmfTUa3PV/P0uWKLM4R1iQqTf1I8AO4QIJyeYVoHPveavFpG/Obg/okY
DLRXiPjUnXhXLH97qYThE9CrbRlG27AQVhwz+0NlyMZ3XEN27cZbDBFH0Vm8R6oK3ejV7Uky2FMy
drRhDdQsD4qP4PipS3GFTGRPRLowNf+39g159K+tuflGjFQWD6eLcBZUxOduHv0CJnQHC4lDQch8
jSJNLFHJGJmdEbVVOF0Vr76VgqbQhR3ZVzb4X5IRxqfSehbsIR+sAB1E2f9tYPRiAqm7iADO9o7z
5jEQJ5t3ZAFASlKqoTCv+AU/kvnfK4oCNcI82OHMRy67DccX0/ddK3UYQkxzYBZI7q73s17H73UZ
U31vIhA40JpxdPdEITvwCNOfA+Jb9TvZlvV9JuXlUhTM7KKaJFQPk+9l+jlZXcfHI3i2Rd3gvyLv
RYdynZYB4oMnwccVT2kxFjHRD2wX9c3Gfkc/bwLCa0TireDPCE6HcFmOl4G2P0Y2RXlpnNVvY8Tu
7ktFfy2gz8NMAEjBWpIepjjJ4bbnuTb5WV2y/Es90wDOww9fwG5mSDSid6D/auEMv813yK4oF2J/
R9mq4EqzSFQXTNwW7WvnkiYjrbXwtqb+Hrg+JFycEUuKG7qIFyK061NHHxrhMH0kvPnXpUVX2T6J
/d1daVaPaxdtfPts+ZBnPgL/E0Plbl3tIvkCFPko3g8Rcc+pa+bhmpEGscNYu+ZQQjvFt3L8kz2x
4iBZAAzoPaKSaO8hpde0MOIOBcMXD1Cuvu7f1NBJYYugl5BvtZJS6UPpzaHl4E81B49A5OtBwgS6
5B3UA8oU1LLrjJaZJpHLdJLLeukKH1bo1A6jLnthIOLw7+Y2uWOBTyom6KQoCSO0E0H1UB0UsZ1X
cWe/QGb1UY7YGCqw9dzvWW++Tqzw+ycAV+yo9MSXdtbEfTg57FCN7ZjX5ZVK5KqLbqXFf8NsMHG3
Ms5DbwdwGwE9QM1QqnawEDoe7675Y+9atMnzqpZzZJV0Gjpu8l3B0A2P+gRSlLf1i1I+UbXHDPFs
xRziR6AMufNHbCt60NBz9TTHwhaMdG0+LEHsMhCO08FBTFy02zof4PyqvlyMdEU33qThqTuBzInh
IJWvX0PsAZMBIFVCAqKR89h0Q4baH94WDl6Inuks/8t9L1OOed/DzqvHOdAKElvuXNQ2PvTl1cLR
4eNWII4RNCwSX/4ZKE3jjQkbEybEMaPTIgNAEgCn0gmOxAfpZcvd3VNXe4WmFP9JIVts07Cu9/wO
n7ff36Mb/Ugzb60pY1Zq70XC7V5QiFIR+LCKCK1j9nsOOIV99bhnu+6Lt1EvaQDcbqc7SNc5lUQi
IKiAq/UCwT5iEZ8EzoR9Eo1257MdD7u4AT0mJqZLUvVvX74cynYq/MAKyu4xSGXBoSMJOlMSuQ31
y3A87yLcujpwnVmU0+ZvM9QkpeiZn7aumo3Yc5uQcHAXSdt2A+dlJ+M6xAPV771g+1eJ0IjeugVL
h2AvP6mtXO6vTM5QAWwRBOLGvkFmYWB2EQsX7orxxtRSsjrVv0zi6HWm3/T74Ul1aTTAwiGrRwS+
Pcs7pfSpbSWd9zc7x9/ytDeWTHZtH71fBkbQFlEH1qN3tHi4MvQghnZ0Mtc/ev5UUWhhUwUG+hFZ
2wHME7KvrwFSdSSbJTjEd5qExYRg+zTZJxzEfbpEW6Nrwm2DNKIDK388FggxdoMjMb2WpHdbAALJ
pzeGg38C7MkwTQbSYsps20ocOCtYsA6avaQaNUwjBahRMPXaSCyQeOdvPoHLOzljvtIvMJVYPByo
dhx4BJoyikSbSAlUUT4W4yOcIpsc+mRZ4xpMdGfvvKPjbVGhxqura118nc3TjS9SD83bygF2/Kj7
GM2zIn1WBsSW4GwE3RKJd97bc19dAKcMs6uUGIohOD00pGXA6oc5cTUm73ZTbddK8VmobgGe7pEp
1oblNzTCB1YMvfw+Qr9/och3Rw47HIBevC/1DEVtxXzLvziUdDySbucV9D5rTrEDEIIG0RkGtcrz
VtTXuTq9Inc6drKN3tIVRFHs3JTX9+CevFsBi2P/nSaT5ArtUZrDJiyQHAOZTJcbpyhNH3ub+ZTA
johshGLl8go4iGtqUefEujIDbov01ttW0Aa60zvpaH9nxd4wyB9JYfxbyEi7TbbQzc1SbRRtgsL2
BIJvd+ZhgDT0/BUIrZKhXAdpKe/Fsi42/MaXNSrMzUDPmDCHXzZ3wYPs1/buoTRAeD4gGNbsnsr9
fXm3udt9UfUyy+JUlKLsdrXjHFILZVoiBJcfFzapjFTLHq0TbQxPqfKCS+bFSLU5beFRQ+eXgi1x
eN2Uy7/lh1YwF14lpYhV8BQV5dSsMLix5roafxTfpCacmYx0rb8ZkTVOP9aTTkaJyJNUNW61w/1K
Q+Mt7jd+Ra91I+E139COSwqf2TjL6r1Oe4U5RA0hXfoGywtnMK2tn9j+1DbNPhyLCKh7CI+Yw2KQ
lFdxvnPwRxYWx9OSHwxg8bJvfJBZnjfrI0vp0BgW+dNe9MHmNNsIgn3jDZ37rXCGP4+xqD9p5eRT
i51pssnzUEeFRuz2lHSlgqlob1CRy3M52TMdEsfTGWW3auQ7OE2+Fvh9cg0AuIpalTr0D5gHUDUY
EP+3oMnFBiLEgoeanHWrzFv/CDOKjlEZu/PYsgKsB6pSHstsWfHWOiiHFPNHrAazmsz0SpE1QmpQ
ZNm2a33VvL5B4UjixH/hAEE4jAg1OTWkIOKNWi44zkHV4YSIgWBDjIGxXY1KDTFBQdIHXi9u3eVI
GscSru7RA7hhxKJThCVjX7BvPKe+OpNaRElU2H2TXv8hnA0DiFcUqeKtCiVi6yuKWaFME8T4E6ax
m2efJQinpqBlPczJkVVw4qf833S7upVuZ7bKwh8cYRafZrkiWfE0fPoz2Sfufqvh40LiHt4MOfeH
W2Ft+0EBCQ+FgTVRN16HaCdg+Y4fXErFdxf/PgM/I+6b24nK+3EGXMfClOVTSeFWdbFsq44ojPtr
st/J0VQ7f1A88MFnMlgy2YY71c2SZdyH4K4JYHlEM8pWTYvq6r6fHilSlVjMdYr6lLehGqnBVitR
ErGC8LfwPlXxy9DWQD0zaomSLU8/FOAHRcQ9YbxSXla+aRDXgq/OdS9ZPi/QmvXs7+1sz6q9K42W
MUkuCb53WwS2yab266jnzxiHXQLe89p4gR7+vb1wBcgHNR5PbxSgz4mWeRzaKthYlVAL3seX14N/
MPKONvvsA+sHwR2rr28cBjtPcdYH/wm1Z9zlfE8U1h3ttQf+CPHNYzMD0SCVnf5r/cm7o1x5Kclc
+9qnXtkUJGOMRk92csxvAt7h5DbNitxu1IziZhfFtykFyTNxXZqa6CTTl/EkuBzY5ZkabOOzijSR
4N068kJnB8jYg7l4qlp5scOaOCzUFncyzq1xKi11g/F+5xbaZFSSUuiIxpine2zXyP1zqWVdeg85
lhDhDMl3VAZiAuWpL6qexjgD2Ksb5OAXXBzKZ5tkUktz0IFnV9VYkXa2rAXHoEb3rZVgFCXyzYJZ
ijCGgV+oPjMXe/xKmLHD5Z0NSaJwzLXklXhuA/yaN1CPaRMGw6IMuVjnmAgb6CB2FQI5j9EFtQKC
AQCZTyHeJcxRodUwocSnRJ3bJnM9E4b7rvaINTcHbJUZWQVO7dQkRRRpJ+fAvLS1xXgPClbQKkgd
XgFGBnfd7WIyxVK5a1caVGHfBN5MBLOYWrtkTTtlsDucQ6SsZuS91V63hh25W9mAA3laowf76+Tb
33vk/lgjAV1LeTISksyr934GPEsMnrmwmnvhUjr04uOiFhd+AAyKWXH0ZUiEmPxcDK5Po5kLHDCc
3n51cuAeAKbyWoCk+zKWQtkk8VJejlf7J4LBBY+gC85F2YNREfmKH3HWLp9qAT1pAcDUZm2GzzDF
S3wYvRUsuOyitPqZ7nMvH3yL1n4u/uedyxZXDyVgmy3fXH0jdg32bbbvZ4gny6sFL1UeFjaCDC/2
+oIpLzbp/Wn+cV7J0QZcvfUo4v4Zja8IXtW8SzoINX+xMYIZboihujoOYjFaj0pTcoxUYICwYtf6
6/jZFrNNKZWgZRuhlY+Db/SDW4J1268zbRwG0tewVIOVUcfqa+aSTnNMdVjbznBV6Mx999OlNS3L
pecMBQim6s3WnegBPMZnqH2Ji5kV6qf1U1QgzbQIYlKk2CmWRc6cnCmvuSkb9cDSMeui6QpeFVYO
Gi0RKlfPNSkMtcfetOePlUOta4gcnHH0h7lo+RKSdUS/7/B5b/zV5aRb+E8i7HPb3TgV+hwParvJ
CLAGwketwX7j319XS8c2P9DJ9kD2JpH41/nVHW9fAEBB0AwD0pw25sb/Eg6eUYmANkP+2nKRubXP
mPCAXFobhJgUqWXX7trNT6qX70s8nM5ExYkNIu4AanIEVUwWwt1XscbpiIP0aw7aLw3wU2C7Rv5P
HPliYayp+zLQe3QCJfImd+bUihivktgyCTOWp7QXBN5v80Z3TwXhs9NAYeKR/lLD+a63xieLdUSz
Q2PdbeRONOvobBsDwzKEp5SzheoPjltDNpMKG8rQH+Cr4s2/BBvLe5oI7HfjHIJ3V2VK+PQHwCzF
VdorciBqnMEU25alWfmsw1K2Ohn0XJ5ki5KVHJ6I7AQshmj67LuqD8+dliP//n95P2nO97CZaVph
Lt9a2Nti++4cOZ37snd2l2rjvuMy05y2rPi50weZwXWHADAHRPjLkC/yyVm0+e24luP+nzX5Y8Qz
HHDvSxOunK+G6czZT1zXVPcosgU2KipAY1N/afF/JigNlNqywyIJzhT/nxfpzyId/zv0H+CBAOXH
/XqUuRWAOnQ5S70M+I7aZzV1EOLQVc3brAOoEPCslBZyTbSRK/RFgAj0Rm7ZIBrWERVPtEpGWr8S
wojAcmvqqHB0olSC1YuX9srlwHEvgaTSdtAh2Bbp9fa96uVHkLWiZ5uLldKECY7isOX9plsi8rwW
A1n1l8ecRZGwT5JnEwL4X5skx5zAqZNsYmD1JlLtCgwG7mgRuoFbCYWMxYDb0HCJbcvInyprMd/T
r8Zk1+T5QgcR2KHZeojGOxaawqy4+lBFS1jHAMginJlD4CuVKvw7jb17J2oA1D+m25At2YF+J8da
QYFgVJ58BKhww07kdzfEGXooJqGU8yGj2RqX6slKeD7kqAb47/hKSCyyobRcHSaurZyfUzrg+8G6
f5HxUZ9snFOyO+/K04rwZeJ+fLiTVbA+K//GVqtRUGISNojJJwKsZXo+ALJob7BUnP+OvAhoqL8U
h0Tr0mD9AG2LXS32qJ7V//Yp6K4wQAZKRyHkpd2GT3vDGFquQl89zTUb8q/8HqR217oh3roNxiuo
/P5avh2EBT7jlPsHbaf4BGpHpNsMbxRcXpXFnyl035RKy5F/iuVjTncJzEN+3SkYXCV657uTFnh6
NwcmB1wIX3GGZUvvzr+rORrjVBbBQ10EOOnCnWQCQG+7W7Gi0NYuFHlY/JhLpM1XvItoB1AN8HYB
CoKRBqs5zhUiHye5aJzJV7FdVX8Hgt4b+faRHTr9/65YtcvJZ8CH9ROof0trQTV9bLmJANyZAx92
grKdfW0n9Hr0o2V4d1MWqkS+AqTWjcGX6xD0LSkr7Xdzjc8q0xsefbzZEEuqczJSqvwULX/obL4T
NyqMBnGgLfXrvxigatpiqfsVlsubANYG/nmqaXK3tKnkZ4mZ6Sd/mmKm8NLb3Q5j6OiV6upkDpbO
GeKwwpCDP9Sx/JaZtCm54ehMSgHUq4Ttfn2A4xeGZIDOF0/ODi0oMOVCKtOlVH4qA0QAiR9rQJ7y
miMipKVcnP5sRQxB7VtW3Hf8Q3yychzJVC5XAxfYC1zbhU5G7Ia4gXUHa6iR1f8/1NhYHwiaBctt
oZ4WGOtaOZiLRVDR5GkxCV7j20vtFV3zbmhmLJj920ydJlGS/v2ORGkvrpkNHuTglsY19ccFwcVJ
P9PKxCyjjEz/piTcbxwsF32D5gVUj83Ifdqy6X/sgDMdevYWT9pNUF5IzYxGkNHwB/ETshLcsEYt
x74CyKl78Xk3ZIcBh54AOc1nabJ36xtFStLkC1SqbMesE4C2IYG2+GT3c4o/J/KsevAYO025jXjH
nvmTpejlmv1e+6p0/LvAMmP0AMfC7vRF/SwBhxexQkzbw7JrkUzLwUnXVexGlzh5FWGnNllAOdDX
LyUXrz8oEihWZxFGGNVm7O3EAzcKPR1jDtesSe8FgrlyzzzvZq9cYB90ougUQ/igE/jUyWEmuR+M
pvTAoSfCSFnm2gQlflQeYfepjSvol5kGA0plM0pKu5t4GpeDo3x0GIZ1AHFclQJUsGGAdO0DpT8+
85THYMhTbuhDtZvWuoSPo4X7fpn/klquBb/hckoRfin0+CXabOeTNRqtnB/8ILQnGz0Y8BYFxCZJ
iiRWhNn/rxR7j5rVtQ2dh0AJ7A2vqXX0ZemU3WI9dTDucwLfURGOCGTcVesFdze8niV2ovMcqM0Q
khlZLDqorn2jcXDFUrZcTHq9vjpzp6K9dutfw6RYMDevwHF1OZfpG+t9LrjDqmQXoob9gXftu2rD
iLVJB5VG4pEVzqQuIa7H5NMzhMVhOLtm9KAC/AWUHWs37rmrXHrFVRrhDhYv+Hp9s55GuSSeXDiP
CJhj+L7Lp6xhZWmfVLQ2x/h/+lwn8+brbOwplXlnNLngyXusS1vK6bOFb6qDn0f9JSU9JLHbkxHz
EtUjaPIieaVb2IUoOQvSLT4b062rMfm5z/GM9f58xG17s5rCVov4YcD5y6w8ozMy1WOEFXbHjXsd
RmJ2VEsRDSzViDwJA8j4HryJSymT+e+8SvrGxeYbIJ/DzShuViZ0LsVvZnpjwlsHzxWtOSrxyB88
t+dLiBEQuDloS4yrOg2Qh9RODyMMoWbmDeGFzyrVT8ivWWhu1NkPtdTlLBzNH9scuLdqTRE2uaVm
clemD4/0gjUj24IQOUTYbAezuxM/dIDD3Vl+QBK61YJZgvXte6gXFbJbOjIOck4Zj1/TBXV5+0X/
OkTAOd7x6JU+8Rvp3uU7LgqXhvkiIRsVQwbDS1NFcgaPDOGjJxoid43PKk/DhOB/xxswcwRn5lMb
5V8ugnJopHcoW9ShAFjz5d6i7fo1l/vGGXcXU2JXu63d8U2+uS7ysjhygNsp1Ks4jM437Kf5+QhB
udEiGalXTdSAupS6imt8Bjepozmai9uxHRGkHu/XIAWHfTD4rlOIGjVe7eXSLKvsBorj/+QHaAYh
t/kkjj/Ds4g1sdsKOtojoqR3jjD/q6E9MbmAKiyD2eZzjydq+BfLpPWv9BfOJZXlstAe6f/9A8TW
MTQrdVFKjyAO9Pl7W8N70wjz9Nzch6oPrU64/7tfOFnjsj+YKwOMhgjQn9oqkKCC8eMdDbDq4SNT
g5CtM3pkcSmepzQ0gQ2j1d0ia2dRFE21Tzzrn7AIvx6UWOub1pBjoZFkWAyvmYJiEso+YNlk4L61
A5pyMwdr4rF7fABpgb+MM+aaaIUvfmAR+gMUBWB3w77aavhSZyIUWuJ7kqpEVIheN4jg9GTHf8Z+
0qSihQ+Y3ArGPoYFpONHq0WVzMwsp6OXddEt+C2pECF3QNDXV+mGIlLMjgE7se6QGF0es3kGl27A
43MpmJ43f1E0T9AORdVp8sCOtB3SBt8TpHctEuOg9CZQjSPf4d6x9ZFEv4ZtCrzVBPgGwgYH7DA6
bTJ4MuIvwfdgXEOYZvXZWx3tbuxE51n1uN6MZH1nQz/EazNEcZKJDx+wwftUss6ngsk/Xcp1CP/P
sJLu3UkVLvnRHln84bFY2tjJDQUbHSWJqH+dqKfJVt1R+ZBvABUCZizlr9cphAMXHLrW9FP8AXNc
fK34i/EZnaY1XKdXbLXCYTD3oggW4yX7PwXtLurUCcjXCGuKAon0Ivnm/PFttvXS/xrUKo/mRr7U
098vEqekL2DzlymqG9fTRQnMAtbaDjn1xmoVyycTk/aikwF9HErK4Hb7CJyT0EJShvR2IrpV0rzK
1+o9zVabs7kPJeTx5nvSYW0rNR+IjdSZTy/gqvtnEWjoWp9e2JRe8ByIFuXw9JuWTCeQ1lW5ByAU
CQq0O/ItZ1KmiSmrSVuOGVd7xZ2DpeD6ABg1Ne845XRDKDVeAHkHO5PIDQQLQZ8oXGuAakVKDmjD
GuvXlIl2d99mlxHPdK3Ze9bwuj/uwRNkNFsaxKOk0iexMZGO0mM7GSPQvIxf25RUFFJEDAwC+8Nh
20SAUlLpj7zHPCc4aPcQNQi0POvIekONZt92acPVT1rvXK2fyGiGazG1sSEmkwmymhYRBXL2lmqz
nua5xV/2WKS4osKiUH8giJwbMrO+1hYCJ/2Z3UboiSXPXQ6nlyUbajDI6idBfkKZaNVizZVkLy9C
9TbhhA0rt0bQJo2q+BJOFKIJRJOhDsaG/ipR567jhY4NfuuXKN7Muqi4cygYTs0oWJekb+BiYxjK
yC4U92hPA+T5INDIYmpCQxVb8C1hibIylCvFG38TINSw6erM2JMuMG2sdE/mFESEo2AZjRiS3Xm8
oO7rAigGHfftXauJ4we33Q+OAWkcdDrTDWY9CSBVfLzjsYjVXJ+z+D/M/mioowYPYn5J7CrhFSLh
fKmt6dvk7WvqAL2UkPX1H+q5jyujb6X2lsN58jhxctqWAFisEokU6v1MseC/Wk+ExW4nb7PbEPov
V1tmJQQq70twox3vouV9NQfGSa/WaIRoAI52zNb4svSE/NkPME5N7boT8jtEmH+cnIz4L1QoOPpO
wj9obXZzpZyF7NSq88cPYv4VxfdUDZHCXnUVMlkoTSTspKNWvnzEcYTjR3LiaWTkxeG89J3zZqij
gdIAIxdwaUVkj22o0w4iRGfXXLpQuQzY7fQ8hlgLefe0rnwJR4EzWw5M7oE+toQoKNj3eODw0W8o
vy8fCWiKExVc1lwotdY0PWeBAgHYD2xAx0u1yde5jYZ//nLuUH+QN2T3foYhAmKIcOwwjt7RLxl0
lz3XkMG4t89M8zSHmAkbD0CKWOJZk0a0vIg+pxL2P9CyA04lgUEJC8KOF4sJGgWt/ahU6JUWb83i
WYcti6/GjWhqaRHZP+5SWKie9ewRFg1SY3qW91PsBZDc+YFZ/Hahhd7Uo27yT/EsczTBWShG3jr4
HLhxq8z8qI/U6Be59tAjP0P5sCoYn/ttHaupb/iNsCseFNS0M7WTYgYlajMwsY8kLphrH5nidgQO
nPMmxECgjiyBT1lCr4xOLuYOaBdBzFrqt1FCOgtmRgx4Bmr1prmqzTinjPCDSu8Up71TQAs98gs3
M+hAXf4/bdMmgS+MRxFkL+4k4Fdf1Rd8JxkyHYSSKQ2kUlw5Eswhh6hrxnmR+emzaiwfKwKuynF3
9iQ5ulObZeByA5rU3OsWjvAL9jYDP+P5JqZqz2MNvfJdxQ+//LSH+VFcQKWjz81WBwTS2+xP33Iw
7vcBIF46awf2mNLr4Bc+nEbP/53uxgHcu2s5LEDR606SS5lqD0iWfGQWII7IXCrHqJc+4dPS/ADa
87m98cB72jGOvE8DwNhLC+6ufyfG2XiA/G4A2PlK53yVsN4z8URsZFPcycJXSc6W7wr4iPC2eex6
brqFxLbtAl6cY5OTC1PNtn94awwfyDAhlJoDrhF2sCB9FHBljpbdLm6khJuwbKwLasU6PYvFZcAJ
baX/pURLtVIKveWpsGXdcNbwV/lmRJz8nW84TsSwU4Lfsu92jqm34KgzH+ZPQz7bZPvC7QvM3Z4Q
pEtr6TRR9z2wYE0pN+xdWWuWbRiW0GIkvNu59jZ2dFOhS5ATDKIg1kRx3H+jhjkGqtiaFuYUqmjP
vzkbu/4VPYrqsepIj+hk2DbuF4QxF7UPkXAINST9raic50bHglZF/orfRChiTx6uLGND56gQhAZP
iD71SqesWiGnce7TMjplXQcEKATqsMBMjjTsMvTmH4FEQNw6LScoDjdo1UuZ5FxB0VaMhmhMFJt4
EWmmgYDBuuXGm6DvTsNX0A0KaMCT2rphrbl69PLIaCO077O+zUcGluBFoc9V5xOcMRPXz0M/HwKb
3NMIJDj1LiaDdwX9kXk81JUPZZmPQL+gXT3Czz3dzgIO43n9LJegLbuqPQZkyj3IZmW/NtTjllyG
UbkQ8Eyd20ENbWbNSN9KQOpy35rge5TpHCUBCz1hKvfrOPHRb6opCgqPSmlDjCzMkYuucAAoXjXE
L0rvim9RFyQtdrr7cWbYJE5XfC76dxrYPYcb7aNJyEhv2+1aVRhWWtVvxB7JAUf0LIXQAMqbb3h+
Ck3lxJIFQsOr+/8JPPs0TDLZn6EtjNyEK4vdt52iwml1UDgvPqWt/2MLxRSPG3PBQOSGLv7mbLP+
+YcSLcCyOtUazZS2EK0fEfTaDhHGQI/fjk2APyyj1IYYgXyN/604JHI+yWYgK+aOyXJAAVTI/m3E
Uoqf6P1kjGze1vcCzlWNrAQF9OIAr9CYUPARWn6LCLa6wE/pOUaLbOJTBbE+uGTzkVZwstGjH8tW
WBopOOwGLkHIrYY2nf4KDtoQDn8cNB9GHet01k5LPHLeB2nfSUYHjNBkkH5IXnCFFAwBDMBhZpbG
cReBfWmU2+n1RMa3cqmrPu8gVL8WH9TyDlss/i4T8y2Do5e83rQTTmD3qFb+5SGY/Vhc3dOpvbgi
S4SftER3d3ZJ8Y7FF2mW8GGZlHEEQgvHDSyNA5NzUib0fNTPC/6yaMge4jOH89pv3cxV8TImITF3
M354YpRmTGlyru6HVVh9a8PYBn68yI096GPo1QY1h1SVQrmzf3CYXiYajzqlzfjhF+SM6WbouAY0
EiMGi/b2mBzAj9RVJXZLQ4SeMJsfZFg8+08RUkQB0AymbzBJR4ogrBXPYUDZwVkaU6FbBAML+v4F
HE7QHMSEbMTvw06ukIiJ2pUc7KY7ZGnKtx+2eiBeaGBTfksT/5TtuydDKpb57XhVEMUrAw5lhh8E
yXKx3MH91pjrcDQMiOwPZwg1kP5jRXdEFiilX0XnxAtyx9y3ZP5WoeRMoFA7YwjnQ2QHHox3GL6n
dlAZZilXhhR66OYDjWjZla8tyKB6LtfPlJYR2Tq9pVA4RmFaZNBCnWfnZVD6LJ0E2YaqCLE0r2vD
Sn5ZcNlLO4ycEsSDvDwNyJ4zr+1spdiqRPhgDhNBvDHMQEy9AhESdB41NYTK3HXd9XRF9TBjdEfU
dF9oSU7nWs0Vx4/i4wscyGZIZBgFnU6Wkc00KJbyhGUXFbBVR4lhFXjdunT4507PqlsoYAsmT7Xa
Fv6pvzeLJHlmlBNq1Uikdo6TdlDb2DyI57/ThzA1U7JtapgvxCOw6/k3Ke1PGTXeFn0SHjsfSWYO
XgOxHGpiaGqkoa0Mxqa+clQwDOMXst6DJHi5zb5M0PMyuGBSK4RFvrFVg0kFc1pqMRVMw6LZcBdG
/6IvcFKz3eGHMOPFoqg3RhImm8ZJF98BuTCL4roCCEtTmk85vMYQwJaoYxGoteljlC3gL7OQMhj6
CAkyyK82wLyliWHIY3s3aYoBUC+2AJV0fgoV2ds1VMk8h85F+2QkXoQEahcPd0DS5FOgwE0tKUks
uK25K+RPn5QjENGEgr3sYEwRAKv2/mIb86zeZbMxMSaeHJIemcocJwv2ZYk8xshg4cDcx8Slj3do
SdltNtq7XhMaYyB+u0t7dnTjrGGIBWrrcnghGS1FUqCmus5Y8epX6M7vTOleAc5VNPJ2WPf46X+q
GfC7ytg842+L
`protect end_protected
