`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eyi8awNJ1g+09H4uyqBjpOQgmdL1BMUW8g2f1WNdLNBif40R3VL15Bg5mVSjEhu/MrZVqVV60ym7
8YxbyNqErA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mlf9vrU8Lh52SUEuxQkUpz64J3SYRFjQ12n4wix/sw3oTJa6muxvidfpdIiVFJ4blIkTQkMRPkbg
fDj8h0sF9+AKTeU5zhM3+ZU/fFdbNIC0Q2X8WMDlMi49K1LWyKM79UpzEDtbS4ALqVNafm823hPC
pUb2/Oa3db9A37SUNYw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PV9/3mPNbClKl+m37NsVrdnraSBAN3+giH8XQPhuM8SxY9OBXQpcetVIGg2Y9Br4Aw7LX4WOezA1
8iP342awo0MzDnKqPYSHvgKVqPJKurlCaYRvFX9+eUrO2LxjosvkHoXMyUkwk5XErqQ1mZqrE31s
IxEWyR47zzTd6YIoocBCIRQ8C7HYpCrAv2N/6SgQM/hNe+cV6gsFkwzJlm+kjCCne75M+/GTWwZQ
wQD+PQjjxKKRCPix3sPi687M9kb3+/uULywesY5HeOPKyWjNBFFsu3eoMubvAhqTr0wBpA4Dv4VK
xFaC/6YExubulX72X2hNxb6tIopLxFpklSzmyQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q4OqcZBA+jABGBs1mOeVt7TEhR3lHLDumRAKZ4H/7m2lbjSg8Zd07QvOOn2gvb8hTRrHKDiqloSl
wwiFYCd5QySycSxIFUntNs11ACMa4pe3x7ZCtp2WVu6uWnqiFOUfs9Cgw6N7oOB8JDBypVcBcsVN
O+s1kCPgkRKNHtN4Ckg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HlYgvM8J8iKqtwQYE2GwgmChXC9qyK32U3u8iXxAuoNo2MUM8eJAT9Ng7m9Tj2ZxuL+f/3k7ZH0M
HhGTHhmk9oElHVUSc3/k/UmjjzKYd1EtXdC5qnnYxSlGsd3IF6x6seAqRP+dZvQzPIkLgL+qKNBn
3beL+/WVj/Um/2BXqISRR9UfljZjs8NsHx3qnkCcHerbHUlITZ3EYzHlciVGeFkuXSwZiX5kVwep
nWjwluDzIB3QFWDus5PIk8Gl/Lp4GTQUhvKgf5wFR0aGCyZSX8FeCzW3XBjUNeATFFeZZoRr50ah
zYA1lP+Ok/XBVBvAeXIeMwAxIATzNohyn/LpkQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11888)
`protect data_block
oYPjLnMmyWtY93MY43nLM5KXPPTRwXlGRboAffPj/pNFdrLjHogz/Aihv/qTk+udmi1xhf7YdEry
EUUFX93fLWwCuLz4hsTxlex8blvxgPTelI8scwKXVlO1fpfmcmha+WwFRK8PwrVZRXF6IWYNl3hM
eVIA+VA/4nFB/geikS0rQa9OKnJVXMy4vkGnMis/VZDscxiEGjrJywS8xBqKtVWZPWKNFvisXlYp
jTqqdQAkrxBHZCZRlVyLJ/4VTAg9yCuB5Bw+O78lsKXFi2iJzAhcWr2dpa3J0Li36HVCxJ/W+KM7
w0fAflbf7W5WPiMaiSPWP7ix41o5IlM5JJpDjwMypPAScNbW/gmy+41J9ZnUKMwmj+t1wiSkA4LQ
NdhEscZTWS4XdIlHvtrkgsGBSqHnudaty2oO5Pmryv01LzMOUgIHvGL11E/l7ghdY9IlMKyYii+7
TJHbY7TytCZgyhipXZVltgIZl9sMimyAapO9HYpyxOggEEXJXbWSApBXkBSTAaqIk7bUJfahqLNz
lH1H5P6BV2T2+HO4rfHBro6NyJxlOF6eFAjc/BFNLUVVUyzwD/rapL1MbtgyKNMfnWG7fxpqdcNL
KtAdxgQ6xGFIo8REANju+jYIn4jhFjHHosS63AND7mlPrufXyrlZXKqvwIIjGmdJHpHWbE4QrFi7
8tzxytoXYR6VqA+yuctFKC4p/P2VU+4kjCjlEbMMM45Z7rDm0upHS+08pAa9yiv0ZTOShuiZErvu
fPzPO3x/NIk9avbM8dmrshBa+BBU0OwD+O0QH0NLXRm0Tip8ZXA0IifbCj7VV3EHJbC8Scnmu/xT
1hBh9qO79M4tZxe0XL4cdQkfEKlSyidB/lbJpG6Mc/aMAZBFwrvJcwBA/zb4zGsae9A/LAkQBaqT
9How92+yxqi2BeiUZByCcoohZJYKtco+8WNVQp8H6P9aR96vbJCU5OHRBFjPNOit4RGXq8CBe84/
kCt277nr4Cn2FPfyrak7fGoC+g3PWL2KLpqGqO9XtyKSbGFkJdqRATJFo+SmmmAYnroRZzZxJtpy
57wDe4AfVihiZm8k6VIfTx8Hbji087QcDzQZepgtRMvpePNFDi4x00ETWwSeqFxjiJEZMrukO3ct
yP6MdQwpYv/l5Gi8NSlijFUU89XdPzHLvKAzq1MSmEg9Ej3TkrHtSqfx/mGQiR++UEDQ/W767jor
/vP5bMlclyvefjF5YP22pjAMVlHu/rnAzMOwBgPrJJuM14EXL01j1H6hLVr6UtlVf9py6sdMw2y/
bMfjew8+OhA0Xf+Yi9tE0xBcqPh7KswwTcFqmRYzth7Jpcw6RSf/Ujggxjqtrdys7gCo6Ru3z75M
14wS2Bw7QilGoKt4WJyCac1py0GgiJoLeTKAtXqPuo4RlhvkYAV7h4PlKT9THR9IZtZiRG8cFa5M
p0m2rBonRmiraar+2VIIPSdNayxlluufpbrkzfa23RQnWXTaTalDKoe8Ma2M8beNb4agKc7ZSjsi
8P3dKaxfQTburyB4OMWOzrYAnYajdEe2lilY0zXRLf1tV/ZA/Vgat4c4vTB3K/S/W3+kd8+Xlo9i
DBGqm0zjUpsfi0VZ+NB3gZgDifGFi62Rw/zaFSJeh8+pU+4P51KwdwcxdEDaNFgV9xn5VN3rwf1b
0Nk9HxYbxAPHZbmRlylF68qEMA9XoJKbW5ZZYpcV5qmyLgtiEHJeyNCaQZeDxeFA1eMrJSskJX4h
o/DKXSzIVeCnA9DI77vtfSROTISuOat2tpzLDwsbFW369GqpUBJF7UlGpchG9GTkwCSbXGTNVjrO
30G/1sgQ+gbtFcf3WEavyrCn77kJY9dPdRoxxeaBZBAcFx9lq6pGwSva3jjrPWtViKM8/Ybjjpz7
CpTyxWPv1TtaSAddibrZCJGRBhI3v/iDXIs8xVB8zEZ4rVRhmBbgspD/ILFLPLTIwT02E+24QYK9
jRqBfy/gx4hVlUkweaJmyJbOsi0lcyyolqf0eULGAwlqlThOS1XJ0oiCAAZhl/rw3YZTAWG7Nsms
SXTH6b3+G2E9zRTmBoEhPNqmUXKXyPsfFC1Pp5fHTmYvkG5WRM0qVbBl8kb3pZ+dzg8BqNt9G7e2
Jh8Kjlfr8uZkmXKEaLGSlJM/lcBUUrkTfs9mmvR0gRO95Nj+v6Npq91L1zBFfcGtvL4pK1fwyUca
gF4Oa7pvNb+nqkrNchHyMQAUe9RTY6IN919ar5RtY5cXtSnp5O0Q8hYUrQlSwvF+tPrKL5k54c5V
qKd/mvwvVEe1DPuco+Gy8d2DGw1BedsOUhlrPTCZqoxjio6OU9+BIvcZxh0HGCZLufbthnI7kOAb
uZXLhQ4fhfk+fSzm1+JBpzr7o8s1Dm0s5quNgBuFZ6HSmdAxP3h1+wFRITj1e5Q12xXftivvteNc
KgK0ThcO164FHSU3cxT+g9oYXAy/MVOHbqWvxzNO1HZCTNahFVw71AjyCrlvyobUGx34otqPa5Dn
PT+7gEoxh7fjeb5hj6/CvdenNWgXVq5/tCNQ3swbNMnXm+ABi9HFKp4bh4Zh+maJGQE57yEDlXTJ
ztAgOFDO5cbv+u6e2ZzbsbH2JBV0XhFbXaFFC8VMOZZTFT6xDT3xAFsHo97WSiOo9ZOMu+cla+RK
/AreLeMg+u+gM74TWeIvittSKpryxPA5MUoFm6j2fBmsT7VtWNF7L8S7Wiw9K1p1T3o77hX7jnkN
ootTlatuqyb86cVTPpt1QW2zqu8hU6qtwFvi0Lf1zGtqspqv8+fyFCMB3Mn4oIgglGLarQl6posa
gb3SzBQwgj5Wy7r2c67GQ5aeS1lCTihYK0FkJ+ABs7R/ijrIT38ktk4dwEK9diXIhjxC2jQwZzP6
6H8eOYVB6FEAR9rW5XJoJHcQzsOiLSGU4xDeq0XwiVIm5HfvCplEtmAJfc2hApAR6U28nawwJXDF
BgfyCD/pnJ5PEF/R/4o+RCD6SB9OTLwjo8rGAsdRx/xgUY0fUsJF1e8k8qgUw9NqjtrzJkroWZf+
q2M1LRD/x9TECPEaGGpRZY0sYZqkYZzTrSsp5pY4QdeU4RdvJusFXTfVDe2JINBDaqqXWvXbHgIB
YcnLZ8ZkfMiZ4P9CSjHdXF1iUqa8HI7mvoULNRlUVJhMhy+3d446OArl/lNo1zQoyDBJfUH5M/Du
II535pCNJJ/6rVBwXIhu5WAqX7hTg9nA207GRsEkKkIm9TwOE7uS7u8ekfacdk2AAeZIUqbpcp3a
HntjZPYYo2Ahz8+7eSaro759uOKCG+G9RCBkFvDrc3kyXGS4fkXSVtf5W/O85qgPaNZrGwRwiDo8
YrCm1XLSOgqUhYEtwwmralISJPHuDee2J1koKI1Ur9t5BxHaKkbfTlwkZGED6BfvnYN4WuBsr3Zd
3CIdJ5UW/d8gKFjMeC8zxnr6VB4XiYQxeoY1eq6SulI06vlKxKZZ0siSmSWrQzWFLVLoA/wJkHj/
C8GOYCSDFX2x8svsQYi3XevaKKHcSqKMdSaXLZY1dF7FfdjYUgFjgLTVDmqd5xib6VuOP1ujwmv5
dNQ6oNl3dNOwGF1h9lFTqHdxkKc87khNCxeeA6HeKLNiyRyDA5B9WG3Ja9Abb2daAIxXd8lQ6JPD
py+58Vus7RASI9AUIRJ+Q8EFCGEtV5Ia9ehR0wHFBXGyLgUmYMLJUqIq+n2582kkqlKZp7aKAv15
6S+YR3Lq468zocD0K6ZDV0+1CF0SJ08AFeIZBXm0+8SehRHhrYHdEIopuFH5FR5c64mEdTAyKDWf
4nPlKHnDLrWbHvdfycfXAc0Mk+JzDU1oUy5/P3ErxW5jaenZYMppQsAmVtEjPSJaEUg+kf+W6w2z
OuHHo1cKnRg6ZZFaB5+V/Ma3uDdUp15zUSIk8+K8jg0J9YzGI3B/m9a1i1dQu1g20G7nOdamplLK
ceOXSmckeaiaIcPSXfK8YWBte82hO0NVo407M7MbdW0d0i2StdutWp/5BSXvcI9qgmhOSX/qaKxz
GhPRwI75/f42UqlYz53XM+7ixPO6R5iCaQ0b00np5L6J40AI4kTvf3wE3gnOmyeJqGbvT8RVDBui
TwaU1Nvux9O4ESGqqUkKGPFL5VIN02ABhhBBIGWh0x6BT3rfD4PrJVEOOcCk8hsshlvOcRbNYosG
ID+PCTj01H546u3AE+vkuWbQtum6eSpgrcUH3bdRQ+vu9Pg+KBm9xqEl4Cy0fMcZ/Nqm7wcvZYyW
dx9jwZk2KgvPsYKFMT7DwqoUc+z0o+aI/V68sUX8kCwR/b76oxVb2Eae3MC74nkkEY3DxvQVnJzQ
qvrQ3Zt4Nz1m9L9uLtl0wZ+rX932DsdNPd9TZYZ/hTu0EaDIR/72MxBG3Nj1Uu1Zlcg1j/eDh0uD
WkMOGz4bHlEAwmV9s8lDM1uNsg5I93+Rfwdq8zZxNib7qxKvRMlFQpvAEsvrijvOKG109SoUxMMH
mHPo4ZwtcPJ7vnm+0EtIJ2P8HCNOdEwb+Y8peFbe9pFH1/Kmd2xW4Crl4pw+tAAhryDMgeS3FxRp
uOsmxhtEpAYx7WqKFqgZC9Lo2yWcOAEdtuuk1yN+lWNRK5CJ/2tJQx+Aw2qxNP0XlQlPvZVHCHGs
eRZjC53oXxRQzpvEtueUP/rHRkPrbu4Oyi47u7+NV/nlnPcpM38DUXFGUPl5VPI2tqNzFOZhZQbf
eqIFTIdLfsdxaME4UjN/aS9YsRB7XbvRkgkRY0D6zBS8kJl4LGt/R3jCtA1it9ZJnR01abV4OSa+
nDpdlq1fwfvF9u+XW+pxDF33PtR7ZY+77UeHxFcNBTf7IXIgbRTmEwtjBoCcgvY6IZ2/EsHcMVBd
EQZ3vzMoONewxBCwLIy7pxxJlCBn/Tw4renx2RiUbnFIBgYmhT8ke5bXQ8wtCqPQPdvGVRR7cuP/
0ikVPDhRgi2QQUN8WG7HsSJ4REKhRAPMYdqFJepnIwitaoBrRgIkM9RHRozu5Fbjz/eoPo2cpm7c
DmZj+bSblOAuvExooFccifHCqvien9Exm9iIqpEzCIYAauVYdQUPHk3etVU257fi70oASYtiId5h
kcnCWX4NhDayx0adSx7djSg1QJQFyb1C+FAgfC8Qu1rVIXJbbV7O00pVPtE/We4oWzQuFwcPTH+g
JjhjURI+IqiVNIcuB/0r+gMZiLLnzVm4FTpRKUt9UMFTCA/Lc67feiMghcmgzyA5QlF8QpeOBYgd
texcOjMVm6e8cwoMAKEuO39ZLuXr5dCfGu/CpRw/QAtz+MKBVnXoMkXOJHc+MAckzwjsLjemdWIq
PdBK8yg5Pgqr9r9i4FBhWIktCRTs2YspAdBdUbbXo4NDvXFma7WEg3zbYiweSQp6SlUqN5ngOQ2l
Vlwnkvgpaav2MfWWpfZculCCetVHTceurlNtedh7NDxdrZ3Zf8d9EHRciGfokjJa95/a1SmpS1qy
o++B4RTqd2AwNM3HUhzOzWtE2MIAcr8WyWFztrm3Nt2vpiagOpt5T1NmwNdT2iiKBVvImXnycaZ+
ivXRZfYtMknPUCFGtxmHAB5XpxzhfNZ5RyZf2ge0xwTXBS3Sf4cRQ2H0z6JAdVRSU2G8Q+cip+B+
RagPbqKAkLp4u+zte3cdnMic6qXokUQoFslaEFyvGuQE/JlLhCM64AqM1p4QC/elrUJ6z0PIpX5t
G6cXbvbXCQDI8azFEijeXWsj2fVJyWiC5RlqVvdfZI+YJPRAH03/9H86lkW1u7UgVcKCB+8s76qp
K+cKo1j3WzOs78PRxNW30ojp4RpFtJRjajFC+k1PpMPR22+eF/6JF2YRoAJlfNm7HPem2qIOcpTk
OVMdFcE8mW7uNg2XoVRL4vmWpMxrXpSgGmsd51iOggyv/OVp2znGLG+1sshq5j+2m0+S2cHvCqxm
BdaeVDi9Bz8E3mxJ2ixZChqn3KbV6uS8xhmhTh8/3AdwUGWXVjpKaoX4Y+HGbbZl2Cn29Kz3gy7O
mu2zDelwcL4IKLNP4ipupsU7VHkbv2k9p/2brBBhl+M08TBov3azjclbXSLgmnxIJ6HfaM3dw1cW
wlbBlITQyvtNagzLXMLmj7mzENLQ7gmss1/wb71sqdDocJKp0MpYZNYHPbqD4mSG+mmT1N0hXnU+
7fds/RY+T4yKUakyXA94Pb1XG+m377erIvLzUIYQ5KKCCp7xZcAelYk+Wvm5erTsxXbVj8wcDpUD
2lY0plup+OIepVgcscGRJ7JmIJ1qgUWpye1gW8+WV3/ZrNb/z1J9b+6qjvLqK1Ft+F5vIdQ5QTd0
DSQAX3QNuURIL05bhkWh9EpXJtvpHUeToovXY3jsx0/eIr7NnuvpuFpu1SfehZcHSKDloBQ8wKJj
zYTygmdV5glvNtchQmQ5oA80HQvwLfw7Fp/frmLOYpuITyQPG7+5NT2LNA91beYi6xItYECV28Vf
4H7C2cJfpgTNXzpDcGSdWhdWuBn4+gdJA7Pg3f8/lwdyYUWSiHqf1Hdkak0bQTBWCVAka8HhDKxs
3suBBXO59mMcbjntjw5YlQq/p7D01leghKKwJKB+7Bko+B9TXkxtJOVqvVdgZz1yvijuOVOVQq9A
uGglFwqPMxrfp8uZ3dNHqDOlY9DohdIRt1joevylFY0kTDu1h5cXs6A1iS9iFvZXGepjftUrf0V0
QdeZBrLAUiBz/V/IHus5XY2jYZ6DPIWRh02vnvz5HRWdPiXIOt7Kkuxii0XtsrRFMYmEXQl1Vqq0
V84Kefyf87OXhAU4ei+MazbGumwUZPEb5iS45dhAdYuh3uQdvEqjRKS5Jbm5gEpIFi9BHrkeBZv7
LoaTr7qHIhdmr+AmczK5oMzBGwkRvUuM3ExbuYxyD6V9eImGNDPb+ZVbpBJ0Rl2G/2XDltRF5mvZ
NcEAzt/5Fr8JrH2TaKjrC73NER/Aw3Jn0qD1zX3zfMg2J+EJpAOF/cVFPY1kHJ3Sb3bQ1Y8D5D5P
PTozvOo0NphEe9tVtyVChHSHiEIp0FurrEtS9XN4PxCze0RXOVsLPAV3lVDP7ZYgeLZyPdqA+xkw
0KJcTPs7ZRA32cBAhknkg+E1C7sD18fGxH8XWEpPjH8xVpsI98lBSiWpP/H5qUUmpzjQVlakA2Q/
GC6JR/AxnJzQBRmxieReDcoMnECKrBkoJC8bL0o8hVkK0DYcbj3ICe/LfK8dTy1o6mz1icroTzqh
yuousfWFa8Si8mPwV9rtmYclKxY+bC/fd7ykU82mm4lgqCEMpxIfTXyuDRK9YT1FfGG87OqL8Cnk
yOyIuVlbDzRxvL5eef0IRCbOHEOWFbfB+jdDqrAV3JRd1Zg+6KMc7Ju0iVp75k+QlGZW09a1v6Z4
0bvfXou+G7JopL6LoaVh4E+EWwmw7EdW31PgkTRxHCj77Hn19e20Mr8o3EJj5MUzfZUPDmtxwInc
zZae/Eu6TXKnbXNbeayIgWNbT973JR/hUwXoLK/RAFrhVDZFpQ5sn1xWv02TLI1V6yygDi7XxQiG
qEPOk46hKcy3/nhjHecWzfJSitbg1WbrqioEpcTqaXWForq0KSQib11XK28zm3eS4Qgk8VGSaS5Y
H946giMiTBW3US0Rzwtq0mlolKAIufXXhzKOiSiUbqVj0DUyYRTC0UVz+h2X/egroafiPosoqs5w
3rhOPTTRCDcTIDnWxMqyw71DNEY7ttilFDa0kDnLUqUzAD8OmZZuLZnk8B2Bgz6MWlYNxdwo9E1r
gvVLy29T8xbv+zyH96IQtX05kj8YhzZLf3F7ogapkaVFFG8uzcIS7SMLLv9RVVJ2FZjsIpGh8qLb
OADecyeuepZ5m7SGLqAL8dFL2350sfg8gKo61mR4A/GWvWrzvfm3ixcBq0j9cFgOP1K56vulPfOK
HetKyKl7qQjMzQzR7riSSBq8kSNF2M7E+nhHy3CS3lQLEt2S8gcgcUr/UIDwxHZQAOgSqSzwi+SP
Mg/QZodwyICSTExSf6hmcVCcQxtSXUT/XTBCa6q2sLKuRyWDAg5SERxhLbiMtrvi8qjvKy22LD9f
RbqG1Wga3a1OIFaMJIgqs6vLDLzIDbaxaFEmZ3M71UzGK7RpJ18+eOSWQZOcG6pR5JTpD/kpvu2N
voG/k7/MEN0EVbuxrcPYtgq+vAe18I6vM4dL25p023zpbAi1w1QdavphhwouI5yiCMQSj1AYSj1x
k8cbbSGYlTBi/2YEcTwwL9ALnirL4QFbk3jWLGGfUWW7yBXhhZMMCvxIrCAZQvJRLUnya2lrr3EG
fZm4h8g4GVx0eeqnkob42+WF8JRo9y+tYOyyKg/3SbA/y1qN5/bSzJqOrVNJuxidVHCrVB5BGmCY
ix2vLVPGYBfMK8HeZcfKdk9E3GTJi5NWzCdmZiUM/SEOvOsIy/Pnvi1FN9poPOSqX5hYAiOn+xz+
yPx/CjS4GjsnssA7dJcZD9iG14cq/AClaMGtACY1lOA75UWe0tIHrQIK5yf6/n/QlROP7xq6E8zE
SYlgByacuv50ICP3iQTRV0qfmYZ9su0yvOfKvEkGS+9uO+SVCNCxvaf9apRU6j0sevBhP6G1hVOE
/5zC+OzNWWG1GitECuqT2uo/V4Gf0qYAPus7iJbLWY3wFjopa8zeoqq4YbA2H+69FHxh4DrT36bc
mHqoEezoVOdzzWLrisE2CTqMjAu2vDV9HCqqT54qFzTiW6EJ2vvgJvOH7AN11lxFRkC+OEbrhB6s
Bho5+PvjByi74TPrHH9qAzekTpiS5UzYWMcULFB6+paLMYLv5RCYc0Amx3mQN+zRmghAJFHVE3yu
uyT24rgt205ClAOqAWTT1QiwRpfozwDsfu0wq58eI7sKt7R+LZXOSojFJ3xwGNvt537lwYFl5vfS
WckcWVIhDiuvA2BwXf8ZWK48hUM2o1ZXourZNHLAHKAHbLEHCr7HjRVPV931VYagKTlFWlvE6zeu
MYhgMM1CqWvApcWy5DCbJ5KyUflou9Nw1CbLyScRx4/b52zTTGddwRmYPVOMWoRVGs0stYzHzJ1+
Oq1UCdTWa2wWOW7z88QJ2Drey5/FhYVgNKDUcsUNToaOmo21Yzhsej5gLl5LFmX9wyTj66n2s9Ft
VRSNF0eOJmjUO6rPcpcpPjC7gffQmpvpXxLt9CNo8a83omRQ1FNPAMRuFvUis20rKS7i5DI+AAsA
OGc+aD3RjpdmMmO2QC3co0imQZSwZLMTr7eD75HXYPMp2fmUxRHtYNFwm49sfEoNRPo+lg/40Kpb
vC2glOwhWrAHW0tWO7UoVEy5/goBRhiS6M7tiCHefvPR5H9MSilBXnFZNn15znxTrLp0LrIJPuER
PeY4QmZ2Z8jZJIaGktJ8CWqRiOXmpZTfN2urK9t2Kvj3MJ9zAcY6J1watn898yFtf+fTYdhpGeNa
TMtBqQnHeRFux7O7FcV8tsqfubUvThF2N77ieSwSqEFNiCFr/mDkyRla/JzLdeFUQ1bVBJ+SRJ30
Mtuu6YGe6+wNNa/Lq5c9bdDhKNSruPGFVrj/ctEVD+44JnR9jWqbd/QNfDkV2cOIzOsSXS8UPDgs
37vTtbGXy02qhuw+S5c9QD6U9MoUX8XqhOSv6HNBkD0PoJdCf8Q1FLnZZ3S8A5xoxr08gKR9kaQ+
HbdGvp7AziOZodhSJ2H55snIWFes3neCU69PwIgTGg+WO73X4RlGPi7iYn79Wb56JwGGGtgKbDNx
jvUSeabnWvQVBBk5ip0FFjtx1iNHXiOp/11GX88zxnbhrFCOACkpMTzKkG64r+9wSZs/EnhPObdf
Q9G0m0tZCig67wN2HgNk2Ka4FFKmmehG5hf/e4uEYmREpDxs6X1T78fFQuTXyz2ALKGLdplTe2O+
Pe1RHr8rQXntAbczGfD84o+8QO6p2NsgCs/X5RaUDq6KqLCSLVf4Lk7+dIHsQG+toK42ath0Jtpj
ACa5v/6N9trpPneL9yAvXKKnRzcL6ceCYr8cY4NcawbinUi8+QOtuESNz0EMfSYZ2W4kwu3uFut4
2D3YySpp2oBrdqQBujZnokygu0WJZ1u66RFpazeBmuYfGr+mJddCB8sftCagwKvwyeVUJQFu43Yi
R4rUpyOgbNk+M0mxRb2IUZYnGAGV1k3vfnfRx59Se5huZQEyZfLZtr7qXnto+RgcF199g6d/j1hJ
gTCJkhTccVYKpHU00sdQ3gHJN7buG8SCY2pfRm2RwQiiXTAnBeF65ZDowLHobKV4EfWtBmKGCm29
th6At6DoJxjclICKWDMZQ9QYNL1h/A8vT8w8hWgWsXb+4GcHHCWUvdvMgDYqoaqWQsSQOeB2A5Cl
QWWB1/aVx19P2ykKIJDylNAcbExM8R2++OT4F/gCaN8rEH+w+/jcGcwrA01htPcpRLKcsljyL2vq
kxeUINciduqTRf+fQ5IFp0/kyd3Kqq16TcYfKA8vPZ4OEUt5zxESBPj0uvevdf8cr/SoCAkthtj2
5T5XduD3SSXrqiDjh4haVa2Qky/JeQCwY9VmE50Zw8wIkBtxWCvo65UDeSr2GmUIqE3XYC4iNQw4
KHoumhuFhW42fwAFTSAP+TzxAWotA1pF/m7hB9dsH2vvRrdTrqwSd5IAj7S30LVIJDMMAmN1sbku
mrrZA/P1mkF/wjwG7snwFiI1uZQg0gA+mv0I88JqhWbeXUkG2QoLmrruWYjVhFyVVJ+iTZM8yHMI
CrOUeYeEvzHfCRSO8jOFOP5zlnM7xNdcr9Vq81E8hXJ1btZjP0rQfqIJNetHVph09/vPZSeXrBHB
/tqFEmPW7wS8TjYNaL/WR0PbMTYnx81eA4R9UMtcaL4WpRdjzBwl+RZ1g5luRACor9aAzR2SUGMh
uVFTNLT1/R95zVmPAwf+stCk0UOa8uZ7EkKGv8SDffmAj78e1BT1ztKLtl+7enP/SXL1GelmKd8O
7YeHYnYTQ0BUN3qONJ0d/ea7DsbRLOGsun/9er61XjBvMblcnj7kBwAPZe9JsHCGguiZTtRXVe/r
vY8MGCItC3qeE4Wn3IJT9dxjwyPc7Vvg6ejm+k1e2IaUNvyJlCS9optRt61BR6zfoeMfdTMR+Hdf
0Yxsj+3H9a4BB52ZrNkhdCEm/zUAnNtfbO8klj3+IjjMN41DJoEjFxnnezrR5NkqZ5oIBOrGcJk7
2drCfgBtM7VLy1H+YLxRauiyxCzM2YiFzQnIhb7JrpfS4nfNHUANJzWuMZKsEO3ikb6BoTIbLKH7
vOjcfreghXH0zmky8MfsFthivoY1yY76ABVOrY2xcYQZ4OHlqSw1PRO6/zc6Rt3Orua8YbA5Y0BQ
SdalS+CSSxGb1XG8KTcC6Inm3qHrs9tiXTf3hp8G61IvlDpsSCNxyR77lb3eNNl3nQ7HMrcMmPpc
Kleid4iWGJkrjpsJ42bo3Is7DxxX1VUbKS+4jKrJM/g6T0Ou2Jv12MJ/aQTGBApe+xZmDCsl8fp6
yhFRW7ZqcLhO16b3q95X4SUnPQmVaWauAACctB4GY2GLwJu1m23yQYv+9AiKRZp18uf8+OssEB1z
UfnvPPBMVlyO7LqmS0jqV2LVYkVHHW91wFEhWrG5b3FeatJvP/tbeMU93ssfAPS697Z4KlWlPtiy
FXmE28JGq92fE+8JyjfDfc/8he+SK2yzaNzOWvJOucoGsdXXGf+sciW/A8lSIisPJ4VmT6t9zt1J
RwthqrwZQaMnpkgDAxHdHrs+XYnVVikPPo6D8ToYpFC3Zv7sKXLIGaAt/0nkWX0Shc9iVv3EArj7
v/0Ff/fkZF0RN4FmV0Pf69sY9LIggMSlIdtLPzcBqVWwAKy0QmT0uj8wEum6/MvTdmc6b8CAyrW/
BaYEhCjUUoClj8HsVD2x16HvwSeNCQC8cbnnBZKuK87W2tcL8jtpadPOeLklWCcwaR0ureejPKrV
JaeF67IQP/eLYm6o6Y3PDkOflC1s9mInYaG4ccbxXgst8l3mE+2WcaI8Tspm0zt4gZOP2YW09Lkw
XIlT4OWn/K3nDtts+kV9HMIPXwX8cpRgPyIqxeRqm1QVcUFAO8Z5YHnXDQeOA5mafsXaKptyIPVu
G/VVVQ51sptigP4WRC4CSzOcY4dZhbcNVFyJk7HeH4w1f9yvLZma4YoY8O6dKUUwWvu9ozV3lQ45
FIPQ9jMtlpzLrh7gTMU+23aafo17rkJVcJq0PWZIgD+PJmYX6WslmsDUJ30XFRGX4s9ZSfnFBj4a
lixTTffRXR/x1269Mur5+/gB6NmCw0Hy3ku2QF3YldxPpK+g+gpxWKTIihiLUXlxzTdfIwHxoBjH
uPCFdIWJ7h6cEv7sY8QA+ta+bI/iwwGGq9nO0osCPMn0/q2OxxBONUWYYXukKYDnTVZdz5sY9yB2
DGN7KwDueDOnwKkA91uLuW9n4N7CrhtgSmnofmOJEMci3WeCzd/fkaMhbDKnd5/dluJx53Ywh7l2
0fdqp3fj3ZCOw8nqsYHhnTWuv8YjCAtPwIEAWSIRNiTCiO3xHzmd9zzfJdx19nqoAlWPnvTIVlGg
HSiAgQcvZye1HaSVMj/PWBuIkRLyJEAbjFqZPqJlzVF9ZW2C4eT259HZE0+6X9HPMZoK6b0vHNrJ
5HfZsbMHHvo745DR105cYkfRgUodsHhnje3RysDrFeH8b29XwnHn+PDTFQG1GTLjrB5KBMi3Oyyq
47NVM7/UjHfsyUuQ4Zllj9qXhdMIAnHxiIRXiWvKYI81PWM2e7LYK+Pro4NkwqXlFx7sc27iVYkM
s8HuC9E1jayPqfGLU7WWxI7c8jM338IqEo/ccRpxM0NR17qk7dGFLaupX7md8c4pW5JoI1WbuTjQ
k1xWDfhS+uMfHhyVCrWQDHo+0oFcIVGYrHNmpKfuo4uGVPZ9ofwbUbi8J9jpzEZmx33jL9YooNuz
zvv7tzperbLVikLPQQhaEvV6RiV8X17zUpOn7JcEGYYq+IS4dWkmcNPlSD+9Rj49AvRf2d+stbaf
1Wp5tumURwIQQXKVDr5NnxrKerB0mwmiGDPXakW9oZkTfh3UAlOP+xnkRYRx7+V7+UOi022qrybb
rflFEz1nk7UwbP/XFxS0bpSclrJFvcHVdzlkzajDFS4r8oH/KVSnsahCUJ46kopdTUWaVencRfpH
8y/xzIiwS/z/JGirTIwcXPeRfxZvNOpqkeUUVAn663dODDD/QTNuF55sRSCQSdEcaMFzjM8J4GYj
TUbvJgRyfhOYcMcp0rg/UTnIliBpFqIbfmkDgzc5AP4v9jkqeAI9eJtM0dcyM5x7LZQuTmc4+GE3
ZSuOB+x//nwR7sLR+nBoqn00E54xwkophbfo/XpYrauidTMluifhDf4WvhIriBTRB1I0nExeJdrb
LYZ9x2RQMCHkRo3MhwBaEfejvc2SAPFTsLELf9y6R8A9kcmAihp1dG/U2tpCJNOYAfGU6pDG4BGF
aIGuMKpgpmAdjr1ra5O8gHMYj55BD4uTph77sN6lkLWNns+o00uUSHsLX0dlqebuuR0qbQr7/uF3
Z7Q6pL0K3745MX4rvPiDQIEZc6dEf2kBmkAMKqTxMXlnNYeIQj0dX1zByqG19D2P3YHax4L4a2oP
Qw43E8T5I8PuPDpa5o7uqgLALRIcfnRgStk6gA2KzipPzNji0YRL7aVTr0A761qQXQih+g9zWZkx
FWftgRU2vs3aaUS1iKWleC2/s4gCmg736vV8v8jYADr0xKDzafui9OKDKrnPSdcLvRdGeXVQHhfS
6VUuh5wo5UbAtwEV7X4BLx4RCyAjikVB0uYaDmMWCr6w+1M5B9Ilej3l3hqap8/svPCR0yu7Yq7l
WFiGEcgGUQ+vcyjtCAMUEo7T/25bR0zGVaHBz98+HXs27FZYzbPmvue1HkTg/YrsC7eBZDzpWE5i
uVizhE9Irow7jQumnkiEck6GExLqv/yO9NMgW/jTq4mPAkInuQRe7qDqiRiyunQ2Ig041HLdRevG
5PU8a/G1GqSn77SHQub4t0Tm/kReZx5ZqwMgKxN/x40pjQazu9pmG4VYFSxvnYj/mkqGRxt1Wcm3
Gxj7B0CmRMyZfQrov6rC+GYeHIGit0WWNmjjWaFxlRzeGrG47zlxnixI48xyHwe3wl6V37X5QC3I
y4vYRpDTYn6AVfZ3Wbosxl9Z+4QIcFttEqhs5dSzdjBEYc5autfPJE+yiLGYOLYDL6GXDBHkpAWP
sEVfITn11zQ/0z69Vm7dgPN9gTthlfpeRSKW3bRVS+FLgnHI9gUqbBuoTtaz2USu/voixz5BdCKC
jfmZd3gZFtBmxBqs8Zv2tfYFBhiiYV42xW1cSe7Ceru2wIfbUiM6YNAICqMvDENhtOp6JiBhsqpZ
Nz1yGyz8BS7elQL2Nja7in48DwUOPMAqvXOdU82tRaU/Ww6hJuWJ7nNGNgWvEW6ioc4wl2X0A+qp
ybN4fG3NIPjV/+lDEb6Oqg2veFaaUth6VuuZ/js9ewo8kpF3wjcBBFe8ZF+QCeTZDtTM5rXvyu/x
kYHisWaS4KTT1+FdYDZhK1Yw+GqrWxpD/eXr1YFPD7x2Ft6P1eudpMHdiDI+mVodXR2ZGWnfcVd8
Af5yOyxmiaYOgRZNJLUbNcGrncTwUzd1PIgjCtqMS03yfHiL6T+4zpWWVY2tlWhdiLioS+m57VrQ
P1XAT+Hxhd9vkWrJ1tpYS3khZuajlEs/JbIW1d49cSrFNh7olwAU+nNG+1AlhSv7uaptiON/Og+m
5i4910zC/52mTJUAV1HkTniJcBzhS9JLAIgx8ihqk9SVQ3OpwVSHhEvaNJLL3B0oJWQ7t9hWoRhH
0Ls9vr6+Sgg2/lmNPwNxTGgS+jSEkx98GPz5khbiifov5UoVrvpwqWmSrUWNULfRwMINuQCGYX6K
y8CSdveRwP/yW+osU57L42U3BtOu+Fvgoh8q/u0x2JQ02tS7F2GeNd0ILLUpMkGyXeBSeyg4tfF6
WHwbTSAqh6Uzfg0rhHLeOVp6zgXSr4Uz/pMYU82AZW8yiUs+B9+dKE9l/MP3xCBdo9ujK4wdQjIP
wmBOtkV3zf/TyW3WW5644bbMPpu2pHI79QxSC0yD7ubFBbyEbC6Q+yFzqEa0u+p0LjKKo8BfEaJq
BV+50A0WfIygwewJjYnje0gP+gGpwm9WUcB+FXsaeB7HzbB2+5fTT/iU8ZXRlLD/xhlmHaeE7ecN
l81uQo8F1lMx+/O40lGALfWWtgFH+7Adnyq0TYhnbe2PtJ8jLgXJY2vzD55Hp5LuC2+24XHusQ2S
q8p3XOxoSkhTJP4qyJNuJRs8ojBRNxZFHtIn+Lnv/W/yHkS4CuCNUXUM+SepcPI5UkunOOMYi/cC
QnhVecPYE7tOli2CovdqOoM3k6h8iESJiY8ZIJC96gt0V9+ECP48ZACdYrwUEu+KijZ7ZMpxlycZ
aSoYHKoXh7q/RNmjL2q0g4bZZCQluxZdPP0iq22S+DZ8AwwhzE11laKDMUs/DuSXytSUBqI6zh08
m5ESa7V9hCKP/gqO5u3MUroeQRmW2zalhHrYkeh+z5NrWCh0T+6Y7GN1MsJXM1D4fgugGG3QGBSy
weeQKmL+BnN7SLlgPWn69oZ18bT14XTCaVQaEpTKWHCVUIS0ijFoSt/elBUcdIo3/ORbYMfpHLZ/
lw0DbMUk9FIjlPrIpXyVFAkeQLgpmVrZWPW/vLxISfR+LAbuuxXMpmq5WkbhztCL/6nxfEQ7bR3L
MmarX+SQ/auJty9ZSgQaPBQO3EYWIChIv6JrkEfE2zDIhQg7sLFroVKgRwWC8/tzUW/NNNsMs6BW
xW5X3jthym9MSrbO9M41nmzLDG7oGnSV7IcN0HvSyzs=
`protect end_protected
