../../controller/src/common/ControllerTypes.bsv