`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xjg8AV2JA2PlExLYsEd/svxeepWxmGsIVTUMyH/IxBun0XWM39gyApD5yi1906KDnEq1TuRNPCA0
/pxmOHTc+A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H0aFelE647AZKiRMrUGit4KAcCc50nhHxkL4BRx2khsBUOv/3FSS8COchZbEIAFBTfDmofRV3q6h
FsH/L4SNnRkWm1IGniu+BQIZn/c+k6+zebupL9lSX98V4H8DVymZcL2mKB3nDNaLEsmokQl/Nm8T
J8/1CtUNmMacgsMCQJM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y0Yq2g1/K7T95gZF82spoGVZH2L72fYmSmEyVF0bY3P4bdPc/KQ017vF4NICNOftsUIpbxbXu8bM
yW2ODHkTxiJUXAVA9RVIgv88EfazVf/q2bNav0BQW1F1Ut5fXpYTrCGZPjAD02We5a66LcSw/BOu
zk1dPpFwNTM75bu6nrSVwQ8IkJHZY1DBsfpTVl4YBCc7DoNy3ytR8ojyR2TinqX1t50PVSYb9Xel
9tcwQZsCIftqNADlRLDLW2oxG3OtLOrSn14mQdlQmIsLVd7c1ZuWFroITfX0AKozIXQkM0vEex4u
fMuZwcV3uY+BeL8WPdwKiWfcPCKFffxCNI4Zcw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KKm7ZuMwo8vHaPNflK1A96zuX2no33mKGdNppXhDt/Whf+z5ks1/K77paMzb7H5K0jaTB9OGTJpc
kf4ZEBXkND9FbV4rod38K7u5J9hvaygWB5mh8Sqr9hHik7+ahL9Q4RQ255rtdMtEn0u+h9HL/BDH
cSGhLPdFy9DV7fCVeFs=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XMZ3rEIcTIo/wmgIIVya7XMD9piySienTVIDJWWmPbN6ap2aKCRg1rI2rPtu6i0ICcveQkhhd+tp
qv3gUWWcg60HdoMn2BvoWlMpjQcTYeF/7Iye5Fe2sM7PVY9+ce/M3lCJ/Jkeuuh8LA4DIH2JBVu3
/IipUqRxt2kaKaKG36dp6W5W8yNieMsfNeOR4Pk5p+c4qJdUzq3/cIIcXV59vxBAGcf8NZAvT88P
KRjWuO0+jFdTBonjZZystspBkw14yw/z6xr2gBgLb++d878qqymqzwu3L/c28Vcezc4rqhNZlwcS
fKeTDgqBZ9cfB0j0LtMo1Vyj3GINSPyqLXxDsw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 998320)
`protect data_block
kqVgxRhwMsp9NNMVKoiFVVtSoW91wDXuheqsTM/WJaijQykA2SPJTdTjCDSLDTwTlODd/N98lAAD
6fwkipS4A051pMXHj2z+9uEIZ69kWW0GppjC3TQGgNHUbgTFf3CT9MQ4+8oFLN35Ng0IsFm9Srro
rF66PYO3w6j0TMX0s2cz2ZyV7qJEp1f0eWT2tFUSZJF7qCEHrjMo44JECm/uL3QDuXiwbG7hE/B0
MkHn2MKcLXfZnRCLmKPHbePjf/PR1L6qWUWGg3dtZmPXCWLZSt9S2vEsyF+Bw17ottX/HMv7VPPT
EWsgntYVpiHvri5K/LWHxN9ie4z4cInEGmIFiZMymvkulzyneP0t75VErFuz1hEGMUNjWzVlS4Lv
4e1/3EL0SKUI0qRreu7L3OAYsprRDjxVptkYYZqf0EKPtcOHXgcpS7sgURy/NfCUo31c5qK2sY5O
8oMqEDJ7yt1dz+kp5JmW3m3pT1XMxTFmlpQ7BLKXOCMQzsSVVK3nP5gSuY+m5jFXWbMn6W8RozWk
jc1P2aQ13EjrN4RpEOuBErRQPNV17SJ2AP9Kmzqr6/qM4XwjDWGF+NoVk4ww1x7NwkwUVnJqddLg
XYH+sc9+XPJmfktmTov5H2rStjH6kV6scoMCcWjxArzSCAqMslfYozwX0zh/fDHLSr1Z9z8YPSl9
LWtQ2HlhZ64a6w5jiGCM0ETF6TvTOY8d+SNkAjBl73IYg2LQ2FzMIVtM3HuM2Zn1ZPcNpeI/8/0o
mqBc8JmVZqRoJoScL0iJqM3b3bol4Cz3bsT93GQG90qssLPjPcw8ad0Towe8r96mgWV7KqUOMeOd
Yraq7Qk62GCClR9SwtKxDcFdo1g3KIqiBz0SwW9xBvwHPrFBZwp6UpQgMjYjqnofrqjfdbM5m6D1
Lo7Le4r+vEMrzI+XbSfOkvTilDGauNPRVvl1Dd3dT+hxvXIEMpatDV1oKpPWXhfqFO8TpNjEDtEU
q2NMiLBva8lQGtIZZ6YQEYzbFAZ59ZQC6aI7C9aeTbVuOYhqFGWp9NZUzpjt1hmb29oQuQoLwxIC
xij5dw3q1DLbXkPIspuPX+qUoET3xcuL9842NkC9H7CqZ5SP+ubcwIjZEsSUQE+X3I5kDa7I83qr
m1qhUgO4lSwzdESavyJKn5zGLeBAY/M1vmWEkT7cqJ+xzriSYPTUdmMMBHz0JkGzeHKea8xb+QWa
mm88X1KyB57Di+xc8GPr3eYKypj2zM4X5dli0le2bLHGZ+5v/cnHidheTO9KSa3sRkibmIbjFZoO
Gj0ej6hJDum68WE1j5Q/GJ1TTeXpwbmylsyXmpC7CGMJBFFGChPY5/zJyjFnCV5u2hrT5kJ6ba+G
/I8D19HoJS9SG3ZqaBi+lzST1iqhp/J44FxVayIG5YMGhItnSnG0VKaS93Sm1PKAQvHwSCdOU3bZ
g9L9DucFHI+5m7gsmHiDxczK1kNaxkqs3lTXBYCdjscg1g8lStD2zdqGgcwk+OAjc8+x17/C5wXO
aiQSAwKlg1VhSdUD7AspNnhgW5UKr+TO3IM04rpZQAp6vknwUx34M7cI8gU/Vy1sPUeaCyf9hBHL
o57+KdTmXNv/0jwCQTrUZsXmccDbgnI53G+PqJYwgBWINWKaZj3rixUt3V+0k/U73P7XY64QmkjR
zFfD/iU0DEtII8OE5IDjTqBvy3ndGnrDi16DfoZpgpjDNQJMIsj7c64z8mKLJuV3TTqgyD7fmEKa
ksn6uLKuga52ErZHLWfivOqgqaDLb9UAMQJvRs5jM5/Nxqp67IWGwfw5pl8e7qNzpOFjQW0bKLjw
Lht3hWjyCl87a5eYEVke484rLD4NFNEK2AornEsg7GAvZk+qHSPehWkXTg37OVgUDLsfTiekn6xN
+rNKw6OrZc1mFwwitrpmA2IQoUytpgWhwZu1BqCWXef5PT+e5pAmsw2QsSQQjpfFlLqtPYn8At7O
coI/q0ed7tgYniajBg5yNOhu2qR1kdoAODcz+0doBXIGsDsAF4fxJi0bPeG+Ah4vAQGA3cZzLvyQ
UqrjXMUeR04bdpleUhvmSKf0gGjuVDUyIDtQc2OTZNl9WVQGOHsWMQmbpmnHrlPESgqJST+CWTBP
jeufm1qxAbd56Q6rQzLCmi2fnihXpLUriUr1sdOVxHkv+nyMhhimhaSNaMQN+pH/bAgurObPy+60
c5YfxryZoZaffFr79MXG4oVwu7DVkHB2BGdEnMSfeLTKvrlLC1SXEvLOjXgJiVuD17hyUBs3N8Wm
WQjSDlijjptDXksCi67AUsQVwRqdzyLQyPkF2pPwhUNOwKIKs8xlXpDE8QZ64PLX6HK/vki5T3iy
prDp1yeOWxz8YS2FBRzK/AJ5ywvyUtNu6GID8aCes4RQUuUwI3WjTzm/MUqOTSnyy3sitJE5jg26
36yNx5QkC0ODCOwnlvqZe69U7RYJUuh45JTQ+ttksuzD1hNGA2BZSl3ZB6+hUxj96i+sGpVHkwoD
SqF4IKpCAt/9fG5X0L5Oi5dYInYSYQQi3G7VYp1ZEIKvs1rMikhlY5RIagG4NBNCPP5h3jKCWpXd
EPfpM7i1BHJDo5lkpP7gdyidKflSEbndLgfOkSPUe8uwb/EWGQWZdnouGE/no15NLP46/l700XXk
hv1ceERrqOhW5pDUgGn/LQt/DwRr8Xa3AldEuSgDyiIuqm866P1MdTChz/ltJIhRZHqcN2RIyobv
Jv6jwoLaa0wUpT+vNAv+Ye0qba1p4TKJFMKS47DP3BOV0DdcgiAIzVevt2CIb9YvIvQ3lF3H5wFR
T6C3D1JezYibo9VO+ncB22R4xZnEAfP+SbkhN26jJ90vA3LdBC9oY7pmcq1holo7VSlom0j85kN+
yH1ooJwflpxW6mADUApnqdEbOq6cKxaGdQlQNvibfJP7i0MLOljnAC5UxrY76dQmTz2lo5jHGvQ4
Xm1Atr9J85oMRvUA6+33kJHdH1KvVP99OCB1YJQo2su6sh/7RqcT8Co9qIrnGkgacUghxduFWeTI
JKqIwdyBkhCtPNeIX6ETXrjX+0nCE8v26fcZWjqcDFywI5L7Ip0BBa1eGQqlAT5ndnYmclynaUQD
XBPND7YUGR6ZVghrOK89RtOvymGajFYsuGpY9xoGbH/ZS9L0ivdjsUUyhq3bZaBJOn2QKyPqzPfk
+eCyddA3cC61f5FKCBCfBD8cP4Ud8sS/y8LwAuIeiPfhZ7yv9+bCQhYByOBfgVI2oI97+Enk7/zS
aJBk2fbCGsZzrNYPoXpDuz7oKl3TRO9oJFyaUN9isuNDvlZoZcl84/6yBuR0HDNf3CCIXwJlsvmQ
SdtK+ev+puV3Iw5DWDN6yhgwMzrmiPvAu0CuSRKGEVMxJR+Ss6ZG+0haHINgAjQLYwEPSk9O4/61
zH4VYTGxnpIkC1kC6xbM7j4E4C4CQrZyOvCOZyTBDRNQvquwMn445FL45H9uB/49wVZzTKAQsgkZ
BxfiXuEaVJTntnADNZ+hSydi+6D3J8OMQdMNSf3fQ4TeiScXJESXTqBg/R7LdRFKhcFFz8Wm/dkm
ENky7MAPVLas/m7H5mZHAH9jxJRR0Bf7/pvZ4xqymr5edodN90a+CnVHSF4iMPDqUrhqunf7FIUC
teVqVOz5XJCO5JHy9bgbzUgrm1Nj7HeezQsxf4OJwL0heQOrhOtpsdWsZgDvjKO3EfoYx/0mw2As
7wLdeT9wAaJsxR9iATjyKdg2j/YVFnPvgm+rxOByefyoRLycC2Ku3PKnFkBKFQTC4RLUv/Sp6YlI
PQdX3lHogxB1X6wigMe90x0AEyl41yuzdQZVIey2ubhYrRN9s0bSHybSqdyRdPfoWtC2KLJK9HnR
Yc6DcPPwEbmAl43KgoK8B1JNzOTep42IbOnY4k4NN64hixB4s/zRYkWp8h7UeQEE+l4RvZ9e2YXL
bi9IezxmM9OaK8vmW7tsNrQ+vVCCT/aqIsLDdMua9Qn11zRJCPTzNGZ3G23htLagPW8uEQJ7sLl1
7rkGRHQjzg1963wfJT0WWN+1vUcBoo+4RJY5MSZC1BxXCIRJKJP9GWVt7oldQFz/MDsykyH8IVDw
ozaqS05N2R0EkaPnY4SOjjovoMgJ5DIcYqYs6yszvCIUZtHfsEhaGyAMKBH0lG46hHoguVKQ9dYN
2WYrsfTsZr+MXqo0g39rdiBCYWbSODTrOW8dPF4FtyIDNfFVHGToMGn8yZWeDyuSSQHh6A91sVcv
nvvvguE4DWFARuvSx82vjK/xih0MmGTsLhjVJ1z986nF7h3LKtP/iYAI2DMQ857kFuxQ0g+sSKCJ
opCQJKHOiv2l7iDLO2ff7GOGYeO8d61jP3kvBUOUZGNWSnE1/sC3UMeN9CsiAwUg+SpMKNmk1QsF
DkHLo50JQZPknzhA3m4d/ykXBK97z/v2KuARPn1ONBRupx8HyVGmogDeqpwdpJIu0pVRmxDVyTxS
zkmbmZiyC0McJ9j5wSg1fSOR7EQ1ce6wf3Tw7jmUaMRrFM32htJJ1EjzZEW75HBDmNLXxU/Nilyc
/PUeQgGWxsQxzZubhcZ2fqWwJsrSSc4jz75/3h0x7f0hkvbgsJJBDDWc2gm5quNl42vQtqBrsgSe
mKxvgA9fVjX11KSxcvjQ3+gq/UF84Mr5klYlGB96iMigyE7bpF2VTyZJYbvjcsQ03iw5qSdg2slj
HW0GpVCSqWKEiNETai1Di4pD3vxEJKWxF7MqAmwKpGpWDMFPSUWn0akLOPSB21YLamc6xuM3kGGS
1DZOxFxzzUG2K/mD3eJBi/PZJCSj2QLr+JtKjBFy77XoHX3SvlhVEV4AipyK5myelAGY1NuK7tBp
lDoIkK7CQ8XVB2EYDXVTmeRjk9NhvTADJ6k5NOlSsaMKqkgGqMordGvWnLXyuCMtGmSnKETolBUD
inDYN1wMsfKyBmo6igGy6Kxxyu5ZFQQLE0pKXGcuAJmJqt4On2NozR1Hycah6Et93JxqBQFldHSo
2xcPDkJPlaREakwXQprlw+Xms5c0QTE/ppJv14WhcAslmNoWEUNuDFzJEjhWdwOtjc49Cm+JhtCk
9qfSYzXo2fDGVMxYlhGX7NK7uiVVHg0sdgHD6zhhIoeNfCB/YNPtYbsKCVJpwhXwX31zo2NK7/6f
aWtjhc7u+N/lqceysK8EP7cJWz3myp79np27W55YaYDIFC5TXGRI4dAssG/MDrkR16wkdcZ7bSY/
jUZP7kKVXLhX9ksB7zT+derhVggGOSIKD2+K6rQcOZkcTr/REtfbYqG17/U6e9pbMUnDllrwQHBk
/gkm/wZhFqsDhniVJHNQQu4w9Eg4YRAsp5nymqLNmK/TstJceYyR7htElcDhXkfrtIr6aGaPhHGw
MtLP6vcfb0LNq6jPv0eUR/UHLpDiqe9YRkXeBGqqar0ctxYEL/FVx9Rjy6X3wPDQGBZJ6T1MzKjr
L+A0q6np1vT5e5Nkcwty88El8DswUrspnj3O3ntAHb/Y0TmPxBOPFR1Vh9qTHDUAbZV8VV9DfGrt
GITgCfm2489g6eutel52v/4ywi8zwgxlxmX7NMe46Fs9M7WK5Yab6+/LeYeL7nS2gqQ3s27M8iiL
xEuSluiLBjBPm4jBIni4JQVv72gz4se+T9pww/JDHg4U1AnK6B/dyurTArq1xe9+VudP98GRnuNQ
CG5TJKhWB9VpbnXqIJBCtAxwZ316C70zjcId1j3RT93sgq9P+JCH1gR/AzQYu2L5mduLShWCt33I
74L+2pzVjnLZWW1buFIhExP+sSk6/aUc8xpA2B4LMmjtUE35sIUcalhayFPm9hHCtHbrloKyc+F+
qGkgUG0YZ7nxXK6QiQEPkkAQUP3xKmRFtpEQlxe4SS2BTjtfCNJyA3XHoy1F/LAb4nJHd0/rEJ7S
w/ZuqvtM9K9+eeGe+R6S7QhkmojqFFjnTMKNcL7PlmJdYDncYEVtWYYhZ5kjY6dEN1NjajzoIGbL
yFEDUgu3ALNIOFSoYcdGyg8eMbNMYBE2yyx07ySopt1gM/Hr1TFdARsL51WJZUlxGZwgbFYdGZzR
OsrqSxxy4yaEeaE53psTC6jLUQAxR7RtZqTtsJl16YBVMF/w7q66nSD3JgXlmgjZUq4By4Y0jOIg
LMzqlM+tYYrZKaSoTpjqSjqs1PEQ3sHpoVtpd51uDPzM1WYV/pU63+/bqw0ll1Ym1XquVT+Rxhs6
KZz+CF6aCAIRoTW4PxWEElF+SPDRhC5ILKIEigWmnb6kVHM/Ag6CuMY2YPJGpZv8dkWPNeQ52gko
IH9h9s10sI4mE5mYRUuA+yWBM7R70l/3hqeo042tgshoER+GYjTegaxluQ9zpAF9QnDHS9mG1Y86
oechpgiSKJK/RTCN4GVOPhQ0FCfTSBe7cDlr+poDurRAYbGdcl3VKejPV/I7I0nzLDkzTtEP1/pG
Yu6UCjFQqgHgjXwOUAI9Nn6+aSULRf5riBJTFPfcwSUPIRDfh+mqqixv3FgcNVLwwYu2sl6pQ/u7
b0OVVrwtXHELhPCXwDiNqBMI3X/3DFaTaq0oHBlczd/k/tS+CjG9vBO8l1rYRS7JA0+CCJGFd9i0
TqoNalyVPjGkFzbfB04PWkqF0naDCVW6B1c7Qs9UY1l7sfJiPOXizRuv9XaXY5qjF89ioaAtVLhb
ug/mdKg+CMTJ1o4DAlGVItMlbdzXygQgEnwJcRGKRTAT8YJ54uqtCYA8SprnVhArh1cON0NwYjwY
kE+cAp7OPz0nQ1zuIgQDBKL5fZ/DCRB2uDgtSQjhbWG/P6Dci6ylBHP4RioMXQ4K6rQmYp3SSxD5
UagJ6g0C41BFoC19Jj5ZYEBPbLrEau+Ay5SyXv+vtX9eLf72eaNYvp1JXIQjP56d1fDC3bZ4gpnU
j0ZGmCtETjJ19khlmuCEZRwBGxDiOxYqYwjc6zTqUrXDEbnDWIEs1ckU3K4Fg+gPRADJlNp2Xh5e
hXR6QOLynQNVv+UqUGni/IUD3khSTdQt+WN/10ww82rl6liUhh1XMbI5kmjR2mx5HrRwXzyRcZwZ
fgScFZLrjERsifpsNNVJ/hJK4qMqAVCjTpA8x0X5UrqjGdlGs0zjDgHRb6jxuIt1LxWquU91jpGY
a+o1OWcURNbZxekaN+aivPupxnrXsRYvFHDPtzpiS229PM3jb4NbGkdqIpUsqeweFL1F2pnarXMi
c12PbikPg90iA1u13QBfQbQhLSdw/A5nahexZqgfZddpHuU3jv6C6M4EDGYD2MvorsPkSqe8ESaB
tLwiDOFcsAFgWPAXnFYykPNAOpJDjXSKLyRp83wPrbiIN8aCYF+lYM9jZAZqszkUfrGJWRRBEuwn
CguH6cgAk7hOfBEBcBVj+wL+/xy29j/NYZORsOXZaF39oTAdr7odsOMsh9gnj2JaZlWGmF556Z5i
7GsyiRUOMdDMs6u7qvi1Dl9U0sdIBjWceo+sy+BW1uFvv7KAGnGUePjYlQ3lvV4niDTIhj/Ws7vN
sKdb5C+W2oOciPP9EpIJO4XExvu/edwVexuHHLlDHsqBJvQGEu9QOs4hTIMb48+CjmV0fwWCTFF7
90m1ChR4RsIlfGC6FDgI5GKbHhHdOgPus0IIWxKw9eVQN6aaUSKjdJVUonIa+6/Vfp83kNe4Dkxq
3K55fSSm4dufrlpR9XXoLXbz0hpOMr9jlPdYHONLO5G9cCny006PswQn3idTIksxpbLwyHMRFCE1
4kdu0OqFbUiSc2nfaalqVQ7SExxFhUyRVPHnR99r91SZE/iumgZE6d4DhYds2J8AmMWmQ0rG6hLU
PAqKWl1NbTt731K/fOpL0TLEVYuBYqkP4danyF7j/fuYVp5wRd+ZFBa5jtBY+aStOH+EVrVLOvgh
xEN8uRRCZ7UhqypQFML/zoxYZDa8lLc1j0nhkMwbq+Txw+S15G1qeUvEBWk9m2VoPPqWklU5hXQE
9/XLJlCNg2gTz8N0lJklzrbJ5pw2vSYK07qZjyt+yfkpTy70N4o0fKEH9NEUyOTHjwRl9CHBYKSg
qpRWSLomlVGwVz8ncTB8lB81c2SAT9l5SaE9grKqP1WWIMIrdquFZqhv2BfKw0mtP3UqPatJ88cs
ZYdxEbSuyB1Rrj8A/ROi05nJ3FCzinG03r63khKE+I+8iiZizl26rFhj9l/bwPvKPSLm6VIEFM+o
G6dd1kAnuZ3sFQZGOfQjMHI4YWp9pJAiKYnlX5NjZ1S3Vi8Fuef2Ui0OjQ1LLB/4GEa48f3gfiGA
jOxJC0G6tOp4wicifs3F7K8MgRU9Hb1UYQMvu1q4HyvBFgpRUsoR7UKEL08UFJVniKpgvzBA8isy
w/1QGN/GtGyosaC49uxxieuolYLpQQzEd1rIQC+bfR3CpiQxpESm3oPcA9QOIbHnnoM3y1jqNliH
CgHWezl9arE1hdkiDPwV92wlnuwfslLaLMuNXJXboPYFalzxhdgvNw+VdYf3nfSBGWWQ1KLEeXGW
iHI4ahViY+kU8/QAc00PbW3Kv378hlnray64JNnBa3ko1iB5kxVYblZWu573uUmxv2bS/wso5Dh4
x3dvN6pv3Ha25t1reIyufBH2E+gqlb55aPVwTDOmufcE1Htbv6VWbYBe7owuk2CisUHqzvY8ujsE
IE8PqgnZVpFvpg8cSWXk2tXmFtjbPC+LS6wBlyjJOZdeJmB26G2JOapCkZaVd5UFmSNHto1kAAaT
ifAHuBErEOdii58SqHez8+9li47MsiwaCo1p6L4rZQkHy890aYYMX4ABD7YmJWuQ2FuIrRwofKa0
YX2unHgb2hcRzYcaumf67aGZmwH2SkW/Siupoffu1rfiyqF6IrutJ9wvEVJ6AmLsgzhTXJsGhJug
fqc61E+ZiCdPzWI2aI0LDG9Up8NtfGjvnGfqDlUtz6dJFtgddm7E3O4BxSPnvYJz4iMgMRxRedcd
TeVEFq8vuskMFh3mogpJhvveajPSolrFcHAmO9TWpSM9pdItRb7w7Q78B66xJ3Al4v6Qj2dd8OP9
jzCS7aLWZfVPXAIPJo/gD5oTtDUBMd42lBB/mVPr1IVcLCW/LPofxnSIJsVvGu/9HiqmxFBhjwou
O6JJQSYFQu4u+Se7qGMxzVxQdJtWyMyVG2sOnMnQleSdchMJJRsxr+5cSLIyhgvRUuzXhg7BgMaN
OsHIJekv/pYdo47w85ED68ztG+GCLlxIMTqn7JxOcljVRoxVhRPSWKrnlPbnBez0NkHWyoJO4J5j
4Hk9uLMd/DOyXBXVSLAjM5SD8o4yp5Dt8hW2TPpKGEMa2YiZ5Sy6WSpQgtwm32hXRhRBTlK44E7j
NT8IJQP7V3Q43S+0yM+mnfxnKySdtbLU7vf+rukjpHDdejWAtJvazSMg9NN1uM4nvk3T2dZBJV1+
kBXwvk35fAnukeKw1uhEgHkE+or5SahnAazvdk5TK2uzCLtdx+AgppmZWDFfhzqdxeaKVV1NqU1P
T3kt/97fvNOqtI77GZ3AStI0HNoLiz93dhwI+DYMSFRwLjf9dmOS6Ggwv+zkSMbh1RHKPWqffxmF
e4y3xY6GHXVuJ7gsiK9YGTBQfLskABh0jl+/EP9vAbtbH8ZrJWF+yQixUNaXfZsAqFc3zpK0RVdf
SaoBr0Mpl8yaEI+vZwlzsUNHxmue2r8mI+Ndhz38Hq0RcRhSwzxHCg007ht0ofAx+C6GQ2swIZkb
fPAzC2m6VLltiWpgtN7SfrvxzXnfQXpd0cHH7iU0pv+u+2xbl/z6aNdEreg18ZJw6sb+MstTOlpV
29dRFqH4NO2XsgjqaAzsLxFCAdFnfP+fiBxCw/auvKdnlvS+wzt3ZSRGYcuimVkOVJESMftw7rgG
a6uhlvs8PPqGCHTlno97nmvsGRHqgS7/qycn8N5FOszYvmFrH2asIcevk3S1Fz491dyphvI57D4H
QlDJ071vwAgdmAO7yqggTlxCjgApkas1jfSlyNk889yRoPHYwD4HXNK8WqR/p3MNQSWVL5lV+h0o
RRcY7XVSbgRgiz+Y13bqHwjL82Q6tlVqoNVg1WkVejf8DhGM8ChgakjLQ1jwFWq9PE4bSh8YmbTM
/kiVJOkKsGmPYYNeyeCmprfokCQXqOY0/nEBT2b+tPz2G9TjinCjOZjen0LhWMMGGuiQgR+o0BuQ
ulOJIxqw5k0+kV2M0UVJOlSMgGWOOR0LsB1nrK5XFMj7bSIILhyy8L/BJavv4029GdAOfVCzH7lJ
a2GCPNyxpb35YJB7c3SSYxoVtBvy85IQxM9RWZl6JRnyNWpg0OJbYiAztC/GOwWomVYs/USnwerh
7GwFxAbidjjPqQbdKj52wk5ZC/22Oc8w7oM6JeIPM3VScj+paJofMpDNHrhKBFF+7OXnMNGPvKWE
V0FLMqsMINPltFFl0axh/1jKaQe/jCRN/zxQw/qBvjwMMx80Jhz6Znau8QetARR4AypWNE3mM4Jg
+o/FK7n+yMEIDYHUJWEcMcnrjAfhtHKAM2eLvPIX4XkAZteU792mxKpLr94n1xZecVjTcM909Xfd
jn/2j2G0Vt5cDuuRpREn9+OFa8PAg0zcy6gW4fmgDyYWSDNiI0YxYZIfqKZfBQ+pTaKMRdaXPPDi
QyUpPXt1xpQT2PByMcPLZQRzt7bfIg26MRz7hcJtYC/dFFWtKo6pCucEfyb5d5FQ8VB7Mf4RN7S6
Kqn5S8ybTJDbCVV1jV4p0KUyNgi1/yb/hugftI/XIfNksKlHm5tr0PN85xEp8sZ+pi/MDoCNZ9g+
R3Ks63vziIXO52bh+RjfJnCp0EMsnikZGJgwdHaw80slM9hO3VifRY4FC3fiWa7U9OZYXNxsiHaw
awGOw/hulEI2ylWIt6iOoi69v5+jtUJWe8czSaVo0fREKZRlG25wMsgrpsY1V1Po8zr9ZxK2iQ46
JUu024PfMuVZ0b7Zdeid5QCKtJL/W4OxXHPLel4lGHL+k7d+Tacvk4QCjWdLH4k3UTqY669sWF/X
cfinZGAGYaSZuMrZ0LZrNbocBMkFZm1clPxLQ4oj8Ru+qGaG7HhwPPFQKVJ1O8vHUwfIbDJRXq8j
G5jE/Km+n2kNOKPZtMVFCm+VcAUIzVrePnReW0quXTpSITq07oTrYR2ASykGVlgjEHaLUdrfSaU9
FGwKgyrC6uKVUT0AoSouM/nQdDf+OPkBMnEZc1wmily9iJzio+82bvKBG+GnuN1wJvEcJnemA0et
qfaTl6XoOPN62XU2KmvWYXPv47KXGi/1w5qtypUD6IIa/Rk5ETc7uDF6yWiI/EhoUYNXJZxiyQxH
DMyLl3yRgH16WoO+nFhoP7gAu47ieg6ITnpJeODP7lz0GtlXxoRo17URjV8bHn5LlHogbPKQdaOI
rDOYHQLBc2v5x/vgiAwp6Qsa8CJVNL0oeiAv0LGaRWopUV3QxVHYzhUyQqKsTAOawII4LldGx9CK
TypGg/uPWRiVSTBBuYJtPm4fXb4ZY+5IuALu+pnDliBTdgEtxLCiaL+fVNzK8zbOA+Xi4Ix0bvrK
tBFfIN6mIdMmOMaJVOf6YHq9J+coD9RDwYilYJlqLdvV1Kyy5FPHXz0M4nc4D+NYoNzM41mziDpU
j5Urb92WKbexbb8zlmR+UbhIlxE0Kk1LcL50Z0iO8suxlhyhPhwXe9OTkkPDcReOYQIrGTp3THjO
rHMHb4iPrVaHlQvZuyEzVk8CauWUU3t9bDPtj80cnuU1EnBzQsaKQ3wU9wBKTiVxlW6yPQ2YFKj7
Pu6d8hH/ngG4xegvGqDlY65OFqKtJBRsGPUE4u4I9MYyydW87bHexQHNOO31Ah8D/1aiJuoNLUb9
oOSwzohL9R83kflPSrIUWt6Wh4iwL6YAgqQQlzm1UYKodienRJT0rWPzVN4Rj7yHRq3H2OZYooEV
BhHFx8qu7PrnzR+zbJYvLY/OgSlVhodktqW9a4GLmvIYrdox/DvCpITE0LMrimbB7N8ogdZdX9cz
EwmFSLLbIF/TraQHLP0id2AwbyzFuRiZzT96DK9eINRalvLqWBLCZ0yWuO3gQ1aK5aWU/yXgzngW
ig3l9YjIDKQc+z7AV/Mb1DLKGwLiSEHILSGWgWdJwZjjT4N9qV5GBgk9SUImj01L71YLagl/j3tB
idALCUNzmb8lSHVkM2Aw2f1QLhLEDyoIga3nY1zzPsuH7dgybfhgHh0ewZv3VVyteJJi6R7phbxc
8yMZ46YMUnFRQ1NC7boAvt1ouy0zDDScyb7wsVg9m/volMhnFg1JyXwABEnM6HWs7hZFuKwi+j+2
a7It43ZzGVCSD63MZlI7YZ1q8148cbmxysD4yC/QByg0gqif7BRUe1ThwnxpfXP7mut9uklMRoll
zVS744RQDUESvVvsWml0hNMuk0wjFWGI/u1RZGrvl/ErSGGadPyegmtbzRdD3v45z4aXjaZQDw2w
k59QSYvdcQY3Dg2BBH9fTtU5r3/iz5Dz+zzVhDhHMePPKue3m6qnTG/ttYfeO2cyHBaUVLpAIrKE
H7dReQIL0NQD13Xq2whon5q2M0siJeXf9eDnDAtbPzyDamoigZe+cV5pTQGbJeP73hRHDDNabBDx
fdPJJG2qybvZxwqvmHWTQRmirXtz+HvAUyBNuzgDGxi4q50TpUX4nYZPsHFn4sl1DNiL0iYp3Oin
OEcVw2gkibOXkZWgnd91GEfWYCZQchlXDSBe1TUNNoARrED04AWTNGfCXy/8dUxXdqt2SvxYIID5
YKkKcrekvDWuZEwBbJ31HdNxQQWVKA/xfZK5jGdfgGyySv3H942ZNXJGKAKM8TVAkdrQNJZ/OakH
IEK4vwDFYRzoOy2/73JVc92XXbkn7yQkrRE4a5zCfjIRhnuTnk0AsjV8VB0YWpraSX9fbOFnyodA
Pi8CjChXIE8uqIgv8EoEYL4YG0VWXJwUx/dNY2RZN7Lmg0rfciEnz5UO/Xr5ISk0mmDU2gUwU6wR
5/bKQKLiyiVGtPWkj5hIeTCqATpa0u1iOHuHOrDos1fpTwtiiIPymnUxQ89dLUQ8u/Do5D1aiJCz
HfddN+NgG30nc74tU4NLagD8GHEoGBZQ+OHHU4i2Buny+My09xGtqITyV+yQMnjON9aeIRKhtTB8
qBPpKgpH0vgGVJ0M1WrnQshh27ByEh90Ojg8ygzgqI82Kw72yChkdLdJ8X6V4Ve/lN63J/6I9bmR
02LgCeVCyJX8gMklHo7Q3Lr0HnBM9rTIgOtKnZfzihIqiBvxofnX/PbEHKQ8mbEtnjW2xFLmSQUB
Sj+Bp2aoN2NYpt8WPz9hZx2O0uGuWlEf/6xGqtotiY4XZ/82/3BUK+T32lcCYOkCP6QdOZ1hhAIx
65wAHyIa4GFhaT7vQD1Sez6uK2EI3tFd+pEYz5JwPLLgdpbp+8m2wRvz7SMWX1Yap2NkrmKNro6B
GHBWgLRJ+UsG3vRUpwrAisSm0FDcx1jAzRvJ1LLifEa9c5fHI4X32GOp1Y5B3WU6V12DwI3l1YGY
PMJGcqDjotmv9WtrNQY2tvNjAg8fPvuLiiz4CCKkAOAgXGqR6KsT2h+nKYlSLbAe0w746m6KiVh3
RBbgZIOCy3CwEOCnGI1ZkHpFBsae2llZbRQS0ccJbRErolAks/8lqbdCjq17NZRvazssXQ7JPRe2
/mR+pBJDLaz5nZfcF4R3AY+SEjusAt4oH2Anf/AJNpDm+ZcRHDghuO/oYslABsk/AaTRQrQH/o5O
y3rd1S4hRNV/thRzrJ7Z+965JO0OEUOqFGKPGdVsV/KtVDx1OGOebd8kl9yU3bNCDqR679EwgaTv
XsZE1E9FjvALqyLJhOREvKhQkgEd9QEghafvT5KLhsv1ZBm0/43QMBcLCeHwT71nZoD+3/zUPfHl
37KiKtximjZqsbD7yPROCY14Nm3gJIgHLYbTi3D76YL7X80yE4mcICOrRIX8tRtx8CSkUdYSMHL2
5m6HESznSG+iEJsr/JkYy55s/A3zkQKPkqbfUwM1LRjCZVDKO4jz0ksUFXqxf7XMEv6Qloi0RiXv
ywNtFr5PEMaROXMpB7qWYdFVsWDZuJNwkkPYL2IQu941jGdt2lgjHCRZJcWqf6QzHwOCde8vyvGh
8awAthxjIaRNq5lmgNHjLAMeH4uv8OWHoXe/hIZlgfvoPyjIopprf3JtKLHMx9t2s8QT413vzgwA
tUfba+9NrVdIjFmHrTKnVGV4gPYhxhz+D7L3fMn1A8sqsxRBWcnAbP9caFz+FYfIOewa80pAVi0j
BMfGzrYdv++hccttw/DM/fw0IzYoVTf23ZP4pEaB2vyGgyV0rFnvt/sXhH5odM/bXow+jAYCfMQm
ii42D1UkcToPIqX1iSjCXXpGjp8fSijOIq7qMUoHUHzMp0xnfQhsi0uQanlRajbTTojDJLrwnjki
YV+AU9PHi5j8e4DAqiq+lw+ChAXTYwiS1FSJf2/RZ+d/CKhqVQFzGKWrip+kixnMk5e3UAzRuEDQ
uBGrVRp6IUKnOeRekxLrJ2cL2Rslr2YG0meUlx6Av+F2hBC4YPVxm6t1wbakZoVT7gzJzz0RT2CY
A+afIjrI8S2nsyGEujUJRsUTTbcrXSG3QdfOuxb3r6HnUFX2ktU63ztCxjelDhQV9n2RBoM5m4dr
i/U48y562VYre9YWCL0v2snWOiFgMlil6yirzivhX/uFecNTaghrDZwBbDPXPrkazOS2boWVRpNr
aU8XDnlqymMApV6l1owIuMiGwFsaXjtVweNhL7ucmAFjqi57HfgMJslFQyO9ilEW6bcMY9gGxnxL
FaxYbQUp/sY5ya0xAiqSGlqu/LRZcqsn2QBVKggeFYf23jcTcmtGlExnIeTmyQ7JYuGi8kw9I+IQ
dGmgZ3O4xADwt9H1Y0UrS2fKxJrRfL6Ohg2+zI9mWaPF/N2rS4nCzgF1vwJK7jgngQsBouVIeMjh
fLseh/bKx2yngXZXBtyDvgHixlThHW7A40UZyh6nZ2OoR1tOWpMH56M5uRKWzNd584QRqWcsyLlo
k/aZA5kc1pi2hppJosTS3s33S/cL0XkHf2T6YdGdRgaLSS/A/MS+VsYQmX7qHl+40osn+ED/lZZW
cMIG6eI5WqlInuqQMYwJPSAUL+LJHy9V+O0WcASWLsEJ1ZzgVSUcQrPFbc1gv65lccYSJ8NvT0KP
MFVaGn9/gThBzhYn048st58zSIjb7gYRT53yTmX3ITLajgLSSyCRJyVY3wfQf7F5EZIozYC5NLKC
MlzQLSlLfhJKcDnNMHaQFoXKcwvwEv6mgqPTiolFaitIVLE/JTRXjLUnMTVu6ZdjTZIPx/C8Mj93
uSDbY5t8M2gVhZVO22zvg8SdNL8bzdGB6cWHKyvNzNOZfKAzHheWLe23s+rYdxXtP8r1a0uNPGz4
Ukoz6X7kYtwrh0ovLWCN0GPxUXvhAm9VJ2J1fAXsR6EwQZTpi88u6EQns238eDQSXrRdpZ9bbfky
GM68PvbLbbt9ENOP5p1XKb+aGpkr4aH4VV4+MjmTJ5PZMLhC1ybjC4ikvgCze6A6nQ0AARUAXCeY
Qj3eGT7he2zn1/ZaF0mMUFedUeodGjDICpBZ0zj6M81VIClQnH0lZ1IUWm4YzaV+jTIj5/Nwd7jy
3B7XemaV4QKFjt0xuaZgWVVXN/CLIJZnH0JtnRGlJwBXMu5+unS118p397jaTefzDwvUcaVX8T/F
vysE4knqoJlGkBZ9kpT/JrLWn41n+Bm+G8jkxsoLJLAf8tYuaHUqifoT8sncbUy1eIKpmGHiKNUn
Z1dDF317Uv/WlSkWoo+qWw4biNFyNrCehV7S0UyBLComQHaD1Oz3Q4HvlOij2b4eCLzv5J56acR9
tni6TXu3fZv8pvtw3bbZ4xNn0QVQCSACKKLLwlfZec07IYukpHygzuV9VKGXNFPEhTcGidcCr3HM
rAvYKgRy5grAvj2K0WQVx2AwP6N0YBRsF9T06YZ5UefYJNoRrt5LxcPENAvUbEjONP9NmjrRUjDp
2AEUSZa37qsuNpYXm54wC2Spql+/jlAE8Mg5L2D6yXKXCrMsMcaqFGql3AFg2goBye5d5U0ftg74
OrkdXMktuTqZG3XhDrFTjxf/GV+freCCXgk3TaqsaLQ9gFWFSk0a+/VI9voCBOxXhGpKR7gArgZZ
/ofKFFfVAJXdOZtafVJr4D9MutYpBPUVbDrRXpjxBlrFRw0saUwZIyXH4hlGebO/hiQUrDVdKgRM
SVJOZ8hWbK4EsBr1NPvbpt7277kRXlcP4A04bHnKYs2UG+gZaEkI4JlpETyoFeX21QYRElLfnuLn
S5iolFWU1yJD/rB+hkWx5q0iGIimXtmaVY9+hHkwfKKqCAFuQVQ12R9WhhMpMZFzp+jZDidEBiki
9LqDMaoh1pr8C4MOo/NNiSlPw0Q6SfpT0ru6PWDsAExWBYOaqtgxZrAae5p9jTWy6DINa/toXV28
1nVHRRVi87BxRc4Eh8i4od8MEmLceoDQiC4g6vyUI+BUH3agtSNJ8GKcTrKIrIrYriJslilSB8wz
KlgZgaYcy6dSb/RQMRGBY9x52El3WrxRfsO8BfPrUuZJrdImxVnt30VZsPLJf/bX3wptA6pDzTVy
VTGNF7EkevjNYVqNIW4RZYMYI7o5MczvA4xqjqGY7NF6ukdVEa4jdQAlYXivE74OKnRA/9gfjgKh
KEQKwzK2yTSUG39jtH9U0u6M9MVziWOpKJr8ORk/oyh+mab2px/KIcoCOPf0pD3pZ5T77vx8r4kZ
UfVZLRs9SMnpffxSNWFIuNIEIeNl0VHpnfiZANS4Y14bI0UTtD+zZN57Twh+MRRDcylEPX4+xAK4
xfEST4SqfsLcoRk5v44mgf/2NvZIpLI9+jJ/3wyiAfzpEligU7yj8y4XFbMnavV1QBOC+rsKyMuD
hvlKsGHrTv2y5Rj8R11e6LImkZTFXD1WOnbDKQ6JdN1jyJUumvGFcDjTcEhENAcJDPUxkp6sGLSu
LIoQDxs/LxzJ8iu4kkOc84dNADH6qQ34xleJyOUPo6mM4DGumETqxPr05Ltl8KYyUw5RfKbdD4fQ
bvh3tJa3ziy+k4VYfSkz9WXqpe31n8latqNLm70NzmzdcR65bzayRiox85Y7pOnpuMAwds0r94o1
V58bTYbYz9iHm1K4K+3V24YcrHv7FGwCA0tDBOx/y1YMVWh/io49bLSDweff2RLgT2QKJLD4kw6P
1a8E9cB/ZmFESeLVx5WDpVmYRxr+zfUKDpwhEtYrlMxg1P7F6/CxtJ/0c1dOjCGtgfuPX9rSdLJS
vU3xNRaYgCXp+LWZEhpjKzfStxb3Oa0aB4620ohHy3/neg4qDwSljQDWqAuQu3vdnTVcbsgj6em1
G6JxRqcdMDtfrpyFfOLglAV9KPo8AjKlRzeihU+/z+F2RlJ1YAIXiw8WDpG03ofGhCJRhY0TN97b
qsaj5wYTL0EM0gUeq9H1sC3K2BJHRtjzU/uhl/0dnLc3IBN7sJIdsqlpShG1BqnJDkCoUwpcXzNl
T8SIC15ETLMHohTn7YBrgw+wv0Z+Jj+Iw/Anak86h7KVnc7ZWEySiROJ4xYol5KdpAL1kn++YJKP
vvgJ1NNc7zPMBshi71/D5td3/8fq8euVzw8943Uq8S/To9MjnkBFRxQc0lX0aAQ+ef/kAA9Xojll
yqGF6rrK+fV952Jo5pupo9IARlLxAMGJ1SU6wTKjyRmmb2v6Qw6mPIQxND/IWVVgGW9KODbfj/AX
NyUQTo9TSsz2eT3q1xCzgc1RzdLW+0wXrUf0KLF7f8vD4G/YBtIXBhQub858lVZF9JOK9+AlL4lm
E/JoqP09/BwFPNNF6v70yCI6SdvFEGxdKTU5dwhcUvVFyTbtYT3d19h3oAWcHxkeOMFeYmLEvCXz
0x8h7NlpHZsVPolt+p0x734T2Z3o5vMkaIc66GyzmRrHDuNDahFXEIg0l7c0T8QjCBQ46qvOLkIM
CW6AUj3oAxJClssp9AB/O57cAXiAQBd+iaoqJILVUWiEF1rSy5lBMIxF4Zln+HpiOyolDmciexP4
m7CxSGQ6lWoio3GRHOwOb3aX9FnRKC7WXF3CmToSJ3D1Q8UAjiF9wjuv5JogQBudrfFJXm3+M1Sr
o9AvW+EjqX7JSlNehzddkqm8SjsS2VVWLOvzEwfxTJtVwze9Tk+dU7rA+XXK5uV/h2mA1btM5hUE
C/K3CWJfbSRRMXewqMFssilqdMBApzh3o+52SMasV50FBVlgYC8rylUb/l9/Q+IRXjTQNr2zcJVw
jk62lLbLiHjtEX7Hi1cEjuKHkdaYo9ndeiHR72wrwPLot02omrj9mHKGK+kA4BvfJ6/DTDgdaVtm
rFkzVw6nLS0tHql8ZDghdQFqiSHt9Oi16R5vqTVanlfNeNDG0BIvGt/N8x7dYZhoJABZ7N7M0xQo
pOYVBR/4+vrIVnXc9ZC+gW3h2/3b4kgSyadcfoSBduNetB4zedztsCp5rZNKBtrm/7eLVw1zIdjs
XAuhukYPKJxkYpIeLOaHC+3phuCW/syyUO4JKXvrrsGPUbQywabLX/LmyNSS0snWFhxZj3og7cfh
tX7aBP9Vf5loPNoKXwRyCBSuyj+Ks4+7vT3Kra9JhpLT870s5Qa56ToSHoo9howoi8cJzwndinRE
/1MC2h9FJni08CcPjmmzMl7p2BL3q29+qdI0QNq+RB4+lJsCnhb0o5x8QpvLOnRN8WpbXsVLA0Gr
jmS7VciQ7gJNBTtGZgXcK90djseWcOu1UukksQbUh92Yu0hVn2PE5Wyjf9LT9t7r3Srmyv3CBW7h
tR4ypbN+LxjXsIgNogTvuNv7ndK9b9ypVQzxQBbb62C/3+N6QLRypDMWOmk5Qajz1rPSZmKCnjmL
VqH5H+nFF9W11geCn/UsYeoGq35q3FZumDT5ogM4il0uyCP9h8CaE96SacUAsKNyPX1m3/X3LnH2
H+Unc3jQqGgHviRPPUwSsUNpySQibmHjgFeUFLA/yW+7x+5BdF48gsZoWw06zIKOBIcgleK+2Gn6
TfjuXhO5mwf4QN+oElALlC1U8VQSYL56Vi+qruyTpb1GJ21vt2weQMPlxGcefAjX+SKJEY+4g05e
MSQuEVtkx95aLUd65RIOzLYJClCgNiKJVZEUo4yHIBlXSedH6ergc8NYIZRtbpE1HUx6t7nKccYL
mhOuREHd92VKdrxb36kvosEkillCx3eba6UU87AMfWu7ZgkXJXI5iwdx1yELhUyOltkCix++KZJ+
8GTuTHKFQ/B/hnsGVZEgTVOEC+Sq+JPnZ9JAHY3QdkrDio3hZN17icumFD6P3flB6UZZidhmYGVf
VMTsWfxW+DmTDffrGDzF4HsHHTcjczwNsdM7pDZWvGNBb8thvH8HWTe/JB4HhPRylIJprDvXUHlZ
r6yo7os5dWyigSCKbA4VCVcwOQps9Cu+mA5r57qg1KP2YfR4c+OOfQX3raoOZIrkEliOdKc3Fa3L
5w8e/+hLyBAPRYcNm+w2Hdmg4thhkEW+o54TMa73rfNA2eQEW0W2zzjQQDi9Geu5ZuKK8OeJMnO8
bq8wP+wFIC9NaaAv5fNDlxi+bQe0ZON/dD7yKZjhZfx8BWuIaEvh0OpR7etsSBau3DKbOBbSK7Hz
/PfvmuGW4TDm0ts/K9dK9RygxP0KCeKTilLOBVnZ7/Yvyud3QwxD6zwTQ8i4BHkqfoyfCQKYePJV
ATNCsYeD3CfVd5H6Pa9k65kXbLNhve47LQ30GMLlrn3Hk3M5b/mGe314PmcYisXpkA7S4yg07UR1
OknBf0QfyHvvAG3db7xDAvsp921QFlVKyTGPSVsbKjczoN4Luu+fPidKq75rPWk6wL7EYuATxr5A
Mmi5YxIHtEiYTyLXL9ehLMWjXVhJF5dBx1VCB262dZgH41s6VCmxDgdxARU81zy/aES8QaxLfDum
CMfbIWI5jVYJn6702kuXXa8p4J1IeQQrs5Eoc0XQNUKhf64JnVBy3r0Ql9Ki7tsy5PO3WEpWPRMP
d4uxcFUATXPvkrKjI9+4omDFMHN8lsa23/pfXQ50EWsDUuNefGZNWXwUYTU6bLsYBFX+rdyBRnoD
zLhbdwPkZBB5nSmVeHVzQIt6rX9PQpqQJB9w9+seKtkTEw3ZQo0lHNG61OQNOouUOdMu5pqLYY5i
FUQZMmH7+LqMHUF6gvtKHt97FHX5gGCmkfShyaAief6fVDeatl8gMvjyICbqGRRHVJwPrtfkF4id
9nWQ2wKVJMC4cXKWI4VVgHCnTRj3IpR5mJUIEeEWxkCxiz71/Lspmi1MRGZkCBW2xLfXWkOC3m+R
Zd39b3T3gPsXA+CY9r4wkzwqYjpvEdWiDqqG/i6UXo7x9oDKZj8Z652qB63KvqIrV2fcP+1yZSeG
orYgs/+MY2U7x55oZObPTv2qmogzy6zeZCKwD/2Dlbph23d6vsevoZn92ADS1BqhPrwwhvh//jOg
Kp52rD+9q6Fkmeml8i2LBk2Z8WtT6GOgqTr5pQvxSDSB8ViBQImD0djWE+ob2YFzaVQzEePOnxK1
u1Ef3FuE4qC0zjdEGD3CCXdGT1XI+QziDHqnq2y5pisCG7k314c3B5HBYm2LAtWS80s1pac41Cfc
Dx//e4xQBl1aySUOsClko9eVZpHyCbCE3/Jwdv3MzR1wWeGavGLtdz8EJMUcm4HGIaotAsctNiW+
cdMWgMUvw3e0L8fZKBHUlUDSLXz32xhDOlUzKjC4DLH9IFza3jdzTYiQB7IkSDuJouqVoTOtyqxp
ytbBkST7egATsxlHztLuJDkW2IXkOfzAespJnLOzz4gS9/qAOZjTtzQgAOqahtgJXnUxNCNjoxbz
Krc0hDAn5m/9vIIa4U2sOMsuwmtK0RxoefqjYorOBGhzxazwnvCGGWgBg7nDqFrabSAMuXdHCy1d
vDji9i6AhC4Yu9iIGe99gKIn9evyGJ0sqpkHmQhgSv5rRjmtNGCZSJ6lntOzkuz/anZOwyLSmDjE
13VoYD2vQhhn12z4ZdIFMf/jdPIT5v1QmMMG4mflwffWquDrXxonFKn8uwVJ/thc/y2OKLZt9YTF
ALwW7LZxL4QCXT5l4MCeggPk/Kcovvt1tIV8J8GbBHwPxBPtCZLE5vMObaU0WL681/b9aiYmPHKZ
LkdSxsapgvmNfY0xWU8DCd6Vabt0nH1L7vZstQi8UG1TFoeK5uOK/1+MZAjxNN0rHHnLNErktlUU
eqARct8wGmsL7sSC6VoTGewtOS7G7efUyCLQEb8wy1Ua6HyDOADwyFlDWHc7gFkj4VXk0vGlAK9O
PoEloU6NhijL6lyWgz3yy6Y2nhIsqPzd2QO63IicpXC5gPoNOM4hChI/N0m0e7PKN4XBpUjhosuq
sa5cycF1b7qMZG1gYCYxK1TEnmr5ySeQNJTiP5W7tjYkzmJZlAVDqQ0W3zyuj+PC8GfFEaY2NqAb
SO+HJ99/tjrW26a5M9/apOVw99Gf3lcJCrFyd9Lb390FaGgT6um5C6sKyf0iklwMHVXemsru4b0L
RUQRK5jUL8gwOcr0ig102qgHJ2HEhwXgq8qy4YficFo3ed9Jd8LKnhu/8hUSfnkHnI8p2Oo0cRQc
8Hfyg1NX/JqfRrEbMu0c4H68QLrYVPfuweCpy7APk/chikiiRdiz8/Uv6b9vnJLCW21H+E8rhZm1
Qs5I83zbFUbDNXhIYXcGtlZjanpCwLV2w9Qpah7Y71T7gzBhm/KAmRR0jYcYkJbbazwjplqsiiWS
XIFWC5F8KAVj5G/LbVqAuB/hiOfMpy7qpVbUUIf0CpQSzjR1K1BtMwTmjTFLm3yKFMbTghsT4wNO
cBs8xXmGZsVl8unYEzL59mQJGaXGLSbRpTyB62jb8qAi1tdE0Ae1dmr1pI2/VrqxAIKUiiwfdKR0
KmwZhZ/x8qcWHVErfa644EjO9fsO3OMHXPrqjvIbBxHynYAp27sLTsIVJAMwviiBxjfohPbojF/8
//+75UxIz6RAezYdMXRF9ymNw81VC26CC2fKxzPtX4e3AHdbuyV++iLSPPtDdxywOKeDtTrdcGDI
iGoo4lARHh2uhc+BJzms6hRUmUBARfo8KB5RDZHHjlAuQlNH8lpcsBKe2sQBAIc4Rc0BiT5WymF/
E0g3uHrfWEhBs9dVjNPXP/MCtzKieYQjiWsrXX5vKdtebFj+pfWbn0e4AAfsU8DteYFBIOCglsV+
nTFWtSGHa0plmPjVLxXdU3LHE6jooOaszuQ/SgQxMHihhoc8r7CSS/tNIyXy3Iy6aFTx6CsHXX5V
57H9WjX/f3rI/ifCPj9pyRqB1XyL+aHnDrMyeaO9GEITs4HmhXiIRybSrvWaYwjjoYvj8QbwBCWH
OtjNrAwGLKj1MJexoj3bMX7f1Jcn/jKzw5WO0MAtFyXSkpsb0q5bLA3RdmxJV/xJYuHAonAFGr2R
Hdo9z3xVnhdo38yHk0Nzvh2bEVA4bUW/Cv6RztmgdrfvpmhMLfQ2Xt+yQ7ctaEDU4P9/kibLmSUc
CF6ce+xWq17laC6Yhxv2kuTBrDiS5cvaIyuHPJR+JckSCU2E9ZwJyK9eaixjDKabDQsQANrRF55E
4Zs/X+t3uAFGFbJhXQrRM3UD9xGF3BjIAeBfT1PYNljC7QTYp0ekLF7Sxd4AiUrXM8JcVUNKIAAR
jz3zrrEfJ4+3W1ivKTmu6NqLpCUiZf/3pfYjQ98sqBqcea9Cye9rszron7InMPhiVxx7pMa6Xcao
JjWSj20w3uHALg5UW9TrXqodqhXppOo3DCClsYKyezzpX8vIJVqIYwPpmMFEvDPLptHN5e8shBEy
rTHpQy/A5SamcfAbcmzW5FsQTtPjEcA1nHY16znC3krNHC0XQxBauLoYPlObsYb/SfDhPsFGN+4b
JzQOJ23CApNbF4GMdKBfzNg0mYiGjBvUmSJlJ7ebytHlJ8vlhZUFWHZDUzQYTkF1BewlpPtK3Vcy
ei80lxhTmrVbOC0OwjjyQpFR8xYax7CUpjq1n+lw3Ww61CwoY9Tb2snl1zcCZk5CSfne8rmI2Gw5
o3kKntVOGwtteLb5aSdKA6apEkDbHGx+zs8fMUPDigt719Qcb5xgKP3TKt8KzAA2TRUb3j94QySu
4+m/P4lfCOV9dtxvngBwyxwMCoiGtu5ianM4F7hnJyJ98XvFRnJQ7/iZ7oS9Oy1RF0YiyQmbL2AR
CocBxVqFHWeh12jkyBZd0R4Uq1AjgyrD/LTfviOO1N91/ZKRfMCgpgD3OI6rdbrD2mKLaq7nmFHf
auihZQ3r07f102m8gEhU3wFk0qFFK+oAyAX3QF+4BQ8j+ai+DevII4fdmqRNf8LpA3u8EFaF1AkA
BSz6LZRvIx8CFV9ma2EH4qHvl7ZhPNKPh7VHJ0zJbOHihTvVJEMccJG5EXeEm96GfRMw+28gXO26
LvKu1lnelOGdG2mDs3lnSVB/xTTLzDz0EBGe1j8SOBDQU6QyxAKw0lhjQvebB7JnGOOtRHmohsG6
F4LpL4xemNquIIs6yRSFsOT8pCbLL9XfdxTcaaI0GfCWe2xM+wC9+G+VjkCqWE+UicKQfr0XEdU7
pIP7Av1uDRIeNxJu86giALPIjvAVwxngJ2gYSYUYf9hE1Pg51YM5R23RlGNgucgTgakvPIp4Sq+K
soWDImnA/UA8iAoz3dS/bUaK+83sXuo6mI+AAQ3uIjEI28e4ACScteQ/PtzLzNFONGvyj3R1t9F9
RnYqHOCJkCuXRWdI+GhuE7l9r+v18eAkJLrJx5WsEI2iiIGM0mbCl6Rsf/Q626iki0XvP4lxXLxR
7P89jBpuZ57Q03eP4+po4z7qijsdiQUIae+8+Itm/9dJpVGZNKdwykfHjriNvjf2i1aAKvpqmlLR
02iTZHnn4WZr/GMIRzKIajERVJOG133qy6NLsTmujumCZuB4H6XIOs9pHC+Y2zSz3Uts+GX5fZDw
yDmf813CTDgCdR5dm+gx1JMfe3t2LJuSyWpEG0jsfVWCUWNctQc3iqfQxNsCZuWlGfxy1rO9Isv/
rMYg9hXvi13/cTbgmAzFKrDXbWTYxQ37zhsnQNeIf6p1n8ga/LcqtZ/W6OiOixzPg3lBInbn6cjY
HzbxybAaPQbmFERPBH4YgZ1JfluPVgRKk2eJZThwYLUWw5fFagV2r21Mj2GcBVPP9K80GmTmzSYk
+7hpY+G1wwn2PtzOaXtZe3pZDria9A2wOfLs93exLXH5BRcNrC4yUAiIjDSu+UHUF8gW1jqcgz1Z
wFL9wkE8/NqxbjXEZ8aXaq1HZvrCAM0eFLpngctC+69yZ4JQY3iyKQZDe4nOMA5L55lkx1SIzI5J
tZ+0ODIFHS4Tapv293R96asf6QEA6zzixBqTa/CHwTE6TPD93EKpjfNuinv7qF9lcOO9rt/WYCMr
66CQ52QVNcoNJa8Hdjp0hxvW0RZRxy4d3p6IS1PFq5jvvIgoNlcpAeP3nX2ad7Zgf+SL9yJZts3Q
XdpwgwSWzvk5YNg7sTQjM+e1bi0oP01+NbqdCz3kmu+7zhPlUbm88+saB5Rsl+LuVtOD9+hWeSYZ
+WDnXVr/+lZmuWH+PSPlcvJROC5zU7P7FgMZc/Evo2THid9x8EOkLwdWi+/NY1HVv9RcLJiM5Nk0
6Dr/uEl2bZRelptQGNMkc/pl+KlamVYJtfNlHg8VJgHCSqtHurAh87G/8skHVtAtNsr2UI0OQx2N
AgPHP0tGGtyirrSHlW7EYgzk49M8QssetXwTGsp16yrohWIePgEC5ui9LE2ehUUgr80UpdRBTE/P
KYlv4CFNqFeMwGxopIeTfTzvCJyWw1BpdA03atq2W0yyTJCAvuN4RReXdozGhPDtqlKHJQf5YkFN
uzfOC6JhdYGWRT2UzBgerK3WkgZbYn5QU8a8Or+e815zTd7ualhxWzHMFKYSjZkGdoXrZfwC3LUm
3OnssB0lC3hnLOLXZdgD6Qb/7Dp2pgJe44DhFRGsAs1jRruFd/IyMiKU+JNjW6BJd5hBfczp7dbh
4/nY85gm13rZvKwqLDUhUSvfNYnQ2Iy0n274unbQfmKJ7mzCeVdc57078UB9d51TzyA4eqnV3h5a
zwRb0JiSG4pP/TIDoW7yd7a7xO3KrqNXSbe5gH9pRcjgZeAztUzdEY1G+0jdNExEgaikOZttEbf1
pw+J8x98S5SquDI9L5cRGS9DDZcU47L6atKH0Lwv/HKti1L75TVbEfyNA6rKLUeyv5rVnvY00ndS
NMcwu1uYM+bc4HcsAVNKEQCk+B8ZJbEbuY/G450suEpwv9C7RsX8XLM8/hQXTuEo7+XWD57+5sr7
ir9QWXpyeVQysnptjOwXZ6FcRI0g+3v+P2M//CiGmG3RWwSe7DzJzYGADimsXhdbk1nGGdpUpTUj
GzikOiRbdVrXymh9AFLfj3j6QsOMkjrdYfuWyKkSLLbjvEGrEhLhb6wThzJz0+ddUKMKfkJUUHKn
EeiJU5BCwWKIAPDsk8i+RJ+WWdcd0AXqqaJCXcRq3bKUnPrBV9DElXepLCFa8Dntx6y+6z9Z92ez
0fTrazBm7LeX4s0cgWSQnnb+0Q2wpkFZ0KaJ1cM+MptMvFjCk50TxXGLg9dc4MfBwz77eI6ADg3x
hTNFAiKRd9AMutrEeTLW1gKZz7/sZ9P3JliGI+mpjU6BJCGDMuu/bR0p/kR9HFXtMDwNydeQ72Ep
NTDMBlNXmhbx0bmj/mj/V/ua2On5BKHxVWgD0WXt/cmUzO847ws928eTqILSjAlSWY6jXd83+k6k
R3VtHduO7N8+RV/ltzH9IqMlKrBGy5yCYmi5uyaCudfPxke8vCsaOZ89lkHAPLzZNaNzQfTltmxd
LMPNVTp/ysgsmgmpIOUh5cYcBkiOKtBZsDIQpMjIzs2+PXRDlb09GFkHZgFsdVWyHlndoqSvTwRR
P5huz74bDOpSpwDBlWZrKQK8CUU7VG0h4ExCCycAPHOPVWs5uyVeXAyHfr1/49rCb/OMg99FXAit
/H8zdw3zN+CmKJH7Z8Kj2mtbkkKkJj0RfXQMB4ZNYXsE4jSIsyVusarpBI9q8NDSp1XnNzCCJxo5
oOEWEEUyt5kgddjCcOBJDPUuc7f3Tf6/NePr2RkmXBLZzTFRnkOpjckBov0fDKzLEh28qyxgiOf2
dAl9I+LHF6ybwKJctOkB2hxhwXYsgTvvV7y3emIToWoieQdMMVXIfi5guIgpyZI3tn7e5xnfMfhA
zJycrG2hGQx+w5KoxoMeqkJ4acB9EVH/RcfG5GkBWXvi35Pi357Lb2SmWpTXm4CgS/RLO38+x15C
sDiRVeLgseF4Maelpsmk5UYhEBU0SSBnldUSmL+9zOd13ATISpLRfXkb9Yz3nas6R2Z2m/L5y/dg
PuAkmM8UQbk/srDE4GmJsfJFgBWPgggTOz04RMzNm152VoadnwJYBWKjPb+3eiH5ZyImP7NEB3s1
XZoTRE+NFHDTONxaTjS4B2IaZMRC1qyAnY3Ld5pzb45USYXy8mD2wusOvHhHLz94Lj/1vNTHvYh0
Coa/NsFMc4xByTeX3QSrSHtLyOGQzfJJIYZPnrNwiWoRwDOByk5pBI2vnB98zh6W2sfo8X+yFuwu
DLufEtl+Fl80hYsE1PUPlLzIrCOShVy07qV14Hz+PBxki+7MQ+XM1Otjdy+SNcwWroGZgLZmOWKx
r80S6agt22wpO95dfx4TQcLzxe/+dGjAMZB4NhsSl1qKFUxcdIR+8Uw96K0LU8/WIQhpfkzJRsT4
mNHXCjFEsW5333M52Sg3XoDTzl2IsNYyL8ScJKfbDz5dRqMF7Jm+fOM+WyptXYBu9pC+TeoSYVGZ
CXLs6Cd/rF5lQ1+jRF0ZBww9+y/ZmDcoJtHXVVwDsKSoPhM5EnOM1NeZENnU9GXeHyLTUQDk8i8x
YiPpkktIyAZPhm6EWdjaYs89QRrn5p88PmjX38Tzy7Z9w+DUlFYRnDHTEtKsMK5LeqQoJ0zFWKIl
x41SnvmBaTRshV5YPrwsKKy1eWaa8j5mmLDnrLNsEnL9JoYNi1zQg8WVg1u04bOnEICNKYkdr1Ch
7NFF+hJhWN0q/sw8Wo1flGDyjct+P/b7MANe39BgeYoqDLLx7Y186LbRfNSyq78tAVZl824md56D
y90Bg4TUmo/fMQWhDTFYHUKDgz1g99gZPy3mKwE8s0Y6RN2smiWkyzH/jALim7AhtGgAwSNaGrko
iPKuSV0sa1FSDEwLoaAa72/+u06+sqOxzWn0wSJkG8mals/PoYdRNT9hxtfhQJ/N4VPM1Zio5J1s
BAjVM5Pfc/Gvk7HYbSO6HV0uHpL9wYFMUuo+XyNWjtxopAF1PUCY20bopea30/hpEfRICjwjoYiW
Lxbi1Q0jRNeyIXelPcsi0KfsRzrxtya4DZgwQGj7uSvbrpdIJJyOD19j821qpAiHVFalROFQyA1T
7bCP7ud0elqSTvzlqcCPEhAHDMhyX0OcT9hGkVSbGehKEST+IEeLy+ujubi2xgkVx5g4q4yTotVr
PiQP7XatGizT8Ff1G6so5xov6eYsBNL2U2s9e21OoF/gOzsoSjm5sXjhtl1/PgQt0dED5NWbYmSF
p59oPT1dm3/z56doTPgKIXfABwagBOBRcPLrvQ8GRnFuHwKWrFjmhBz4imcSQ2n9n3BnjpwnhDZv
cGazp6+S9LPXMSGc/4yxbWPHrP3u7RSWsezI8F2JM/k3AO1nQ+7moxqSLbgQrvS/FrtrgnQAYEdI
w2qJ8oJYUuaNn1we5x1kXO/ytfp7kvdxPE4QsYDf89jLyTxuuowiKE0UoU79B06r5JOliXKYn3QR
QIJgRsluVCZad8PXKgffcwI9bOaer32ycURinkTgyWhirxr22h4XRFf1dCR801lH5pcJLMDATL7Q
caekBXrkOYMPcdjt91maX0aPIi9WJe8kS8LPDU4cC8EjkOEQdxtSM8INCH7rw0grjHjKEBiftvaT
zZ5xK5X5pcsVMMaAqnCwXgT8RKZkDDBpIkOTmylsNVdJcaJMJU8wUX4GU7GcLAJqUXqVNTb6tmXY
J5/AEKUtdEGYS8fF+wvNBJudH9LKqz5fY1h6/sHpaGzVYI/wUOBcDEF5kLs5VJ+HQWBEdGbc50e+
yS9Ebr0YnuaSAVBm14ZsV6YcdbBbEwNyG7xeGrObc/CT0SuRq4DJjGnLaonvLqmHGX/WA1H8C3e1
YRautI4nphwdlZGrF+hZrmyNbiz1mtk1djnf3Bk/m8ve7cTcNwyHzf3iEeWUgGcLF5sMoSOWaCCW
h+JJKzmURYsI5Bvyfn4NMQrahmHlZI9XXgd3DYPCHaRti06u2Nws0Tbon8287dl2aSh8sUXUE1J5
I6pCUjBZUK5oQk0AakeZ29T/ig92BLnEPRaoeAwL51CRMcWsxsWjnPhJnE2s061CeoTEO8mv6srW
N6CfhMA/flAAtavfwqKQYZeJrPdattjA2ZncKyNajLk31cs1xvE0QesbV1aV2P6jrpFxazD1xZAj
/H5+QKC8jBGw1fVZyuMimbbvbEXZU0a+0GocD5WFbeE0jV6qwwaLdBhuxHyFuwvaAziYISREq6HA
IxdH71BntJN8DNHC1Rssy+HfTvb7RDpsWfzkg8D7G9P6H69OJGwbpOiWcBk7X2av7LmLsrIpwHF9
JiRGpqR4v6Gpaii4iJywFvA5F4GeaW/G1wvDFgZKYTBU/5XofQMJKnUtCcszK4qdAJON8kDf2Nc2
2rry17bbDAv5eIIaFMmD9OPoG2p5/Z4agCzsguqmRaIvsBLBFDU1bK4T8rcRe0/etsdS9ITTGqLs
Af3jwUUw1RqSXQzwImwi9yOvtKRTZDF5sTs7scz9otTImdtjPXPNY9/IrNzgXPLANHNEHJovNBjS
3iWWHsT39UvYCE/ZMP6RkCXQOj/g8lbOv7pxXV2h7noygK08MjalYBT+tO61idLkv1k1KGilDzkg
a2bQxkkcHpSc7nATlXUrIaHVPgzzgoyy0DAc105F664Mpo7Sw6KgCTlrIh0Xi0hm/mRoZttZIgle
5MK3HgzV/CKiUgI24n+Pngx1UPopNR7Un4CdX6TcDEkHt7iuMLdCp71cdKoRlgr7wTOU/tNXNYXw
bpgXWy5bBgeJbmErtOJMJHrD1IjU40W3m0xrF94WgU3zXXtKV7PGydiBJ/FjXCParUigdMa060sN
FUzSdPSX/A9154ZIMmmVWkeACVGxf3LMFojXxO1Gh3MJsKFh+nxPVWZTYduL7RuwrRNJuScn4q5w
i/pRyAaTLe5LQEX6WMMVfUtSvnTX/oKEYiDXRy2DPGIOwrQtVLTWIq8rCbXHrPpkyeQ007x+DDFo
0LLxsw6HiyFEk0hXarhAtryjSNdSW52c3eU5uVxcYRZG6axxhABSejjVKjb9PSXia3O1srSgiPP/
DFKzVEiPEe/1hjjShO9JZc9k3fHCnHGIprtLlXpa/av7SU8+y882AoomwM/+8/GKsNlN5M7SkiDk
9z5QCcfTclkSN5uWFRa08e4OfViV2Y8Rmj9eyVO/CJgriS0qxWujaoQJ2WSrX2LjBvxo2QUA8lia
EjPo1zTLEMUOUTGHV35E3dqiLCaa6bw+V0JJvvQGIYsRAzWcWFA2quiYihIjoKaxfaxVjz4QzCni
DEH/0QB2M4Pwp+pnN0FSabTA9TcSfjHXhv1i+pZjjloC+RWepu/X6rTLdXVMv6ihS+FQ57iAJL8e
3zEnTEUyPLTX+J2r6txO8j1VS6pA9DRk0YWyq+lcAm2e0MbLPyf5TQG/mLjwCpIDjW+/CyYVfTiF
px/VnsO1qZ/Mx2Pwb2ewwV+Jgkxg3rupvR59acazNIpzmTVIy3UXx0vDvn6q3+54GHucKTEcJx87
/F9960f3abtcap7jelpUXqceN3SIlx3yLs0XvYsnqJUC7uj91K+/QoG+IoKD4XEQAlVa6V1CpgMC
Ev9IR2Xvfg4QHV8jg7hBXbOe0zgutz6aJUlGR2RhfNUp1u38n5MDtk6lhxc9MVki5Fe8S8xUzo4D
H0prvASFjS1YbOAFLDI3V//hgZ/vImuvjI96mNRz3u07voObgqm342M39M5USIjVIThpReW9IIMa
kn3GvRriEuXz9c96vdeDCb4PwhNFTS+7d0jjcZZ48MpLdDCG6BcjIDvgwvu4+0kHrH3IpxrW1A/J
HA4iolMHKJqZ4KvJtwN9AC40nSXhLwrl9v1TJO0P4VkpS9HrM1L1iEgpZcRoXz9gBEo22sMl2koQ
seD6onwl0WKx0sSahgd/bEsHz8taYcOkZXQanbTw99FWr2HkE1/vMw9Od3+7Ne1/E7myBzu7dxUa
tEHFNNNeckRmMX1HqrZFLsxEgOAGW8sH25hQ+0Mw28HuKPxSJ4LCy9LaFTGrW2gT7xguI0YvV650
LEQ2d+4ZRVkPvPKKhXmh+Z0Ny9Q0KcHS/w80PSMWicZfLKfUev5ZeZffSxFECI47P6anELRIOIsj
UjjbIQQs5t14NsHlWtzy4cEmmxRR5svJODsfl31hf21FNmijM0w3aICPSyUfjb/qyW7Xeq34IJaH
+i4XDYRZ7+YgeAuCuLc6grV5ISkX9eaveOPzKxSZx27A4FkQRsRe90TbKOZa8fnis0JtzYo9viLJ
V6LWhNePuLUvh3KYsdhbpeaK3OfJF65YcYJ5vJ+Exd8kTuxYzqe4NUGlmFUj3KC4eTtR2DdpFOAh
IVHOzxK4/fyYx7d12JhudGqwiz9A7DNeTQRRKxwB11vmVCDsZTqys1dfY2ng1In67Sy1QPAQy+ZW
WF4PJGwC6LJdFbHhyOMLyt11wIu7cP05YI9mNBaAr7nN7c7oiMbDWHqz4ieTO7lc4kQWZ8toY+mD
ltg55RibeT2BzVWHSQMI+qzWIzwsaC72XmVISw39ZXLo7EWJb/oy8+67QFasnXOAZY3A/JKTQXfm
fZlNwk8vE1zjIy4TWjpI9mAQ+CZGlaopCGVfwEJiXLNKcUlqnEdaPG2U030Y+Omb9dmG/8KYp+Cs
Za5yXt/dVoIlJ5zvesl323lb0CyhYXwYdPTyj0Fc6/NEPeKlMK0BKdhEectsY80fxguvHpX8jGfc
bIYRnu0o0JMHSiw1nbyr0pYCKokIw2xZjBz3uj6JXVqmqZ4r4DKXNkCA4i0sJ9eBy/xTBqHmnqUN
LCqBTpy+J/TzvVXqWfceM5K755svZcxL9R31EEE8m0nF7P9hApNJ9wdggYhdIF2by4P4ZI5YXFwC
43rGSl4b7Y6M8KT9Fuah7hBzcg+4FLNdT4TgnPiyggdc4lHA4z1l6I4YMdNWzH8056SbEGID3ofi
MBI5+2l1G0Lj4KSxppRAopt7buZJv3v12M+RmEUN7WuC2mHYciKvflzuZuNiEfvsDUlcDIQXNd22
OLdbU/lJd2x6pkfR3/oUTahmdPIj6+IoYENKpf/rIDcASNrc7Rq/bqkcoePoJf43wmsI+62zO25C
xRGehR/nD25/QwEuKh2Z8Qlk28nvTgi1NBZedW21XWS2KYaqY9iUXp65eLvWMcvAwzFHCVB34dej
E5NRMmsOAOIuBwOm6sw1iA20lVqsLEFoBwqSXPOGKhDlJKwziJtB2fgVRdQlC/yFohqO1OX4K2UG
Tj8zzTS7QbugxCn5NF4WiMW//Gr0RzzP0Xu96POaEUpsqU01Xofc8Bl7s2JZdjMfsgUconrdSjU5
6kyygKD4syC8RUgdzbdJnnam/tTkoAIGI7qH/Bh7CkBUpov8DIFQQ2XvN4JfeORpP0vaQcTBHWKO
XjHF9FK/gfzqnwbFq27eHm57KkH2/qhMc+RW8fVVEzWBwC4t/dNGT0ixinR8EurVu+wnYJIt4EIV
gMRWlf4k9aTRySZ6s6uR7pOIapT4HLX3jkXf/fTtIIRXT0yv8ZJKtpvXmHrNARL3pv2eUl8wzNdv
xyw541xOOCDCQpE4w2ZFIminkOVKsAFexvbTI+KGRSUgAQ6YWZB4mSxwJSUIo63vhcXGu73cpgVv
3vZmbPmkYL9JJVru+wtraRnZgl9hOX+MLqqiX3pHBmRR6pJcwk+vSU/u2HHRnySAwy4RInGk5mzd
cC7yyZ2jwh1LlvAvb4VOWxp0OPkqxTj5GgUYWSxWFc+vMUzDJ1yoS6mbZO4CNyxqh4mqwK4aypEz
b76AdIJckeZg6UH/mX5Z4DYpwRkgGGZBwdBa7jVx/KwZPTezedn7xPSzb09w3j4CoSIcStX691jS
vjaihfxTc1Xn+tRcfsuzpe2JDsKGCmszvH8N0dgFICxonG8eaHPuHIuSGClo+bHoSWAp81Vt/ePM
gW0VlJUyVoqXteqA9aFPKr4fQ6PHIjTaK4tef2kp4SIJolo1P4tlcfiwzPFMiWIevc+9iUI8bPUa
WAVFKGo+0op6OhZ0e4IllTxiE43T/0Aky0A9DgW7bLYIx64Y7VALEZVc1X+1JCp7HOPAtxA0kkJq
nLQbRcLzwED06Li8TEBE+W9Ongy3luj/vicyEDJwK2tD7y28I2zG1yHYZ34YIBMnGyQSDlEadcst
OevoYSbhgRv3xjtRLL8RmRmDFyoAZ1qTbYDkyGjRoQgnZZ+tOiT2ne2SUS+1VcNuTyYzKLiPH36z
66O4Y9HjmRBPfZGSe5AfJvNEw/RbBe8SNDmiO57IujiRTC6ycXUy1sJK8T7YZrJF/qRqTUidOc5B
k5IMVlvZ5OCuDMtLwz/ukgEPTq2JaVdWmsBuR+9CjPi1myI9x+1lCN2uqP5krput0qJII9ie41tj
5Nks/gIQKSmRZCSoGc9Xa5vtFi9RMfAtLh0DZMCGi+kDL1GtbHYkeRwXACHybmysEwI9hYTWRClT
meCmHGsYsLfNAtjp+TpYSCbpD05xEou9v0XlYr1sExvsnsxwJdokTw8gv8L7LoUoPIL4PTQwLTay
hEkQ51riElymeHkT9KPVNOKZZDzgIXag387eGtvdV/0AEtHdjB6vQ7eBM5RNZpBdalh7bb3eXJuz
n+C//ZdU6CvM4QXJPjRx1tlF6oxEHfViGRSTqxnY/wUpaLX4XxVFKeOMnMr+0sNATaFFQfiLtbgy
o7rdjIz3FmBX0BR9jJ3AQW9T1VAvuy1E+V5nufnCR8uZao2aX2PKwuPsZFDjCR7xxpdPqc5WYy3v
yMTdtUQ7C0DmvtdnEveProCmrSkKpNiBTUZGA5QitiCT6mF9w0TO5tJLMcetkFmOOQpGOSz087yq
q+AiKP99wBFc90KnQ7EIsghgmlKUThfgHD2sF5c/oJ2jzxOHLMqlEfCFKaC97PmXDcHgsFnd6j0x
ys8ryonldyxDfidFNslfmJ6U4lysOEdUjwQhOQAKJttq3dM+TU0CvL6hzMyL0kBcom7IsrHNxsSY
q3eo8tzyua+fPRFYTYzjLdVpOvmmCGFN90LRWBoF9pbQHKFvypTTefwNnpYGH1ljXmMg0oK+gxkN
8ou6ht8VrTa1eSXHtNv1MQWOZZQH91VEM4OS08R++F3bNHu538izi5HjHWTo8Iz1lFfOdl3c91qp
5N6qsoxNf+zxO9yRG5SVI1iEyjwAzPyHZB+zJFrUgS/a1aYLxZbyP0OW7byAtINvRQBKEE8AgTvB
YUOb7tr2XjpFrkE0KuC3DEkNEFeZgNUkKLMtsX6kDw9QZs8Gakj1hxczaa3QPvaXR4263q8RNl75
o1SkkPlUIBVAqWizxLMxzo/pFd68/czlX0PLbY/mFwip0UdUnB1Ad8Xkco3a/z4gYBiJL/9GaxvX
9jUi+k+nK9xTicl13uZI9vVTIhVB3Y3ZbnQSOptAOMbvIVnld+qrdem80aFSIAsSRy9IXsnShU6C
wLdx1mTqWXviNlO336XCjXAnfwYkyvpm+TUywUNT+7sFjMvkjAME41EjKIOlDMQdefWXW2lWu5Re
xuPUQCeVyRPT/WW/r/LuGOB9Id5tcHh+BOpCEehbTxgNbYOdRNLTvXUEansk9pVfKZV50GNzVE/N
cJQwe30pS/QoMYUXXyDgbtK1wuC4fusZig5af3adPyhUiXIUW2W61Jo4c1OShK89d/mdby1OqT9K
3rbdA+gyqqR08T4RCwcimryX+J98SrQkD+KGt2jRyDpU2QCuNP1ukIMBDBcMdJmedpsAgZZx2TCW
4PJhCNo79RUnyZ62jHPf7mjZoPNQOHM+eFOuYX84NuQ480MBcCd+rjbX6TfY/kWDLY7euzBf95G+
lV5HYBVM4trcWxSKJKAAvH5Op8MiN7SHBkqbG6IJy9BObUL9JEJ9Ey6R0EDLBnO1ol7q/nbFD1ef
/pPXD066EoD2FIGDoBHCcTn0PcGFsNxt/PzjXKR8sK4DxfMnnDprLoHDPvgqUtpEzZBbcBtQxkwl
/xdSv6yjFnwKfdz0CgDoRAPf/NMnerQrUWHi4tXCSezwgSBDKIDaR/FNUuw/b04KNtFCwd9puowe
Ov0uRzrmt48yDvgPs52IS2I8lyK/9xs+NyynrHEApI2Z6+AjeJN6NoF0Z3B1kWBBOeawmPCUKvJy
T25nIxCTrXCP8y/boFcng8fh8O6JDWUXqhjvoz7G8AjZYH3BpM0ogu3js+0B8a9rglrfv/6QmwQR
OPDQU1O0z09/6HQbTY/FkPcoLs9whIRF9oo03xPapazood/zl0plgXmu6JHCtNLW24zAERoJRKXU
P0ZZL7HvbbYUbhyt9yIj6ivucgqBSNBSLATstZZqp9/fXpKl3hTpPl/aDr77A6k34b3G5sQnd0gs
ba335tu0yQsJYyp/JAqBRzO1lLlEEcRAQ7yLM42mMOnS4e2jvUUby4C6snE/Ulg35kXt9fdUalyk
PVU9FMGndDas97wlR4xsjPQXoH1ZWIpV5JZYdCjIe4wkK0Kn93VTvbuOQxA737e1RNrRZynydQq2
SCuQ2Pj0IkafGqhHPOs25QifsoLjQLGoBvy8xI0/USuB1rqnQJH1Yagbfzo3UwwNsoIgbj3yNeg8
6k/ikeq2ZV2B0Wi+nVqWfEhJv9XGJoX/qqaZQ554Kz9LKj+8Bgn1spT3u2iVBvfOmGHYroCOqQ/N
7AlDZoEzk5w2SB9/d0hlTtqjZyZnCUGimQKGJ2JWdrn2TpvciaLEeUUckqfRwr0URYMijn72vYO+
iFrCgas5Eru2/xmOUA4PNKfBJCPMWsDDl4L0ED0LriVpuJ6KFdCcTPz4I0RcbGDLCyfnsFvf6exe
u9arHEYs6+Pua+Qqf5Szvrs8g3kj7YOsi7dbPbBxt5Yq6ZI1TbFASybVdX0DJtHCem8LFBBzlbEd
TZF2oXhTIUU/Yg57dXdS6pujJgxd9Ptb2Y1EXljwsmrAhnCFglLQYZPx06pNUjZFi5gP1toNKOz2
GRu3czo/wdW/VFWn0moSeUAc4eGqoktqsEVU9Ad9x6pj5X/3ZbujjfL5p2inqCtNb50EIAJv6u6l
g4ng4Obd2cjqkLF8u2SvRTmvmlzu91rZCSuM80QdHcfFWiPlzhT8icW/wTnF0BD+bZchs58PeuZG
/5R0jYjVt4HsRXUqiwDB22MTrXLM61p1Agqq5SOItmsoIVk9dqJGcIV3iBzvr+9hN8CC0jQpIXhM
1S0NCoVBaDsO7jgkIHS5pNMlFVzDCJybJqzVirp6MEH5AQBAEJMn4PKc/AT5lUTEQBQ5xaNBsnwr
V/kANRjIb0xh7270h0MM0sukJMtFlkEbBznfTwRN5kyCzVC4KibPJALe/3CZOZ1gQbP7e5lc74jB
qkaipDoBTKtOWlLw1al0Zz+WFEEmGIKuTImCbfqNYmyW0R25Rw0UcYU5ZDrxiMZHDb0VcrM0DXU6
IzQ923E5UUWRmrCmxDCuEwuY23n9emKS9xT5dbu/j0H49iLDRMG7ifJVdULOW/x911Ju6hz5KFhq
gXWByUmMAIRor1WVZLArvYn5U5FEfy9PtBwrqodpAjP+lbDvnNTlxJkpUmaMtdKv+EWqRdrhTmJp
cXSaUUaBRkazEZQrd2zfhZSrBSSYEFeqDM6nZ0QcmzOmhizyt0NAq1Q5E4rF4edn9bqhLclRIltr
HcHisOpfamuo5wXzTXvZoeWdGD0RKB3zmdrp0PjGJ0zUHu67kSnE9sk2ZnTo0CDGJs/HVUyiz50U
zh1gtRvatDeqVXi32Jr30YERcYNnOXLMql90HD4ieiw1h8xW2HbVli9DzqUQIz2Zc69lNnwifS2Y
QP2HfWP5XCbs0jYfkoV0XCLfaFBgajbdjF3XSaXPlEZcMQvSNGz4SeV62cIbA6eNNvY7C6qvlqef
bU3gqMw5J8An/5HkyjoaV58l7v2VnVOjnQZMf+pp7/02HYT1qbLLWmiru9H+ppS7ygd56Jgm6e6e
dKam2g97c7SPsqIKHuaZehtlI/MH7hIQOHEo6SoQ2Qhuj+dau5stuBz0jM3NqSSYOIlMpuDxiXOn
6TVjT+VFR3pfsF1ZO1sckTRfQjwklmw0dx4TbVI9lx7TF64cE3ozx1Q2+Ef2Zg5j2vnu766HmUev
/y9HUik3kVJgv+XgkcIbTDtwF/7L+2R7iyE4Ue1Xbk7j10njr4mwMyF1m9fBMM8FaaF7LB15nOPH
bPz+9hOlG6znurzG51QU2aDvWMPpMN2KSjTOwZ+QmqYu+fD0FhqBYBhuHeoefZ42Y8vKJX14Ef1R
EawseQnGUgKCzYXEMZztQy/Ro0oP5Dd5J//tu4IC2lXoq1FeLqU6voj2rc/KzA1WXuFrGGDjTewQ
Wy+ldrbzJyGv5I7t7Un5QYYrhf9JiqYpVW5/2/LvmUT/6+P6W1ApFMfSUysBNnLvgHOr3p8kEDs+
/mDqxJgb/dFZAxUWK4O5FhXb+WlObvw4aAWEl++My6/KSY9HCrwNwzYsyJtvInbbb2VbWv8RtmhF
CeX+l9/sAgz/EDfRFJbOy0qFXiBfWYk0awWO7JCerUEQTsuKWW7HV3QoxdwDGW/lUYyId1hqQNoh
vojyd5aMhEIOFuLm705naRlIql+0lVMTmHMwd5VpR8AmzqCVRn6ZX86fvLZTO7WQzHoXRYeMgeZO
bMj7aEnk/vdgoFRmOQqy2RUIajpwOCjxrLItiEDy9Iw3OlI4kv73sWMOy/wfvB+IUorUWgaV6U5Q
G3Dss9LU+1K8lKJ7MT2CuRKxAVcYQAD0U1+fEdtk8tL6CpPBkvY2iEeOpDW6Q7SerZ4nn58gUGzA
5lEr90+wjiTMvqgZC4JH+5ZFMWG02krXpM8B8s/gJrtXZU5H/BA88zF0pKCb1hKObBjwDeulBFLK
4jlZCAFWVkuIbPrmwE4mRLnDw0m0sIo4QF1LAUzT001lgrGqCzZDwR2bPNZ870UC9/GnDChrALZD
ELBp59Nb/95Ex5HviQKindio+M3lAm8oGchBdT2nlPd+jtTxhmHPOolNkVHnNEhH731IrYJU9pmz
kddk238oRnJIwMHn+uHZ1hdaBv+p0ml7cZudvzYeMYvY5rvmVUKAoRCNO1jZcItSe+YPZ+BBlvsR
t/IoZIWdJFEmpGuc7YDlViSVKbVVgt2WqnPUmAHbe2b4tpXaVZeYUbrx+Sb7EItC5Q9D1QKuah+2
YXLD2JfGRPisUaLbpWKX00tmkIuKM9PmQvmm5Z2VWxG1ay12HltYrSl0mVSBkGm5NAngD3yamdKr
jCTtrJ7xaAp6GbWzDx02DFINx1MANZvOkVQe49ETKYfNSqvEDiXcQI3UxyOQIXpvUzXMNwTSyKhd
IH5PUnWcsWy38GV2L8qoosWab8SFi7I2049x6z0ajyQSfYrSkKZoCPQxKzRkfPPWXQQj0AHM93eh
Xtk8brraiPdndzJc9Hzr0/tzRvxQxFWXkxnq1v6TNYbZpPpNf1rqiZ+71AFK++MTY2hiIqYQv0i+
MG6I2Pd+QqcbV4Z/a53qMB/CWjQjU7mYFXx8nB0nEeTrRnPVL7f6Z+tsKhWNFhEHXuOycU4KXWJr
UH2DkKwvZZFHKVYTm5prNBRfk0nowaIJH+D9KOhGSDu4l+3oxuwxjZF9w3QpyfA8eqyYRydQhltH
cnPfwfnZNuUNBmGz/x5t8K8g9seXSPaPOO7eXyLWgHyoDJ8l/fhNwmX3B8MUGLClbuoE2KzETnpq
KgtO5CPY242YixVo2n8Jq/zkPfKLZXDWF9Chu6Z/7JqT4Pax3R96QgmWYFqcXZWTpkES+TeDLSIu
OgSofMkj0C8TXtUVjtaapM5R128a5ErZ5uUlAKUohRWt2/XFmZBcKuxSJsvqbuJ/Bgv1lDJFZdhL
HobvawgF795KMmQWzP7nv2cH1z9U27iOLO9MzCXpC9GW4pkU2hz9RK2G7UxflE0epGCITp0HOxV3
gAhQtrFF0IsSwI3BZkAIXxaRDpMbwLqgOqycEGkB1GtkCBQ7eMbmFyID8CQIxE4cLUZTztxrccv2
DDfmhWSjsZKUNCL4YUGzoftD2sLiFCppq4JpqFKfgZ9oT3voUXiKo/ieHlw9v+8fPWKnHCSoLccL
0A8NRapgWu+/+lLgRRDhn9rfhYSeEQgSsyHxxRBpemZMfekYFy8cKGq/1Z1iORMMJ5in2wgZxT3M
0iDQa9k2NnoNpeEVFCa3iGtn+nopRGpeAOz4g7aaT1O0Xz74oEpzjwfetq2N58hiG7sFzFnCZAlH
k1w35JXi7/sNu4rxhbbXADFnsrowW9s7n76bCOekjVg4bbypT1ZhslCrye17xoDAdk6d5OELDndL
EGzhshFnCb6DvFbuzfH0CyROYnHXu3zSJV5p+9wuAJ0AD+vQ/JcA6lLuxhM4gDLLUObCso7B5EaE
HFE+jfgcnBdVpvhdiSwqZHvBpFJq5V8RVap8mtJj+rZGtku0m2d/tXg8TCYojCmT+bBtKVwo+iMU
pW5AGOSnTZN4lUB21pRwixypjmgJWAkIHAJj8WLFhoz8MWRoNxESN6o++6NAxO3m4OhybU70xQFb
AMmwPnWGPNp1Jd1e0tajHCiqxwpZZzT/aHBhehN2+owjt9bQHuCQMVoXnjU23hoFGIN/i3gi5GhW
BhLtwou0tcXG0vyJURSy1PZvpwG5khKFft7fYWyzb3mVzU9ttl9J4UwgnXUI7flj6YkTC3bG7GcM
GPpJbe777uiRkSBdQSuBJ0zUIj9tUP2GjvSF6/zRa9T62vTGLj2dX4ULoBRWIVpGCxCBS8HtRe9p
1Hh7aiif4fuMCA88t1yRFgl81aEXkDRqAecQpVmndX9QhPUnCn18BdauYJZ8Dne4dVdSNIIGAjaA
cFnurLx0nbRMm3eWQfDZJXqK6UblTyNg07bjWIr9HbVfBlo6z36l6J/J9zCEGXGBt9mK3e/ILeNF
sWHWrNCZX/NBtgscuHsfzOU6fyIWYexFsQ70kn3Hvf7mAtcto/RYKUZYmDZnQYmWwryIgV/eoqGG
xuzcrMB2lVK44wQ7OidFayEVqDoS3eOhC+OiuSET51wlurhBcKCuH4hskXTVgeFAHzWuQTM6sf42
+KLCt8EPbF49EaM2Gf/yFNV+dIF7uhOXQcYAINhJvU/Zophu6LfhbImNSJDQeiEtVRSl9McB1LJP
t+JhnA/fdQDNEoJovLRhujn4W0iHT290gtqlHR/1wCCi2wFdJR2EpAZEI1bNh7UeE104BE1Gfqtk
F0PYhIcndsJ4LgBKQMxW5HJWK1il33LpLIOSbi9p+3XlxyU8Qa5D0QzAHTuV2n1yyDAjTlkDVdtU
2w1BUVuZ+VR7ZoCrN5zk6YGGd4EdsC9mFBqzxE+dzh9EHnB6FZH6EclSiYsqdvZuHGJfbZp0F09u
LFdEp3iwnxgrGD2t3b163UZDGgbGyi4CI76ZeFo0XyAxfmh9MSGQDENmcil+bFUXKSRONGYk18A8
gSf9WMRT2RBDWzSjtVv+fI3wMaQqCrDR/fdnxEXLT3MMCws7y5t0fopEd4chkcnKaYCdARixRD7E
vqT46XPiU6p4XcoP0VR2dORDAL/Q3t94yaDOwpA5bI2IxaV+JjXhort9G7E2DU2/r8pnQXo70dGn
8dhHMkNaY5PYdgAxFSW+vfQWfh0W856HfnXpsO0F+VVCAwUoXQs7pHPb7/TQoGBU7VX78n7jZrBV
7JQiL7UbzvkVUXPoao2PV7BXDIGCjJua1Bp8Ti25vuTcqLoNATtKCm3rphQk3i+MI44E2ZsZkk7X
sVjgDT/7GKMPmsW+MXX4FaUQ/XKVkxsuRy4ni7XK/Sm0WzFFffRGcy1vPBazwcQE4Z7laeF2la8H
hABfNkYlrgvogojRdP9N7XmwkfK0EX/MDcddDTyL9cQs93uHyMQlc1/GDTX7DtnEWW6qQJES4uN+
oR4CGuMpzXueGNLMhDqZkUrhz0TLPmtQXIKWEv8zhXJYcTkauZPox61EP53WL3hnU/B+WdOEtMXU
5VFhft56pQoE+9vvXQBSn5PnrrItajintk9nzOOpT6YY2FKMoMz7fTwnOh5ZMQIxy2dYaIaolGH+
HyAEMsJFqMD+ynj4gIIOy6UZnItrujgktJIn8ITp/WVZst6TMnsQBiI5PQcPqgqfSxhxRmxEcYZb
lJTo3ktLA63/DVuZryWQIJndTEo++5SSLtTA/p12V8HiJo8gV2gOLSTO0SkdzsaxtncgxzZf769P
2XVZG0BHASSA/D1NTtQYx02pIfBbwrmDUzH/ZQaiJxXhODvmuQhGvxh/AXJfobnPHmHi+PlP92T0
narsL162MbwCU5UzsZRxNY0L/Mk0ug2vdwZ+Z14qUKTSiaYM14T450HFL0eH9K3TFEp4pltiVXpn
6Z3PY5wVzc6dtHBPcwmFbAKQ4SwKIfaRe66fCNWivAAE1LYdg09iPJ5fb7BixtT9OFzMSr0xz4kt
kEMFmEugSsLb2I7LaU+tu+wUbT+mEX/Y9a3Q2wH0TA7rc/gYiThhxF1zmuxgFeP6QmIURPlgB05m
cN7pzoO4yQSI/M7yk4IkR63hAIeEJxd6s57M1XwIb0yfiOR2gr0wWYPJR0CiqbXEJSgHaTeNNMK5
PBoQ/0yIvLfBGD6Rgh5OVeiQqqz01x1FpbXff9ecjwNX3AKsNZyF5POHiZfufAUrFBM9XQnSFu8a
iGKOJCGUYowo77p/ryHSXH71YZUmoyD/6ntPRsMvcZwElNfJYcfyxawE8XDhLXbKZOkMb+Lm/c+T
UuG2DO3BWQvPjr1e6KZQAjz+y3TCWrcS9W6abLfp9sQZUCfFcPOArAebXMreAD1FWmFbCMqmkDbj
CdWdZGcTzXH1g2G6Gp+44EvdjxacFB6MSvQoeFNOhwnXM8C4tgUj48qbO6oBJXwMv3ZD1Rhwq8Wy
C2vUrP/2bNPgYeA0JY3nmzDJAvry+jqCJV/jSqw6f3wPHs0xUoWdkYkxrJnk1LbBqZQtfr0agK+C
wRi+NRZU7xWi+cH52TDYa2cbUZMi8tg6ta+EYdoL6gjVIp0cWtqGPKZa1adRT0WoXNwOgyVjYE13
vxHEkAvL+kjZgGKxGTzLMY3Y1SVyYxQolHG9Km0Nhu5NTXSlbmXiaQrKD8Y2T8i2Y5TDg+lddcxs
6D7fGjhQJIAMYoAT2LcXz+ElV4a4uI3lQXfw/i43Dub47L6FOTawE+2lD5kp8LfrLtJZ4MtQFzHc
E0vM0VIKgYeWcYMZ7y80N+xDggWe7Ahmu2kn1fTsUCajxehH0DEYDGzfq1LgCIkuxrt49zjtss1g
L3Vg0aklHnnYUd8lpUKrFuiEFA8ledEWTLrt0ajmPbCnnF72GdsV5pX1/sQa2Ir2QHhU2mi9szSo
Rr0MzQirs6klBKmsZLiWjm22IklLG2nYnhCQU3XezN13lHzAYu9oSSdJQ1QQyRns4QqJoHe4cXlX
vwcNKEWFPJ0P2vk6yvkGdGL34Bibvn/cor5wlNXkmz3Ri+oDIlsOqEklEN6tzbkUCZ7L52lUB9FQ
AWJG0f8CHDWnU6ebUWI1Pjij8ijHHmEpI1JYhv7x7c9nwUJM/ak4VkEr4ryuWJc0dols0alfR9PH
favv1R+B1Ic7IyQKP3vEYpWfEoJ8BUGOZaxb7EzZrz2UCdAspNlkHwUd6E4E101Lhcma6Yoi5gax
w7118iFxiZQHknwSCQbvb4bq7CUMhikxNRBvUH3R6rAMHUQPMTeTveMS+74IuAB4dIc/IXLs0VdD
CgIA4Z6rJ7L2ZTLcesJcLUD5pd+LEzivV5J1FwqqIFKaY9etu4rcic8lo+YK43tv1I1+Tnr2dKhU
NC2LA+ug41X1vu7WDfOZWcvhhyB7chqx5Sxo2L4jGHIadTiQ5H8PZHmCUScJ5/Kuzdp3dIE2k26T
iaIyWp6an6t8fdgFHmzqLNUi6/dTBhoMmSKLwHzWrVO6RAKgkbTtORh8+jed00AoM9xSvP/vLR/+
I0fqpd+3PLiTw8GXsNlJL5mA9MD409kzLLutmkyG/sJwb8zlawYVC+f1vrSMHqxxuB7okUPEAXp+
Lyci5O7NhYHv2pZh6jMlhCNQvdCRFi6HbWfUXwM+ZpJHjS/dxre6fxgJfYfziUoQvdMB5WAiHCOh
olgcfD+6GHU71QYLfhr11ZRvtPROuJUOzq0lLXCct2oh/Hn9DwqZBH+xG8R9Tm63FQwF9SHgtiGW
bsEp4V+Zyc8inA+vOU7S6F2VA0vqt7ZA9qhzS6Sl1a9PzA2MSDGrdBgDdMYvofkWd9IABotYsHd6
Ltp3EyZph9wi5OpZm9I9De/7l6cZkU7oZ9BujxOs/exRL1H8UVhedMNwIeJkj22cxFnqCADrbgGk
t5e6E6dWDmTT6gB7dSOdQCxmh48a/QXfwrK76sb/WHeZrGf7Q8a9bBX98H7itWqfMwgqIRPUdpYE
0HeTshNPTyILn9obGverB8vt85G52F1ZIBRE7iHzAJlCw58On4BTf4amWxi2c1+5KF1hhy7VufCy
setT3LCOMTQMQx+rocqBbPrfCZYUnjJF+YovWiAYLV5bQ7VanwBUSBdm8xOpB8AgNxmkOteHo+D7
wpVvgSE1ZZRoOwJk2SprsfcVlMVN453OHQZamZ0ZmY/iXKW7+/LYAZDnx3WaO4pJLgdghjK7OYKl
vBKqlGRIBLzGoo4g4oIs7axA1MbQL6k/+LS67joIS/VOqsMJiFQGLvstYLd2mu92dCshj9QAJXEd
OtdLbGQf727/RASuveV9nkatFv19RuvI+MZjiXYG3qhqxviZRilFn77ycroVyv0rPr+Gy8Ti+eit
WvHQpLRMxws6C3WVhZMgmJyAy3GkRoHz55561qv01DFeyqCX+CD779gRyIOhoK1/ykSz3T76vwOq
hgeLTfG3FyXECG7b4jssfU1O1CqKo5xCIy41Q42f26Vq+D0ksNRXbguY6WITM21qYCU4mHt5aBGr
61NlBN5cdKnUiqWoRz6J26t0yU9KBxRm9D10wNrWyka1hvQJaN/JEPgnlP5i0Gi6S3bbzwrlNeup
62KkxmvO16/Y2KnqmD5rifgaNCvQwpN6lUtX0idXL+dPDz2KCsBbRz7rbHVnTrhMvqkQb7WpErgo
IAGH0XQ86pqMVGe+A0/tPm98DsxZA7w91lBRdzm+G7FhHDq11koiFcV1e51VtHD2uoaJVkPQsDsm
ZdmSB2WzqwmzDZ5kGw12AQb4B0Ln5o+m7lJN0G/voxK4bDP30GwoKz6YxbO8i3IZ2n8VMFoAVic9
8nDFhm2oBt795CQH9HpxZFL1E7lnP6eBSWAQ7xOtRKJfgoL1Oh8XahfXAs/3Knqg8BvB0ef3HqT9
yS9nKO4AvHE1Yn9t1pq2nuUMRJvO7tK9FVcLdq02COiYRV8zuWDlbh/D34MaF6USWY/VUBI1G9Mm
HqyJgorD+i0O4XvEFSNwEN0fv6Gdl3Vhr3t3v7D8KwnB6psg9KY/RfWUVFOGrEK24Nrm/zlhj2wr
YgDJ3pdAydsHRcwZ1N5gXYBYvJ3Qke2opLkgs4vo2gHBMlv3QEFX2RkJqASJFB3IM5qUXLDj1LX1
LWRsRm4/BHfx8JvlagHx0dFwqDV6mteuTbQRKG4uavzifSENOvk1zT++EZXVwInN5vMbRJfZCoS2
1Jnk+ToGuyeMtznc9BtgZl56iYcQ/34b6t2RFecp2f06dmw7PyLrK9rrqN97xsssrAeTBkkDoGnU
GFo2tl7fVgn4T7TQ/516mL1Oyu/lz8uwMF0/x9iFhaU/2VOwJ8lX4FBOB4R8ITF2kv63fJ55QYHq
O+V7J76UouPZjsPG16hh+KAAeTS2OVdyvmbsy840JmpzfzcbFlHw/nwEiuVQT6oW6p5gU9pY3KAc
XP4sycIZKLElrCsQL8pOp1rathC4D36sj7470+mOzwGZgFSDnU0ESNToWRhmA1BzQalmKtkpo7Kr
iXADfTTPD9NmTha20T3dl96pG6A2+kfQIlCZjzRcDMjNW5oozE1yySZzb4zDvGkoTBBaZKVhcCYJ
Zk1MYBQwS9FAqMa0gzjpxyLZiNsLdW4R6R4AvbIenJhc94k8fSkoW7LrRHd5tQo8ZKeqtP6ukBBq
oh/hjgaARrVgJzqVBp2/dETQdDsHTN00rLWeZeiJpvxYk2Bc5ZXrdswV4IfOtxuiPVCJXOUFp62G
PpFBUPbo5z10vAcOhbJFxNnvoi8+LIfY1uA9w/MIRoO4QWwYpnopKP9msdqgJ2NaatmV8F4zK2Dg
jXXF1yD7SR91NAJsYVbrg8/IKW0sMfsFP7qzCyn2Cs6oz8/yCRpKAy4ziYoja6G32mBxhHzBVj5T
jLhQnWxG4nIa0T25dZuiKH1Yh9s86CJ1WNSaUUp6/LBMxZkJcSITKiB5eodESoyqhGpY7n/Ci4B0
umsWM1tLN4IbS+DDxJodSjdODGo9eYYaqAzPa/HFQEUBLw0BFdVg7lV8iRR1kkA9bkFejpNqLcHE
0cxk4JT6bfdvD1WTpLtHVglGkYnbUZTSUQIxfSql35kCbAK/J/AwTlyKkMteckyfov1XJ061iOYl
5T6oKsoHUuCqdWHKlHg0j43wGUwFC7/B0YmBX6Jtcipjs5z6r+v5GjFY+gUEuRzjThoqnrXGuFt+
fcJsFvh+GHAJQp+0fG/sJ4gJ9+u7pPTKNxumlyHyYuv6kEXU1lIWUJ1yx5u0MAxaCb5q1MVPuUY1
TkiCBoTqxEvaVdkNPMYwWNmnRTRXQj4wmKXKVsd+/VgaFoV/UqupFaB/HyMeohw+Pf4CJiJ7aBcI
6JDwUXYl6+uhORI1mkxebDt1+86jSnzDUJQHQs7mrPClAH6Ximdt1lCx2oHIWv9elOvU1FHy7la7
v/tIKQpN/wUDv0lcGEE1w0O6+/ZjIxQ7l0qekQ+xaCMW4M+u8hE96bKum6H6xWNG+/MN6A8apyow
VnXNifIp+2fy+QdblY63quPhmxmrx5OHL0nMuCBeKCOb2m1BAELbeUOvMsTjdmrs2OVKAMYsq5nA
rxOVegHIcsIhtzc8O/xc1V88twqJMn4Sv+DUNxZZ35OAgCsM6WGhOP6xwFoKhZSl2o8Rq8wMQtan
h4qp8Pvx/pmJbmC5yOTGkzn3RGy4djPW0Tr58yBDImNStpmEnvAPsQeVXbfIh0Zfi1Wv9HNEzb+i
NwbBSOX9t8uAFyZXSYMuFQk5wPCTslL5qyaNyI1m+WzqBEDR4ZEGw7Z1Jy4fXLzmUPFePdcOXZUJ
NdUFISS3B5vODU4WFt1aoyTeW0puY0ZkXweFNg5sjyDEld59JlhUSWEeXxHaDjPf6oMVohwurcBu
epXyodk51MFyAay8uPNxDrHAkP6jjjodXiD/oflK4senwk5wsWMQNLbiPSSGBXttlqJK4B9jwoTa
KTWlsOtH0tylH0y0g7bzuCYqO1mzRVyY+94AmZcNuFH+YEOfR+5Ga78ld7/cs6AybfndaS21OdbZ
ui+A2CpfAcYUzJSG3Allxcsdp1iAxIq4LxFgQdO+jQ8UFAGMoyhWQeEpRpIESyO2cUmEkXEgfFyP
yS9sGlskCjVEq1Kb+aFuYvZFW2hOaFXSAi/ZOdlm2oDDKjlofOGbMPUOVB+tB2W64E0oygLoKNWh
AmvWkISO1gtKD7vEmb5xkCJuA5uSQAJgTI08HbAK9V8EX3qWuLED2bOdYr4pBNEWSieSiU2VMG/n
3EikbeHYyEf6j3/jEw8FRjYg2/Ob0niSz327/EIxxes3nA20bRT3xmDaYfAjIpxf8eiLV+6OKLZw
KVXwas/vhMzNYrC1o6fRa0IXJNt3LXDb9giSb2utaDA8ryq+LoHq31795+cq4mGTc7kUTaiDfHxS
qMo6opwm791Sf+8A6CiqLLe1cacSeb4JPfhYqYk4JMwTBuOx9lXKp63QdUhfifv5SKzof+Ghcb1J
dVi699gGVhP78fcCvpKldNPxuOB63Th163QEZPfKqs0MWci0o6SoLJn/fNB5i3FFd5VSv2Tttm0E
vPqYGcbyhu564rnFGNA01nwNG3Y9b67XhZMNylUmlmloLuP97Ghv31Xl1rzLGsq4UczYxWU5tIug
DQs2rLsdBgjnqrpsIgUGflj5rpqzFYrA7evOfT8ZmjpJcIbs1PG0I4SzTnk/xamibif3meYhb5QP
3OF5Rx2vAsSReOYWmWgeTL7YfqQI/wfbTybRyeFk7CEQ2jv0b4aXRXFOEVyznFdjPDplnR9DITlT
QXFlW8nsNP/1RFmuQfJFnikUBh5evYCiQZ+9tgh5D0/45Bhc/d7mf1UbZq8FnCUS9zT42tLunCWa
070lvxQEGAVvGogGnxbZ3rks5IgEAyYffjW7Z/M1C3Ci6B2Ah/II7KxXW4RlbSS35ZDZyGeiEsGs
ekAIXZCvtqk1A0Pn76B3poiTUwssTU4mxyOp1dU8OIElzIXLsxyqtGgvw8me50/3aDUAypEOSUr7
qV5B2DDAWzbZg4HTsIR385BoeUdHrKbjAHHkNY+Wd4WQi9F9jc2K4OZjdoDtDDQL0TZpTPyvFvyb
nsPSMVf8S6Qo25i+rgeRWAinmuwIQnDgBgBNO6/jk22DRk/INPAiRnh1GlU5BF35CyD1FBioQ0jr
uM2w6+71gwp9GMdANcLJjLzYtaw6sT3Dtsf2+bn0P+/pIITLaMm1AaI6Jd69ZxRawbdojshOKy1X
DCKyAUJ6aV23QWQbagO6wU6+8FDfFhhKRawwcBzhWJclR0orXaSp+CwAdLIZLMH3iAfkDBsSAaAg
siqdZmNaKCYMmyxBmaXW44daaVpJurdMdULzvgWj+CjD04SiWU/7IbOth0W/6WBSikRy0nECp8k9
rCgll2/S73yvfbENoN+r+Fhv81ym9/hqPqBwghHGlAixj1HwOQaoiIkXftLExQykkluNJVtSIwRh
J2eQ5F6hAWBQtwXVnZ/b3lwTZmrlbgYp9k6h0ucKFSFm0zVFbx0pX5zsDricDUVtl3lZnI92RpBE
GBp1gGtFKDFk3nh0o09XNG5PpowS+ziMPnJq8D1q5HkJr0B522BKcYlQr3J+8aPc3ZO3r5pZB2/O
49HytZktq0sBIEx6ALYAuFMQrExtKcgXY9Dw7O8xIkfnElbAQdzaKEDc6M8QSsA9J8L8IWkU3jBH
2YUqVDj7CECzDf12bdBaUtHeszZv9eiNq59IDdQbM/RsVlfFR9t391nAej2Hq0PedJzROwA4zp+w
bb8QetElhYPUgsAt4xIybTtEyP6rGC7hzP9TRhdoTmk2z9pOWzMBISm+m8clB7VqnJ+1mc5wBiVZ
u0xJLxRfn5OXIkJy7keDhfFzwbAgQi2FD7c0c0eC2f2FQEnXn5byvJTp6BXroXFsVqDqwInN34uQ
Dg0E1KGwcSFYgiGIT3yApLh1jmOp1QHRObiGUsLxTsoCKn3y0A+yY6QsGnyVkoXHk89KgHMemtU+
GDA/oV+/wKr8GllD/GJTIvRhAsrk7I7Sp8gnKBi9fMeCHKpI7urAnKla2qXbyB7Yw1fW0xvNQ/Ma
faG/H32m4P0Gly1nLrbua+ChRlOCsABNupfmu98mkaYr55cjFQEt98SB8cIxQitNhNxcuGivAnR+
6YWeVyM/ZABx/C4M0oAxBASVq0/MBwgJoiXB0GGT/cOnMlS9/WPapAw1dBuKWD3URq2NXZLkDBwT
9gnoPKUSWBsiUCfFHV1AJuwzC5fhFhVnaGQDtToqAKERYiZXfqkgHGnR6UX7EGWz+qdBSHhkRu/L
6D/aKYon2LgnZNTCWzA8N/ephUPyz+avrdzb4VN2K+8ZWYHa8lxShWLoC0wzAeHB5EvXuiiCRf8V
x7df6Gss9JeS8EjwPLJKoU8Zo5um3U1Nd5K0596xy8mLP6jQ3LbrxZHCzZekSadwnp1vGx861PcR
d0mq5elx2pMzCt89ySJksrXsAR0iYwhPK2NDeK/nM5hZuQ9KWprL19kRNDm859BB01FzhqDGv5pO
1ldagU7YMPSw/h9Hueio7/N0EdR22XxJz9JlwEwOuMDEj3Xj5NXMpZl6abCPrkLCIabkOpTBpPHD
aSORKNAtm3Du08d23MJIVIj8zTr5u4y1vXECmCwBFy0swFFp3+2ei+3ZSjP6Jno/5XmUCGiyDNFb
Dz+h8kMH8Oso/cprYksFsjlFuxLyWND3PFsze5I66llXbENmaIkVaTf7IxxIFHQjqK14HdIBLFdB
S39NA37D7kH3Jzk+Vhu04OIxI7JdyKzcYtS61smw/zMpFkmPIkFgiSp95zW4m8EO2ns9NEHmXQcY
ApEC8cTj8jp0J0pHIWa011RRtSxwy2c3A56/oaIahI5hyPfC6Sv/RsidpLzjSzF6EjX0FSv6bqMB
ek7D8IGwOMSKegqyU3KcSAOxYsRP+J6IEP2B7Tqnp9RF/uXvjY9b9C0XXw9FJyMPI0DTdUMrxAOv
DRcxOPnTNcOClC3CkDLFXxqYcaLAuMpHQHRYvhR04jShaNSR820Pv4sHkwB+KPIcIjXZkNCsRAsY
mOEbT1mQUQVBFOgRSLZraavnJNaFoOts2aE3/7mlTR2iiL3k39XySpAaEgNfwQi8n7MfVSjNj76r
tphnqX8S3L7im4qe7crOdOHIIfUFy5o3QYjwtm4TrrPKuC9uYNTv5P/zXEvP4j4bUS1Egogr8IA2
yI17/Q3xev7caHH55UqCNSb8Ewm/n1afPttYhGAG2BA6oytHiTSqhKKvE4UrFUbye0yCQ8+OP2b7
bMIS+FgVgkQr3fYAHXgQmWY7bajiay+V/dVI+DPduotPFb0vtFes/JmR6or3IGtlRWXhf+4Zeprt
zW08R7+oXp11hB+FVJC95HghwhQBAsO+ajSuBzJSIML+Ty5nbOXFd7rBaxrlnoJ5v3Cb/8Y5/utm
IjJO8gAzGFjDnZ5gUXjdKRhwmL3bxFUSngjax5HNx2J4DnaHpIhSEjFv3Xyf9u0iw2MMTHg0lAKF
3uiAYCeaLe3KJaVyndpazI1/jX4EBbbfnbGab17eN7sATj0biY3A9hyWPPhGLKqG2xQkWjMwsguI
XPsXqva++Es9OakjW9uS/8mdjjEvOlfeKCt+NBbOVCkFZ7E2BKiweJ2eQcim26GLrGRP4caANZyl
Wa8waJ4QJ6PXaEjr4YLR6dL5XiTJVLux3rT+Y4HHrOVQUN/tvvsmk3i3dSqzOTK0btVpnhomwg7s
kcXsy6e+5l4gsOsQ+W9TJcHqxz8o1QtRMBjcgkbB9VxDgYLikr4gFOcIbV6LFhYbuHqeh/ZSn5Zs
Ob7o/GeoCCxm8I9uWJ8sjk43NA5bujSt8OwB8uzOOOztMiP5cvMrEmIU7VgjtGcxCkM/lFqT4nOx
rkONwMfyoA5d+Kv4X7MJdCeY4PkIY7sR7ZCOFjFZ0Vw6y+afSd6ae718HrnzIKOVgFDNRQJHU1Lg
5vIOZiAsuZd2woyPuqHqW796x5/iinLXkwLlICcmAXJOWWC+LsXAT4CuWRrDC84QVAH0IHqleCDp
NoXHxfxR7Pib8gw+UnVjQZy7Rwq+OBARCarav9iSWkyFVNOVp59l0vvkPm2DRR7JBGsRKecUXXON
gTZOJy9QYFeJFnRdEtDvo/nlBrmdpKo2v6reci4+Y8SYQQrEkK7CQXkY2q5igDJfLk938j//ELpA
fBUsqH4TTpU0VTvjCYIJ68QvxSXAOs2JeJjuNV1yzr0NG1nJZfFVcdfq08H3zxFuHrNYyufurVYy
2ur8oF/E7uwr/xnSaeqwARqV8MFHvo4Avb3HAAl5ou3h1r3X7HGgjNZyiRNOm2TbMJ4fzWfl+t69
6tP/DdkVEB1n0/NcLrfTMS65B8q4T5FoNUp7g9FWfsRkRpycoA0qLayfpHAaIO0xa7LK7JFVSN3Q
tiNe/bPnZeJMEAjsrT2y5yK1avNMhwEb4I4hh4IJwo8qQxSkC18X0W2dgUYO4mkBzeucsvieAs2Z
1AmflkBiPvwHRuJ/tTAT5Jf6YrKup6f/VABW2Mx4l6hrRtwyW+NOgRIEvcCVR9YsYB0vStKse4Eb
asKBZz/XHq9KO1dvvbBD86UbfUey1DnbjG+SG+sct1Kv1liUo2PckIWv7f8yxxofWLL+xXkczvUq
nnWinTohPe80+5el8w3qua+vDS0CL0xftvI6aZ7ZROyNMoT2Zyf6YPbn2mq6o1CYv0ucG4fWEB1C
hwu0cOyoWnwIC9SYi7jpO4EZ1wj02yUgcn9ed7mEUFktq6Iz5aNh3MqwaHjDMOLRYzz9d0HSBRFC
ZRxfBajBGp1v5uqTAV1yEWFyA48dGtWrK3hjJCBqHreArQwPMqIjBxc+FiEkvo+leEMn38xAWA5r
JM1/foNUETpMpj0lEJzXZrOY3Yz3bE9Z2y2mw5EH1iin42xnpehhrDx+B3jJxFm7Z5wuUPEGakY2
ze7SJM2R0Ty0x5rWIe5dVTTuyhnUVW/J48QiSYETRWcvdFYMf5QgkHAsyiOkUtdSRSi8ANSeYLfI
8nt0yZreryxbeNKmAuPC4iR+R2tqaAVWpd49xYJPgmqXffD6YihoyCHXfGUPHJZ4ctqmEz8LNgFr
kr8F4EPI7kC41pQ+4zB+5yo/ncruwGAjLyYT04k3wVZMR6N4FdSmJgyPOJ+SVBvIt8nmiuZ70non
uFdrxsb9ZgAM3PKJI76LKGouOF82iHHTmTOsO4DAcTrIain4bVVkKf4p9RToV8wgEAY2iL9NlX4M
ci4R5+jpYwLd1UdbP9nTJzwd05LN05OTv23/ngGk5pH2DjcVP69cQbTuJ7OUP0VKLQ0F5HPEo9bG
97GXvz86Edi5Ib01JHJOvrZP4LSOgr9y4235evbxd1+JIfyo0rRwkgZRewXJHpK2LBfbi5RcOukL
ejTRgErr/yxHcIMgRgu1zjQEpaH7C1ULXS18RL98GBSQ8OWjPDGfmhR2K4nNa+i/xUTaFZYiJvRK
CG9TvHYIdEA5l3Q2K/b9rbaV9fAYXb/SESc2FhllZWtKWa2w313Pf9oNSU89UamUvP0bHu1wE1ep
NniBjYjB+hJ8cBvv0FXefAy3QHiabUh3HqdGntJhfb8u6r9AIjP/Q3Vhf2Z945Lf1SMKuOrkxiEi
YW2/nnRZ8QMcrDZ/jCf2WhQ1jRojpETOON8G0oZDwY9m/01T5mUSLLpdpzU+Gqb9hHUJEZo5dBLU
ymHnni1AvRgtqxXKI5x/R71dc0BHI/d+Pcgd0SqRzkxep7fh5Y3y5XnRcq+9tLq3QaIPEQbKSToZ
h7rpR7xMlqqATDqNRo7a0qcbUCNwAiO/+x2xRtAybhIZLro6f/Uq1J4v8vo8eD3myRyyWJ0qrqQa
xvIyZjcG0pXFKORVeYk3eKKJUMkMeybSgUZXaPlQySM5rQhUO2enPD23OPaOZXgDM12x9uTUHIkg
YMfj6Zxc2IFGA6KgPLh2PLjDKFouSJ11L/rAo7q9iR3JClhDSTNVOFT8fLos9RMNKIxF6bQpiqZS
Ogun2FlkYUjxp0R1BnEy7Mky55XbPJsYndka+mKldgfV9VVQXPTwBGLKWDKvOlWFxu1UA+kEpmDd
u5rG+EuTjG6mNUZMRFT9DZ07tRow+Quw27ynt6NAe2zBa4Vi3syM/KpCaWhAeMZ8UvvvJRpRKMiw
B8Hr5jTQWJiCMjUo0FHPUO2bsG3+Wdtq7r9rVKMa8Uvu57rqwQTG2fMoI7+UU7UM8ud8gXlty1sw
OTrSPaJ33HKI4y1n8jRf76v4/o4cEE6b9/9lLKpGlqW8DpX/WJNcbYKde44SxHbUTIv4WcsMgsmT
2nJMHQYAMKWN6yntXALBiqiJtvJjOPyS/GTtxWpMBwpD6A25V57W/+eEq/pND/kkhfopfKzp4XnS
UIFYNDCr/XNL1b2qnqi/m30uMUBC6L1ywf71IAfrGqEeIDUSzqfa/3b1Ie8Mhj/7Bouh0oZyDk/I
M09VVuFRdvovXS91Qu2NiprBmcmPF9mjoGa/B811cTh2nb4cWR9ZpVW4WQGpiCQN2Yhpt+OD1q9Q
1khM0NUkIpZ2kBJlzg3ZYw7b1hTxJ+OcQ8R27dKVUdFwjJknQWjrGffzPO+1MY2zRjflJdrE8XFT
jNElCn7zwIzrnfynNnoe41/LN0TpmUYPZoMkO67Tj5zC/hN8gu39ic1XS42aYaQIyCMoThf4TSqS
2zqNyNzlFRfl3uySXyVqML7CugodJuuzJb7B8/TjVYV32HFsoQ+mUb28UH9kTCnxevO3N+hqCMCu
ZF8UdXau4x2wHJtScXOKEVjzieKiYwuxyQcBYe3S0rnp0TsDof0uQrlb1lVISwaLutzHgasWxFeN
XWGEw97QpU7avs6SHj0WFik7PoDgVS/wpjj0lWR5gpztlJLMDSEhKYhuuiWNrT/wxueXxrQdTwb/
4JA2RHmZDtnqD4LeFWQnfVoVa5OreceE2bMyzDqM9kIAPlvoat52G8Tv/pZZ6X+7+thii7s/YBIK
2b6ZGiJp0tBAjPxFDtMVlc3v/RCKVmneo4tDHPHJMHm7ouJQmySucT9htUOiF7shXUsznUmWu8LS
YGvmNoltsV4CpTBvRKijZh7MRoXsko+zcFfnwKTh87ElTX9/304K1grNQoZoLivO77e89yOgHoiz
mv1CZpDSsYV9HPQqAU6BUY+5FjYY2vEsFRmv7JfUBSVrDSS8wJCzPbpBXikUfe1b/eyou4TOglAA
/OpxcvOpQMhFNxJ2iC7NRplvWAMuzj4VP7NMHVuLFC5qyP0Q1At/3bY5f4U2Sn4Xmzrdrc5Gr60a
q9yiwr0z5eluzwnPi3+6aOGkY0kLfrYjcHyd4ljZ3/3IH6NRBmxzDwfXt5goHdUoHS/tkbpVKBCa
exHORLa7Hk5SHDlNqs3L5fMDPQz/J9WkYX8jZNtMZs4OF6kGwWZAxCqP/tqToHrQJvLiSeoK/iMb
Bi2MOmVjF95GFKSgtfDAzYDvfDYQWbeSCX21Id8o4DHCmkJVXHfI4HwDhC/0ggakouElSGOtfhLz
1KLhGQzSWm6KrSQTiPfDouneAbV+qTc0MuY6J3V1jsjrD0hA2d2rGbj0OZIDzF2Ipi9VizwRMGHC
2puMExbsi0lQ2SD4tl/hiqvdagifxFARCo+c3iIqu5XYuo/2sEI58rmYyYkSmEjXnOdaeX2jba8f
Up3pzl5Z8GfFo3A+REbZtLB3hTWjm9lMB8ZQJWdoKW3tNJBtnPOHpeBRnOA2zOyktBixxTNm+OtP
rzqINRLv8YR2nlWC3w/s9MjB8d0gkQAbO7onKjH+TFH75w0HYd9S3SrAmp/VDWHalYImZlbqvVsA
7OQGNdR7Vz0UcqWxJ/OgMt7fsLB2DSsNxygbYvoz/Rvj9yZTbF58tMhbBy+fRYU4SFhIrhMG+DW5
lpsGXaBmnobLoJCbWRQspKnvQV5RevdaYbKkjYBZrQUjRkJps7cuwySWoqZzsEkp46OARDttY5HE
UvQ26ln8/S/NaoqZw1efIsGrLufodgSaNZgbf2OKu1CMxnWW5Mg88Am/jW+IYnePUwnJeRy6k65R
fiZ1hNyPpODxxpFClDtw3OqEM0g9pQwP7Y8i1GpFY072RCZ7SZs5TU10uwNfIRnMLw5AsXlod+SP
qyw9NC0yyYWXHHzX/Wsy7C+QyC11XIP3GomaKnZM41ewvCTf6JwWtNa3+wAwV5jbJS07txKnSFTd
sj2/Gjur8vLhyy+8n5vd2kKeNsJmayPEOA70QO+uxktQm/LSMVid3jnN9voVzSlnl2F8t2OfO614
QFCmGWQCAV4hvSToaJePwv8iDieUYvym8/PwLbNKl3FD1n5PaN5Txh+fpa0rR/JDw4V0Bmh5vN7B
LwvmcxKfwW13S4ojVm0xu0UePlMvXtF1lmdhMGUKiImnNOgHTqM+dIBYqQM7g5RyRQugaI+HrSO6
4zeLPo6j+ezu/r/bIOFekhr02own3NeK9qCA/RRHVP9vEc4QOfnAIwraR2fhSKv5xoTyQo0LQE4n
1rKMJ5EJ7qJzh1WJtF+z8vFyiBHQeHZPBW0fJHC2M++7Xvyotw2Ntj+0LtZ0aO0hCUYYpW5BjglT
xu0X5JXOrsZq/Bch8fbQ9d8w7NYYTWGZCHshwBnhNyj0s7ruN8/s0KWo37dHtLwyZOU7BGbm7ow2
TWxJeVNLpj4ussftdxD6941/KTZpSkjhM449q9jfTMx98fxWIuj9PKv4y5sZvCdLP3a4UxGRnwOB
cmNwhMZCm4FghHaIcAvPMerP4PoPXe5lg9THGmCP9/kHY1eC69VXx905p0ID1sM3s9M6zX9exsjp
2QWst9/JUdK5KXWzPVFvwENPQgPf83qN9RFRN4xwDet/qZpLZhimzO3S+fM7OIg3k9if82UA5paW
HTwyNK+lAw19kTDgf4a4QHiqE/3STVLUqj4wpA/thEodS7fwPSVNdJUBQ+yk4HgpQ7k6wpliz0IL
pfH9x29BZobNpZu/rDQT5d/CRXZuWKYGyogProCX90wE3jdifx8M7XghZCa7bQ45plUM0LEUCW0r
epAUgLBKBQRPlu0Y49ySywKg2cL056JPhJYlwBclu/regdSDDcI0eM9/RZFfMDBKTAatoLQSqEgg
AE58NE6gS+IhUuW3X90t9t4n9OBwpFOct70ZLQ51O5HU6yG1F0YpU18JtM+B/sXZu3Xjbl3/6nLD
RvOvNKQHse8Y7AT0oBCzefwwfL7tCsdpmCsO9mNxop/3nUGt2PaQI+MzI/eBAivk+OruH1Aw+ql/
Ttin+NIhP1dkOZU6vHckoht390yUnGFLnnwT/FXw2RsOADKGgY6fNK+kd7560DQnSVK2zKejAUXz
1+6XFvVO8Bz9KPd6zJpk+8pHPZQhoPcHdyZ304IBn8PuY4s200Rl7lvfrVRpC2wQHrdPwqsAeuPl
xWcAHrNB+RibdO9nKp9khh8JwH2H2fVTg4yV6eEJVq2kiEZrtLyKcYDBO8uVN0A4hzVPgIEKR/+O
aXjL8/q6MjYO2xeMDMEcSNs7pGKa0EnMlwcS3DXZQFraEZQpamr6eOPd6gyrrR07mbNsDSWPQJhS
cN4MFmy/uVQDJJC9Nh1NjGbM/DPOYKQ9EWh8N9FpLUVY5+e7/yrbbP04FnFk4D18BUtIh8JBHoc2
YUX6M+zuXQWKqHQt3cP2nlaC9mj4zMGUOO6q4PkG4dfX6ZMOdy8uXpNzg55ciOblZvuE3KJb9c+O
ub+Wmow0XNs3ofyX3yS2MtdbQXL8a5Wdg6BGWYTU2SnaDpWdSXs2f6BQHxMfJx22J8PnqBpF4EHb
PwwWdmMStWUL4y7dRBmkXGpfrCHZKZGvgs2bNYzPrgV4P8lSjV6ftZqFBfhyrrqCCxckU4OyOHMm
gMGKEETRrVvsLjtAyiKN9b+Iwj1lKEZC4Od8JoGnQHFKnnEWTjl+RvsR6uzPsipSY2x/fKTPqS9x
hra7997L9r8DMHOQD/Sih4E5m0DOEutReESLFlvuHb8lyca8yosXchizIAQmaqnHKSDowo2x05z/
D/Kol5AQ1bMMh8w8hqjsg1hcC/XgMnlm4FymW3taNE2YubGsZNCjBVanVWCvqUPIWduHr1UCOfuI
jHUCUPjEQ9c65tPWv3NJOofdRXGIRGB4tl8X3ZBb8yZmN4cluQuTlgeZ7PAqz9Y1UiGFXbPxkAAj
uhcx3iU8qI9c2MwX8ujMLoN/WV/WQN71kIsFYRaYV8gzhD6KGFyJc4CtbuGVuXqgC/XMmJTC236h
M06J6gaWwRAGG7H85fgDkQxZBPTPsm8a17NgeV/V/ueBDMGtnoku7/MQLkXVsqzlAZij7OCinz4j
0bkgnlWwIqM9TFy5oHaFyL0gEi+e8w4iiyvwxkP7a0JPWxGNe30CuRpVocYRzJQhJXlMTdfuGGLM
WBvuuVPFHTOAxlRuauoWXJGaevJZUXD+NFhFLHu4iSN8xsiMsnG4XsOKxlSGjqTHuD2fuudy3rxy
iD5oV77juXeO1mhdJMVtL4nKpMUX1jwS0W+DPZRwDt+hYqMshfU+8rAPvk/xJVWfmUZTpMdJjG4X
KKfaXsH+s9ZEHHzFcRNOTQZfeApwb1OkMbW384lrMMoQUHGjmeVUWFwdRugsctJV10l12xVYa3BK
N7x1FOQUDl4/UDj8w8pRqOJuYiV3G3AiM0wnO8mOr1rQNlFMfarwv5MmFPJHz/lWHKk7xA6iGi3l
mVS5Tpus6brZYbqc7XB7fb+FeujfxrBngh4H0JKFyR536zn2uHSnq1Of07g9Ud8ZJ13nhJs79mBo
2fATrMAx3QA0jrM+U4T1XADkjQmFu3aKO/mMU6LTEVMjzQpiMI5wH9gkTmghX3OnuBuZwid8mb3d
xK+teLIBfWI3T5Gm2YyhMLU2Gm/Rz+Cvi12AU12ap6Mb97aW/3yW7M6a1TcIT1CDHiI1oM8lZYsE
Kt+PKTP+1f+uPeLA6j/0T10thiltjC2w//j6egLIZDLL51W1kDNvcIDRL/e+Qp0U2eSh4QbQ2FOW
7dg8M8dd+eFEI/+r+NV2oucGzQtBv3FKXcZdn7NIQV0TXbIn+fKaleas9XALozPqDoO68FQ0eczK
Cc8VbX+j6HewRTXlLneY794wwCYPA1n3o4SfEHSq3xAPUAgpRanT04cE40PNWOGeEomPnGgK+9FC
pbusxLiym4QeGdKvYy9D5zMXGOmZettgHWKpOKg9MG/5ckteNTaGc7VV87uZr3uTq0ldzCkpSpfT
b76/AZh7jrx6INqlJIuRdiEkP8zM6LncDG8TWLlfTWpwEY2kLT1XcarnPH9tl1fZAMglzgssPfxR
XCW5NCqmEctR0icziTJJpspvU6Wsg8Uj5DAQPIT82uDoLZaEKLP7lu5UgVgyCssRR7sw84FMxbYy
KQuGgar5ACTyN2rLDN6rmg9aJM6HTBQuSYsw1gzTaWAwYOzjHWtZkJbv4A9sd8AnASGckd8YAh4i
Tg6qRwZL3tDO//I0xy1B514P7W2qgm3z4tqXVHlRcCZanZLVBosRKLsqGDJ3veIL/s7h45slcaa1
u9hvml6mTTpT+Q/0TI1YjSkHX2ENcPJRolzqpIW8TDiEFne78fjEj742dT7emJB6naNhMWoGwYAg
4xvi4ZRYMYqCmIBaCXrt5wWxqcO7S2b2Obw+zHb8Jdc63eSfvLPQjf5SS4y1fZE/PzR/OIAN4jVA
ZSgAGaZ2aBe1u1I62/KLv1BrpLpis/TEONrrT6bZGAAsYeO6GxrmP5XMAXWAb6GAM1fNl5w06d5I
nxh5e5i4jRb7JyHCdERdiILAQTbYqtEFqc9F3HMzU4S75kbWy27QMF55oPkfmst3XhcgJWTTJbBC
frMkM3+XAcXdBxkDDgjPeYflExN9P/GdPabepyix3q3ws8tziUKQQd+xkgLVrCau4E0PuSBCOdnr
GVcrnV7K6OQXWknMeccGpUbz1AKcM3Z9CmPAnCQhRKYtm2JmdYAgUBtGIQApIdv3uyddkkxhv4JX
xUyQGTCXF1mruwLy+L4CJGaTtMTBncTMN5I/zY+qem7zzzTP7TqTkUD4PtJ/nWm2CY4R3wr4mAMy
GZfj4kFnkigZ6zpnsGzllcalAW+COi33ffeQWZp+lo1wWGkhaEBcKjErRUFVXVzVZgR7Am+Fa2nP
q1Sh9q6aycBhihOgv559EX30BYhixsH/C0jMS0TXs9XzBw0+aSmk0G0PBzyCg3ppNmNQBKyeLRtN
LixjNvQcBO+h3FB+WrxDEu+eVL9Q9V/n/c9TYiTOAhcgEbUn+YetKPftN2NrDDeOT2LAfA8/X03f
o/wEQabFtqAJHgWuFZxf3+EsECI6FcTwtpYdC70pkCRRVRXQjmnjdoOlDkhqTWzq3OHVaVARm0GZ
JCai6PM3THEXcSSYuPwmAQVNXK1+VNGCU1mz9Owp/EhDAeF4isz4RW7YpF0jEfIwjVHHIj95eg31
cKZheFRwKBW+qzzuVdjVpv3kmqNWYZP7pzo1uyuNeSWNSqGHcvW0zBAsijpdLni+P80crXUXFut+
AH1v/QxcLMhbpKWpmnCsORKS4vtPMcYYxekfpxUdXAidSsRLDsarbAaPv4EKb8AyPhm5RnMfjXEt
uZ6u/m+H0jhgfMSUjuXv0QBtfIuQyDZYzF9tv/60pf96QcVc0q3QNhdSWOfoqndlqZk8/b9Ojjey
o1vF99mdbRj+qksKmFnHM5hPPP2CG8EFUvz8li6jbu3ZGNLhP5V8IKON6DZiZfc+f4ixVLWq/mro
qEJjI0Pbv4xp4QmVmrmWY1g4Atxw9zjH6FAH0f49EnHMA0XdyR8RJKlfx4IkKI3bCovkX0w59Bb8
hV3GJu66bLCy4H76vTfUTmUmYzpov1u3F4gnPVicT0E95RhpwGJiWE9OXS57KhHp2I/nMJNG5+A7
reKje2XwW6oep0LpOND23CKAHPXtIUQqe/QXMufsPgK68+KxAl0MFeHIO/HDAVaW9uloFOGOtKQS
+hhUExSEOIFJePQhMJwG+++DL78zdaJNYn+sziYKbWmg6vhlHWR23Nys8AMS6+/WJ8gMJa6Vcasf
uvGtl01GQQnGBh8XBG1slCX8VfhGoe8+QlCn+2i5BtJyCx02dPFIRztZ/1I/YaqGO8AlKr9WMtGX
HEMYpab4+t05E4JcfU8Y4CSMOaRR1T3QhhrsBN5Nb7g1UAQ9C19WIys8Q2Vl+b8W94K+IYMIVajP
hHghKoCprcXKBmSAlKBGyswzG0CirANKfkU1OOtJdY6a971I3atF/2OSKqCbH9P+wjpDxvkbS+am
ABPAQFmmhbYnn/190wP8Z6xu6Y6Fw3Wpuxocd9TwIlIFhhtmDS5Ddkqh1Scn4bJQ7aTbmdlG7Gaa
im0K5M25s3mSkG6KMgSOPuH4Dj8Y+LxAy0AzJcqW+84BJhu51+pz1eWGm7EjQmtrt0tw8hw0S0qO
8uIX1OBMcgOuTsft7LCDScK+yUcrcWdwPKfUBd/gfcuv5qdgp1RG5v+Q2oEdQ2t13rrBB7vs1svo
N7Cn/P7S67V0D8zXPi6NbOenkL1xfggmfOxcht53v0WQG7IsC2HypwPFG+yaN/46zk43raohyzbc
RG6yREBZvbTnhIxuThzmb1LWErS4hTuYx3lGhxg8GVl/Sf4a+Dol41Y4KilmASdoSnTUA1gWOV8x
zMvso6P/PB4tFpbxX3unEHHO4INy8wiVoYQvGSKv0mLZd6WiimIJoX8xsSyumCJDQQ0uBGqV2qJB
pGqhfcU0zsuzjHFzK+4e946ldmIJI5N5oJhFWMzVnD+TykEzh9kFXm9PlcIoSOTa/HW0yZSexV8N
t/g3jDlx2ljhVF2VVA/X3S+mVKcGKFyvK2VejQC3zvs7nZm9kpBvAU3qcSSr+uX/5U8wRcP9v599
UdWe6C24uXFvTQBGTVPELhDrOHrQcFzRkRIkM5RjDOyC1uyF7O1JBYnnW9xmtoAe8n4hNJDnPdml
o9EW/4FF6GgSuQ5Sim0CJB1uKQDxYYCxJmmL+4Mgod10obanqiTrBHVnAXtVGCRuPO4LgCShEVbz
O6Sf7Iw4LfY/8vP+5DzLKd7sVeT4xA8cUtCIaodC6BWb7GvNXnqtvml+0GzHrOigXLA1McQ+vWAg
vSvtiFpTRNemFGT1xo/cJugVK605s2Mri14fTXI6OO2SsFXylZMhCA0jrjuQ8vWWT/vZNJWy3u2V
N/7YwJK05vJf1wzaai3Xasb0Jb5blLxeNLXX9MWar2v7gASbxW4128DdpXANIwZswMxEMyfcQj3w
yeD54UY8wkF79kA0XqNB/qLZcbvZ2g6iLbGtaQZtR3xRrGzbeKdJDwf7jDBUaD061jGmCglbZB9r
Rg12Q5GUeXlZzEYyh8S1L4GFuirVCQkvQjOy0ha4F/Klw+jPNbGDXgMAMoH+Mi7yyigxj9vBSPKl
WjkX7HiF7h4yqmRQijFhD/bCh6l7pxShZiLKUcpOijwMaY0jjkHTvHP/EJtmyovCP4c7ZNZ3j1JD
hPc1w+hmlbwZGEO25iMo63i0EFWW4DPqQGiKhWMAQICJ8If/iDuFFf8MwX5NBUmaM7P9HXaoTnv3
gg9YSrv+R2/KYEYRTNbX/uNW/5g5XRZiDwLwrL3WS26daJAW5aSGRJCseN3xVTb7NWX9phLXabc3
SqxjQK2fk2s4vx36BLsEftTSfN4FGabgC8MppCDLaP2nER9B7UYi4U9B7tKJ67VhyUnNIa2AdcLd
xQR+R5PHHMCZJUbI5ORmqKvTCarkZbwB+IU4bTUj5SF4VqQ0jR9DkTDWcZzp5mV92suszEJ0rDmI
koZgIV1FssXW1GmK1jO948xstFl/isyIdKfc1Pnp6BKHzV8/uyV4Yv5Ad05kT4VpTB6t36QCZdMN
Mvhr50iv2+9MZi4Ay0lTgDF5tkflf8yEj6zs/BDPFYJuRNt4i88XjYHMrHJinjFcPftqmekMPT21
5ZQcql9KCQmX3RcjWCr+UZbzo5OHnfV91Fkt8zUss+vHoNkRNOkzaPzntf7nAuOo0Mr5CdqGbje+
LluAkMl+6rf2B9UBgTlicZb66rZmgQDY4wU3Xnnb0JjpW3DZXGMX6+fhVYl59cY9DafKTNYUCcax
CmWFlnncclztNQnL0Ct0RLh/IlyhARw6Lf0KtDayFgV8P9aMlLMe3eXpYKcgVArXvxeVNg10dUSP
uAeTgHMPweFzfC0pQqG9XaDPT/Wv6+Lgu+wGDTtdCxw3IlsTMKiNfKrY9SDKsQpJ68mYybEUGIUd
2X65jPNfPeWkpFxWmvDk7d9Krt4BJj+CQh3VABKpWr3jceVLxt8qFiLq4UdB4POKZRVi4BwAt9CZ
b+l2gbPMYp67bG40uR2jYq8NeFs2lAHcWlzjPitJoVGFj3VrLXSFuhJofCKwsuHc+pMo0v9Gt6kA
9bYHDAKBz5GBE9AQw+DY0TnPoGEcsY58Zj7PTW2C8KhINpK0gI7v4uAHbOCqOiYtBpIDDyrROAQh
ufBeQljMvEYd92xiEf7qwJacCeTvhnLrmbbxEHO58e5uL8NAR+Uo7CDfp+RFL98/IuqzUll2SulX
KqQpzWsL3lSpib3lgRoDrCtz1vBoLM/CL0FsGXGjsT/oFcJGUcbSYq5S1YfvEWmQs70bB81qpNsI
tWYDcNf+v7Pte0zBWJJuLgyhuNIctVshv1MDJXmYrCBRQE0n+mUfXVbJW9OOzuBT4zG1gLivdWpl
DC1Ewzq9eLvERH+et5iCbui/A1e21m6d5E9NtBukaB7CTkAmJ9vFoX8qTP7iWoFlBLg6BfP5pJL/
a/K2A7ONhM/1i3jwOKL6N2xzh22chj30cmH7kmU7C6HFr+RtYtjlmib24nGP/zUU1AFUOEtnAnkt
o4b9PNnEvtXY7r7tQ7RT6j2rHVMI0IYHJMUmKvWnVWQ4My0BIrivPg/qGja7Dp8EmfpeswlqtTSl
9J2bq2OT1ao2ySFehlFonXGO+7hWFfFPGDm3ywT1D4LKNQvbwDEa/WPO51sVqtiYKnFn2/Onld2j
48w8ILOrBHDEfJn6JOMEPeT/cN4AGGxwDIbHSxYnEJkgAspJYztaFFsGqLn2CXcVV4XQnyyQDSFE
KT5dPr1E/XZw9S8WxiptPMmDPpvO9B3dEvjfkNRk+kJ0TsDhqV3YBHSzOS2XUSiUuZ4kW4MLTdWf
tMyJVzh4Y1xqGGpW4okMNKohrcoQzFROFsHU6ol2svfagnjB47bcsQNuvTZGRW7f6skbF0KXF/Xo
ZnOmZ92PbSjWuuDoxDEt/OUgn/ZvCGGYx56X4FHSqcsd67hvakUM53uPFmqEZvqJCxFZAzUAYcCT
K/nw5dZXpjGgznq+fpC2VQFWIk3nddwrIU4SjqZQC3vjQNG2X3Jx5nn5IRKimVQNwO9+n0Us3DHW
WQy/JACdmtxxc+ZJeNQQy91JMcCix5LALbta/nRMVAIF5ncqXZvf7pgxAhCzn6WlMec4YXiMQOGN
D5A0kAwYCL01QhxByjp4YVooS9K9qPJdZRQUYrD6dUr40tLb9szXtgVbRk3/MWhcwcgnCdDbZKaR
YhD0lQ/+0XwvekPBYc6N8AGjL4xQZvvcTaoo5qvZW0zO158BaEHWwhoT8iuVV2DiNcmeJS0ufkPd
R34qviotam1GeuZ4zpDcuggfOTvHepiOWOzloiSMV4cvstg4KFqPQk6wkJU0heXfUXuEcHwnHIgI
VQyfblXOcxgEdMy8KRkfQzrAM2oR9imVxCseFizCCYfsPr50x56bt67e7JHbLt4DnBVNCsn6rTiS
ZZIIssjD3L+yCjOANUNMtAwS6KPdgaWp/0fnUSo0lhQ4J9ZwRb+VQWRTP56FWMwahGHK206Egvm3
Z1ZW8y/YLw16XC5fX+OSDOG/OKGK+0MaRY7GUDX6UNiUQ7wkbJDWWKhnRfnnoaj6Xmn+TikQlfPJ
8dwVMLJ8Xq/n8O98M+MnnmP+isArmm/KfcBC4Qoqo0GL9UVNxLu8UEe2iRhVCc2Z1HEkFTd84RoA
f0wBMAhFTnRgNi1sewoMMLgyP2Cg23mjWO4nsHnSZRMK9vrhMWM7t4W3wWGEwBuyFKedkb2gpAUF
4M3Ya0SeKemTWvhRqexE2ZdTS9sm0d1pXLclWZw34FhOAYJImiI3hnOeuimO6g2CAEORPEN8//ND
OUMMTY9NpKz8bKyH7jpFxHKk0mAYXTI2YPGYPndfIps3VTnRp3lX67PGZSNBLPKIihE2mzC+EU8y
RhX8X2FUZwIgea5BDqCPqvcFJymBiYd2yjWAfACAvnmAqaC5pT4mX2ZOvfG8kNfWmN+qpCJvwXg1
U+ohj9LIZqj6OHWGVrF/7OiZgBXKgdyMW9F67DeLOSwM/KZwPw3Hhz7MmqLoADhXYWcT4ivE2Fbo
e6qz10F8zDTWfttdn6LoaCGNb/eN441mk/wG/y6P6SlP/A/QMQZSv7/823z2XdvtRU8usHw/GphN
F9ud/Qr/ij9g92B6N0GkSFxhXyPtmI/PwkMjWKtXKMTxlNdCJbGbc3wd8Nuo6GAYdqka582lv+yp
BgKuQp3nAjMriyRolOkKL1Y6EHppeRkDN8z19EHiHCvhh6F1sIHLw0pW6vlp9FHWnvzKA8ah7r2k
gL/Bg9BUDQt8Rwg3OGDCYPnHPcRiTA0zjF0tu1+pN4hMqjymndI/j8UwKCebqwgoBLjPb4YFp5Qo
MDC/JOTeB86jsT9cF6t+y+ec+iOfvQUKpNHtaFlqLI+rbtjihYfR9RA9cqZrnUxNUFswH9CjqvAR
uvij+Cw/XLYp6dqrVOvwBdoIq5QwN8u5BJnq6kIP54U/pEknyOPGIXjo5P6pOF9gDj5fHuctHjMd
mMc9ey1Rn/7AMYUyiR/zHvOk5TNADY66EQ8JRpuxkM8bSMuKNFxj4kC6yi+6PDQBhsP3/P3hjQCH
cx6cI4m0dGcxIjQin+BqgsWR1TShiurlH8AxagcXXxA/1HBZCHg8EB1IP5vybPA/b8eAk0cj/2bL
1r5L1e1sH9qneR4iSxuPDBImgQFnTN26z++ghCmjaYYs0++xhFLduuZ4MazP78jURg/1OgfwJaVn
s2qcUoYiM6E+SfnxOzc5vXnAgU/x9E91RC7okVocGo6SMsiY3QNhayP1Wgxt8NmXdSIJvkfvangb
LtJkAZ+sOcEQycfL0T4NFRhlWh3lJxNNAfp2xwAo5/iW7ZOhTO+vdTgKTOLdHOFAWRSXLiHPLob5
MwbYA81c9SzaN6Yp7UGhaLNStIQ34U2PzEKgsNw29CJadrUgxrZB+5JCvZ3Ns5P+mSN5IF4SUOBz
H50VAamJJxYk5HKoKfL3sdb7dD3MmjAissLa7+emyDkFobsYCmgICakKQqQ/eZtm78J4f3fmOw4q
huzzFxLu2in/EOottqQEC7+CgavIg5zpjJjD7SbgjqU9ey8I7TLoklQTTGpgEwRIM+ATB2PWcvSb
aM89miNzY+kHwYc+pooZjTLn23DbEfA6zZwHp4DMrLrKO8AmvX9y/Dmx9VjDpMEBSIeKTpwIctP7
GcEf5jKPeG0WkcTbfU0ylJ4PsTGv9nh6xodpFHQvVtPVBFzxho7ftFQlkXxAdYxxB7RnIRDSPOSO
nwPVAarN0IUDDShsfN/oqbAJm8BTrBwGe4O9Yko+GFcmXUYjYwyXKASovdibVgOJoaod6bR+h47T
JJLHdgtPD3oV20sHKVE8WNJ1N4Fp/v6ZuxuH9mC0WlPFOboAXqvvTMb9kJmJa4HHXHKLS5+M5OfX
BD4dbW/Ym47eyP5eFM8Vev6PdA3KJS/+A5/d+HsPBdH4o5TAqTJYfdq2cVzol7tElJrhXh85iqkm
e/5Gxb//S0n2GGXYJjVjj4OWqpFjxXbMSOEzF9zdlMTAT9QtCGS0xsr9F64hhYYUwlX7DZlNa0RY
1Xu7r2MQozyHyd029YYddXC4ce3BUPEsjPVvYRu8eQGwx/+ZN/L1+lJgKGrTfd32KQqSmXIiNHy9
55IBkx9E/BByoGr/g5x4R84QhoVaPl4b5wcOJ3c/Q7sKIuMcS3CPabqEp/jDRBdgV7DlIc1/ndyK
jDHa/soaY5CpTWdBNjtf3mEwJGkOhgR0lxhLz7DfClWlcfnuEfWnzEyXuWBhdpQfPtJPooa8G53R
5hbEo6g46fYUhmJKie/51NY0ZnF5oxCiICqcC6BXKc/IV70//k8TFUmDuZ91FjWmT4JL88q1TwhH
f9TrUqkvatap0ApaqI/+yh2Q3AwgrcympQQQKdbuiLjvP1Tfxllr9rsppHg4Cp9ncRrVEyqIvoC1
3n3cY1hVPvMQAu3kn+DN4esdpC/Mb+vk9X7IhQSTOD+HDHFCeJjiO2u9wzYG7oH6SWSBqQ5G6vWO
jQNNFDWLBI2z2+6J3/KNDFAE8YTKJ9f7m3qQg24/XduoROTEOFuzliPNiKFl8EzDBP/f9xTQnxOW
F1y5P5g2rWLLICurGH9DR04y6je2pgzJGNiqjjLdpJO1y48f7R/7jZQEMmYxp7qhAr3lJAKCyobt
3RIvD5IawxfYTFXEh0MpvFWtC58xGevsLk635eqv7QaOZabwGJhfPDcg6HC1SUMxZggULgn7kDdh
/hFURdSwwSOnJHRqwHDupE3v2bo2CJkqbtRRGsVQUBiwwGFVsOESIccZeQM4ICK0jQ9BtvCn7q3M
UjT0CgNG8UiDIvBJ3zD98Bo9qO50InnI6A70Yy2K6MeWnMTZySNEACo5u0hgOJaW+j2U439H/pVM
o5KVSkGHN5ZALx/yo6u2gBrvmB8HCaTwllqyvn96mAgbUtEPgr795ljMFuxLxOOzVR1TLTQ2enId
hLvWQSlnWOrXKUUkiTc/K1sc0eCEwWb+YxMct6Cw3nJdDDNdlCdO8dowUQsHdOBvhwk8EoAdsuKL
vxx6rY3DJdbhPklpW8mVBvVL6TgE8OQbWlCvEhclB5fc4IpcC/dxCc230rnBeQXo2t3rYe6o30L3
m8wNVxTRaiewd0TR9X6YqzgdQz4o4X/ICUYxgyo3ZIpFzOEg5RC9XLETRRe7KQWAV3qCW2FmJ/Z9
KA8p7sGD2PUquRUGkHx63VDlEbczSGLjLMlxqv4llF7uRNyumI+J+wMpSpkLqNaYsT1tE/gCs/if
gE/7ZlY2u3qEyIjcYyTUewA9RR6TrF0sZ8OKfqI3vtrHYp3a2ctlJ14St7WAnh3HXrXr0Fpkc0oO
1nDMPiBKdSO5g9P4mzfuCN/87XaqSDLwp/wy7Yyrerdwwd2iwVCqyO/+D5v+5ZcVb+X8iMD1uta2
dZXj8lCUgMqKu4fKeH07A5LWkrAo03pfK0N3lAow84aAgx8CCnTEKoDvrmSeGC0QZf0ytlCAEnlW
/fdjems5I95CJS1uvAUnPRVx7ey1SgFLsFwu4E0CkRDFSZBawG1Tx7KzocwIWJHTBupyNsMH0ppA
9N+2vCt1JuuCbhU3Bw+8PCgge3KP1BzH3Lm6xAgS4qsnjaYSuX2/WQTG3xEhJJzw6PZtjV7YLHr7
zYxF50WEGJAjpgfOlCQVYeUQ0zQt7EoIyn5jp4fdMQNNbBbn6632FaqdxK5GOzqrvezrmAPQnjfL
URov6D0MTJk6gYoBMSQyhRAdqr/LGCMSkH98VwQHDnlopJiU4qzlgBGwlqgm4UjszwVOFMb8flGs
wsh6tnvTkOK/e4dW2aiy7Z4+PnFCbGgMfKlhgJdUj7soihi/OtC81fjPdnNWTRv6SqZq33fI6mMr
OmnQiUGtchfH4dBA0/5lV90R8Kq1UWgT0lxx2vlxbvUqvoAyX16Fr55Oj1RhuY9v4GtqV9NkeIlA
TDXpD00hESEq4uqK+JcyaAEJOjQtPP6NYXJki+kFJU8OhDQy2ogaKdnySJQQcQGWcWyv5U8iU+RV
LzBJiDSLpkFLniDdqSBM+pByWUoZlp/tVDHSOzYhQWeLUE2BfkJCh/pJfl3T1fOAlWeuyAcfugOi
aoZzxHSShGDZUdqCPWK9Fv24r/9yqjTMOivOUEVISXuivho+1RduGL+Z00NiPOdpPvsX5SlBN6bM
Q8waAnKSna9xSx41x0u+HubRUKnGGYWvsH8dBdKqtfvHDJoTzKMjqjNvSpz0w2Jdfk2NR1+MSDyH
YI5R7jEWQdZhp19sFk334PVe4GmDHICWkuDs5aP/UQh4n+SzhQJ1DM4nalf8Zuzn1g8575brTVq3
l/4f2o3RZvw+RwwlGE5ney9Kk+2RZHg7DyFXkmQOTQbe7x1VH9A+y7X5C6CI6DwAlFPhNer6JUWV
L8CSAca/4n7JxXWJ/j040JHn15qaRkjEgdTrN5d/kCffdAooigCnh4WRteymPfVFdPmBixfW0ekO
sBSrlGk2qsWjOWMd/5GG3s4dOaw5gZK2mDD88OiqWRZdhljaiFfJHc9tV2IlzQDQe/Fr3JJ3vsHq
pFmBKCdt0bXDeFzEsS6TfRCbgaAtmvZ0QcwCzBrOvJSo4ocEUTScLFBpV6vHAElPS4VEbWxi4Rek
qDokWnisy7OQaCuUB2tJJrSGx+4XpApTKjyMgMxoTGmwAyRf45684X91bTQGn2woD/DMMlJRB1D9
adJG8H5D10pqibK4BOoJRqhy+vyIMvxNtZUNwztcVIHZFMdwQyj2JaXk9w4Q6d1XpjpehC2q8L6c
0AeoNeOBxZdurxNrNCadByp5i25oYbKGfS+oLOoZWyBZwRO2t38/I09TsWE/nb8IkIbTAfHJHUqC
CvB8dFVkehqXs0uXu4DbjQYA2yyjjBjODm8xA14X/zAJ24vSyvgg7hdVdeAFG5AF7anaLW7u+ZNV
vaNKhyjzQqmh1A3aShOaAhbnfioNOh9JwHR7GLkNxqAonjYzf3LUuMLxsqBGOlvDSvt97TyJJiaD
9tkwg9AXyX8qzCUqwmdT9nCP9yparnsKe/R/hgVuSinmmnNXRafH/roh9R6NAczF3gyJWPcBGy0l
Fd0CMc+A+zMmQfLsyxSO3SIN5rdt9AX9Td7IHG6nVadFJeDgUWNB2uRfreR/GyksN7RdHCDDg/N/
8QQNrswaGqYu91e/R7hH8h/4N1Id9VXiICCA8Bb4OKYkH7/kPxIlUdxZgPJL9dq3jJxr4oNvyNJf
RMvsjg2Xfac7X/95YZg/10gZ3f9PZyOV7UJtuqhAlsHAHoe3aIjndPnlVqLcfhLd1Y/EzvZ99Jib
4FbFHYwBG27fLUHmjxsfqgg3rclSQVzNzpQ//DEaxAJgULoIZe7XpIfcj1ipjCYpAZt9HOG2uxCP
fgGl5/jOR9zNuQTlroPpW0ljz9MDMpDMDHhf4nnQv2+gmLYzS+vijCIzaQC9jf08W8yPm1PbfVFb
YCajK1D8IQWzZHR95q/YKTlxoppagbWfofcpRmeLKTTLE+U+anMeZ3074/020AjO/sYzu8UNVfbZ
1qNPDOJM3R8pIFSihS/W/McD/69ArAW3c1o1+oe9ZRuFhXI6cD/7BW+exqAF89D9kw3vyflTzMuO
AE/B5mh/uceusGTezc4XZkZVwRLAA0pdUzrMHcwvWDWeEFVCXdvFrKfiZl+KDmZjgmN64VuY3Y6u
x2JpqxkWQo2XB258rjOnrfu1Lt5/qNUzNrtiFKeDhUln8qD7LRCRk9hHyXJsfKMWYoOKiTYug1jn
W6u/zeRlYen1V3KLqnLC+EiCI29LwF8bhpibMUqKmUSkpB6LUeW0kzuPaCXodQg97VbEoTk13on/
Rs/D5KOpwMOq8l7RQx4cR6cXYEkdJ0x/rcII0YSGkY7JG2NtS12J3Vl9Vy5SUJmCMQ5qy4u1IHzv
GdqVP9fT+ccZksErHnezFDbfxrgEAN2NO8Dvfv9Tc7w/SuuewZ8M0YJIZGuw8UaU7OiEAoJmghZd
ZjffxrT1v1ARy4r5g6ICTle2rwuYR0/RlVEIGsDIrUzJQ0ust+lCvWg3HSDSxRELFOGKDrIFSLys
ePtqkNTnDf0QB1u1bGxQX95BfyubiyScqnbPpa3ZyD60D92FvCUBbf88l1lQHD0o5uRj9MZMJE9c
gFP3RxexMtNVa3qDEj9P4bV6eqhRTcjGSIXxmhPCt5/sBK15Xc5Nt+HJcDpg2betrF08f6Gt4z24
gle7H0+ZaDpfpZlNeWcq5sHhJuhCycnKnRA2y/5H9S/tpLH65Md7Ysi4MAtE4Rm8vhdOawDC3LGl
uYsS4u2ZjFkXiXwlW8Yvetx4Jl/6VnqBh6Vpc6rgjfqr4guZGENqQAakgNqNP63G1uTyKFkMslBw
MoHPnb4EvLYH8E+hB+QRf6mSe5fL9NPI1hSKVB+tDyZ+9tdw2mu6bx6lCNxOhCy42G2IXAbTfhIn
zHVrLHB50TCzR2IXaoehOpArAp+rTcfzVjeCwE5O0Cl6uyYp9wzsCAoC2H2OMJ1FAC5bhgHjVHyp
ppt0EVVRYlLjQhFHyWMbilr0g1gJoSUC+gYfcEimNF0pSAEtykjTNNEJYDnHW+z6R/7qLe8YIvw9
lGck315dMsBY+fV3HhPMJn9K/2L0JEOLrbhJzNGUYg6v4oQcSts8JCCKtq27//S9Eg4HTWkv9rgu
Q5aXs7wWNRDY19NS0qzEQrvi5a5DXtB1oxPVhJQqT6SxEXr9xXdbHKJufn/D/t0ByIEoVD6CY2d3
MSsOgeIKosOTMrnFMIzDXEEbY4Fdl7qipvQQkIaA6+06794nrr++KofKcol8b5Xh1Ho4MjiZVVJd
3stO7JX4CUR9gDHqBzZ8Ihu9y8sNgb2UvQrf2azokcnI/QuXAvG6ZXQwC7AV0M6O/jg2/UN0iBmP
Dgmog9Sbp9jq7wCIhuurbphdOQyIXWtNGmaxuR+YTL5StIqrQxJWlX/H7vTRMxrUzzPwm3YrnBZK
hViRmNdBOLkMAIYt1F6LE/Cogg/zrC1J2kmnsCx8JPA4T5Z3OY34BqoRwj9uIcetLOkfQtogMIFP
dLs1jUYrMICq/FBFNT+BF83Ogz01Fiod2tLLlJjnQ0ofQuv3HyHmu0CPKvx+FQOISGfLVCVao4SB
fJbc19tbP5JUpQyerPeQ/mrpy5zdZmCklwN8D48LEekSUIAPvdbFSMrPkzZbkrGhP1hvXe3+3vT2
n0yS4dRY74s1MYJR/xrSmYeDRELyOQ/uq1/ECZWi7Es1jHUQ/DcVqlu0DBHo0cUhhQmB7zew9ZVJ
xPyxeofYFjV8ZkAhZOhW0LwcR7WZ7mGjVUu4wB0HVIesAz/Mrfenf8vidFY9fzjGa5iDzgRQVHeZ
F4uRtL+dgsva+g7EqTi1s8eXaxpBl6W/MXuKDMw1I4+de1w53oYFnQjHEJ0lnWyEyhrrUEyiKyxJ
JHMkYDcqalR7JM+ymVikhXRTXMA1ewTws3jvtFg2cq+eUtfJAy0/07XQxowE18Qq8K9LZ/ZAo0qF
5C+qoYK7qTKaOOuWz8niuZ1kc0qvi5H9IiKvSNU9fN05ElL2YgubO2vlVnQXz3R14l1Tj148E1t0
jxnhbDO3JN6UvLFq/zfpK+Z0dQMn8V637dxtii/XglWOLULss/o1ue9MoXGqgmM/1FLPK54zzKFd
QeU5wkpDIV5ngxqKJ2aLWlO9n1NOf0NRNVqOMCr2zqJS/gMu50BnKZgk4tpKYZBQnf4iJDiK/nJ7
oTjTO97sVrxgmOis73jQood7FDziPqMjU56c2109ojygdiLsLBfDNApTH1gZV7tMxPm6/OjAB/Tc
VDkuyiByge0IXH448hV4zClRndtNITlSgLX0lw9xp/SxNeg7dEHJ2Zysme+ZQ7KchX1a8DsQFnN1
2XiBL0Obz01OTKy/5oXliuDwKNQtVf0urBLvtKkjlcDJmo+OTQP3HnDA2NQ2ahVYaWVVIOhITX/0
7h9XMzJPdjt25hXKh8gbKOzzoSorJ0YZZ9s0gTpD4fkHZ2ZG7xTgcF/WKXM9hTkSL5XSoO87HeQc
ai48pYcAr4dVfXVwGpBp/k6l/V/d4M/BI8xraEiZ5kKKuUUJaYcm6if/I3rvTBfr0coHt0YZq1fv
L2JXiRkHA9pPqCQMizJd+JO7nwz0QUy0wWzGRHOuv/sUVym0dHDWhphVfDnB7txC8NAz5CzKWnzd
1Mi3l2llvJtgUSFq+ZSEIdoSyf4MVmJm+5+chOg/d2PT4xuEkJEk2KbMUhQ+9PjGmcq4r13orEEw
Q+AL4aGJWcGhhUD0n/Lw964/+Z9OzlMb0+LrChTDjYTtG6CtB/cJPLD5vtNX1Us5pHTA5QMHLoJ0
OIP4sCCFtyl319Mp+nYLoCPzi3gEoWtTjwhp6IvgM3XNXFbNQgb01L9zFD6e8EutzLBKQxEGj6Q0
Cj3nZyNSCSs56fIpSzbD/ZCmofYsgMq1V6Cv7XDsEWNqgOOHQwVNc1yhFO9D3PfJN/oblV1DDzIc
H5Hrefqe1WmF9kfMhvXC//XHEs8+FtQpD56s8vox804O3GYnwnYs/4+XlealOxwnyQqrE4hlor3r
ymGIXrwII6M0mTMylgKgejxou/1PDNQvgtBtjidVBTO9TM9UDT15pQwNlRUStuYehD/jezhA/jas
El/wYc43XIW9aClXQ8EruszXJ8bD7nQMfaAg/0AfRwPXDTZzhM6BczTReWTP/67NElBdVAABoJwg
5e1ji96AqwnB6IFx6TSXTQJtVdAO1AOTU8XyWnWqX9KkX/jSecF5OMvvg/ALYEpP8EqoaVZDbuWS
ixussE3L+8q/4/orIjeCOXGDUBKASdnm7KFcoDh1hQrrQ1t0cmsF25IDVhBEz73GlOxhSZNtPGaP
0Q7LjwcmN+Vn238jf02FdZFpbJq0Qrl+jVIp6wCFKVatkTd+kiQaaWHUh1YDkTrysHpsLKteDjwT
bf329VmvPI1YV1DLA6LWj7h/3D9p4KR2IE6zKeb6O6O6W4ZW72lY2uL+nqflD5fSXfA0fqqvya+2
1OtBdvXYgxbEp6OnaKg8Kre3FLhA4b+8vGtB/Fr2T5ICuCnYZIs6Z8KKSJXGJUk5jxRdvzTDtnSM
Ne6iabpF+I+5AAzlg3LSf2Y7XE88i0Z0BGwK4x33BP4z597ePjmoakv4LAj7K2SAMXnDdbSngtHX
Xc6PhQO8rdajYqgRxUSvFx3snbaafJnt8Fx1rZstspMBwx830Bh/JLiQXtI0sqOraSzs3ykX1ZUX
BWlbudFGD2RASLyXaCYZk1b5mIep/XBcft9wBOiu2xsHt8ko4u3WiuI/xG+9xHsP9EqdAkjISrtJ
zOp2dNv1zPXe8sRa69oxSA5oNRrtLdPhwNbiUrraLke9B77j6OVthApkrQ/R7yEO4qc/Cq+bU2Sv
kW7EL9OO7Y6n0KjKUfE2Uyq+UU383FyxoId0PD041uMBUUbbDBTvw/OpI0ar2p+73HKah1BMjv6k
+ICKoiWOm6vLxyJzrnvrUvoixuxmZyhy2q8UM++rzHGjafNk7P8zEzlRlGMH28NoM0yp6UR8jGbg
a4DSkWmxBQkgNmpAZIrj/Vl5FxibmzyT4O++Qtus9Wmj5YN5msx3smAXf4GYSy5FtNGcN8TWMSD7
9nUSZ9Ftc44i1nUWbdPau00hIs+KK5zq83dosc/FPb56fkU27pyfYEDOI66wfg5z8dEok8nB/S+w
XkzQyTSSxuMRn8XdbKjtQyLIqY/YUV8Yhxw3prcueAr23AxpDJJ+yJxxm4x3uXhYDB1GLxPzLVPX
NVCiKoqHUMypI5dtm+ZwZD6MSNaeEqz5uZOXvQvqGos0wL7Q1PlXakbbV2Njt1MFIHo1eyrYV8bs
7Gc8jkv3rYZCcWo1GRaJVu4BZL6TLRGmYmqHbeNMR3wfVLDGWKtVMheQzA/J1I4pEuCf2x2s9pD5
mFK9ZFnCkDIUwYe95uy69mhpOVHxVzUrU9Crkr8xmrUDZwjYJoh2TX8RLdeMA9cM6rMbiqJpILX1
77XQ/iWO/2SUyCWB2n8S20R2Kflsk9KzTmR9KPfp+3Hor9j3LFNg+ZocZQOE/IIFQPTv9Bakj+aP
xE/mci48GceR8M1a386hVkDz7nr586DhrBZlDPUF8fyT1eMzea6q4epRQT9ZKwbktiogLQqF3+3T
xPiHPizg1j39EiHzSDaywQQC0CJj4KrmoXJUdJA3/M+L/Gb6FXUr8JYGoCO0EBGqL72hkIM+YM/p
Y0jIhSjdOFRzPj08FG1KWoAxmK0F1VVpdU8+oRJYlNtV88kk44uVYf+UnApbz3p2oBkGLfnti06e
0pJ3tqz2H4jWJq9tSvDHPB2vDcizJbAaSqiRg/qiiaceXePtQ1OEE8He/l85K1DDUqj8EdauVuyI
ibsa+mjHRjnrVDLz5IK3o5thPqRPjyjsmtlM15CuN2S3WEXquOwAG6NbQoWVnNq1NOUabq6JbmxR
QeOhxtx/umW8gir3YfTxeLUrBgC9Zuih5s18P989LED9ihm1zGZ+wggYc59Wr/kFVfAkBPwIYpM+
GfF6dWsfOW1kkJitsBPsR3Z+r48P7U2LuE2FIIPmNQyrM3SPeHUJIrJHQeg78yDcSVcnbql5Qo0D
jq1topZKTXTakOneHD+34AMKkZ1U99+0Mmh58OfeaUBOe7dR0MYBlp1zqrdtEWc2Bt81mIRrwhGX
vBYLaI4bwzQtCYywmpM3jSrlFzjdtqF+bvRhimlOQ9eW0ld4RdYtBLhgc7orEHYO981tIfyorhvl
im+kF0BxWGdRq+HPz2enNG4sXePrC+f2C7/lkvjrYKDfGf4M4Tzw3GoPLsunLbTzCkFGheJsRYke
BzOjCRo7/46RuRm2xlgtF1sq4QDyzLlybZkyhBailfcpLTbg1B/jik7uaOV/QjNf93EnbGMJgtQu
KUbAJbqnJxHXUfD2iIo6epNuhmRtjiTokrXZpf7m+/+a9IdzC50B+wBNabIkRBIgwJliBpfrcDFH
ieF50sgLJgXDmjYMFkB5cEkwZ2flO1IktKbCVMSDfk56GJHDJCtyqryJH2uOrn7VuMtTxgbjLNHh
4QNTGSB/cgXHgjQpsXfGQXgQbQEHZaXHA3GffT3f+oPSiQtteaNWvpK5kYMZ14eVzV8e4AhxikLq
Gwffuv+CN9qHJFCA2+eOiSUm9DXduALHGEg3P25Erk0vSU7gdayZb4l5UCJ9sFewgIoW/5nqnWaP
eT7gLvjsWD+aGB3ZgmPmvAJQvgaMEF85HysWdXsgIqNHueMLPslPn+TdYphmnqpYAnskjbi6c55k
wU5ovJ4VV2yAAY4yR94MACMiZhUPjRqPQGw6sNqMcc4jpN2HC2SuQKYA3gdpzWyOgDkGJmhJxFKH
ApMw3i+k1xq5OCxtDQTTRDV2TvH5pI/FsTm2EI7+OKf5VnwY9XL6oF4+Cxk+ynC4H+4dHenQyla+
FxShZOm/5blbtxrslJhxTGKPIqBY8nTiMv1uNz826yrCaLiEeFeaxHi0h1ChHXdeFiuP9ydy9Mjc
VyTu/HVLOWeSH2zLaLYwzSHJldrR7u4cFeeDVd2WAfxt2+kanXP4c6fdslaog13R7EbSkxSansJt
2uCFgrV7QD00/y5Rwd6cnnmSxHKFz9StOdKMDeQCoOCG+TJrssy+oJszYkTmI3pMWCsG4Shx1fWQ
FHCAUoE0KRQJT2PSTw+oX4uqPXss9ZS61Rpo+cwa0JKWOVQwiA2D+dnATkRcrzgscAMCJCtB81NA
pPllk2R7Kv7rajdDfJ5hKJSiNCxOx2izuqQKpfdrALIsFG5hO2SxlbpPy9iqypdabXo3iFBaTvQZ
c2VE7DlIiSZIx4WQj17OKLIJovVwGbe9Kix02gOzJNTtx14BhmJEs1n1Rm8pQuNluwqyIF6KTMS9
myKjYTsp3wQ7XCu4qhFSUmnVQfdMUGyjiOHNPKs+Xb6CjBqfXK35aiMGCu0KMIV4nSUjNkFu8RD3
ReQG3NAQ+AZPf0Rp35vj4JFdrE36qTwjXZk5VBO1sWT/+Kk+k/FM85TTQsCgfNoGunYCBLwGfPWc
J/7TKYYHyFrWNkTXLukzvyzTtDJC9kZlFnKEqFWdtrsg2B/E2wcuajEUsNbPjcAZEz8UiN9Qvq56
5lBkWbKRCuagx5DswWQmLDO4Dweykzm/LjXhUadDxIty/vf+hR4UMu3fTecRwrGnErg2GzATttoA
YxdGFGljtAi5ZE+uusChhXhBtU5Wvcom/wAKRLedFbYtojw7cLY00L6oM7G5zmrw8/Lj7P8ebjQt
O9ltvyOMK0hX8Ubz0miPeJwZKw6pBwUypet3uetOeKqvOUe1DH6aF/C0Kn/aRCtx5JJIxeuKzF3d
LumQMZvNMbyIyI7+NQFdMBEO0YvubzFEL65uLfmas3ZEMYp6to6JFQZScZ7x2F/DrGnjqRbuQgXu
w0qBAWmBfXQBxHCrniVGoohmC+sCnzr91tqJ+XggiDPAzGjnOW4LJKUFP2a2le0EedKxEBpHzXHa
ldN8zhXntT1TxtzbHz43duTHOaqAIPFVn6Grcapq2BPuJeN+aeFPZaMIYi3FuW+UoKtoufBwvCWQ
Az7XJHcYUov+vSx6rOQup5ZX+ZqlcUKT2o13oRnZJPGfy/RI2ARfP7S3sx3gM4/KKe79UtSEXcav
9YWA/LMC1vBmK0kngHeMwjVM7M1cjWUjnc6IUqHa7JYkylNgEQw2XtvUgQZZq6nYGwc4iA+J9A/W
I5ceG+BkxgklAXFvwdqiYKBKf3hGoKLYC/iL1r9Jq1mum8PO01ReRhRQsOuJLmtfpUZl7ghu7+Ge
jLQ4qrzSnXxM9KHWIOseu3BrfcBKhsG4srHZagMlIZOVnZ2g5Z6J8LV3kbltCsmCLFBffAvxTjnG
a3MfQMocd8y8G7QkL8r6ybK1YEK94QhDi/IvnHKuADcK08tWgu6XE3pqoRzHQY78MKW9VeAQwb3q
0v7gHJPJI2u/pjvZEcRZN6M02S8d01iL/XMChhqJeDkIAl9UZmaVV5uVs/ussO6Lw+xBLux7hq8A
WcwC2XzZ49c4Nhq4K2K74uTY9pgauJk21RzVIMoVPLTZf6/9fWFK8UvFIfvcBJw1/LBZI8sSYcGK
cTmfgGbEGtXwBeEJUBvCkAIhtldqZ2Oi5hrd6OZHZSqZQYU7hjXz1uZXnSszhej0oAwoAdyu9ozz
wBiriFvESdB4KPn+KCWzTGwRh5B90dhp+I+5UxiOsv9DeghFxlXqNFlrHt1MWVlYp1u8aTn8nWDd
qLmEvLM4VwLQB2GpHt+/t/Ia0tXUSSopavHMi+t6vhh2L0Fq01Hwbe0ZeCgdVpccs2BKmOl71KQ+
BXgXzxmDti0FZi7jpx7bc/mokcmWhLbejvMrDWBdAbZ0wk57yf9IOv9LXKY/zi2KFM6J8JpBi9Vy
XQixnXpU6Dpc3h20CiugDET1zMwSGWugUKIBO0zusPYX4fxPF7xmEHwRVoVOIY+GEQEVX6qgvMun
2jDymeJ/jhgS83DHPdSs2oTgM9NOWPfAK3thFraayARy+YAOw+8ezXC9UZihzRvmCPW8XtOc5d5j
b6CZVo7ElmPc0IWYMbZt0bDu5O6mO23GZSPCdq3RyT7U3KVxJWS6SfmGeolc3SE0HOx8lAj78A6S
XGqKFUOnG7JPOecz4jV/2VsEwpay0tEGcKEmrrzRHrFSXzVpWdd0/GkiwrXlWHsj/RGm9p+8c5XM
MQb1LzB/1BdzsTuHbl8Xhf6zf1hsIRJ3aQxXzpfubaPjUcDLGsOSJBc5GF/r36D0B6F8uoNlSVJO
22onepBtx3PP8/oMEYSgYx2w+5qzOGzFnGSRGU0v2Mbt/vnHIEB/q30Lr4hgnU8OwAwwTBfdC1XA
axwW9pb+vQrM+4308EdIbTjfYDLEoVLe4vGRuRvn2cP1MDjm57tiSRVpHREtpmkT/mPqwiwgV2PV
9xRAyuCTWhYZc/6geaFPtXqw0gU3E0gMRTuTYfvkm0t1pjOgXID/iPU/Bf2SjrX6mzgvYL9RLXrg
eRGq9KvOjOLE1hQNy6Lby9Lh+fYzDq+5Vp4GUPPBubY8z89Or/CPwJ78liRGXpfsAf8ZWqRAIQ9i
1tkIg2Q4LTtuY6eQJf5eWSq+kMqP3Da2/F7mfJ4xEjhzekRUwUD18jz/8cY9H+o2KqZNW5BEMUtF
4p7a7H+yM7GdV2swDF84uBWz0JSR2XhIx1/8a6V3JPDc8KuDEUriXY6Bns9/CDTFqEaUWpLDx+Gu
LfkqP8apP65zTJiBWPfoZ/iPa0dx7KYWsSA1bLbXw/ANNuGRmEJoqT/XYf3NQJAdNUuqpNFTsDkp
NymTu5UddUAvDMWYjuAGFMwDDk2b89AP9knaO+B7sHHHPog4xSYYl7ri6IEwO7Spe04eWnAvNjeb
QdZREf45m0aeKKQY9TXXmHyX+JEGwObJ3paIkRsgYmoYXQT2W6RzlfmR5ZuyRdLkn448BlqJy3v6
zQe7NOaQX4Ubs66edZlFdMwTMqqMjclIu31A3MxhlOAatREDfzpTTqfp7TPlKjQ3B7axJPnK9a4v
ckwHaJ+ws7X5GGJTWTGEzJqphyrWUP2vh/AXLi/xRaYmAHBnTL+OYtQX9OHtNxC4uITK8c2FaZ4T
soYWOKYKo/gf4GvB+mtwgtP+oXbR+bxYVFh+guuKYf1HFLyXkITlBq/Hm8ucsm1pgrzxtXN7SQ5j
Bz1JIV/B1P44pqq8Y30NnkkzLNEagY0jv55/dsr5mH/Wt1Vu2D4/589JSAbpHoSM045EBul/OGlH
972+5KLKSQXog8ufac3ZS7WjKoEHsDcA51G+/lJIiJxpw1vw7XhECFwWgTyZ1O1+5ILMVhISFHm+
2S4Lhdb0zIUGwZfnpL62b3Gda2IKKnVlVibSu6eAyD/mPXMmVK89T6QIXn8E9TiVqu4ePA1fkxDn
DdvXAjR34nINjkea6ppy9oms3o/MIGA71m0oP4Erg/5v681gmLrt7YZm4e0Um2fYQRTKbzEMDt8H
WQxhCBEFxAC1nYmf/zXdrTzkmpfnU6gC3mzoPo7/whG+L+BEDH5+ktcBzBBIUIo0NSgxO2lv8HbV
o9y6j91RB6ClZ2JOIdIANgvboibPhMGMarkSksMu3hUHPMdnvx+nOKsAD2KV4GJc1MgoqcAHyxO6
01hf7UGFqAkgxXarYoJSdz7JqrhvDV6rqpYh3dHQO6Du2blwUzmMZbO98GuX5ofDX88n1fDWbms4
S0Jbi4aUtGO5Jb+5SdSyAH40H1Q9rSiMK/8da8G7GiGPDcqyCCYaV+jGYZvNWLe2e1d0usH6DZeC
uqUwBOfcAF9XXlSq12/295AhLNlWglqMruVwreU0tjQhM7dlWe6PuvlRPHPgkXDWXsP/5c6bfNPZ
EbBhwclceCAmHMN7b+5eCR+444vhPWLe7rxQ1PDWSCHyAOP/jeywe0feqXPwSDm+MtVRHoavMoyF
9L+XsiTwnY4CLE/CnxKeAGdCWkFCjrUMlmve/p3FLh6ZABFPHhiXFpt+XTko1hne5vEiiN+igB1H
Hq3gBkk3cdXUPsQjGQulouahOrCqWyOnNVRlnb37wpuPjAhPPEkDdRr5Rdsh2wuT+qJOvfaNVg+W
OZtIbPgdFe+UEpv0gGXRGBEd2PZvSIRp7yGOS/VG+WLPcu0k1pdbG11vbkKrMezYK0XlA0j2AXba
KmXivUrAOBCujSXBG8qTeP/i8OQMiI+cVksZNYjZAtsdPCDq5zTT/02EuelquKOjhYIDxN6d5p9z
YrDOM1ozV1c1E5lpTq573F9D7M/DC85ws/syVClb/28/ZFYoE4jMSb/+CaCOqlpxkHELvqFtDSBC
UgZaq5RHZzQlRMAHuN6m3IJKOR3X0SHymbocnXgxjNec8HkaVz4nkvMMsN2rXwezIh6JJy6eQI9C
+IwIwL+Ei8+oBeJLdNUdwTQQ9D6T2W2e4/MEgaIO7Gi2d0nBmqtCcY9OlxMVpe7ck7yXgT0x0W1A
ukr4k88MqTZxmP2pmvJ2wGb0vr0nPXQ29tbGxeFmFhLxVy1rkvViDaBTEsNSSQpYx1U8jgQoFY+f
m8yX7zTzi+2eWqqMw5FPHByLiPFnPfeH9Poq9hdEMuRi1/VYMrJuqQ15mOUCIT7f4ciOuj02aqCY
QQCHaBaRYQ8edMBmyWdAEjpefaSv+MErorp78/2LIIMza2pQULUSqfkfnxwhSyO2z2Xk/cEJd+S7
R+oNjTgKei5cVtWBd8N/05xk146TjnA+sFTNDV6xlOpEH1kV0XaFvZ3roO0xj11uRQKRWSEv05n3
Nlox+UZ9Xxvz+ArULBPrvs9pCC+tLmVyVeeJKdvFvWSun4rTUATBuh0bibqMygtTzTLMJkJZS1hw
I3nKjLzM1k5mQJmv4ANRxnrPUh1HKGMWX2G/hf1NYQEFvbDEFsdz7p+GQYCtBEaguVH3JiuwrFOA
Y1G1NhefOb7mFbqwhV8dwzpc9Bug91KCcspYX37CAY5bPC4SPMtL79Kd5pOGTVBc0sjKI8GqXv5u
MUxgyajwmd6pbIC4GArTwKnPIaXIGS4f6KCpew1UPM3BxSL70lWxDwH6f9pHuAcEbdG668K82X91
R6ZMVqjKkv58rErkdoScogdHBOPLCa0lWw/QVYHoAmxtxgGktCDD0KDZZwIWW/dM7hkB6fQ2upOD
2u4xyZOp9YbGC35AyvgZdl4vZKUXECEf89iLIg4lF1yijhERnu9wdBYROVkk2VZAlS4Ha18ELcEX
4AB+RB7qLdvw3YEENx4TpQNCHIll0u1g6QqFTS0oMEkrRhr7gaUvLhTlui7N7B7TPckVxPFSYbUH
YS0S7zUcKT4vHEolSAjPLvxUvIIC+4ZiKSojHZD7v8Zg/WzeW42GDsvbXdQ0VVaaHoIJ78XHa2Oi
kNVZt7TwdwGBJW23FgjwPFN5S9z30ffO49ZJe9wgimNag68aLr6dCFgIl/MvFxhbaBNu3/tgjre0
kEjeJsi6c4JtGw3cRbEMRC3Cce9iZXmWVdAhDHrqmgTpua3fx/rwxTgPNZYxiDBJwvpH6+JEeaFa
ov5mc/dU8KIQWKsUTJlfNO8PpYwjoT4CKL7iATElAB4GS7VrKI7oxjnwb6wp/vhnPtMt5JoqY8WD
XeTQOH0Pp0TWqz1mEzUO4cEigp53UmACnZ+vgi93smol+EQbH0Zucg31+8yufvzAPnWOkSVybeUw
1eJ9SaypD+oOZsbwSacyu9x2y8jS0seldLEr6KPl5yCwImvBBzA0/V6nBXR0k9G23IFCwcu12BM8
kQ2sRKDZ9+ZloCP7hIWD0tnquPbtHzN3HQ/q3EVYmiV4yDnzW7ojm5ocelBDKELft/ePacJucQWc
dRmmSfZj4IwKUJdjVMV8ZTwQKhCfA6U+KPa+WNWEpK75XTAbyPHTqpKWPZoAXgIuhwoC9oqMOOKm
PGR//kZT1Uso5RbETvb/xXmtwNqL2DIVIFh4a8ow5ERtMZqD6mR4MhN4LqGUiAlC2QXdbKuOuxHx
J8FdDj99KegHC9qyf2cJL+03mUqRoousjROQ0cK74TESqYYWxaGQDgt3A4dJvuLRMDg6onbQ6ASP
QA6dFTNOE6M9llzbpH6AAW264386Q9TGAtZvsvmZU5XQCpR+j/HEjDN5yAwp8zgeRZHH3YWKhRbG
ADs6gCcsY3Av0l6cbCcU8iaxQAWn9viHbheeB4nYcfotp78cIjXfDFIkdKkH5uA6NkE3+hClJYlb
OK0jNL3hWw3wpYHW0QAQZJqVafkQTlTAsw1X1Z6NAysVNyo+cI5/4yYbFiyxQXuRnSSUSgOiyiVU
V7WU5yHHofUoYgLyzxYx2EvxwtKqgDhCIrVNxdE8PhShhHCSFgUArbZ0NI+PXu11w+hCJb420USm
5/qeRD565KXqcA3xPKsytM/PgP3qxXECqnIACWKu7LXUpKeehUgycBXrxzZN+wJrfOA+t7XPdXhj
BWTQpBOWBb2mwDt0uG1dFckUn/QtUMP+oAaB3lltA2Rdezi698gyQS9RcApmjgWnYD0EZgDnHEv1
rmUmepP+veC1UY2LFmrQGSL8PDDn64Ss8m689b7hXmg20RhN/Tt2SxgRCh+hYrH/NuXCIDJDUL3J
To4+kuWvLb6h7cfFVBjjS3IE7k6BmKMS/mZmSUwR3WS6F2p6kh20vpZRBu2auKmn/c1uJMmLN/GK
p6HJ5FAOwxULiv9pHHL4LiDCug4VBbhh1O7ybr2RrIleIzsf58f4UC7ZKPUFd+gyXW5IQUWzDsG8
e1xtzTaKRK9TuBJSzWLy1PHVv1NuuwllNTXLTjF5kSkECrnZGNppZHjaChjRmc7usIai9g/bST+O
VK3F3M9kWPrIfXA2ZKElsULFNbPWtjLe2zaUfpTvdwU9qhQlbqjUMbiO+ktaVhFL9vfNmrC0uu55
hbDngkkWHej0gvA4QZQc8jB7iRvFEDa/i5Ldohl1hX/7E2ZzY5LLYnx3x0pKRwruV0WTdbzq09Iu
voVwWez91z3ExzYKvkePaOfJOa3hYa2Xiw45tO27sfKOkbgjW2jS1BdO7eVQGgMVOu1A6QgJJu4T
48nDJq+bev8Dgy0WXG7vxdPOOJ7ucJ6avBc37czRXZFDlNx/2b62jK8MbtVEaK83D3NxteZug/aY
HaklMZcK/AZQoI3p/EtnJvdl/i8tcf9lkAlEJ1vtNtptlj4hEph9WsvPMd7LmKj8yfBU0mhnU6H8
kqKIDHvhArFo0agMOenSnuFWPpD87HF0up3TcTw+X2UqfND2hGyx14g4MBCVa5pbFz36fVn5iJBu
1pjZTKMPiC2jsv4IardbIt4KMlfa/gIwF4E4B1ZlsrQ8cCKqAaWix5xtyeN7UjZFqXIXo3O9VRCc
ZEwGkBT3SiSt2N6cTgzMrTjg6Q4uETgNFihh5jW0V3Xcx+EsptRGve/SOM5mIbaOdsgOiJKf78iG
NBT5ybmFv6m9cbchTQRPf2+D7yr4RxmuKprLteMS4rdwwqrjwslHZFk4kYFBy0NV9aAyQZKcfBhE
6DCf1JZlroDr+wFujfzWpcaMHEtxC3QCDGYStmonrEF+psUQjECZcGlGf/5Lk7PmWXbOSCE2sxpt
kT9UoGlSS3Mkz14CYTZ6muw4cOQ3+RX9bsgN3AhMj7aONiK2mhZyJjphclsNHEauZXoB9YSS4q5f
O3CzF1bal2PojJCaEJk84nCHyzaRPu9d8UoQl8GcSfjaqU+baFXDzzruBI4sKigVOOgE4cwzAbdJ
Se+BJK6tZh5GVF/AWjiiTpAHTj7+5MeFZmmxVpHVdGOtJNl//d6HZzrxYZS8o0XALh+V9K0egCrT
/8I17LdMippiWVgKYWXSs6Wix58qJouEHwPjazex14wmo95NeVqwB226SaZC428ZxdNuDVu90rG7
HPSEi6omCZqkpQSRLfbeK6l3LRumaaWUOQE1n/uFOIUwba4WHlOeDY8PdI2wxfc8cshvpFBIDm4M
IVct19YE7VnLD8mhvRDwk6FSNvoRhb46PxQcecdQDrFavxoPXG6OYv7g0wrtaNwwjww5D+aUhh5U
YbV7H8ZFaFDGMdkYIiWvUmP6zctebqxGC5+jcrZyoubeeire58GcGEDkj87TUo/bgiIkhzBYOaz9
jllInWtP5Cxxc/bxRbcERx0DKJyOx2qckA9Y/HVc4BZE18qypJwFAsfTcGPruyKJrch2Z/Ib9tsJ
Fiv3S4Lcv/pF78Z3WmOIg2cwT2jTrzyQCytgTkEfZ4fDoes++TyD+eQGsFmgs7AdwBU+b3NMQ9ru
qb1ZhZ0IBSJIb0OSUd+/yu7fXn4vZ9s2blkZAHMS6xFkgpwjp4lP9Dw7yxt3C34rMUxaKnHOuNs8
NJ31wtEtepJ2fp5F4R6SU/TzLMjxmdAWGNejUQFeZid4TJ6+8SlcWkpiJaYQGjJ0kwWq6Pn61p44
g3V+HK/YU2npICljCdTev974n91GpAc/GIja00JNM3sLAQn11lSbQlY+TlKNnQVn/z9l0D6/OKod
p2japYY+Db128ovk1EcyP0VYxtBeM/RufhpQhIuKR5NV9TOYQwUO/N/i3A9BqNqai62htaObAY3d
udu4OxUIudxuvq73HHQgwP3MDn8Kr5O9WIspf8YxcRE6dXn8Ybnuj94rU7nOcPjVOb4pLw225AOz
Jp/O35BIuu4ik70LHOtENTsnH8G7KDNxdU57NE07S6dRmlX1FTmfh+5N3h9Y2fPVTY+o1JQ/XM9B
0+Qaq1TlzwnGJ1fF3fT+yyVjyGyGralDBXnEuPoaBdbiNy1MdAvgOJs/SfNBATAgGhITVeXqPgim
kaNMeZRAbQW5jNMSXxW2AlHBZZo2yLMg4a1aR2oWf5LW5XZEzcdnYbny/8TjHDlnnY+Kt8WnbpEd
sxBU4+MXxoioP4vUM+5cWWuMnqjrErFfWfOqGBT8yfyc3AHGdk5X5I9DCirPMLTEngw0DqhWqJXG
LMGq30uRu8NORXbUIpqqlkz8gxI1lS8ufr/U+XDNaVPkSB1JvamZzWh+SIqZJnyvWaznPf5twdbo
O8KaCgmVkxO2UD40ZgU5RBbwyFqoh1GUCyRI1PnUNhWFdxDyFWBtUwihJQ5SqG821rrvAxg+eoiP
E2WweibCpmiI10dJetOKX07BB+wgB1rr4cyIPNynHN5OmYHHnLIe0reLpL8M5Uz4BJX7PnBxLDYK
m65LKhjBQvaKadGPE0BZ87cYDtOeGt36rJwep19p9Pp9B+imxIUxYRUFCLbvCDRmBx4+VYKogRNE
TNKjt9DL72TdHzwqqTT+XlSXcEiKj4U+UaGF5SXrO6UyHOgL+Zor2tuvW6EJZAVoxfMDDH+1WfhK
CsrXyG8SY1mJTzW3mFTVF/VhOROSzvObPwKjO8sP1NkBvx6sjyFGJG8+Yd+iZIHvxB2TiiRPzuG2
sC6QZ9TXyd2/eOfjGzdcO6909/vF7KQ1njhCTAIiq1M65p+AXnRinAMb6lknC/zP/HPhBHsWjOIj
hgpsaM8Elnu7N0I3Xn0lO0k11W/nLVMmTGrPa7vvbH5M8iInqoNxL2eQc/TVgJM0Y6lSmqNWcPXF
twsfNe+4SGNmaNWpQevsGOYsdAuPazqolboB+12jF0Rp6QHUpnm/qvmhFvVo+7XPHvEynj7Ts/dc
IKfeNOBI6Ye7IHk2rUcsV7JOdrHfZGAIJizO6PgupoekBJdWoQBmXBcxH7/LFq/CWUZtrJ2EUgSK
vDAhB3BQJKVGCfGtPFEojRdHdrhYnrQigeM3f9qHeJn9RGyxBj1d4U1/RIf0tdrw1qOt8kRsQBfH
QQYU7S94sgXQK99wjAqJqpjgPWLBXw2AXut+w5fal86rG8jwhwhLoFGPzzkYgSD0iMAptWyTzPhd
TUNigKGuQUn+eyIHHMCJmN082cLUlT8Ks1TbH6z+iWIAnUa/ug6nAXWtRUEfzoHKd+2DQfYz8EGt
hwQhdBX8ee55MPahUpSunre1gr0JWr57W5LleTlO044dF6lxs4yBIU/MWIJpD6C6Bz/MnrDJdMDx
FVsxQpXdxJa20J8RorxyizfMhFqOz/8HLy+LcybfXeB9XzJHKsknu6w/rqlaKSxHG6zfSaO5Dd73
C76LOioGNDfS4gJzL558jW9GawkOtvL/jkYGYt4DbuZL5wzzvGBQnH8FkANQasG5RUf9+4vUkD9Y
FdalHSYal39n2OhyaY8dctiH8DLhbe7Kgh1nxvibueY+4HRmdAuiSRIez+qzZuAXHC2Dj4tfeieX
2NYjwOECsmAROchwl+MP8T92CqhURITDtZFB/EpfaD6GgIFJC9nrxaULIVJ6wHG8f9jDvKoo/Klu
aemxyWcUbWeLh2s0HTXdsGQ0aAwnha734/igIyCIbT9DQZ0qDg6GpEaDeLr0FjACSEonNAkKpyrJ
M1b0CUZdjS6p9ikSFVjBUaGZuz21K/c6UxaLqzlKSEtVZfFL1G/TMbtmawk2bms7UA2F+efuvUaJ
9duwXf0+nfkpxUPinlLxvm4Sq5a/0xPOt1QkUqwKPqLusZimfZcgr/lLcba75/7H+JChL2fQPDpZ
IKF3bRkYv5vsk6N52AN2atiuEHBmTX9zI8PykNWc3ZmzrLz/B4rAZopJxJdf7rHml6ceheccLHjf
oZBUle0J1Cz6yh2JgfVxCWNDY9fxz/YlYSDf5O+YvvzlXTvTQoyt6+J8RghkMVlvrGbwDBsflWQQ
dhUdTnBM2duFVm4fPUeJcbFNXg12xozj+6mNYz+mwQ6UiDQ/Wzfr21uEoKvnEShBY+zzrQiBO8wh
GvnU2mcpK4JYWWk8/HugNHfr7Edn1X0ZIbsWM3xjLN0HCJ7abdJYeJFCRN0q2zO0FSfipUfMjcN7
PWjqoBdM5KBurEbOgxXQDVQPsBvVIoeew2NDs5usyguFyap6qWKtypeyWClUKrRixrujJCPdsTvz
RTiXONjuPaE7mK+LJs30xiZUa6GSObPpnH0xOlKY1OZHPxHG+zm0lpWNVM2KFRDqkfq2/UcJ0fPy
/B41t88aZuf8enVAVVMzSYeRmRHuhNOkV1FLITVUh5499VatX0gHYK6s84bDyPZ1pgWR/A1H2IJF
6xJ002WwuvbFAMu2DHWVwF7mi24mhSBy1fMv5QVpdKUeFCXSSPJCKUfgSA5upc9Co8avWPTodKNs
+yNew4L//rLV/j1ADFhw4NQVKB/GbUHqEmMIcBXv1cgc+CdyPnRFEha0w++imYhSpD+pc9yFJ5pW
WjORshzeR5jRHTTqjC88Op+/ZD8Z4gi2pJMXwfe4hMe9PtAKAQLrmpWy1Vzw5XvQ/03GiUKdbnFj
oVKshnXe8ABirM+qEE+U+EoOKmyL2jqFtrJQ0YrexEIrNDQDO/WF3vboAR9Bbry7dHD2gXf7ehei
lYIGe6pn1g8GNqYWC2dBmPjt9dAicDwJF73dgYNiJE0yaoRpOveRsQhWKce2OEFJor69ZAQRDEog
aLIZPsKo4y9SEl7X7maCxm0Gbr9tVXaXgcZBr+EB8isDoZpdKuGYPsoRr5Z8YHwp+nYGjlemMk+6
Pv+WGezwKBj/A5t8SucQhBgpu67JaTP3z6+5T0S1eh1IaaH1fgkkYp8X3eOuIJc26a9jVw6YjYU2
EKs+WU+8xoP3JzvSmZk7HRZBQHXvuwF9IyaxsDLt5jtyvJ6zZYDFl/dUIJ+Z9bj3agJxUK3naVvl
6buOojudHGV9wAhOuWB5hTCkkhczpeaEzC9fdnB96z9a8C9jU7rcop1TOK5vmyqZLPhh1nYMGnlD
fJIeY6XjIkTh7bow+Yugrx25vputS/2aH/9gCpTECdhFInRaK2M1779Ejuf7HOQS2ejI0Ddva0ER
ANqy6MMsceI6pqthlLoB51Jp9UWNcFwG0rEyFIpoyqU+9+KxhjL9PS62OD/ik3hAQTUk3stFasah
74jhmfLih+sVOOHAVKnCMkK2N4sy2B23ug/EjOb2tKn7GLjXRjKLhJr+ueJl0OG6ppLu9AR+1nTP
TVVI5vjTNVmQG4ZXGfnVzAJ9gMWEdeS9cd8Nar2nzHGbZIUHJeNyz1ZQkXwbEa/4eDmUTdNGrKab
eByb0N5HfN3lBKQT7K9SElx/O2RYzZ8gqjTBg1NUzRr5qC0OoP/k768TNWByljakICb3OB/fAqa0
IQ7y4x7ZpulD8RJ38lchAZoOfkXyZwR/DI+afrbYxoCT2lzuU/H94vt/XX1Xuc7h3J9baeRCnXz4
DjnaOCwVTZ7NxI6U5I4Ad0WrcLnUsb8H/hYHt5fLwO43bhyFmoGeqHykMbU7GST0WFgwzjbQQlTx
4DHZm86qkKngYjfHc7JDh5jQrTapL9+FjDNhvDGbrVU/D+tiXI3JbV165fArnlmGnGhw6xaN0zzJ
OM5e2AO3aAEq2jpfWbw3QwagqpQdteY58g2AHd3LTCjPpBFI0a/aR7+xGK8ubuP4Qp9Ds8/sBYk6
z94/A53uKIUyNj9fXux1hrbYj+OEJqj+Z3BNsZifa0RMhopcsySHqxinUe/ze9RGRhOUUtHlhXI4
9ABXcfSQ2q47V+GXzFp3tijvUgFsy9w8xV/iwM2VLBiEeJsDC0Hoze9obIWYKQDNwwKH0J8T24xh
t+48VaeX//cUGSPp+Bc80Qf4rQFQjbocbVv3goetodZuUEoik7pDDGgXHKQdmemR0jb3edrxOMF7
ZsvY48Wd9v225M+nTVbE5xU165RTOhmyKcrl5qCHctydHuBQTo0/JCqRracJF+TEoXQ3gPjWwA0m
EmlSJAgbQT0girekFln4sn7F7hL63MB8hPM03/Purl6hT4/BnYWB4pPAYspGL6IWI5H6A/4tGcet
S6QFJR+LWnoSZQ9UU5H245JgipO6Uiqs2U2x/ni6aNH892HVwSvdZgbgqsnwdGQ1mD5JL2rVJljy
E1OZoi5gvWXyTyeBshNZTH8rFjaEyGzl+11gvNkkPbZUevJnESOyq8ZbuZM3MQ5G1F92mP85E1SS
jOfnGT2xuxSHytwAztX79BgTw6/BR/Q3EcT2OFkY1+Xd6ehUsOp/yMhUVEGH5Iu6Yn8ko/tDnCtS
FsnbZ62znI1LUMQ+B354UiGGZa2dIQ2fYwJnfQRPSqR/xPo/6+wo5AF3NcLtdnD3SCdjAMXzzXra
Tw8Al32rI6fo+bTFBRl6v9Cb6+gTLFklPiaHGsGlPirJID2LpCAhS3S2QjOyVCvC3KYMMZLU02pt
Wyaf6Nd17/pEvjkkY93zV7vm1QH01z8hN3Dr1YsHy51PYaxUuO/aIlyf9uB5qoGY7Ml7eKwGVr4L
NMfEsD17No3I0503QAiJaffKZuhLsA1aVP8a++VoK5tzA/aIffqt+cwO7zZgJFESbEDu1SCTdmIk
DnQhG6z9/dSf/E7rJinz29bCxpmLbYLBNYyuVnZY8dIDutb5dg+NDidGPjQ6Xn6uYlH6Rp4D+VpA
ROjWAxppWiiL7IaaNOUNexXdmcGDe2f9xFtY2mEXj+9DaXM0eijZEhO3rdAp4hqZ8Rs9jkja5gsh
Egg5Pnp24UH92FsCwBlapvY4A0xbE5wPwYAHiW0Tvf/b/5CULuFqQMK9S5eBct/GQ/XK1dIpyAYN
4RwtiyvSBgmUZUbRvC9lErd1O1VK+AWxDHggV1oDxWzSN+O0KTVf8yrGaWAMefnSHI+pHcs8nvfY
JFCe9t1ukR/gPtEnhOEkpQ28byWEaBxWa8fnlbJA8Bgj4DLYMRQmWHAc67IYwxRBU4FIBkEQMGIe
ziOVrf54cYlLGDEF++x3pdHgsrbTW0czvBvl2m4TvxBvlkY42fXmAELTgupWZKxcVmS2vZGrA9u6
HCRpS/3DCbsBPwjQBZ5MehstyVuz0IVufvzjO7QvxOHvo3jzp4NspdZ//FjqV5WeJ8ujLNCcK0g8
frYyzEI13rnXt/EM+kd5FBK+Q8YmkA+BVFN/+kfQjDPi8MI1R/7NSASwKJYSyGYK3UenM3+brV0n
e5Z/YSeYgJzSlgXUYCL8qsASETRg78j9HGS/rtyvDt1bYj16cUdmr5yLh/yAMHcp1YXx1nwahlfo
pd8xKDCEX9XOcrMno2Hhzg4Vpolo+jJEyzDbDFYFe7RLyLu64stg85bs3IolcBZHPBmS+yBp9A1v
tgk5bLxwkM9aDm/RHyHlYxxCdrWsi2j7OHLey4rZ1VQMpxFnG9AVdsjtlhqHopB3CpBWSh2kZGIt
6Bmo4lqX68sCAcHV/tnDet6yjMtgAmdnD1Ia3YpIPzyZrQC+rSNgDbINoVlR1gABIapgglxa4C00
clO1FPHl4mYM7kTSvz7l2rxyhrs0P7PD9lmkN8T4VHlafFCKIR9N4IEGrbTIl7X46CJWv5daLo7U
dxKSpK6Em923G0Q2k+qt7sqXUiTYdrdzIGr+5Nj89wtgsAi74swSDLszhSw5I36q5ZKGaz/W7cC4
hCKygtcYhqr2cMWxmLNKvU8vTCmandMkTND1ccPfdA9N4jep/kV4oS+7LIb/QUJIJHTLMOLLyfjw
JhUAK2MRl5+t7ZJGDG0HwUiiqo5FhV/a1b4ZXikl1HsiprOVnppJe7p3b7oiFlWzRIRkGyBBCQw/
E76RnKDNsYAPSodNY7W2kM8GtBc/mhPnRfi+VpcFShk4xSumsyP05AFvYan2VphQQSLnculAZeAd
uU3VclShcn2r7bL0Ud2NdzZU/JdP+Bq7MV1S8lNLc8/TAUWWbUHeSKnzTTRRiLtTaQ6o5g+tl2h2
qGKuiKJmEQv3LkWIwwFPjtwTy/TD9OSXbyN6c1RGe2LmQd0TSkyXAOVMF/Y1KA61KGeG6Z5VBY6t
RKEXG471fEZMxQNRm3m4RDRAlUzjadPcEKaLj6dnncgl23o2W3etL9YszAu7CNgGmVcLdC8XpKOq
JAn+RTtR+CRIbDtrh8xnwqx3sCkEXTp1eMPaYbL82DktEksvVoHEj8HNQrLOJBdTypPDX+gDtUMG
ny4OUe+Ohnf0EBrrT1JIEHOIW/XdYxBEl0IDjqSsasSUDoGZwhskh0SZ+fWcntkmi67cMprz8mA4
8lXdlcYmveCuDvgB6QX8OP/EfAphdbD5slKiR/m2SahCKdF4O+v5dqHBUdk5Jhh9Z6IRhM+kepvB
otT1Qqnl1cnvLvJnGSF2Ji00ikCxY4BV1ut5Coxg21YcCKYDnqEsjPdRA9jgXoCs4hCvHe2In0Fx
Ht5dZV7Bp2iba/7ytnMZx9hfS6gRF286UaFoMbZ/vaYD4MaFmgu4FVsfbWAlhFz9/np4ZPAfvScs
imaZb3LaaWZ4GHOm4uRFot4ox5UuRwz+pV8MVGuax3VN8oMWLQ9tZk/rMOnX6ZOuZDaUkg3G8yop
JPQQPX+1Q8zYuA1E6M/y3wkbdyXOo/1Gbe8/XkrHoHCrCaG0itN2OZ5KX9dd0HVGvoWYN7f7D9j4
5/RFt++r7kGPS5QVaDoDyLbrqtyg1lsedsqdifgpmTwDurlBKK9IYlAb0mzLJq+P6ahkwEyqnL/R
OdvADIMoM71hv9dRc4kRi3RXY7GL/nhJeme6tUpAk+4HAk3UZv6S7jbukXdxGbpcsAPo9VbB/5Pd
dHiTElJ4kY6FgoBkcqxQxoL3yD7yuKkZR49VHolpdaybSoRP285eDgm8LLpZwGS8ZnRpmD9EGOdu
YM8Au0g9ydV+W/34kKEpr/8kA9S8wdaJhp7O/E62lbWSc6GQ1cGRy8ccTKxjb/TNY2TOB/uNKNY9
EH7YWsnD7/JRWXPz987UfFdA4JGByUubLkV25rQznwZM7ymD/0iEb+G6mTPahQrDrJh0bQBRuoPz
AX3IlnEF4l9eH9s1Z6SyR02mjuO0r6tToJDjg/tIVL46KRfwAW02LY30ecQ3MIMAebmO3w0BEhGy
V2K5WvIH/sFYgZT5YUgJw2coaKOF4WTjcZOA3QzHt+e/DkdP6UWaPahAhYibGgZ6sgPOh0Tyj7to
0QV6g+q1djjIKJpj1/HGHsyBTkbedSmw9WCO6MLCUoBhY6Ro+6zEEdPli53/BwRlfjBTeMBiDZuu
XwDQVBlwbwfl7TDxzrrnseDGNGcCtgqKyEbrkMOVa8/19GJsIO8hh//HGC0OfvPc96maMagw88hC
gWejzcZFWZheZ6SHuVwql7L7ipZUq5yoGFC3oTX71vOEXxHXaA6gRyodCWAYDHYt5VG2JOj9Ovzs
H9g16qCcaPZ6rSwcYJk9L0NYLvenTrz4HR85r+aAXrUGJRQ1I/OOVI7hFuC8JLhmDt6n7RaF6wf9
0hSvbNO6a3KQT82VStj4fNkFdxXW/xDx2zX+STnmIcaMoogV+FY0ubWks8/T0Aq/kKPMaXDwq5Yj
Zefo9Q52nLX3z/NfLXc+/asaqn+goqzfsg2pgX1Xpdy5ZtopaypFIvXLm94SRkvzvUQH2MS4LOwt
woceuTxCMflo/VSRMqqpY6MfOfYrRs12iiR5ORShiXlOWMF+KDsv7bakitm4DmiKQLBVSDWw4gif
0NSabf9XGAveR3T4QEAgtsFJ5RUUucnowGC64o9vWmR29tteVhhRs6xIKtrESPf5V0RqzcCbGD9w
jfT7sdZZIaH+Ey4xf8Oaed5IYvI8duEYQ1cu/Lun8p4tr6T1NQCyJwdu0VnT9pR+p/exsxsgHcbk
IpsACkpenQcl36kmLmmln9SfKzJaad35QoGJjk6EY6ojagWgtA+xlwPRwymFsuZzem8+5oQCT8dM
Pcd8y0jRA612gNjZs/i0lhQY6MYEMPCTrW3HCcgkBvp+5VJYVGbY4yeplLCYZ5XMTRCz4DI9n6Mx
uyWUk811/sTsNaPHKhSCwV1C7XexXqDM+4M//hWVKWoujU93b7bBZfZDYVHdECCZ1Hmtvmk7tMbJ
9n8Hh1cNfIGiLP0T7Kc9Hwvm9sXCJkJUA7Rx7rlEwiyoyPTjSDlzvzLk3Z8hZ/IAZFUvpgY7P2XZ
9bf3Cyx8wJTxS3UVAGxmg9LalfUPkc49KBhOFNXrWgsu5eCIs7/DVlESvZ6r8tIlWG7qN6bdLyzJ
HPkgu3/fACxlGUIbUINiez9dVXTO8reobcGgOa5MGmyYP2b4DuDvb4zhJUGN3gVV27DYPvv6/96F
md8K0WumEmLeMUoCvuZD4SH9KMDEezJ6xa0RFpa8DWCHRknKZeluq9o+h8ABRr+yMnp0SiMpoa+x
Xusj6ywt7ti9madAloUB+amLdIOsGwd7iKO+IbolpSnhGKt8PMb1hN/HBdSXCnvOlMtydpsphX3m
m7n/J/Dc2R8f1kNDp/yxunAVVFSfCZwBm90hBBQeI2c7mmtDTCX3qAsNSU6xeVozViHHBtvLnwUU
DWqKYCciDpEY4qOvUj0AyJzzVSO8zIApNoP0RFzTxvN1HvWw6wZTc0PHWX9KeEa83UzA+q8mFTQz
d6TvEYMwi6wrvxG3sbE0ZQszrxwanUz7NlCa6ghzE6NtRET5yd8uUrg1JgThA/ekKEWrR7ZVZkqJ
eJG+o3Ab03EfqGJtu4mUHOeUUCummrJuy+jeg+P6vgHjDevOQz0fUKwcMtHItRpDCqm3Bi+RKtBC
eTU9PHFlnUi164NE1u+NUxOf8qB2sclQ15KXpGs+Gy3HpUdyKRwWr/v/m2lS7cBJqgx1IpcGc6Xk
dfliYAmtLO5aj4LOuK+YWAHQ2CPq/0LDSuXF1Ha3hGQa5M9HbSYQmYMgkjBldhuDdFACJgL9EHS/
qH0kfIZaPWjjEyBZDJi5r4+twXJ4cuRA2+7xFiNwP3clsV4NUCUzpQGMKg0MT5mVJ9LWesgCNr0U
M/+81r+an6MYwhdbJ7mEOSEEXgS0xWkolhpaOfzaXquA94Ug8B9olpz1WvQomb2o8I4XOH80UCA0
ml0tzQaBwFYJaWRCZ0w0Oj10LDPrZHDg8hS1rtvq6/CVHDWQH4gdtKfuxFoe2irx/t6CzJkOM0b8
APEW+Xh9gEyZla5IDypVekc9JAqV8kIZRD/TYEwXYFgG/ICJdb5gj4ApYa9u+KpynH65hKUxFAy0
tgcR0SlJskrJcFpvhWB+tXf5xZy9S2Xb9m0i8YIUh2IHnBjofFka+HPdXWmL0ad8Ck9V9I9OkBJD
Nq379z9uqRJj4svYBpTjfOSmcpcTuz2g9InCRIpdmpjBHFfgRQ4RuQAO+8gu/D8L/kobAtaTv9Fa
jicIkrHi62QkEVVADjjmCISzYToCN1TBWbIIINdJfedGUeeQ7vR4c+mIbA5sbjFFYuecM2BBwJWL
B3WggJ72bIZeu22dPAxw97Wrv+D3mkKiO7kuMRdp6yQxsuxOx1VpR6YIRk6XapguwcsM0j4W9yNS
xYvk1SgSrASUui6+yy1BtY5L2boguctvuATHyRpHKT5miZ1RvaH1ocAHiXwAk/qH8wJlMED8fGYu
5gOwMcN2JV2qASwrV3CukQKs1P5ETODOozyiIB/P659DlPtvcaYO5FsOcGmy85496qcEh2EjwCPV
Ltl07TeSGX7sNSdh/rY2z+4xBSqwk6YVGNii74YGMGBr1mLH6//oLGJMDm/E7X9BYjZJQDLhCd4i
295Niic+F5hcT/ESUdrDOolPFiAUMUZRhp09iOQaR0EpVII47rWd6itvCqW+ltxMDk6CCRV4hYLn
08tMJtugTScc9KKhkcpdKa4xTjeyL0cEwseXQfXc+IUPycGmHiBqzHYlKYhFCFTvSeKqVTdBeg9L
QcHolglgzR9gCKOxlLUYjOS3zjY50fK/NjPUGDw8GjBcXgXynee+iHd5Ipj4cgvOcwnGD22ZVvyV
vDlfw0hLfxi847vPSDhBUSILyqEsqbsWcQwP5+ZkNJeFWStUXKL+p8J/4Xls4rfhCAblBpRIzb9V
dotGbdPvi6PRJloSl5hvMuRtrIvfxDS0JIXzzrz2eDrBQsYSbvC/puSFGA7vSHV5SQz4YsD1dYTR
cmIXSvtKy3u/aYDBYC79dSq0sqqUC3/cFv1c9eQV8Sk1dQhkj2+8VBPfZFvWXw+Zo2v0Wn6Kq+Mg
2Kve/4Mnnipe+4G/wc/hy8l2meHeHsM5T0N9z3CILFDX2fk+kpHDc9g3lPW4nRqGb9PCSR0XkNuO
Wony8ZL768UyHoYWvC+v0qH/ZARHIXHMgAehTSpZi445jWpffCS9Em64ceY+W6jEG99Pu10x8X1u
z9gzIEw6svBsj8cueBdFlaXgfED4ejspTw+IxDvLjm+j8cK7E5rkh7Mmwzv8We8lZQwqrzTk25oC
fVy2EOA62RZHA8SRah7CMGhhMrS2UX7XSo0/Kh1OQV5OuOrp4FjGFVoI5GfttHzWb5JDLlXm+J7j
5pwTOaqbS6bqCQnJU86Qy9nol68TYsVfiZDJF4uNlemh2JPIY+rO55VVbplPshTL2sn8WrP2iU9C
il7eHx6BgChl/0tssansm8IcZvfMg776/lkP/QQ0L5XXclKAK3T04ugofpXpT1Jp4J4nTquVe+Ka
PHv2DsD5SDmgijG0Qn4sFVxSsyRdtkgxhZusYzF9VkAFz9pBfMX4FWIIOYuHp029ckA32jCANrcq
FwT8+CNCnEnm+k07MENvBdJKW0a4fgJj7MWYIjjX2vuKEv9t2TLAFLZmGTCXt1AMJr9QtoHbOHJM
559iR8GeDCy2KIUesYJgOGTQ+km4lN6Opsltja0MFsVeKdpEJFOPa8hxvQVK2ns223bh/L/SIV9x
xXDIRa/SCPb4jmO/jkyNpw3A1ktbYb+sQ3wJQtBy5Su56qL5eH21YwSgYjtOx3ipdLGOyWuuu5gZ
Fx0N95ago54CfvMHrJOMpfb1fHyQCAU+yaIAZsUa+25gKL2naWyUFbGBeRn61q50LakLvQlcefa8
mrNS1lGlsatUBi821tYOLFG8W/jV6MRyPqGnflx7spZOFs79zhHpHstpJ0v7XNXXYSUkxMTe1mSX
/6GbUeRN0jZSXNrTlK9P0qwlDGrxpLf9Q9sd0mihDtDUQ5hZ4pbszeBjng/dUuDykugS2zry1cQe
UbMnnn0p1woNvC+F3jt790hsZf4qykegawfnbMCHHFsXOHsbNzw21+5KUEAODAmZcPaAY7dtVA6E
P6HgA2bJsR/9KJsWyn58pJDyYmJSOUkf/BCXbIIiAMqFvZeXtY8u4tuLeI+IygxDFtHmrRUHfTPU
MV21M2tVjq9EjuCT+F/1p5/tEjJftp48YhysrxBzUzYrHRlyoQw/Yh+TVVkAgFl2tcq5Grjb7reR
EFwMTAT716dmrRhKeZwm/k6xG249+5Kdvj1zwC4aEhlmlNJ8+AFBCWoQ8SuYx+2ltf7OQmXdRgWM
8aZuTLPJbJ/NwmK63LVTChusDly8w0eWHNm7rCR16kLg8gNfRv6BJODG6Om0X9AXgW7CQziErrvU
iTgehgIzzlebj0BZ51LPAxHZk8CzQm+JeiIouwWJjm4FCX+yfDGoYQAwZWaLVkS7vCdSNcTw6kp2
qOTQjwkHDEcJ0MktpfOTJid+X+bw+38nZRIQMeuKtVLh5+o2cfO4hD1Qsv2gmQpDq+zvsaObKZCs
0GklewiVggZtaRZypcP8FqmLLxPwcSp1WSWV66zL66Q+D3TjTgCfDmZcxYk4pa2CGrlQHCC+wqeJ
b2J0ubOLThHPjlZL/+QxwMrQFFqR1yI2CVMzy6LHniru9YhcSoONw4o5r+iCRDruL5vIzmqFfRCV
FWBHutSxqNjmJXKN+uf3jFoS2iqnwZD0qtJuhzPF5nJe6xgv14gghwKdzA3j0ke+kPhjgEOXUZaZ
9VbGzz/GRvdlqn0QNA4HCB8JWnCa8mpmVGcyFboI65R9UrBPbFwAfHIHXzxXOdSGrbbyM5AxbTtg
B/8WWJU7DJ/LNxNnvkTdVRNZjjYp2L0xfQaB06mcY/q1gAvW+CxuS4w89qjoXaOVlWGIJ5KiG8pl
nbu4UpXx1tdhaR70AoKm72n4MTPQfngg6l446w01B+lvPGVryYCYlWWRFugviuSAnTh/ckbTA2i7
QSyvDU4wE9ZYbwdb79xUc2YqCwF+0mLYBGdPQ9JSEGQLundozp6rbNOUGtUdiWy6vplvv/r+RBDJ
BTy7Y2GU53wBDhkMpU3U7VF1aAR4Wj2C10UNbSCxCL5l3KaU/iEoJc0S48Bf8tnnlnimK/qC7eyR
wPrthLInpQQ3xmz6TKPBtR+Z3kUVUcobT5ZFm2dSVpeUH8R8uWvGWMNQQLdCu8BXUCRFG2AdDWc+
1q4YMEO836vuLuVtbAPY1e+AC/DnTDJuQl14jbh0eqWYp24ha4IzYhxmYJxDSTTDKP6ZYs3ZObPm
RbdAR99a4BfcyO5ijPZoqI1joG7TSUqy9FlnaNVzuXemH0cVDWu1Yz6cFESf4i8TLY4no1U3oElB
UKvxuXieXY2G4ucUyXLGa2ynS6yQoHeiqWcvSd2qcvGfi2iyxhXYYcl5vLw0U5+Bv05tN3hahmMs
fYUiv/GR46afmouf3qSlWG3p2LACVsFXlzNoXV7qpnUNAtwm9r9dQVQU504yflgAfjE+zbInSfbF
AAzenDsTDoZQZchZfZXFbl3V26gICKYHsYeGRh00ESouk6hycb4YF62AN1LIndnt030kCt7exPw3
t27Nai68tG0TAJgHK5Xv5D2/nPDAoO+Bk8b5FBAT0mkzWQHeZ5eZlY+L3YnvbB9tHoYkquBMnrvf
IksHh1qmv8k+n4qm+p7qzNOxB27GePsxst1vQILoxOI3ZFnThW2u91d8q7dKFTdwCqG++RmbiByK
xAuLeWY3IEMfALPDbpY1MfQDCoL2V/A7cvL30m5hP3KcJKSQwz+wFdC9uA0ZyQBNGOqDw1WHjyQd
bRCG8izQmiRihlCDpcRGolE2ZeWXuAEKMbC8ScR0aCSWz8QiMTF0oDnNrOyJ1TebGMQMIhIub3cO
8K5hWQ7+c21ulQGZFA1s6cb93jQTw/GmW5GBeYd6EHQ9rues6qu+ubX7bE0CQ9A0eNm0q5xkMY47
beR9nVCxPKWIBhk6JCIRCuqrgO5PCxceDabm31o60iqda3BAsiSIzv0I9ao0PYDgOXLb8lu8WZl5
mWYASwrcGoPwQUAp1UIqg5G6RcA5quKFeq3HeNm5lnu2CJl73bAOwr2WdaP8ok8ixbgii9/NNDOh
kpNfvFb1fJr9wRqj5dn3jCSJtvqDr89MdZhF+GnddJQhPckdKwRHmR1ekOsn0j8CXg2NQhbSjSTq
qR0WS/TRjh6oo46kH16AKkookkxeKhQ0A46mBzHQDCBtOVNXZ/m2MZX2YuGtcMOCySH7L8yoaQa0
1u9rCORt78XFEBLYJ8yTALwTVPsApjSaccZeiw9qyklq1jECJf+gVlDQi26x9pSQ9z+5HVkkLilM
fVJO67canzxYzjc39FC/T3LTpgxY+aZrInocyt52GWeK06fZh9zvaI4q+tJJHQTr73gAoynPZIWZ
15aM/S5xFFWtPKuggP8211yAawkPcnVpNus5oRhCQchcrl2vvtTgYSX3zyMacqp97LuYADnkOxzC
zBVIeTYxSBke+Ff+nI8mjFoRm5kCIJz8aD8vNhMibOfj7CniGzS4DyqOLvoT9O12DqN/uxcpf3nK
lzYChv4klBUHOiJHf+XGFxqkNilymvp9fS2n1GA6UVfXEIQJk4EfHWw/Txwr9PCZEpDen6ItEVUf
wbHPxBB1m34+AgIjFe8+zv4ZM6afiruULH3CN7rpRPPFzj5gIwhDjZi5gpJPLPicjOpJfJXlTTZt
Qclno5aMXDbg9+taG9HGXm3iX8+IRTmasGa4TbJMX2af6YJ6J8Cmf2i9NM0vKHD5penKhSiz5o+g
bLe+oi5RgpC0A85ONqSTO7JzZCholV40pO95gLlLEnIpDBWZrRV/6i1q+1Oi6cr1qzyVaBZg+78s
/AQuCNebQWk/XDxREq4cLcurA614b6+BjQqXUBw9qzQ8ZKwXpXv906zIKBqOyi9mHd+/QYnHeX6P
CY2n16cCt2ttikXjoI4A06G7Kg55v0ZoNP2hl0QI35JmFf+o6vyNLOwrTTJBUma0rLPrs/9ISqV9
YnlbX9+GCXzKx1v4eWZQWc97I9N8mFrz2jzHJ6ULqVTaXhuLUGDABkwGKTOIOMdmNyFNSf8rNz+q
i510vvR1psPt3vRJ4yWkwLBJ17ufsUuYjRBZs0XNldgbnx23a/s2SWUvAHL7mh3JAq/eJnSv1GND
asplvY357puBW11g8j76cbw4Z4+N6Wl+z309jM+vfAbuAroz8x1CRkGW5XzNZ6N1yW9jQWhRGBxr
9Bceppg8il38LDnABotPL+eCViMBbjBj9p7lKcHvZo8o2Dqzdeuyh5LRq3D4kjhfy0eAbw168ol4
ybmsF5IJUSLrKuORfnoWFqBc6+qxklKrCuADBf6s7pYjulBa4gR5ZFdGBFVsiFM8pPrzqBEVk7GK
ieHNBWUGPdqtnEU0wpuUwS6mmrXmxKixNiLFmdu/dzy6PSQDbwcrZvC0e4c77MxlAuKMYH6wrBHa
T/oIVqKjyl5xT9P5+tp7G4IbctohiqlVOaqzlVN1HVeSoSnE9yNreYZWbB3vJ5awSRoR5YACGP/0
69YTQt9QCsumP1sX8+7V/eC3Ypp4qtL8at9UN47Ny9UrzkQ7z358cbOutBwXvlwHukLJBibd/4mL
pYr3LM6Fym5Zz2cpfHXhG3VKg+EFk9L83C4m1pvDMJn51zztqLkICOVpyuX0Sl/E3hhSQX/FhwmB
qjA5ALSwaLLB5Sda8uGUgWBts2bBvK+spuB9WeQ//jQD/XJMk7w4jAmZC7+m5kzTEkDoKPx3UnGs
WaZqNjwE3TNbEByQvgITluBRDGZWvwQhJtVVM5cF4ijxMua8fS2qo+MkxT9yIsHQle+aaHd3cIQJ
/Fg3eoJ42xSHwROpWzD0zORXtkw3A8v8/LeExy1kq1EmQLu290SNnE8Oa0gOB6PpLF7BekiwIEXo
l54krMDyf3+y1z2ixc4WbqwAmqUj+BIlp36RS+zkXCpbDMNp2KfeB0doTJD1nnFz0kgu1MXTB67G
d0xnA4oSB/zXLevEQsG4Cn0pk023rmvqV4x52s0I66xVQ8e5fNsJ2iC1OEjbU9vZ1gL2+bVLOO8k
OIfxoXFi70tB3zwxtKH2JlUfHNEZb9CZcjmra09m1xnj53DI6ToqmXm+sr72AxcilVoIQDr5dMGP
CdhD3Z8U7pkU/HiDfkhLHOHYaMj0J/I/TJIJjLS1ijQciqf2s5Bf59a4ikN0i2qwZXAeitDCXsJW
gjQ9IZUJW9Ova624EO1KfnHi8k0z+IycHR9NAC77X6J/94q4KMdF0RhzOmPuvu9N4YuHvXOGrzw0
5SB0CDMl9FQB6Z7nY5eGumdKKDT25QnYPG4vpNE0AS8eJMjPNjCqjeY0aoZDAacpvzXkPLoSAGGK
D3Imk59i6iOmeez/SO4hImxIMcpoyDIidGLuBtliejOcgeVHDIuvSZYjdQXN0GQ3E+Ump7R2oojy
sNnCmXCqzVarZLNtPpc9Z0stT4o3tIlE+DaFpCLFIYsNXaLf6LwYIc7NVlqR0Ynj+4hShfBNNhk+
q7GBNRJi3zTjTn3BMpUNQwsW/eHwcnaFtLskw4RQ6v6uJh5ra0X4YvRlwsRsIFPOrxdgJCHSi9Yq
IYL7NFpp8bZnBYgUB+tQkp4tIRcarUvWjqwJoPKPE49O2KgSRvbBHii6zWGh0xU6JFipAJA3LPI0
jxVgl8cKFT7eBjQs5pYfsLgqdCLY4kuK6nGLrj5IsdWpqceuLwmHhEG90Q6STlkD/nMVUsnpEHRP
B7nnVLsNLvSUdH9DgimanbcMtVbISXUzzujGTr6NKHaRBxj+eU0DzrbCwMyLpeLolOxb1WqMQXoI
/N0apHBeDP29bIP21dSq7a9x35kZFNy1Vil8rJAMo9NpvHCxU3/hmtjMQAEfBi0ba7FL97eONCVP
6kdGByu1Z0J7JwVKendGmgYdtna4m4Me/3hGrx/WyHUV6UiM/aeiZTFSFG5wQmW8Ank3ONJxv8s1
XGw2nz92KvEcgI8UKdyFNoDp8ohUOzXCR8yTEyTl8Pm/i6Hr+a5LYIwaJ+8y6iXAUbxadBebjGVT
i3zPVa5SBzF8G0Hfh8oTBhilgCay4I/mUPKThTAPkDCxJdTw89zkqKlYAreAeEBdswTd7556gzce
fx+7q2XNvLOIKqS0V3WVl5knfbWT0Mnzp96PKMm+utFihyX/TGi4ew6Amo8It/PiyJoZvzZDaw/v
B8IUgheBWzvhmapWiZ3I4G0I0D66xa6hBf+Jy9PhsUdSKYxKZtJYS4fgqDHKOG1MitsPzxcMrOs9
1KdM+fZf5tzZLcse2oTeNp7tFOqSI5UFm6GjaP80HVPXjfWx+HL7fvs23HpQUCkeC7JKwTAEJyQO
rdkbxviKZ/g9cd31YCR4VnhBtnB2XfhpH4EJ8Xb8d4qOjLhQHKw9mtD4GKfhZTLETlMkX3M5/jmG
HpkzYMF/r2uKDMgTgQvLzmaIn6Ur63R3exWIns0K8js3u48tC8eVwXkMQxT50VzZc+qnHra+qF7d
0fab6pt4KtI9hw3JSL7QkUPUvgN1oA+i7bsNWTroooFoxo9gBKbBam7a+wEB0H5nQFfQ8pc82Rsj
UJx51ZMyWQvYpkUWzyGkRTxTIYX+zucAeYUcYzb9Jj52f8QDebP4z8haiDbAbeN9g8HMKgdd8rLB
ZVAgxfBkhw1iLDK2tOm0bBO+RDzDFObFDUcQVk6oHdQWdhh44yqdlLkELqQBIEXFeBZSod96O0kw
+eBvXmt/zFRazs7vmpfYVm6tsF9L9o/DL2sJzjQ9HoonRZCikfAsIDo5SRTt7G8o9re+buTjvqpv
liP4/s/nMT/KbncUreyyB57AnUXyLpsOPnGpZ1JXLWK89GSvpg0YzL7PQJa0yWhYaAlPVzM2Y/9V
1o+H6qu+prRHSwH6k60exxZVN4uDKcg0a7pxVd4pHik3dB5ryTdpnUAnQlQOqOqbbMeZd3vXD0cN
kI6Z0TGQQ/FK8Yk1pm84zFM7rFeyqkzW9W19Jm5dHEB1Lo4LR8ZkHa91A0RrTPJx6Gg6iEmXG9aU
SjPD8K4shme4wF3G8dRSBoKaRW1gz1OPoocRMsVDCI4f02hLAQi7FkW++wy95o68iDJxnKBOPO+H
fL6DaseYAE9QNeQEiqZSmRtSw4HdYf5Z3CwXnbxdpmyAvLVe+egd5AM8UgYVwh8pAMfUCgzAVWBQ
qBWqjsIwj5pN1hFLHeZvtYKOVoKF79wMX1NXYm1CXGkjl17RPD3J1Gtl7ZcR5zaN2O+279m6rt0W
HNxXONniqzX1JpeKPsn+Z8VSon0w1Vd8Zkmhrknf6JPVBTjddo1hB2cboEyl6osMJ4Po+c+GcPA1
ptrX7MMYPw/DmUByafNBwajVuyRkncOzxmynWe1nlzILOyo7VPHIqKDSg7CbTN+94FMwsqgVseGV
1FGF7M9HCqSL3EL1eGeB02tE/SfX2x8gAYuJG2iGvCTNEOXbkJqCMqaPs4Jk0TgO5Pn7nCaba9RP
K2242YjP2agSl7uXLLbFVC9WGh27Zz9w4jAEc/tLp5I+ibPdouDRdw9atWgmI6mxwEigc1v4e+Ar
hZbFS2FUCY3mtzvr0AJMoSgbJIoBkL99SlM9/OyX1TqU0ak4G6xOcAyDLqpvh8p6PU1bJzJBzU3P
LwXCMJ9Pm+G+rH73BKND1QbOjyAdFrIORYkNZ0tJk52gC7CnosIz3a2JsX7p9IU4Zw0spOX2adOY
y8pCDGU+T2vCWaN8M2vXpAEWIvbKmxrT8WvTdQTmghK3j2sIkPlJu02jzlfxG1N4a2WINiWLfKtV
dN9Y3Pi7JjCTutr790bHpogOIPqcN5zXb5t7GqoRU73zgSrMkieGqA3ienFSwY3Ze8dknyLDT8rM
imSABnTgVB78jhxctmfCh78d1Axf8DSRMWaN26qrPXbnxtQx1I8S4TcBjFC9GD0QNoLntt70R0v5
wCDNSWhaqCjvpi6bX2hhF96P8/6JOaqqIzrjzg7qb8xB0IyquaNNjvcSnupfuHIMPbyL4k/TuWak
wzJLEKz/Yepk1p7vPqU+72FbqeErO+ZNSxvqZyzQjp8XbwDCLWsgPi3tKz+GZ7f3b6PrPKaEdLGV
ckEN8h3bsz3SnpmLdJC5d1H4AlmK/9cm70RgmomiJQql9U7Gys34Z8xwFt6tb203terQMSwhEcir
54y9yi4PdVQxQRMRjMpzRGKmwmys7IiBrMgnaLhWuvGaHqCrWdcQaM6NTAcgHlUlDswCcSM2MbLT
JZPFU6AVAM9FgIZ7mcv4K+tVsWLtY2pxQ8XN08M0baKhrurS9xD0DyUMHxclPxROi1tvMOxORnnh
PfIIpR4RKhpwydUtCx5Smvg+W2Mc/TEX6vTxyKx3zgKPOWEtiRGfy5pBLggxd6jnnVVkJusn5EJM
VSoJwBok7p1kVxQ9gRoQbb6qqCRNn5xH98I4mGmH6nEZ8/HbZC6xofmtwLygYoUdtlNe/ay5FdBr
Snw+hldPGhObfmovd51Bwdq1V6QImTm8lI9QmdIea6OHhatKAUg4Et0cVL+A2J4EjEBCIwlC81Dh
GWDZyvc2hnBu6EXlSgXlLGFBUtmvhX7T9+2sXiNR8O705fnj2Pc51ukCRbp2QqbzWZ0xmrU2ci5d
v9p+xJ7RfiqNlimUe7/ucQzX6HY+gg7N+MZYxUZcDUzcQCIPMQEOFV1uq9GpMEqY7dk1wxUcdqiu
ZXdmsQr9ObkZhnf4Tg4qNCx8YvSFO3a9wkJb+wrTzni1vKBYWnQOBLbI4K3z7NLnN+3KBjw5FIcs
WKqUng7wo7IYn316tiFhTCGLzG/avy0wOSaAS7DHOrUK93FWbS23Dp8JA+rHVm1BoDOzRXQpHCv+
szs5zxs05MHrJ+yXjBp02Nwc885H4xOu7os/gApAm6CBBJ+951WsWuTuQju2i3efcqafI7f9ScKQ
4PDXzSlcod6OcWuv7E398u6QW97SviLYa9m8+4A7hCOVJQR+6uiTrSHY8iWwdnP2Eu0rJBA7v1HE
ueVFq16hTbsnafwa7cy/SSEYnuNiba3hT0+jRBJoMrxgaWcEo70M8/W10wsxXN2LRf7lVG6DrJ3a
kByPtqSm7DtW4iZq0ubHaUZgCAz41cLsB6hZsImw7bSXdcYobsOAD+OPeURX6dPbDlNnrfiWVyBb
BoV8Os7Ow0Ns5454qj8EMpxigNHykhkF+vPgKwKAUrAgFiqUH4fn2JoKrvPLkYsmO+yHQwMnhpyo
PqqZnfqn1KRiDTSQ4hkk3jXYxgARPstxBGvEScAGJelynAMWPFfsmdQUn1HtnlaicutlJPSHdKrg
qYQDBzPTukhHFiRqx6APblh+AQvhLp5uZ/MzKZn/YkX7I2wzmOuLtarYSWNrf4EBe/P+NnAVm47+
Qd2k5embSA3lyFDLkcDshNkITmTeOgkVURw0J7NhCiPv3HziXWYzdUrCA6qhCYBSnwYUPpiHxxEU
QbQ5xzMFfMYuS4tc8PJSKQwljZyP/rWVJYuOU4pBycM1AVf6wHv7nCWrK2Ux3e4Q4HUGzjZS0UXl
9NLT0YQqvAyIFbEVal6mkAIY+eFsJ+k9LseId7j/XqTlgPzhrJWknmsNQa6ipPB277U3ZymrG5Qi
DOiCMbbEKqIzx5OKfimHsdBwDx3VBrvzapnZTAtCYH8WExXRaMVy5TecrWw9XiA6mZxm1fx5WhDG
TSl976FalBR8pESn5kPZzGfGuArla/SWunqLR4Uv8kla2MptpIr2SdONcq2q2B30n1lDCyzyxMgy
49z/Lgn4ml4RrGwTm9jIEctC4TgsqP1MjqRoeeamiuNhuX461sn54FQ+wfJfB73Fur3UNE+CCKES
XJILztLTCSZTsxJtn+wzIwlkUKClyq89bsW98O2rjrhFaXTqOk95eCbcBobY642D4cMuQSVqop+p
lFjtcNaF3uY9bRZHLEr7fEqWp1gJD+6oE8BhTuxwe08qe6NJIHOMStehsBc0xGVsLMTf8OEM0POB
53tAJFBB36Kj0Dn1+ns/L1WcdsjySmCgDQXgaWyWGsZPptG6H7nxsqUMy1Kzz2AJN228xsX46YYb
Np3yXedaht05imVRlXPktrOAInzdZ6LOMeRVYEDth11GfQnHnRK8sV21ZVRg6AuYHQXYw9noAXHL
ZRxT2b5BUsPqkOne84dpE1YqmLmw3sWXGcaOC878cZKeNao7vwomyqwH2b1685fSco8J1E4FDDUX
YRRmFp0mghkTtCCGGeYWsf1sRFwCiVlcHDifQQuPz6tFb6t/GUkxlNifyzaEJMRDxPpbZmw8Zcsp
fh/3q1eyoTIdmTr541yG1ds1ADx6g3Q516UMxcIpZEAKDCluZ1PkMTwwLHRS1ao2t143azzBcF+q
/ic39Bmm4uu+QJz+3rynaGj/zg/iTmtq7rFYHz8nd5NyFlwu9Nm1wZj6A9iiBX02KmhNibAo7tV8
Td+VEGliQmfIxnbUBnC9uLBu2C66M0yzH8ZijV4Vz5UZLN2MuIC8HhD8lT/MQu1CY/8aWzxmh333
MFKOSeQoesA7AmChLYKK3UsCUnAAD72llyAPn7Wy9T6yIBYtpdRGgBvGu38/VlIHIlf8gPGIOYyu
EXQ6ytsaKwzqMWt2qJ6fqj/csKh20XCfdOyje94ixKNsafNHGUest+zSge0jqsdLT0iqM1WL6Csy
Pc4rBPDj9vlR1OTohgT4GuEhIylSteF7YIJRItBnNqm7JRtpUFONk39ulFQhjcdX90KPzg8lQUaB
ifk7DkGZBkklDhF5hMAzuVdGbQGRI9n5yCpUWoZW8jKGP/5kBBaoR2F8EDUhwODw+kCii1N6wNYR
AUyqh/NdG3K50qtUNu8xQF5qINjgK42yyDryGSRMpMB1RT9OdQR6jtU8CwncSvAzl1MsRBhGHmVk
hs7GUmhLAmo1XSgZxSr8TFYvLfTjWTkxN77kikepE4GeRZ56gCdpywU8GuHDgimTvyrbvQt3NqQJ
PwYPX7FgM9PtKEozBQOwNEULashiaYo3g+8mWM23Uq+PkAB4ZpA0BfbFcfw6AH0sRswvILbKn3nu
6NGJIfxp1bIILcljsPZ8sZ5FgIrsxTDq0ytciN67ooa6OREhE4y5nL0zU5JLhs8GDFqb4C7e2EdD
dysnYDNWBjgtgngFAIuHDGGJnHnRlIzhQk9U0214rRvT7MLsvfH14lOvQnkKDwh7evv2a8grxZRJ
cYQGriTJrfnbJiYHiyHYzfy0zomKc2AOr30Ji+x/ohyJXpQ25bqEm2Gq01+SgU084ScwcMy95wSf
BMCoGUuNdHrYSCAZB+heUqQ8g8+v7vUGaDPHltdYobQYpt7PMu7jCjoqe1c0LarGqU82/m1F8TSt
xZG77uQEy8bvmVy6tqGxycUYdl0ukCHFQtEf656rmEIQKVmX7LTW7g6eIi/uZtQe0vJ/T8ZdgiHH
7K0AyMUdwb06m/L1CuxwwrNtA+lJWDgCwiRKg00Ay9C1t0Sc+2jGeOtOYYMhUDdSrJZXZ7rROy6h
O7kjPh0ymGlsRZ1zcnpoTgsXgAHHdQD6qrDoFhB4Ij5+Aq/GTC8brY3lsxiDswiTQr2wdANWyBkm
0BxdDJT7ybAgBHB0hVaPthf+cwvTv9n0VVPsRxeGCYU8Xbal7f8ebDRMG55wXwjtU57tSfeJiWOI
ynbpbs2M10pVaVMX5ifEsHQU/NSVldUXFpjGVrnoBw7VioqIBHzD4ZFgNABduiNX56Yv3nZyNTmE
eSR2wdsrvcVvnE6P5nI4H+KE4aNv6NzDU7X6Yb4y1i5CCFafavpFtFPZRnBpys2G4Z4b5dzxhDQ0
3btgAU4YQtXIwLyb5ZnxJJd0cV7f4iGkPhXJEO9Zu+kB0VKpyMDyWu8lqVChgprWCI2fkfpL0s7K
jCpeCi06SMMQNMnUiG5sCH0Gaq7jP3E5SR0LButVX0D7DbM6ArwKZ7PVhhq8e8ZlmMOa3AGKppo3
gUVRuuF72iW9yan2onk3CV9rdUmB/Dz4iBCaV08LecXnNEqFm9nu7AJ5aibJ4tQPr4nA+a4/UKi1
MBmPBuMugyBIiTElnmJjqutkVmcWwMKeHFvdfsxUd9uV7RNveYJ63YT8mNlP8nnk8fG7uJJJIldd
udvyLynoVF+zOAl+Rd979Xu1JIDyrlUkT3vtuo5buddnDx/z5kAVItGr1OpFK5irngs/IkuEODQ7
8Pi5zT9AxYMdajoCjpGUUu1pQV2+MJ+LsaZct0KsH2C8yB6tXLhzlTdMXD9pZdHmKwk64w+rweDD
vIyHVmnd4TG99I5vPrxVgNUscAGWoJ3sv859mRFMvzHQdOGvUyxWF1ea8PDONaLv93dbSPkGvo82
ZZaBEsXhe3Vj3OTkKOn12oaFvTjpIMmSNgT40SMbw5iPeVGTh2+aAq9FLH6E9+u6NRYvN1AmyvOA
27azXMry7Dsu5C+cinicaA31dfySA4nfcuyPdARDMxgV560MtXipyn6/pAqjffmC3murFP0tdMHK
sIclvb0MAvD0Tp3PL0f/GAyolIBA0v8sF/E9180bhk2UcFSEmkiU9PvTAmqGu1p3I5o4fcQD8vUq
7lNQ6J9Ba3c1rBMk3SiTUUt/0DWDH2vnanJ3OJrbRczaviEatFUt0Z1BNIOx4G3vB61N6pK537Rf
ucNzbKnH9ZvW3dgkr38GIC2WUjEksrh7lit9W+yz90LPERx8uLueDkeu3c4NZaA0ykbgzMq0P9ko
9ORtvQ2tqfKVl0HdkfdYy6XdMbNUKkH6BPKO3c+n6ZWopy5Jmk6HEbq0C5bDr0Q0SxBYOADFX+0B
myRGlVR+bVzn3hH8V+KES/v6hWJ37cHLpRJoGELOxBJpfwrrGtlaM6OlpisdfwjzxbWfe0IafwFQ
kNeNo/Ua7mwqzvwYSwMpbpWG71zw1MvkZGvFrtyiFVRqhf0RsGF21CGx9GXcGyZz9asRWXet00lY
R/SR+U+3uHpjFE6KW6oajml1SAZaYiRMBmfNH2ia42no6kKh/xEDqPfWgxxQxiOSJM0f2RBmhCAS
7t43tncGJtOe/Ndan4//kmOS3p+CbYLGiEFKGAOlZYpwvHmMowGG+516R06JmTMZW7+B8CPjfvuH
xog7SXtSaW9P8tg48S42zB75AEfy1CWM3cE3g/LWu1QhZlClSZMOozaFUfErJGjMe49CZS9bgbhC
NHLVFO/rnVcmeuKvAFhsg0X0fia5I3grSWdyQ0FVipFR8FEt+tHk8gqZ9MPV/wNzTbHY2RM9CsZW
7wp6xmcXMgDuBTDTmfMOblv8seDFqQp2SF5rWeEnhDXCJprizLR5WWC/cwlf4PsBQWMJxm37b1Ls
thDTULsDlh+AVOuc7FZJsjSsEmza5/dTltFwoRslxHzSZQlJ4cPHqEw04ehsWKNSrguEPpW+BtHm
6kr0pF8tqG1gyMEnC0kjt09SJCPBo+C7v6ckI+thcyXScJ0Z7GWo0n/F9ejG5EWHFG7FLdFE5Ich
iwZcmRYc/ybkqC8rqEaBio/2HjX2ixPVU1XQdQZDqa1P7CUbt5mI6IkB5oUWZqFlzO0R7v86aL52
z7+YTToYUB8x9JTTSrPJo/NH65qDe96ovzWU5XdOABgLcLjiFSFw1EGwdoGbXXajY2Gag5mhkMDb
/+CWSbQx9p1ZHKYs0Y4ckUAtQI1X/MNfykqAulx0xQacx44HPizu/zOLLHCAX+cnCTeesBt4qnhO
6Wr/kHdSYD0WIB0kK4xCHpCOvk2ifIa+RI4usJeZhhTpYpWYxrN8NalI1oZ+DOB5MnSjLx2IGIBJ
6yL9EkUy5ecVGEBFZaWTfG9szPW810laUPPpyN0PLBJ1MfeRU3QdngiRSNXIR6cNdxFDpj/wb/Y2
nUWABOXLSV5Dthw6R2ahMr7/FJyKoVDtGdVHAk3TGULCBjMKPtsCxML6AahulnTdzINmfR1gUCEK
ab6ZOXApkyNsJ33QrRcOlthG4Zbg9/BvLETMHafIrzyXjq1Kn9+jhGNq3cmhZy8JA0qLqsrTLszT
hYKYAUatEkT89FCzHwdZnMtcWHrqS2FFKl48tXAQl7/pQcevrr7+4DE0HPuWbjKP5h4Yl2xpuf3L
m9ioE+CFZLXzc1cvsTKJVP/nkqNg34p7B4CRjt2pVObxMXnkylvi2994NAuTK0m+nNw1nbK/tO0Z
Cvk1/GAtunCZPRm6ZDllZB5PV7/hRzdhwk81hvFlxEHrCfiDSrl1i8W5T1/s35PEbdpft2kn7kgQ
hyZqUAPrdu7qhf+ho6REtJEojajUv1A3iU0fCa9QSL/qQze5WioUlqJhKoxAM7lu/oeeIuQEVfrQ
qH+nn6867Vn5fgQEJWOMPgFVCNfz8X8uvJKkW4ANPcg6PDFkIzQy+1+O1CxK6H2/WJHTG/WEhXul
9/C1CCQnVJZDukBMCU6oXDMzPb75d8Ff9m+fqpjmwfGS2jzLzlSwk8tuaEjBdTBjXmsfNuziT0XA
Nz5UeORZRznOthMLIRfxOSPx0bv+HDAjam231oJ5x0BdLdNmzaQNQTQE5+Uc4PTIvqJgEANieaZM
cPF5BROqK8U9/5vfMUQTCrVH7VirTsixBlZKqNuOzouP6qumQ21UeOLJWBONSv+bjEma1Q1mcUum
WeRZOTyR7A7JSoVoODpRs9XjifNZaDjRyDc2mOtxnGBN4bS/y1l13U+0efbd19ITUhVpRWIsKa/6
KRNUnvRbLLwSB5d1KdQBx+XTVAg7nGc0sMt0N+rF1e0iSB+/tMQDPfdFNojD1Cgilp7/9thj/BeX
oyAA0F1wXYKwOdxv/7dxE8XdnU/THp5wD4N7uv0dsZeBXY5FUxyokjwlCixG2e2TKEm/iwBNVqHv
qxCAIGfbRihiz7Siit0cI4OeDeFpyhxCS7TxkKQOq6JVG5P6qxYFBMKWa9A98jWHxY6pElWtQNSW
1KFG7NVzKlUIIWoHtY2ItK36vHwcxhs1D3YpVXCd8+gbPkwVpKNOdRZctCzpTnYrby1TMkwfwAKj
KFF3XVQlkqcjUDDvyuBECa5qc3qM8y+IMIDfMdD81FJ6gvHLVJdUfhKlqabUgbjO1ySyLmfctW39
sXaLt5E7Yef/FgQBuJ3pujHEryJOmSs+DNlzdj/dInQ3fiu7IHeYnN1Go3oTNdPUbE3EigUA6hFh
Voa7IsIs6k0F0CamMG5Mzxu4QiQBJfe/x0NRmIw89Be1EoUtbHyKOzu4KgnbBjpZ2x4DdPXGR9hZ
7cNwWfhZo50Gc4w2C3HKbwhIeTL1s04HWRFCqwYGlm85xTGXXPu/wQKIDIAJ7gCSLtImh8w02ea3
OhXu6t92U4UQFldJsizFn9gPjIWRAOvY3oBE82/r+2BKLK0wtgglWUMSj2CZlSeSlHNmmosMcneV
ezdO7Jh5AH3/IxnerercixDHONh33lvERA0mr3ba+/P+wjmBr5m4/IFWCk7apC8SQbnVz7Ra9GaN
pC3DTAgZbwTyqeiwfR2lNLl76puZYU9Ah4WVcHyBobk1wIeHC70k8l7iHVErl8ze4xbF5FOswEon
vwk8+PyYlXepfxuHwMO5Wmc6KqWSa1WUmtek8pQ5mkMH2fzcDPvA3vRFWozIKrAOkwRZhmAtNfpw
J2XCeMCL8ml8FVUcssf2BRlFm+sJwGam965BDz1mvqj9HObGr920JKI1QPie/iR8jO4lGLdSpuyW
7erK34l4BwhSkG9iMWN1Cckq8MLRBHbK87N9rEDgPR3DJU1Q/AZqRAtduGBcwlp4uPoON7xMjHQ3
IGZu6kk2R5IrSuxGPgO+y4REQ8mshih3KHCOEuE8i9d7vna4NO8zZymVpgNk0Muhbkg2AXXwsUpm
NfHJZqK6plnBUVwnIlij+KymwvNdtd/2yV9FvZB28VLogk/O3f2j6SRqIpt2guVuxo4+rt5tVBBu
grgpfFLo9PW7vPisQgAs+1sEaLAhJnwhtRYx/K7aMce22KMyItZkOtVovBQdBy92XjFgXmgn47ua
rZBRuOr4I12FiEAEkeXnhdIUMZhMctGNdV1Hw7P3yQfCPlYu/LpL74IBjs0nVEbkFeD+3rRxgxCK
FfWfDWVZM3of8GjaTlTbGejqh4u0hZe/YC7izmJ2onrpIGJMwOEDKVTORo6GA2H4cfScAdu2GxgU
jTbATWO91SOcEiIto1KZJ8A6GXKT1KYNELw5czaINHPf9WD7ZXKO8/1vHe7paG6V51A/hMTST7N1
S+ocnDetWjng620TNWl4msdB4dSRJ+xaLkeduuZg4X+y4CiO2v3eMhNLb0UQy+MU2BlSQufpTSjF
H4dUUEHUKrKLOtiVnagfP232A6N7A/JEdAGardhlkeuplG8w09Q1jn6RbtKgzBVBUC1U3dogYL47
xg9mqjvQaIWT4Mduo9Pc8Zyw/F2QvCy+aE2+QlAqzMOHEqZ596eWka6hz42fiXyS/awdr2hdmt27
j3kWsAA1wmtWlYObX7FAg140xe40Ih7FZ8XDRDqp1qjVkodufZPmJHIUk5LW4kH6n5GOzlBjb7W+
mqqEeXFdHZ3sWzkchlRRDAIGdo21JR+oN++OOtpnLCUy2ZVH9rPjR0E84JY9oiCf+1/ZTizJrtg7
RNDK4BJ3DH0n+k2cKde6Fs242E/lVYXEtBxWlKisUO0FP5X+aREUE3x+4JZCnilmPK2r+9pB0f28
BgTp8fOTTbpXbn0pRZGoopX5T9l40wUES2Ofp8JZNd+HXomd2MLw94QCIDK3AXe3veZtBfK7lYN9
4sH6H84OOJ4vy5sBHvPNDs5l2PoXuX0zCVLJK3E7lKTUc9KY/1WNr1MaAa+D+b9Qd/GVYrlW+182
wEGZLJHLqrfYnNUhjPVo//C0/e70w3+gzjPVrgS57ghGD5ljXb31xGcUpKWjDvC1kwiwue2sOYzY
cCiFAOr8T1jZ8N5B/S7bzWtOpoHDqgzVpOR6GOHoHeIgFStuUo++nd4MGnn/SQx/8O3Dt1+u7+u+
CZsuVQ/Q5+cLR8AK23Ah+I6VaszBEojum+f4IjoA0aa26mwiVcdsMmTmckhcX5JYTRIQ5M/z0ECT
bg7TK54+N68FKPy5hDBtpqei9rYiARz6QnbUH48R9hPi/+B6ItiEapSaCTVfxydurxgLvsy9mCtA
GOcSZMR+Ql2+0nypKgwMWVOSm29P/ivUAdqkzKJj5PTp/rige9nuulDG5n9ELE4Q+v3AHYbO2xbf
6taB+6M7gg5wpueZi1e+2fYn+xMh5ui0V3rPQSHQntD1KdSoKqaSV0s8shBywHohTOe6SScUxCLF
o9UvmAx967jAjX5/wySMCW0CZRYKiDCOraygLoeaJo/75krux0U0aLTAJAeIvBBMXsmuVA7yQpkx
vIOeyaDkB72+eyUe10ZoVl/okvON8u8KriqVVxysRqty3yOBA6Zpj1mybAKSou+uVwGRpFy3zopF
m7XK2FdUPnejne6HMln/HYAmXiKRPFk7R1tdu/5b+qO8wp2sXi2QYVGqPXOu3S6Gh3Cs1+s9t2DQ
5r6iByyyScHhAkeyDQS9szL0bpDENAMz3xHJJfhouqsnA3F/1eruXyHu5eL5sz8ofremzWfKd9lB
mftfn7ukB5rbhWUvBvek9RyPENtRgsNjeRQ61ui3EFpnGiixD6J2JPmb3FO3EFcOzFUT+dq5yqEU
dG6oyAICK2/iEfn2VFvKon/FI4KNyEOts4AbEvWxw99ItwuURwxNtfG60Rsb9BiA4gBjTQdh2qOU
vuiksDCiR2JTQu6EbXKJd9DwTte/HoC0pO1XZG4bgQrbc5QgVx2UNZ0J7pjjX9W7PIm9o46DS6bi
ZIPrL6xkG7DQMPGzc4AsY1zbCLavljfAg7cDtYNTrOY4Oe6R2dna53cLR4vLS6LAQyCucMFlw5Rj
tEGVwk8Ecvc6uwZ8aNnXYmYAw1uB2vHbXU6t8UJkY2t45oNukH68y4Hq0Pg37nREEX/XloiBRKK/
Y47nDCQI7jncwGS+37kVPEgpbv2bQtQPjx+8Q8fACYRuz4rHQxEdkQr2iGuj0Q+gXkYSay1EAVTx
Cql/vvpIxWlcKKVhbrEKrc6Q0zWYSVSm6BsSob4XxTM1Lj7UsjpvKy+YCRqBdByZV7vt50XA4b/w
CYn6zACsXfvimfPmQNnLQzxz6pxyP7Z49/J/+HNaTxsAMPtwTcsy/DasBRegfTjQr0QdJlQTCDSx
11WPeeBluEe22p6pCmLG2iVn4WYsV9jZSXUU9WY3iSzwTtaG73FCeH4i01gFQRjVFUJ5l4vML4Bw
zvv1QkfBSzIDf7r2TGyD0ni7epI0RfVY3Wq91dO843syt7lLNe8GyPcVKXR+DiP95XTYk9ud8Ee5
waKEEN63uuu5o7Yomm+rfkj1TdcRTihPNV7d6b5qYIpGVbLyKhTFj+P/lyMnkhrCUrAjPlWGtivA
vsrfXMK4g6IYsOxf3osNbfD/Kc9Dm4FRALzF8FfKvxQ5MQtaZZphDVKfFpyM4/9QrMQi0/Po5sr7
btWr6ClPOI+91Znpz7PHxCSBwKZcZZS1Dy420qiDxvvBgAi41rdB1ojbj//IYuopRjHS8roXyVCk
WX9QT9LPQCsZu/SejtSWtqsdYvE5qaSwfHbShYEL4ZHHUrsqBP5mLACqRw3QYrHGetnHMeQkR2OZ
av1RumNUCLG5c7VV498LoMCRQ2LtxKCy+eA7Agqg9bOPsqstvnofMSg57+qVdngxCbgZxBnJoxCT
sWUcZrFYNQZIQEQY1tfszTsB2br7ErRtvxQgoHjrq0esS98YQ8mnwOCLAQ57oibsDygBxOUXl1V7
haICKXC55kwuZdWcd1T3mAZkjV06WhwoRJ7xpPMhk7gaCg/SMzJYoETSSkP4yqXvkkPQ0dv0od6c
/Mikh4r7cjSQekVvmI8ZpcF2Pe2P6kF9sTqMUcUnaw1Oq/a6+IIqfwLkoHr+Px4oHvQSpERdYYME
5KMu76oNr1EE/xpYKPk2muBpzXxdUE8w4JucWs6JkoiyUQAgeA9VbGaiABPTZGCjoS1mA3i7R9Dh
60XfN9w3T7aKE+BxS9mUGB4PGwnIi9P8GhubMjS2owFbYqZiEBWLECTZ2lDHnpluNjlVD2EHlvSk
vL6gIt1DHZ/lOQlJDVANCltY64ABE6eD5XYSmPXcoU49Ul3hS/8b8Xe6MA2HOiWM1cnPDrwnd+zb
Ltz+aM0nqSf+32jR5jGsfC4s8H3lVXG3RHiFCz0qtw1QZIsfCvnBf/uK7nSQFDhma6NERYLfct4n
znRSKQx3XxHXaorRH5WMBgPtm62AG9M/UazpsT60Y85UnRY+G3YHbB+IzMYfcDDKZ0Z72jjA3lDq
XZ0jQ7KvKg9qlsKYeCcIyoXSC/Ks7BT7sngu0gQEutQ46kagQtKmokp75R0hWWNGeUXSkEYwGf3m
SaQ4v4SOG7haXwmt22ZId7Pz4ZEJXqMMx7mBaXRkrnNq19L7TY4COc/vZpGfLNgSjcwwTKqQ8lCg
hcVSf2RrE9Q4i9/x4wQAZ/L1y6z3GoYIlbkpVxMkaxlYhg3XiwVeP0XeP1VUJNTvb69jSHeoysme
8fWVcOrmOt5D2p/NbjeG45s6jR9ArE1S71vXr8jzjv7r0IapSdvRPjWcTLqro9zQ9nA2Qzm+Vxgt
RMLMhE/XK3VQTPUo/s390fMxt3DAwgC56K8cPMND9vkt6vH6tNmUma7fRZuKyEknv/e1LLtcckCl
wGgeGXSV4lmevLGECcfHBpOMOG9bCC1MNyt8AQgFi0/mJ5IVJxtQs0VwKqn6B2jlFM21ClO63pMv
qo3IvbYKTdtO+OqyqhTR9n9N5wZdCo8nbSod3kksSyES2wolV/uqx3zSbfAIUw2SR+5VS1Icdljj
Sky/ODb4WuWESzEs5Mzn7tOxGhOBgf4zLyL3iktfv7cZ7VBORaVmUMLVdPs3Bsy7ZvIkuk16DUvj
jT85GRx5jqYs1dMprbbBoRCHRhbKeihJKPWjx6mA2ikRf9s4XeogINtrZ9tHNEj1HcQRIC8QXsfp
l1Jinzd8X+rOrgqccNs5cl/eZLeYM+KKFXcCc3EzU3jwd595HJlE43O41DbK0JpDtOl6YKaj6wn9
xjHYkKaPmy03is3QspyaUqneZDGHdrmlrQKpg0QI6JKxe1XXxb6xkIP1XZxwMphgrdlGqKKeKl0J
G0TYFlwaFepbUisib/eC7/fqzAfoifwEBamsPx4MSLUrBf1gO8nYdhaZ855hn8qnFq3Y0X8TABdO
+CJeiaLbJZSRmQOhaIpsUATO5q33Xmqx8l/WKAGKCNHT2UExgoOXU2BZbrm8OK+hF1aWvvHFMtxZ
TY2zqtbZ6tQXzWRGfmRs2t/SjIUTv1tK3kJoyXyUxK66DiJvc4jc2IxItrXR8L0BaK1Kv6EjR72z
OtPl5mzfuHcSCMW2TiDPvFAAtNfaWm2ot8AMVructMEx+W8m+at9EsMreyKPIpEOzokbV2qcnDj8
aw0NxXu0GPLK3YMorgRe9Tkw6Mv+obnMvwHMHERrHSCpYH8DqRzZTqyZ3UkJ8JJDkLvqqzROJy0A
r1zkEzeQGpeiL/6gyuicju7WVjiyXeVQ2PuLy7m5+fetieXBG34XAFgPUrYGWQNs1RffySPIhzne
Ch0ARTcmh9shSvXaP3vR4E2NsUOcVe5LQhlTOS+E3tbEc3lhU7u/5XC/sqO3x+YjoLvdMVnYsDk9
p/kG1fg8mDUHV4OzBXY6TI7Ze7jTIn2vmXFzgYBxYA2M5S+wD+yRQMxCMX/To016uhqgQnkaf4dZ
Qphva7L6A7KwSf1fngFOUzoUctSbOm1jA4LSS7tivurn5X6S44/iXBx1Y+hZHyjv1oxuPZYxkEKh
yf49wxvPcotQUg0lD2Bwq3UFZVWsCAaHYx2AnAVmGRwvuwxAplWEmoZ0fCGdUoUeiq65XI4dmQdI
FX6mfLPoNBeSfzzxd4ePJBekGnJMHULnmW1S9qDtKxdQSIut2Fk00Iq/Qy+5k3tMZNiDk5jcTfXR
CvsWQegJ9VMgpJ8Q/HM+um1+L8yOH4C+wCs16SVmgt55EUqWoQQLWk27hRa1m/Rs/bx2m+nAAAma
Ev4g5MWm7NxMtuytFQVvGVzl0nSrrNO0CQJlCrzmm+Y4nLG+ngPNujJHxQpSdZj8busUgIeLvgpi
srhflvna6f9Jw/VMWGDVEUbXGmBuC9MEH7c97qOuFwn87oln9B7FGiFIDieaELEXYn7+zpahAPy/
oLyqLAi+VPLSq2jgQfEK3HCOCVR4wl5bnsPHv8fc3TmbHg4LLTKejs84fwus/hqSSNAJeXse8bv4
fPh9rFc92/IakelCWa7+WN8wDhiJ5Mc430Tu44XQKC0/4hUcirJtVKe7orcM501TYOLilRglxqAN
UQZHqB0DcQq2xqsJeZS1FQDoDG15gbyx7i3aYUJLXyGIh0wKNYwi96INou9JX1VAr/n1+BRIdTCO
K0alqXqo03joWKNq0H9pRkn5KrmgpXPimam4ONAOcXUl1JKX7vBGVPtnBLFe1DMDTtjMSeV4xiIa
OUXai1ApveIJFD6NChmGoxng0EMu+vKvk/GP39URvROmWY5GpV4DPreSJzu81hTWzQukWlXUSQew
hzZo5FJkfb1MccXcd62PKT4YIjuGr7Fif6sIy046po2AM4U8F63QpQI1CHEQSsYQanefT8N5QSNn
IBrqii6eZHM+9SaC70UBO7fso8C06wxBBI4aFj50k8ZZj3+l5+nry4DgNpvRarjGHkRMQ/W18RIF
e5LONNRrG+OGu1FfFnqKRFyja77+N6PVwkBNXUvcNBCV2GmXdL40RJvg/oCO0vXmxtCD4LHTeMC0
PqcMXOAvvAh7hiCCYgpqzYzOivvapY3v8ombNS6LNviCYkdAd980DjrLb4Er+N50Ce1/SL0L+rwM
z71iqo/UOh9R9yJrIZbd1gKPQMWpUMA/z6zRemljyXZpTk0yLCdgg7NdVHDGrJKZfC61toEz6GxR
10zcQNhJVaMDOP7mfezLilq5U091z9DmCNTyTZlL8P6Si5n6pmspWK9aGJDLhQJ/thWLe+HZkplN
8A1KqZe0YW+/rGz6fzR+CHGESaz3Tt3oAnxvYhVg3YHEUEdfTodDY4oOSEkzhJefm6zrwcs8RNwD
VPgz/imZttSyf9aVxraL77fofqqU/Sn25WgwFn6Pa4bv6ITXu4NIW7bxx2DkyvfYkdhxpHRc2f/0
VaxXZba95Z+RPgoOfpuaH47an2iNhxmFrdrT4O4fenJmVd82WYMIGDBY0FUVq390XaOsc4Ihur/i
dzbmDX76v2l7+C9PHOfXWosksSIxChwDFxAZJNwJwnBRTkvxGXsX8UrWDHXa19AFJRWVij0BPFUC
z5fzTopOo2RF+sucoWR7DTnOJCIGhOPyLGBX8aOKnrhMBxcsLm8k9OjYT4ToTIRmvG+b3LaYR6dP
J0JcBsKas/MP6bL5wcbS8LcVXZYm2NCqUnot9yCcsRvnaGJUgfpmDR9JYPszXhRIPurHtYN+i9Mi
N0paNh+o+Yg5iNgaNWBdwzqbtfSCJ3DlVVwWNONTOTV47EI22TuRPdZvmaf7qRXy5VA84TNvzUnS
G/s7tpnu85J2KWYNLWY6vEs6Tjt/a/oYfKji0vOT8YcEIrsMCugyMjmjErq5tCqVlBL86P/n2aM3
UNhUUcVEH66m74WACazW4lOKD+R7anfxoYD0M/edwsPWwhcCqokd2CqBjsnyKskgJDot9/DpCXT+
Vjk8AScuMru3DwsO1jN3COB/hLVWaxq0N0aVXySLxY4NCneMO+KEsZ9oBK4Q0yMkZJI/JwekQcb3
iE0rveeh90S+AIozDdVp4IwXu5YALCBdRDU4aoa6+u0F6wtC/rTyQnbfMzKGXOcz5AvfYVZ312O2
M1VVXJf958DwUTSAKEKGmd/oFSTR4sSHUNG116McRePYw9nkwXsLrgHHiqKteLXIjThERt8N5CeP
dY65oCWQLO4ADXIvOXKRxnNYTo3WcR4ev96YNHQw9WAlziyl+NvPiTuFC9Yu7bw86/dGLO9qPmzr
EENhAPu8zS/5xpI+kATW0yb7Fu2I8stxLYq8E1d5X95JLQ2m5eUCVV73PLCOx5q8n3rRWBc+Nt6o
xqmTregWXKSSgLpQT/GgGTRg59O7TjhdQnLnsS0SQA9Wm2GsQV6sTG6kSBa0ORsJYlf4hzlKiADy
rSc90m/jgTQXEQPk4eGysjJ3BcvkqUD0tol9CdQMgnG0i28lJNVoVzs3StdRZG8zUAFryEkji2+D
o0p4bqUY0OMOP3//MsfZQqnNeuxwjilvsnWOsJt3GasB8FP1hntNxPWE+a5+MbHBS6Oy/6R5Mmpx
bCd4pURZUPpTOjE1CvnpEo9HD+hhSimYB5bLqqpGmbcAw0j3ox4pEHDbJ2yOTvPA6lgvIcpK/SsL
E6tJaxUdnozkQ8L+XWXOyEdkGEykg27+vxCBsjkFcdxBJcN8fpv0HuMsfu5rYkN2oSTViHGq0ynR
ohJ4bQHzf3oWoAQy8MKFDXK7Di9wVVPSngg7cowwe4fcSJm+Jvdv2YyghR4lNL/QGxD31gbP4sGS
wb5gKHmX8jM9NmLYzZ2el9g8cOPjoVlvxDctJbpGvBGxnBLp43/kaaeFp54WLBaatCNiOmI4h0i6
GpsUI4mmqqsTqazU7VlPyWvUlNchAQjMlQe7i53x2ef47DG4EkYxAoVijsUp+SCAJ4xBPPkuoMAJ
NkAd/P2XulL75qQfykpUTHS7uqCseUCRzfNC2BklOVJZnGdKBomYFkzUtuhfp4HDfh8W4ZfWljTX
AcOAj34OQ2d1Ftp/BVzC1dEoRaYIwpwrcPE1RI4maOOobaKo+L5foY1UGmUm1BBVMQLCAoWpcHXQ
A14hhCrkg8r1Q5CmnV/LOqYAaTad/APWxYD4TKESjKFsUB9YaYs7SUf2EKSXyYn4q0JZSNSqyfQJ
0jOP9kk4xGnrdhb1ZQzkeE4J+3GlFYiWGePQqfnZhM18zHB4WTUar88vP+u0YnmgDZfMDyb7CdEF
pI5/6eOMWXGCIWCbCDPdJqMFB64yOYLFceVvfynq6LqrNpFBVnkUK54ZyywiC/3V6EH3M9+2QBrG
UUvJqCsJ7s4q2230lkJenIi362yXF8d/LlnguzLZv7ryB11sjsBuEkaKfFi7CcEF6H/6PpPYd2RT
/LgqV9SYeZKj4wQ7NekZAwyM49Ek1GmOAuOP2zHtOEqaQljRISqMTXZHNOWzbRyysHhKIE9LJu9W
jp17LRgNdiXWc/oTOsYdyLEUTMDwmQKWf8jRcR2trlYVbUO48QZE7tJEoFeb/iQQKLiEUEBpiGsZ
JWgtZ/X96+fU2IecoUdfwXEUsByqhCIPjTPk/N17Y5eCwf5j3Qv0Rxm0z8/eSxRq3dd13GH9i9h4
Mm3S6qFouYVdoc9OYF+L/8gl288GCTGAG86ls/fX0xijnQkNcN9lsdJbTEb1b26fI2af0UiGH2iw
hhTGUFd/nme2r70bVXHIs5otm0MNezLQFKTyT0igOHIXAVmfdSQz8DY5EHrbQxrz4NgXpLNA+x2j
JPAm88ZGhw6SKXlk86C1sKvZlCXPXoxPzW2Ao21gNRlKGp/lkYivpQBJb/Omn/O2b/0CtdKJVPg8
XWxBiohZEYtRuBDClbMdbOyU93v8s6LMq0C3UkuFzZcovR6hw2rmtblruMLfaDcStqevg8XjUnMM
JPttqIvpFtX3VOI9kdMaIB7/EEW/0lgekvV6URFCCvvNT1+fOSees0YzPDLGnSQO8gk4QWv3TMXh
95ibLz8i7x/QVbU8qH57v/OqwFvj5ksm2L+Rj2TWQJV/6qeXTfI2sEhOjvKwVGwAT0RNLZgFPGQo
J8WSqONR1A8VJHtAO5OHr0tKT9rFf5WmkhQSRk7RrXBRPDA7+vWyX4kYB+wsbsyp8D+4PaFGlSIb
Vp9C8MsmljyD5PxUipFx5cJX9HP64T6mWIPDTAkbFgEdex8h8uniHvTCfT7Hx3e8Jho+yJUWYYnQ
W683FeY/JeU6d2FUrAXWYmmnYoTHnDHJanjXj3HrVPSi8H8q0AFm9TOfQKMgdrAZXBS1pgNqHU9s
7pRJJ1Gv5dvU46LMpnqOlQ6lTq3lIxe6EhihTT99LD1etBp9C7a5qngbkyoPVYPetPa0WLiA42Jt
TyWLY1zblM+5kq2Sllzs4wy6pANw9n9442wuJWyz01Z2drTZrbkOJIhQOFH+vLw1Rc96K3j/InGF
HlQlhq40iz46lpiEJPoFceymKWmT0npjMGa9GvGnv//KNKaaBtE45ab5ztu5GQcfkkjOrTw9ykwR
1/vozSelTMirybhJ6L/e4Pkqgz0U/EaXrE8x3dSsaKEYtZvxTZc2y1mWQwkJXNiWDHvOdkAgdOlL
FajPX6U2r4L76WIpOp3cErIT0MM85sbUD9LQfy9Z7baaERC/OXPn5PQo4nI0YrlE+G5tAY72Pj/R
mh+PLQfbYAawLJ0VktLrpSPtFqvbhg54JDVBzhA6x59y7pQF9qiG7n5crEdmT+ld+OaThZADlOTe
OkR7tH/b2u2AAUhvkYCRtQgfmIaEB+WKfGR3RqrXdHEfbrEthujMUfCoDflBe47JXwbISIDL4ZZK
TA+0ZbWB37vvm11hHRCH8HJfS6tmlSwjm/dfWEGFATXUbXmzCTzFFVIzX3H5ZZqE+8dBQjoGKZD5
eIGWxLV9wXyk8y/RYnWiZEYMK054bzo5rlVSKa5HhkYOCsEb+lkLP0I6W8DvhrMnhqzamcvPzuxq
xqa/D1Tu02fn4oq2r6cx5dV9R4GG9lobOPzB/A5HfG6xGFYt5zHxJku451aLIkHsf7sAlGbua04z
IOzFd4TfP6oDr2D2gCqbHkUA1ArkyUuuyecV9ZjhjpbOhZ5FvTVCGWYnnljtMUUoFLfWM7bvmAcY
g4pfnjFF744eICe9Vdg3N+i9nRv/oBdMu2cY1F/puvPKwEQIjuQtv7208PM6MAsZnt9bEWwhkbs4
8DjUwjkPR/S06pYxZ9bFbxRUaGbB9VFCBiSErlaRvyqiiNomrSYjlXz/Xpsdp7NZWtdvpTtI/v4j
3XY3vEcoWME5Zvthjg1GwFdN5Q1RUCaZM3GMcPHCBBa/YFHWFGZ39sj258mGWnY7BpVLquaxH9sT
G2tw+KEPDvDtHJD1+ZqnJeUGdHAF8fk2zkesmIetwxPY/OFL4jh8ecRvHOtj7mjSKuCF17mAmF7o
NsnEp5LUfxuE19QyPvfRwEET69T+U0GjvPV9nBJm0RiymNKrofXvLKYUsD4T7zRV7/jDsRDuxnqn
KVMTNzUi5ZDF0Byoj93wV4iUHKpwpC/yocFYGySDI+EY4W56fjJtcMJ183jjdMT/rxWfgwNCauFw
Qpn1iDZQdSu3TYGWaH1In7p6EU5PD/9G7dtPslENHxW434m4ig134mv9DMx3ty+vOaLfLARNIPl4
wFBQJze5/J99Mqksoxx6yrvtJwC/9LwSSrw2p2Oekyv3kBrwr3aJzTG7BoE4a4tDZGl81xaxGgYt
Ggw91XwOY94/ioW7VLoLIgdzvnl9IVZB7pgGLUl3PouP3bWzWcV2ecYQFqRqCoYfCh21ydtC8hqq
V0fsbKy//k3mSii0jAHwLzTl/zJRB05z2LeIkBIjMAqGszsa3BmLRgJh8WsxO0hpebIfrv7YzgpC
x6n2jyucpcgHuY5bIUqFoD4fbnQwtrB0LLN9QgKJGndnL8TX1VsVe2R4s2HUMwuJloTsR1GT9Pvo
GCHXtFE8bYpdOcR/TieClow4DlnNHYz811DLtk+dpr99d4lNhhr8Ua67XFpTYDDzV1HEbF93sT4V
kGGdqea5WiFnINc5jkoWYgyKXusCfZzxGYi0YzbQ0Jpv/WmNN3hGSGstP5G6swgGma7CDTklfmgo
rh+UKxSi7k8YrwLlwpjSfLUPZVRbibhColgd0YRs7HxNaluC9DyUOkFaqvi6rVhb1fy7skEX+BJI
6V18UnHNsDEDTasZvxFXuODID1sHC391j6CZYgyB1l7jcu+GS6KO3TiSoYWoY9i9Jefh02cnq3Dn
NXhEfJZcW6dV34YlVOp2haE23I/ZGePBzBspYwPXsXLLmATogq8UB7ydX5KVwG23WnpHZG3NBx6q
jnkz9mz1ULKaTwj+hXKDHiFhjdCKKmYlMo07m5imCnB2IFDDoGxA2qXUIVeWuE5dKOOCyrSF0MAh
SgQjcX/NhwDjMWnxt03a7BiAfKJgf8ww2066ocmT0KLpJ9/i1Wra6xNPcTu5bFRE2EjpBXyYrctN
44Q8ouUnrbKXofn9u4sSnYPX0ReDX6A4oaLvoRN/C4o4RjCw3Jiey3ehyYlbx2ZhEWrWs2QMwLVd
isRJm87ugvLkOQVT08P0diYGhRBGA0x5ca1hNvmZFXiCPpdXAQCNceHVdSP2WQlh68Bdy5Qe626O
3wqmHzEv9Z8lwqbWT+BO1MYMe4FJWhFR+lSBH6fUX2W5TvnOR/MJYgh32VR0vSnCEfiBQ7aT8lmT
7S9HUkSVStWZKjAj4vFhITYuXjxIfNILwLb5qz5bLMzQaNH7PbjYNG7TB/YIPefOt9jixuZmpOdz
32J+dwnWpFLG0GOAQbctObcohHkmynKyaeHHo7JuoDisfn4bo8GcsO3ZNnb6bUwpZReJZWbuHT8f
kxN1XTetK7LHMdC3sVLbojqbdvGdR4i8yJ+vWR4bBAz8Jcn14K1qMDGRvXuj4xel2l2Btw/IqKfl
0TpMcyBfAFs9PyTBB90gq/6a+p9f73+MZG4QG/yLYOeskXDHBdG4QLiP7HbVBxORKxJ3dhOGX8F5
Qnu7iyIg/AhrA4U5q6R+t/2jUs2bUad3Hd1AM7SYUhn5+D2VGMCKGy04bJXgu8wJTt43wQ8+cV6P
rIqX+mPnG/X+1k59rgOsCL/e7EosMWWTTjq96cK6t2xMftbYcq+40TKuzXZ1KUR6P744w/LwfLdm
FsxuWOMRxcX0Z0f+b3WJMAPnVMRqBLS+DY+W41vfcMAi4WEVz8Wce22VAYyceaK+7xOnbR6ReGgS
54J+crypEhtleWuwMI2ZUz+BzNlBcmtmcijMOAY2tCwwsEYjHfwskQ1Ftv4zUIj+BsthpcHEIFMu
aXLT+o93nGUekGWyOKDp2p2odcd+bOi8EJzBPra+romEeWXA51x850qlby9s5Frj+noZxh8PtmeH
aeN6y6RF+i18xrlZwx4lvj52p9bTJj/eXrzCHkxBGDVNx7R+JVxl2td2dbEcGLuIGlygZL3IkZC6
/q94EnGT0iM4TIo3Ijt7ZDOZ7jlxQP/Ut6TWL6brkj0LJ5Nk/UB10HtnXPI2XpTFa4O15RT+KgH+
+mB6S3MaRxtcILmpONdGhJ7HHRQ3XA/6LRBbgCBLTbsU0BEM85NjMUyKx2Sj35g0mwjJ4IC0BOzB
L7IhxShq9vgUdh8aAHeHK7uO6yZ56UsQ6uBhC+lEBmOugkpcPjETQ/l0Uc4mV91XoFF74Rb9TSmK
hCRJSg9ezA9AcxX0tdP+rSoW2eDqxDDnQzRk7iFkBLHzGa3YxzOQZNtp2Xyuqy+RXAdaRwm9oYcf
satUYNHOUcg33c+nJYfXif52cWEuEIep6CnEnP4TSPtwqrMTL3tJw101t2twcejSYvuBU3BjYq6X
2aQO5VRhH3YJReiLEWsHLg4m3wi/mQmsXlmfk2x6LCa051adDkdVZXdl7mnuTFcb+ivC+yrekcLU
dM/ou8LdPVwIQzorpK9GtP6hqsZGkcPi4H8rZTzk8g1/MZm5HOToBliCel0afa9ChW7NxVo8DMV7
w1jKyrfdfaC7DbIKUBhVyXiXVvPjYl9aL6XK7OZkQ0E/5Z6x7A8MMaAVdOLtaCTh8yXllWK+0znW
4hahyoYwT1eH0gG2sRAaC6QJbs+30q7MoNK4r+Jr4bqTwCg5P6hU3/e9Bg/LYlJVs2qAdZ4OwMJM
GraX9R6C+MjnmrdQViSTTV0sy/dn7HrS5/ah4epC5RQcLZW+6CYCbe6YkhGKVHnp1LIRRQZMLB/L
dxY1Y/E6i+SFDJ5VxvHAMuex19oMFC6uU7DAxka7UhY4ImjfZ6jnGiTnf2VNpDBWL4qxIr+KIslb
f4SgygNsIDM+Bz0c0K6uQw3tVFGL8Xg0D52CymD5w2TOBI0wjxqo2vLbmANhe7RKqD+8Tbes4g85
H266TeiAn9jjmxDU8CyIgys+oNhYqwiSIg6xDXneDXVO0ao5C1Wu/Xbz1tUQPR4jaEjhCDZbYKni
G9ZrMCXpwxrHZf/7Zgu0SqtNiiiiOaLqwWbEbH3/k2p5l5KAhNmTa7A3wS1unModJnlaROqAiHon
PRbPWmwlwY1JKkVwEB3lTnvZt+bZCzpKncTsj+z0C8/rXSkEGAYrFI/aPTcaP8gn7dzeRKe9s/03
djLRPDHfJPesV8r6+W/jjxxmDMh9l5Yguk8P4uULVeiJaw7O9eLLIc/4pX7qLOJEpesc92QoEBYI
LFTSyX0FvJKIZREtD3g4WUVR79v1x+Mk0MgPNShKllnJnMbiRAHDRRunHrDR5tE02DeB+DRrHNYx
Z/UrFuElf9jnnANl8D5TyL3We2DkYqhGUKQePcXfVF9WHVcwzQneRc1/wRnY2W9BNvW0gXQJSjuE
GSnvW4ZUXvrMntaeWN4sbx5XpK4xJQGz3QsYsWpAAd6n11ukvhMLzt5jCEEgNW7KIWmoSKM/6Rmz
GpYholG/PLvFIpWFrP1CSlhuN+tsLZ7b/tTCpQh88H+iHRWAFtxy4xZAbWXYKQb1F8hSZw4ujgUb
mdPF6JVJPsQ0Kwf/EdUA9/gN68csbZ8vbr0ujSsA78mexOUQmj23jELsgyhYDaVUFxCVghQjQvh7
52egYBAPlKCC/6pX1ay7jHtP9ani4Bra0kt4Xe0D4p6s82vgsWX5osmTuwFCz/4yoAEWN0jtoxn6
YGW0KmnLWQdHcEcW1cTxO4lgd11OHV02L+c6z9ArV2WNrF3vKyIjP/x4Xg95B/06ce+qF4T20hFF
bd8BYha5slZDXyKMEaB7WGVskFKna1KpN4yCce4R/B0SaG7P/oK4YLUf9grH7A9vJiEdJfEuMgxW
gj20vwrFmSdb5lleAedf/Q8KSq36pWFRXS7ZsWNf5lj9CVNc1ex2j4jhRhCSD9qog4wjNm0oyHrR
ZwsLmY5viz05IT/vJUYYQTF/muP8zaP1fxj9K5hYbTS6mQoXKxcccOZ0SFqVsHveLob6FaXwPp4u
+JDe6TsCseg2km6aIoWQM0bw3xOHEc2Q9KQAuOeqX9xYqSmpviXXqTxTPAJJ4eJJsGqgKeFGvYsa
5VjlcMFKPMD0SvfidTSmLj+MiNxsyD9iZdbvumdaRKYo4gXHCYZZQNx0jeUHfE0QXVf5Tbo7j7Pg
n3D7T8/bHxtWjA6lGWBrUNpd+0kWIRS6p/qsbjKYzMKywkrf+2HhdYwQMFgX45aEknV6z5R7k3g1
rX5A6fxoIGkgCRdQNQ2lhd8tKcHzxrsCDQS9/Pd3TpLk2+jGpWSyuE58DgXWVufqs0P4c8BaADL1
lUn2C1CvlGVbKhMdoAnRahfclneGsUWaa7HClIoXWYMRczmhk3G5RYr3rHLlbszZ9Dn56s0hsR17
T5X2TaQmPFwjj4VKawX6g6t2R+1XCojjXgq/pSFZ5RBIE50cyNKmZmTfttl5DXUJo/29XyL7JXGG
RUFAn+b27hKr/0alObMjhItjewO5HL4KfRTlJdRcVEuncBxebVnD2dgku8DwsW2NSMGlpbWY8KcC
L/SlBNYx7TXiFCKr/UurWMNZm3hzQh6BuYt5Wr4jSx9iUKpv7oWUYu83dIPai0s/j+l/omDIDLbr
TXrYybpRJfQj+K5xNbGbBw/RDAU9rdWWKrzSW7oGoe0ksGqIfP+tCQFX45ISabujL6qmB6mwMDCp
edOY7DgOi49nGNoLsy50ZY3pI/UOeY/oSXR8H8VKpKEaPs6YhQv9bxURbEVpc2FgdxCKJ0/wMkBG
CPKlGMa0ag3r4t+lyWSuq4SzUy5reST5+rJpBI1OEWvqi0Thj8wcWf7bTRTA+wc9uS5Ncf1cb3r2
Lv5Za8dpkFL4VFD2727zEbDbKjypOHJzmH69n+8WC5pO9C+CQDnOX+5rAr3bnQaIz0I+QQUfZPub
qZXu7FDuGSiXamrACJGT7+gGsAc2jKnUWPNREa3bpzhyaY25AYLVVxlz9uoRv1Er3izX1DAi3Ckm
D4uQz8sWT5kJhM0jTS27f1mEifAca7aUFYeLrJB56UPk+RCrDUR3AUy4I67fqK6ZT3EH4OVvD/Fa
kg2Arog+NuJhIUK2nuDxermE4b2AqdDtlBgNvCe0E5gOoG/pi1mWKRMoK0KBEvYj77ooNdyyClHi
RfkrWvn67QDE0kBGSZixgK8talDYwv4+j0mb+vD8e8nMHgRJnNI9QRHFm86YAxSlzbIlKUjUE3SO
S1GUMisV0zZWOaJJjNXzlEDolS0cJPCbUMkhpC4Vehn+ZYiDF0Elbevcf6qUrkjsl3N5jX25PtwQ
AjHdjyJz/SKrIQZCEQ9GINWy9UND69nldf0MOjIQw72RrNAtT4zU5LvywF+rIv78+djHiAyWcUUz
K7bAW3p77Ts2+YGpKl4mAlEoWLy5o8kjnoFdFlrRdAZdDZsdGg1+9gnWIFMaK7o7K4bSNtmLIR9x
z6xLqvVtiNdJ9nkQi2Sx85dcqBxCUC/luNaSXf0wvs21gYLYiUxVXBYri9mcrgh3Lc6QXlpfwx7P
JSjroP+v3GVbGDHvV3V50H203NSTxNqJQkAdMF/r6OfTsnTe6rSu9hegdvjldDDursHVg/rYhK2R
9fSU8zserOHrvtvudk7axiQR6YqggCWSCj0s3ob4NK9ruqcW4rCjKMQmWo6YPFx/VvkEd7MaMrrB
jmnUoqWUWE0AunNVrgXmRO0CqG8RYfbidVSOKK4Ad7OJtLp6QvyCLib0NbGuqwrOD3eQJSAo5lHw
NzqBf4klkmQEkSFOQNjmzKq9mfIjy1HXUly61L/EeLJVcpTU8NjoG2fG53ouC1tSUteA1fILt1HL
3rgQ1ytNETGY2F/VDYyZb88PXwjspt6Wn2ES9EWKZGw6whnCklHCO3rsGc+hheofZzwxZRr6flZ1
MUEeTBVbVx2CGAK2qlfCBkUoM0jQsw4HEFld7wQvxzmd63Kd1cfTngUrSm0/uvbtZsjPuwSZliQY
36ArR35WqyWRU53bKg1NiP/psdGE6LV4zSKbJ8l9p6Ae4PGClMeu4DsnXYbICq8eDIYfZhAlhzWY
rAOhlFNabYQiVoGzbaUJruR9l7jWW/9XFfjWyGbYsENAJOuk2ZMZWxJY8y7O5lZ6Bupjn+DdwXIn
zVOibwHlCWik+5DmtvqCZmifDLRhno64+ehE08UWS2I8392asM5hbzbV2Z9WK1uyonyp3wPojDSG
tUSHqkVdcah0EFwvBcrcY1qXon1BJq8MYl2jiFsT7Hu1qKX/3PWoIzQnTxY2ZqzbxPuXcF/R8U9G
RF/XZ6xK+anKoQun/RgrRA3U8rN9E56vqWHtwvq4ualZP0jLj1PQXg3bxrYrhCjzVuIS9sguTIF1
8AeoCKhSrtQyo+DPYpSvRnuCSNyhURgSL/G7zqG9E/54ZXAKQmQ2kVu0ARpIsNvUFcqNw9WLOBni
h6ZUguIGBRxTiqYlizd23cxyqPnTWZmQAX9rj3gzqsEq8wAp2aX/DT0R4tMQbLoNPkgfQLssyJ+L
vSKc8INgmre9pM+4lEBT76+RiMUMx1kv5fqXLyzaDbQwN4rzNAwY6t3PlTsf7xjhBCKji9o+/mrd
YcNJzjyozwuVWbTiWVqd6IderhsBz+98QejZdfQ0m69uvXSNobA5dAOUdUEKEiuBPzF7q0wFihO0
UXQzQkk5sJHPocHB8Y2Iwtjhi7qnIQKVtDic/NIZfw9SMP1wtYJiacAV5e/LLGliabGaw9mlBmxu
9uZQtfpQH+W43GLo9EKAxjRaCytMmWcOWrHjOnkMdzQ7rVGUpCVcYYdhZSailaEm10z/ZiJQQvYZ
4ElTjQaScWBQqg1GEYbL+FZ5vyQrbeRltpgMY9dyMdxDOlYqXqf51wq2NhaWqIatpCJuKj3ev7bR
aDSKB+aNbgqldJjKUIc+Dn3Ba4v5II2g6RbG3sIjhIH8cwIvNA/lLUnsntPyhgxwhxcXqi0qzIZj
n4YhmCZUbBgHs6Cfpffj96ipdhU3Im/WsjWy1MvukuXe0lMalJh4r7uQxjIEpwGNQIvkzfOVgyBl
N+FF/u45RnhgpfaQTAsiEKId1qjAij51U44gtRO9SJCjX038M1KwNNAPa3WI1fXnZ6sbOwm0+XQs
Hbc5tQJ+PofCihDQHfvz5BOGtZX3fgkwYIclO7PuiTdz1/6XiRr/3hLF6OPAdlULkL/Z2a+KbWRR
/8FLnZf5P+QNc8SmKQFKBTzUhrX9i6TbhVnwMJwp6vSYEVVTUWSwDS0IPVp/H07U/kfjx1qpFpyC
hmOVTkrTaQjalbngvM01b1+Oo63Ahssn2SlyYvpY9pLbPW2sLmQiggDerBlV9qj/XoG6E5eeK9ki
nD3wgXqIdF+gdLefDcUc3ixg3SsB06y4Vy6ipwiBdNSh0FbG9uYbblqLZxsCwQKVgVK86cBWzWXH
rlTYaPV/GDyS8X9/3DvjPkJC+h+BZpN6Zm32lGWQ8VOpJHG5p8GvIiNcorVywEStbK7iU1SE5leb
qYUJcTTNxJeVS+yfTFvzlDq5hzt6jBWZyW0X1hRfjcfEiwApds2FfXmJ/YGOas0ysFVoMi2Sr1WT
V04CYycJBE2oEM3qjMYUWQan5M5HejghvyFwd9E7HnXvpajW9qd7MpIc57fXwMV1IaolZVrHLHC+
/wuQfjzjUkrz7OSz1Hqc9I3bpEF7jmQKNSBpn+K8H5pV54NKwEVjPyGmgVHXUwjJcHqUG0AvYb4I
go2sVFeZvp5+gjRHe++t9TY5WuF0nN8RE2K71BLc43gJ+L5sOMApMqBtsg0dMMn0X4rlxxdgWWBp
b1DA7ZO30iYww+4GRKIJ4fDm/ATbAcjnbWD26lQv+tbCrhr8a4G+JF7mliR9tVZYStbOazJR0okj
3NwADZucLMyq8Pib9sgVzQONLLx2w//OR7h+Ke80Its/fe8UbALOgkMnDStQ/NDuEFDgXUIvPuN0
klcSmDXHLoQtKz/NR2D21kn9wDDZEvkaL4achXKt47aEws3FUDvcldWxkYkmILUPwanZc/8thbLf
YNqC9wZkowFsFZ/IEps2tJTw4NYP4VYU3iEDuY88AzXPNltYOgyyphBidnRQtHImv0SyrXRi/lqW
zD4FF2frMGcen0c7PqwY5u4TrSwV/Yz6KAoZ7tPWxbyXm3SVYIv41k/tvF2gBtMBJ6gN8zlzmx+J
2xOgWgBVZWgTgJMw9yf+QQjzx87RKTmMQ8+ZJSrGFDNhEXd3Heyt1BV1WrVLIHQbm8JjOj9F9ukk
IEgLyY00dAOhbrh3BhXikslIJ8ygkhh4g3P/70K61kT504th7aCtGuwmbXy0xmmbKnA3r1juR+2y
XPh0UEf8vnvICaF//H0TWhQTOKm6Uc44AY1HnEc1f28uK6NH0FWKsBgt7dcsxaNKVmaNMhrUb2mM
0IcopJz5R9TetJzAK/QYkXwSBXtGCBIrs3ZrmoGX6CUHcJNKFZlQaBB9OiWRaa0YY+JmDmJ1Y8xA
oSYOK/kHqL7gb8eKi6t+3rkBqSCLeifRFqPSVLOcINvMYalTaC4/cwCVMY36D2C9hYkUfjmmGsHA
6IAKBrFZLHikIdMizVz7LO75Ll6hVYy5w615ifL9pO7UqrzZZZz3BiYsxa655e0nA0fHWz2K85Si
9V/DhGu32Idq/3wS2Z2SZlHS8XZLd4jX6b5AQBPgSHEWMvYnPqjDCXAmt1WHYg8PS1HU69odRW6E
vaIHKpD7o5n89pGnBIruMyeHFICAAz+ZbefVGasfo7RY1pLgrFrDZJpF97/SPZcBZa3K/ArO7rQp
/srOPDrM2m9mWj4ki8wWRwVGCw7L42nIq3LgNsLz0AxLJW6GNLPwwDoZ7IIxX4BfUQqsyd53k+CA
RYlgnVOUL/iryBrWLVqGBb1O3ASx5Z3/GuCtp/Blu1UR83+hy20PqnQ5S2FVJBnV6AX4QmJ8mWYm
8U/HLGW2Zk0mMBEdWDAxqbB2CjMiOXyQcjEw8UqPL/3vIl14S4vZceqTLovRNOKjK2zM4m69Xrq7
AFWhhpF4Q/k8EI1DybDk3i/rMKl3G45n8YWyvu2tzkKrimCZDmnstjbyGms0Bpods0UumgkuUG3Z
61aQSgLyhapoCNA1D5DFlsLEJY772vhDrp7A28n321p9g8HaIvLYDEkCl+HxqKdiN52i6u0PIXRT
EWK4BcoO1HpYOWIzyelSaCpJ4Jf6ecAs0n414MkiRfL1SxwQC1zDzxqVE6tHSOPykhfPQ6kRU/no
JGRaKCnHKF7Z4+QdRIPvCUAUwt6j2Dmr0Zwdrsui5Gu/4otCBa8i4gkvbMugGUA9RzQKwRhhN44I
qH9XnlQX0rBHMa801oOLVV0MustZeDISX0/99No9LBWjBj8uW+LtFj+0+kOaUdyS64RbylpK4DA4
TmL4a77HPeJGuUz/US9skm2qvI2N0k5FQp9gDbgPHV2uefOj6NMtd4gE+uoBQtOdMwb7KUXCQqOl
zQxhR+qbRVseapkc15gyaD0TcozuE8u8gXbIUOSzn3I3Uk5mxAZOPK9tIVsdnKXON/iuocinNdPW
ikRt7COXPyLqQzBRbUWWMMrLRGaDyVwX/osh6FTbDoDnCq3varaaf0qCiuecO0GlDq9LUHPFtaMy
sbQPFJp+mG1WQmW6OyWaryPDZlLsdTUd1cvIGsIjhuE85Pjtb2jmdB0s9MFaUg7/O+kfLIisQbR0
vdvpB812/RuU+ykSBemMM8Eid7vk2iRvcF8EVb1obIT1lkWNTzhPX5TptiOdg09hdkoBzhWZMeCw
EFzcGs34pOm0jEEVTTVDYOBXaEh9b6ptGslKvA+qwHVlxRViWbArKryQbt45yVVNQel81XlKCLeo
kFkp2QD5gZODrVo50+58hAPfcoZFR/gTbP3R5txd8VERuBJF0rfLcw8HsWz2368cR4RAzrtOSD/K
HBr8qcptM4abFX0rEAdwrZRnl8z/W3GCT9p5/D1cYyNxWQyWfedkUDR92kFz6cwjP0dAbUo7yY8I
PqIMBbKgnoM8u8kutV7MzOKB6AIV+p5XYtnHVFZOGE56MoQFCR3YrhJBxgGHGXlPgoax01369qvz
QLjgN9yIj3FRA13WkdtQovQTvM5cExK79zvsz6banb+GdkIziXy+ZvcNkW72KG/VkcOQGAfy02vd
ZGC9fJOpEUVRg5VVTl+aUp5gS8Z8ZK2i5aNejSatyX8I060XeJbcCdQVjGAo0wUwTZkpmnSrxymX
Cn6/3ikk2Rc86/GDfc24tu3sjCftbICLN4v8pFrgw9oNk67cW98j7zrgjFD2S1QLUynqN9oiqVhQ
sBCFvmmUKHZ1lEz4Kip+yaPK6N9VeMFLqI53E9rc+IZkiY6Eti1uG7KveSMQ2I1kpZxrKorZhvcb
d97sf97Y3ofdmMz1bXUoCQf7ZDCy4HzfKZ4adOd9cNaimctIrH0tzdT29vzMiBrL27nQL/LEoZg3
iX2q5biC4vOCkVj9DbUlu45CQN1lNuuH+B9JzDTMXSJUDcJjWeU5DLGq8wqGRrU0ffALB1DBa6Fs
jAosp+WOqz9hlY+n5HTfjJjs0cZAqjbQUCYljfs+5fxkKsavaKYzCylu4zy8V2Ny7QtW0QE2rv81
VPk/W4bOYElM5bORHa+4Eqknue86knHwxIAmBAN0n7h/4O2EaidE9ozyQpUldaS8gwta7fNgm0w5
SUfTvwHusETba5a12qmLhnzVAnN+972qCZOqRU3OKmVbCp+nIcR+UNmrWPZ5+n3z/9shXNFFs+pz
weRp55uHbrlfE3/Sw6zO2vZVgZPb/Vxyxn6w+XpwMGQ5l8v+ZVsrbttpJnM4CLhkRfyVeDSF//k+
WvH84+bL3s3s2D+ueB1EJ+JF50cKWbkFUF/gzWZp0yz6bgQteClwvRVq0YX5xN1x+PQg+qXImjqH
ZoRBHQD7j9WTWqeVV6qyPIELLWFnUCqZc8DpKDlfjKg+KmuplOaTDv0ZAXs4piBnWLL3mNN8l6w4
DZLkmvLKo+o5+Cmir15RrdzA0DYmOF7s6n4ovUywspGQogRYb6d4eZOXcwVQHCeG11i1+Z+TZFEZ
PskfcUI0H/TtppTJIXQNijIMMn0ybdIZq2524PQqey9P7EDYLCILD0vOi0HY23LzmDk7nYYMrp+k
/0MhtEF66G35iugLRp8XY3vsjZ3bUlOklrx+ehiuibR0Cxs6B4O5YFnSQjyAJw7wW57g4MlUmaiR
7Av7Wwq7OefQ36ksPVbPfyp35OAVQXAt3nLnjiwT20dEkzkhPnKbK9jD4rCvYphZCPwjD5qrOxKw
Xwkkh2xh1IzBneMSFIadIdEAXi9ZhV8hpnzC883BZiO5owb0SDVNR4KsgjQQ5TlIrEw9yPQvmhLi
uB5c2pjCcFFbe85oqASvT9XToQZ30Vh/2NyPP9w27U5KnUr9JCtQg7eCGZy8NIDxu7JWELqFAJ4b
MClcft2XX4MndG04rU+CVkQoiUOphzBOlg0pYYs1YemmZlvQJ2IFKItt3dMI0oLMUq9yrzOwtGYn
wCRXBBGPGQXu+QOqzchuFvJfhzq+rBoPRLTf9HtQL5EUkUwqTAeBvYPWfW1kBELiExmSnnh7nBoS
uLeEPKalb3XLmkooPFH25eh6Icgks/zlxSNQpSCPcdZvWAsjaVQUrbqGPiwXyeaywkLF61FCLmti
V3owo+GAKCr5IryYmTkxuEHYYamNy9h8gQC0x8lCu84ZwdMeRmKnKqT4F3EmC4JgC8/aMtjyLPTE
uNwvHkUMQ1R0snBB/KfG4ugYP7cNPJvNEY9Fx1YjgRd8LwVq/k8LLpQTVHsoVzcnKn+x8f6LgehQ
b6ePdyGGa7lq2WlARbI4nwHPtX1bf2p0NtVmOLIFuREmCevqRMwmdwd+yPdBQ55d3e6Hg+uYbEnC
sZMHoBBxa/qkfth68i3LhD0QICYBlQcigb+TFqydRZ0yuJy/6llm1eo+7vSMWpz6vh1h7V3JTjjl
CMKc1BQs1gdFtTVLqmAis/7F69w5biaWRgwEdWfTbW06Y/FpymI4u6FlMVKo8Mh2Cvl5w9T4/zWA
Dt0oYFz8NZzIh1uZSS9/1sm/pxYsAbHOmRq+dNJg4KFx/2OM+lZCsX75wTem5Wu9qHw/zv7dY3cV
oqkCV9rD9GElr7vv/5DzecadEFY64FZiP1WMEpxEHgiYqYM/J7BxtEa+46SXD25CPwzgqOr9rhKP
zrLeuPngUKaIS0+y2bO1yjdQzWFv6YXvvr0mH0eZ31AoY6Ic6R3eDIirnqZop9v4ymM6aYYM3ivW
NtzOkXj4psqTHG0upnJpach7x6rUXsY3BWwP1w48RBoS5P9lEM8VgnmHljNw0XekE3l2HGHb7oI0
tpW4eA/uCP1DEV3BszDR1RaDbqTV51nAxNEXH+xzrDo19O2TJ8CQt1vxpis8rTxRrVdZZ33RsCjI
kR5onhnkcwnIZp/gDNzFkhBT6IpOQGQNfF7/VJwwGYuEeW2key6kDkY9r0tMK8zdzmhlV6TLDDCs
upDQPV5sTbd1HyL7Zi9MJIsCjQOpo4/Ori0pp0wUMRdC9fum2QlUWSUjGw1iz4ANKKLl2EIF8N9d
yXhk0gfgwvwTK9HkgSF2kd02SU9Z5E1yhg5GqZVsDlqJbHHehWJkHYbXqExXGuN14HBvnvb/CwUs
u1Jn943VkjnQsfv+D+ZgbzTJ49B+Zeo+x1TKHEJcWkszWCgq/J+RMg23OnG7jAJuHNDs2y+wsv0M
/jSYu8CC4utXs+1rsyr4tVdWxHkPtKQIUMBMM2u46Whi3Nh3Vc+VCRhFMsSIRbsuRcF6MzDZm8gn
dvSZZTv9sizzVCg/nrmZJ+6cTvF5rTeJhztpAyUWQZBiLmpCzps6XXvbAd8gpL8uB5PiJ5iavZV4
NgVr4Hx7pt2Pn+WAIDpQZqIXsTyEqzmn3ORZzSTbhNTtQSDJMTPE1YNJNtCkzmHglt+nJRaJNLVA
KAbRA6kbdYmo/PxgHAhsVYaZozKtqUBL0RrwEYJ3sO2g8E60pF/2AjhLxSE5oW17wkrR70lGIHQQ
Miom72kVovx5Kmba77M2DY+rVsYJK5ZG2Cc5GOdp9ss+/MzFSZ5q1hE9EcDIdXqOKdeS1qSlOtoZ
OhYCk5mSxf5C5bgZgMOl7kWvqm8Fid0L6nOPM6sIFvnxwV9yQ+mPuTe8A0Yg/wBL5Y+QJOnsVWw1
s0fA+lEGpE+wX8zZD1RxwJLDKMw462D1/DYYtcXP1tPqr0Z93fJKAo6rnDkS+77zLIocILEKkTpG
Bggk1s2cMbMCPuZHykFCGBDspcOSihSFRpecKAsb6eksVzS+1yi3uma07Gn6QoxCXgRUF0KO5kb3
TbNiI2Bg/mRInMS7xEcgVbBCsRBSTcJObOoDZc9kT1eirY13G08TfmLvttRXrEjq4UN/yblcOE9D
jlDBOj+LBfDp/77Ulslz+l5o+yYCaadObLxO1oZWKKhXYNg/S2HCf4zG4funi/CCiyedUBhnl6cB
ePG6HiYTAISx9d6fCBtLBX+RuHRAGATcX0R+hX9Y7LUnBCiOPmSGB+S+0+O9eX5NV6251CI1RyLW
g1gfC7HeshYoe8ED23xPrvnDESNRGGbZcNtaCZOrAlRdUdlZKNKONlDAOrcf3J23g4WjXqTtlOue
E5Pg/2CKLyAVMe0eVvS0zcA9f0L5AbCWMdN/IJnusvClmrRNWtxzuHApFBJnx/UHI8YEOADQ7N2S
cNNspqdZu+oS1+4cbqx4sYdhxj4IX1jcy1dE5AxfQYIWfOmXfJVkeeillwUCzN9WhR9OoiKboksl
y17UUPloJ1+CkiWG/QVA6s7oKBPSSXZEQZyG8pSXy8aJDdTw7Pq7St+6gGqM9Fj+vZugavEabRqo
EnQ90RivT58J/Rt5Ccb42bA9FiIdMt7QUSgfXrLo80JIF+jYCa9qE9uH4YhvBrwQ22yQ9qtIgsF7
XqRn5vKKfpeS6KP1yhqC4pf9jBm4iuFokiJ/Yv4wpU1//NL4+3bYxoxjeGFA8iZn5HVhR51n6Bwf
Cdpc8hiFP0fyl+vPCwun58fCeQZrr3SSvxF3ZnUefxRfZStn7vd/5Qk+rT10cMN3YKZsMjUh8hx+
FT8tI2yqpBaakgvzpDjQmR1bOi+Jmf+cvAGCYdOhTRVvcMo3xRhSDer1lghypxJNpEWPxbr+3+Mc
rQqiqmEXTsdquKXB/abp24ILPLYoG/VRCXSWe/TjE8ptyced45mlYOSQXPBWJiyCzWs0I0a4AQxG
+VuhhqYDEyGaAUeq1a/pwFMSvv5wsuLKRzpaKETLauk9cZbhh9qAaAtcEaYq8O1F6WY5cF3rZmK2
3RcRrx0bAEz839QiBMUgtnC5gxpHo8lKrLsVKnNIbF8JQ2D67RDUzbB5qXRRmOBArNFibNB77VIl
HYySyyl1kU7RJ+PFVJqWLXvGyohe8ciz+j4JvqkNWturOfGGtmlE8d16DsxkuBtmy25uqBLPastt
Mid1iMNLbHoUq8JnYCLsFVH3B/aZjXtbiZbrEQ74oKbuFHBKlV/um+hlqMqvJdAHero7d20Z/69g
ycoeHQBBFIzTtfCGAgdZRbtZeGITaUXQ6NznDUQHOP7fqGC+SkZdXvojiBMN0A4qtwCMfx4ihkQP
mx77YQPiHfMJe/BoU5X3QnUYj+p7Ipr4A6eKMlnhP06BBfTE+wByywIxC+Rw7DvoD777YdEZ6bve
7QMhssQ1+cXsv8AV8pkn9E6h7BMmlwh/x3M/3BVtngqE8G6MC36i+5IlecV4ppB5+I5VZFwOau6p
VzXhCmh63XuRc5f0a9XNWRYW1q83cKM9BDVKrclxASmTykAyJ4hcR+yhWqj2au0qYCm8wdYfp0BJ
90NVIGIXYdFTXSDGxvEMWG/dC8MO5tkAG5LcEb4LsINJ1Q/fD/XDBuXh4+5ytuyLQIIhn5aIJ4c/
FAqmqMSxzkBN6l0jOkLqKCXUQJWjhCWvFdAOTjB+eMKeKvNHxw4b7sAzBpdyrzg7InJQYa5GR0PC
XylrkyV7B0+SbtRLKsr5UASKCDDCguidlFz5JkpsCLLe8d2tLpBD1HMKskir8BG/LIz2xvau5vWC
VhiyDuW7n0yxOsWADvKk2pCC70e9kavhRvxlBemhFIKgQhj6Daukgs+/kCe6bqAxX84OtI0jucJS
DZamSQJXdWL7zUdJEaKq4eojSxyeZNYO6axrJ1zfgNT3N+MFqMyOmU6ti0dfErPAmJO5eYoqF8kZ
yjaCe1+h4Dwj35MbwtvPkYoroRNJpbsymwsEQiAPSkSsf/l/4+ndTnW+6+h0HhVcvKe2WyXiDA4l
C45yMayt5hUXhrGFjjFsUc0KDHpSFq1uK9D5sShnP7cNza4uTgwMXXep5h2kXwrwuD3CVgVjrp0u
jVpPdwYvEF9MsEX71lTD4ffERq8kk9ozaF/v+AZWIIR/4sfTC+ftPxvzaNA+vgvRl8KfZtMRFcl3
7SC1lEBt/vG0hseuZcRMKP2+qO+ez6dBG6RIaJC8yAXmBgOsvBMn6mOoLeUmQvmXdvXu4DEWcNNj
KCsPoGdaFjyFWIc9FFRobkyvNj96BSMp7JPm9mF8S39ra+sTfTPUNCeLtY1IQHPkbuqXKhmtlXTs
Oh5+cA4oER3/c1GBQg2OGRDYGhIdRQ+EXlvoV9GzDtXFhxybBtj/LccRH9MDD3EGkzxJxkxGgWkZ
N4mw241msLEShQo7/tZ9qlp0Ecc7XR8qY5lAQrLCL11KVKPun29n1HHIN24LMMj9PpHpA3SL9Awr
VNj4DFlqyRp0hPUNsUoFcgXkXxfHw47WX6jblJV3UtTDckTSQIvWOAe1OhM/DM2yXkGleWla1v1P
x6S3o3oZ0f/Nrb37J4In8fNbbVjO/tKck85JA7J3CD2w9lRHXjd5bLfoczv+/r2/q/URDXse3Hbt
DxJhTN/6Vx/DwDtfCHREtKjpAiFUNnPL82ePwRXuiMFo5j3H64i0Nu6/hWUp/PFys/OrG2l6Bq+H
mpPv7kJYD//7R9DmJTIbMBlVXWeijqb7SF/XLsW2qK1qu1b5EO1QQBRRrp94XXXCI2+kaT8PPEXo
rH/4y4oBPDXPXSyNLYnIR1QC8b2KMv7dxtKOfQwJI39a/tTqfO+QdUYBLrqgvMjEPaBVY9ctgIzy
2gwvC47pPVJxMw0vHUddtFyRethgtUYpZ9jFwuR4MdukHECGRXxu9uT+eF2eiwEE7EHWwnoLzV5q
qkNb3IyDQ3+TbX9fe5mOYXPZ+UuXbINLLUgvyCjSqzvmv0ipIi+FrjeP/OC8p5Gedv86fMN057az
q/WCa6RGU6LUejYVKS5PtrBs4tVcVQ96Y2+byw2q3MO/NNUkaJAQcj0ZmuSGeSunvbF+VNSd0Ktc
nivJHFL5XQnavjAwVy+nTmvN3x3cfnXSuPKkqjPptn5CR4oj9HVdk7OgjUodaPlnaW9UfdekQszh
ArCuL0e2IAgWNICe/+vjci0zx/bvkadwP0a+pEpbr75N2pNyVlY5LavulFxkZVAeIdZMuXzhxkbL
BhOAL4yrlUJWgeSA7S3OMVvamOB7J5BVKYWeEYpy6/ClmC7CnRqlsdpOPkLBlRc6ekD/55PIeokT
lsrer5TwZizAnIk/GZ441SILaxU6ffB3iV/1jO5l2beTAmrLGXLk6N9RllLwEkprDO88V8KLL8OT
WgdMv90sV075MV8tRRrYQ7XA5NX9JHF3xOiv/zK9/9QwUhNwCMLOrBBZeGa5rn5wQh2dGs8rjraN
X966o6zycRgu1wQFzOwb7FJKNMLox+w58QOQeEK4bpbCZll9pNJMIdJ+q4HxdEXeco9G1JMZvrNP
hh8esI6LEVcJMQ2hjbe9edTVpyXFcby9t3A73u9LbHdm+LY7NoRkOdOWEruYgF4aL/QgsnJlctED
If0ek1CJmtyJ68PRv6VjLzOXX61uchoyn7Sp7fFKztPigjkyCx8aT8pPzvwbk0zpDSJDMxMJyhKh
SBcT1kSP4BlHLfolEnUMy15JonZSs66jEALtcGF9jVJ2m+ZoCfZUWYLHYqtNJUVb30zKadiJFVUN
O2Jij9tho3XX8VsMQbiqLwvhLdJzTVVx4XhZuVeuQSFJcayLdTiNQyQP5gyqLsLcfJ6+KjGbS6i5
ZhLdivd8AW0krf1TF/WjFFn7aHBdmQXx2KEBQF2wjE9vrHZO5l7htH1KI7IO0qxYPjHnFyLnWo+T
jMYjvEQD6HK4QsoH+u4UYc/N/uwkQExD9i907Xh/5GFNpfV1d3bYyYKtiiFgDeADDaOIv+48izYj
BrtB8ujVagOp4EZV05r+ufq/oyosB5ye0+zBlFIYyl0JeSX+SdEhFPKBPdo40Xou8XmlS+8Z+6Ci
07cbICh4dYSK2TIa24mZD8hfssEY7e8mDQd+CfFwy//5gz4fKp8B871FhcDJUkgHFqvkpCqNx6vF
2tQIwj6nKDUYrBWqCrn7TSrp0lDZ2hEQeNibQbpxG5r8J6+y50XLtaJvKUiGDu+TQPouB/2FkUfW
rMHt2B814mJGqnmsPHsxNbxoD1Ez6+c+eY6vqnzDoHC0UylbTpu6kzmEV+/NQtt/u+hTBoeEoOtq
pRsrLzvyhVEHoTv5hGWguAlxOvFPRzQTGn4tmBH5XYCiZCFyfqyU34T2tVkfqsm31NW0OQnLi5Ka
Xrh75iyB18kpnE1L2EwdXugU6Xd7umnOqOf1M+rdbGZzpCMnspNGmZ6RQ/3FxC15QoiPME/l03sc
mTyK/afhMegzVA7Js3B2trVQjncXFA8Hov7rmDZWKIeHuBtmN89yfyyrHlI1gfMoHLKBfqcjd+mM
EoorW13u17SHpB7x8Syeb3oI9ANt2hy2lDalmnQLDSaSt0VyojH2Awc597VL/0J66hBel2mdt0Bf
7f59SHAn+2yAxxjP/P7IysVdmAoFYCpQ0UDYFbgXcequSTdEk6WsL+n7IFs6Of7AlenxK3nsR/u1
n1y93FM2LjNFiUWJJnN9uJ8bYQ+zNscTpjW563CENtJa8gJlqxk/EX3CdmfgXEC+YMerTRAHOyzP
re0DXDr21lloDf9m5ABnTyEsboQv1Hy0olz5r5AdR6W16RG3LqRnxNDdwqIHXNwvxJ4VGmMJI9NK
XZgEpPky0Ga6YuHb+mJ7LhJhkEwWUybjvYpvJ0qWW17En7eiXmWRaT/eS0usQuuaV1DnQnJ/u5L8
05KqTOpW80KkgcDTJNBxiUKWXRlo9tmQTXIyzEvQ4vaku7MvAq/+s/w+dy8CAfk+Ft6IkFZJiaXe
lboTIXxTRi0pDKe+iA7gC4u07LUyUFU0EPvPwsk/SHphCVhhmCOINUVHUy2FYLDdp3fIF/mVfoXg
l7IsuJSDwtl2EPOKsynaqkqTbEkjoLgoFQw+RfnbjBEI4C1+XS6sZggglAhiplwPKuIUwhmbgAdv
Y17xwCvHLxQz4q71Kca53ufxkhyEWQxn+RZ9W8qx+SskIUbkNTBw5naFdjKGPB2PoT89DrrVYItE
ewMRFIkNjXgryUWAFYzP+cuRRtpySNlxVgGFNDfB4jjX1uiPsMZzVImNhfQiNj81sZBkWWDC9TXb
434DOocoEp5y4HQn1+2PXZx39Os03o5VvLAuYOzleWnPyY1Z9X44mZF9hSFiPSySSz6zk2crrpyr
eLSpTMllSs/OP6p7U7UIhmVpavItZ186P1BHYTuXSBTE2WZKssRp/fBbFmKsbHEzFaLVJNadcmuh
25GXTHtGV1NAKLORho8SmkdE6nJ4rBw/Lq/reWHO5CeTI2sUpSfau3qF4/Z/qEQiIO9WisndYrcX
avTx+uvb8AkPN//coVh8dof4x7lur+l4qdNp7Lxn8mGl2BOSkSnFNoUJq+3Y5OYgOA579Iy9b9md
61MmhmXS4q7LIIWN8JWYSQAhwO2dNMdbXQfLcnv+V4l9IORYFrn367wSU/538p/SRw0yIaLTd0KC
OMA2zeIHo/tu4Pk59+7EzDxnO8WAikn0QlGsZmtzMcCqk98rUnW385y4IC4ITeBu4BrZxf+qSBHM
WcvFnVxL67ErjBhVYbhMYIpVeYF5LMTWAZHSqrdhdYbh12ChqibjckMkVlVzOVbQLo6/j7YhmuI9
e350rFEXdGcwCeM5asAu4+enD9u2vSQXo4T9vTxmh9FV920LBsteHtPaMRr/tG+bQ3IHle7kI1z/
WBV5EBSVKqBoXlXRJGzDSv4vzKsfEfg9K2bmmcxrqlgAgYc2z/dSWG0TzixT1mobaZFbW/AOHUns
Dt+b8cZh8n8UlvaJO2fCcQYirsdnUsGoItt4zRaLXn3e/ysxYOO/WqRMqwGRbnPfn16Dmin01aXf
XXeui44KHWzJuPYzu2Hy6BLUHRgtvkkohLJ9+vrxwKzKhnXAI5gdu0rTS2JFAzb+knpR5glWg3Jq
xYWeBbcGfl4zPFs5Fq1kifOQl6pPS/zcyV6jzaxkUEf5SXS6d59VkCu73p8W4EA7ilkEpCW45qWj
mkTXJsKY+PPHk+RyhnNSAURVjXBUhmicz3FWiFqQRxa8faKySRl7LhSRaF7jYVxRuy+60dnkGxPd
1Mzt5UwmvCn0ajPdScQ0svV1KHHIveS4nE30rGOVLGH2oAQlgaFWLjXbQqLBXsCceXRuN5PfaFiF
cHqpM74Pl4S0V4hr8gpPcgI0GJ6rTx+YVUUzVHfQ8gyiJMnrBFvojnhM1/e43UitYCJeXTd9XoqJ
1V5qvwBLg+UDmFJZqIgym03NdyTu5Ae3ahwLrCLUeRwMUxjf50PAVTMORpQzi5XfemnQPnwllQGZ
TuqZQ1gjI+quDhZZUw3uIfad8/W3wzMQtdYqiF0jStDpDIuBer94axtoHyqgHAmckp133nl4hswr
UVvH8CAkP+fCvINW/B/RV34xhvGe78qEJ4/K1JhKknIP5uTNqUIpe0EMVBkGqH6EDVz8q7jHgPiL
zpIV+LxaH0Dn4+E9DaLhAsWsAuToUx7UYgI8eVmREkdyjpzivQAwEmLd30bFxqfQLPrXzGHpnCpY
8XF79up9fLUlczWV/aILOFSMcrtP/pWIiQRd9SsWnST2bSM2qdYogcEDlz84whYzAarAHRV5gGjo
/+S7JcQM6y/ybZ32xCb5RCMsEQp7CnavNysuHwRPaG6C1fH6cWY8dkmIt/R44QMgw7gqlHoHtXcO
dKglVkvz0EF7ReAY3M5lL+D76zK4mAAXkAH6IsBUgO0QWN7LXR2sy4j5+Sqr9GRievWZMBQT6OCn
7/Z8Uj36d1HMQf11vj2+CuTtiJYP7slAZhw0imS8fjki2r0L+w7JRsZLBhoQAZtoTbXDt44DYfc1
6+ryZqMDSLfoVtioGJI721ivZxrhc52y7xl54ufawcD684wkPf1Qm14sPOh7B1LoLFtqmZOee5v9
w9fchlQ3qPfNZJaRo+CXRQG57urXO3+Ix83AlRUU1F9zflAzFb868T2m/VhSVoXcx2S2Dq38mHxd
JDucxLEwQkKcBy1Hz0bCF0tKSdZpEXCJuf2sVXrETkeR4Tixs1HnJMN2gbSJZ/yBoAo0XidXpXNF
rcsb1MhqFeaaiEhPmuQOtwqtlbuY0TtoXFSSIXeQFiU0E4CHx9YK7wTpX6Xbc5c/cjs0JD93SJr6
1oR2r1elHsyMV5YkEjBtWVsOlRFtNc56tJkLv5Hatzo2IfLeEgDDQW3XXfnqGb9qqsh2QvmtR5F6
F7gRgA0IuP4aGmXRkzH7Ba1OYPSc02nyBagIXx15xIVo2c0ESFcRQ9aIo/jGgFy/ZjhGxq/G7aOW
Qw3AcM0H7YoJoWQt+rbor4xBBSbAd/zDqOoyY73WBKE8jeM+RZfgyM0RZzYIg07bfFEE8b2kI0rs
VmgkHFwNP5rPz0jL33+WAg9v3A4OVet/mYOjEaa5CM3L0e+YFCCVlOkpU/RpNXvJcyvr1zdVQnI2
TPrFcN6cA1L4Moj/15wMMaHUec4Vr6yxZuqyi0EC5IbCUu6halGLiAvCmDcscsl9NJB4bH0nv6J8
181CpdT/vdIVdHKCORMYsk27I2GtN2USVqUsqijw2K6YQG1hJd4iF0EE3exuJVHs9RplMnYrqe5E
/Y4vPr8Y0oEcz4qcWWrpoafTenFG5k1KtELYQKbbMzSxyhjH/FSPnttdKwEH8NskQhRrE95F71iY
pnapOLWy8sNEO/ZjTVJdNCUi8xIG9ugzrTv0Mz/i+ueG663tcXglppGeyIbOw03AzN7PqXuT/+LM
zlmzQPX98vY0UAuu8ZoXBnBvXrxK+nwxcNB5eB4SEGCIE3IOKvUr0ItXL9FaHN0SOBOtqzUcUjC3
TskDXoslB2GkEsZL/1oyMOwOW8WHVPu7W+K3Pi1vsk1tHtDW6HBXZIGxG4LbMZkXi9Jp3NauRxon
LggffsSnlzDVY6aYYP1fXR9auftLvLKG4KatwUjbzVjrwYdwSdWnn0MHbWP92VYUCgj0GSf3jGvb
heFNClXmy9iRkTyU6w2x+o4tWUCFt4qBMr7oKis5PQfqyvWMjfwvoo6KfbKa9UwdIJlHVwreO3x/
Rm+NTBTBVDxZAsiq5eotbkeXhfV7RtuDPsDPzu2bhw0/hgCk/d0iOpUpccLDvHgndR62VRI6B/Be
PZrbxqKF+0GL/9/BOoy1ebfAt14kxTxOy9LZhyJJ9ZJF6dAJGAIZKICZdjZ0lBCMu51FSz+f3hN4
wzK8HfQyYC6cDFQzgv3rkKIEeV5wog1U8VivXlITWNfBaCxnaSl+DJ0skFs2EIrTzLb6b3wQKrgE
aHmvaoblVX2kb4hLxHriZbVHJ5HFTCfk+so1n4ktXhH4m3j5AiQpGjLfsfzEMMsVaCsfaDocWl7J
/7QQYd2miBZ6Es8cJUJl2wNBpf0fxxS/USutFbgJLWdsF4pKnRki1NfieY4xoRQ3anbz9ZvFSs7x
WBdyOoEop5Qa7/6QQfTd7/kX8QwRGfXTSo2UubuG0AjVoRt+pAZI7ExqreJkzb2Pc+OMI87S3bzZ
ocpBY82+ElhntWC6f8Ub6kVgKJ5mLagLAJ2QMT7pMOPU5KJjjXtj/C/RwGPgTMXrCe6qsOv6LTqz
8kNowOEb8TA0p4VOcU+Qr6i61DnUuBoOkzAXT4Hq1U+dBuw1QUZN56rINVxISl2QzDfE+esLFr1f
fvhbS8XgweNjwNfFbkJLr8iUkW6b+gwc8DMJsBhqOV9SOU4XRKCiw7uIrXp2K+QemRPnrSyHgbqL
JU0oFLkd8y5oAmyt8yJucefp/gh3h0hj58rklZol6BdBgthCAKcKtyxAS1wZrhOl2rB3dD7QSdEE
wufhUFK/ADR8PL0KO8ANxesEBueycKNG1ITa6X8dlR/LSo9h6d9ijGTKhHovAKPxDN1gqnk6Eyj3
wQFRZt6ccuNKoN8mF2YzJ3nVghgDRlwQ6xMVNx8+Jnk+FZu9DaAD9efv5MjKHSDEtK3LNQxWoqg7
khhuLXCsy8OU+YFNmDMb4Hi60CAgQVzYFgtZgVxaOwChTfqbZT0EJCdYWXR+DP1ANa5dnKK3b/ie
sdlQmN9rtesFTTg9iCf/Yk6cLVQNcmEVOHuiC2VlDn4dZltRpiIH1rtbHP77Hx2Ygo57HbmadMiM
GsBtMiyk/fX8hzOhM+0rgytlorULfpXiW2/FhOgsgF5P78vc7eRdIUkR4MHq6eTPCutJYYe/HOw4
FHCuHDaATazf23sz+aXFBiVBItDiMcDzmU7EmTRS6ajHU+Zv3MrmZDC6SMFcnKlz1OsY1q1bOmqw
iY3MyTMuACJCXSBLSQBo6iK+4CLIhiXEV3VRF9OHCfheoH1rpSNaS0+76ZomruBZt/SfuuyI6oq/
ZANmAQYX4OKv0YRTt2PRQWR5IEyQ5tNpUGdn2Gi+9UBYVkd6pVc51ga/R21o/e/fZk/aMaXlSRkj
IDn1TsLplHkFVgQSpFob1mFe+rfOr1Q9jTgyKX74xftGp/9UI9OJkaYCZRueKg5C17YQXdSKpLN5
IsdsyeJ1JeuYmtFzmggcVK6lyHaeuEpBT5A+CLPRMXZMm6OL9QxxMO9VRlq374Gi9gDkbPmaidUV
VjDNTK2/cO+Ok+NyGuz2B2PoBwdBUehcrTTZLMwfhYMc87P0LV1JEictUDWukGtcPDvX9K7Pc+uB
9xf5nkp8jaYkAOqfX2VWey4L+AT2TXOK7UdQJAolPR/tHmpWjCHcRBevDpihUXih6LNgP5SXXdNr
OFMOZXiK5uCSCCZY4cXRhhe0tNwKKjotoZXfT2kefw+rVpoPAx+TSCQMBMRFv6/al73ija2IgP2j
PzIyl23uOlXm+EE+Uz0IFhWe/gpoqhNAifgQbM9OboMMDRvpu0cV27lrUr+pJVbgU3jeH5vOeO9Q
cPli6Lx7X7GyLBYVF/EiOvpcyJPwCqx3B8Pt58KrrAUoL+vM2mIeNZ2BJxQ3YHu6vqqdXaQAQqEv
nuHAfRqMwYlw2hJRs7kffXxmPNobakShhZ7b4y46Kd6etWxGywEOP3u6dVYzBZ6zwQJPcUvSws53
yCyA9OZX4EANP2nEldFUmKQr/eFEBChLBU767XpaESjfmcKRkomnW32pw+qjyY155ky2qxI10p9Z
o6PZylCp3EtBP4C3ErbyQY+Z7RysK0XC55Eciij1ZRPrQxDhqYLRPU67jS/rugRp++FlkICHWIOB
RBEEi5e8mzziJnz7JuVcZ+PjBkhKRFSlALxHSctfhHAPPdLVfc/nh7FERyvdpT9BI9WMydEX4lW9
FkFs51fvJo1eoTXkPFSRNYZeZr8z7gU86uCW7T0HKk+tUI0+QFKZE6uus19uOvvz2ZOmPhHreAS1
OfM2a++OWU1DZsS+rHzEKSB8I02UG+XzwWooMeF1S/0BaNyTlON7fqlXlD9j7CdPNRozVSNaPkGW
/w1VDa1gMWKdGgsxl3te/972MlcHwmwbdoygIM/vFrSJFyiZkbnrWJ94IqWOVQx2jCpXZNKs/36v
XSWiliIx2Ka8rl0tiIPTJeipT4+c0KRtNA5WuUdTneIw8MBWX92VFZ/ofkayJGV5KJsEprVXRrK9
d1DlYHm2DG6TmZibExaun0w7dDdUAFe4LJVjyU3OrVZcadhOOfxwGZb+Y7fO+1c2nr97AeypLICd
MOjViG2/uMXlRJh+/svbhHuhij+CQCDD3angVjywBvGcr7IWZ+GhdndoiY4fNagHtGga8XRzlM++
llZY6kPl50XRmUf3kmw6CoNlfLv0TiIRG5rjOsfr/JHNbGhcUsFBoJheRUKaIvU6g9+AXpeYZXEd
zzbIou2clElnzyQ8PhVoDSGugIiqZ2Np880IY8SU4K2TmmsAKTXqy2d5yNqidYIQ31ZdXoN7VCGy
0ZulgUbL5Vb6TaCmw+0bbxC998sDLtfWSQOKCGoMk4kQi2ooZaY/NDj2qVqb8wEpFxsV3MMKSuFS
HOF38NLKcO4shkdePURc2ht8/MDCYW2Xh04XON6AaoHK3bFwLyKgTvOxlgIoleTlH/X6Fex1oqH9
vC6idUsN4a1IEbsGyvspxOPxzKwzQ+n3qtPDFoI7WQHMwTZrKFLtUWZxjqRm8pRtrbIc6wSTJr3m
XlxRkGXALV9UizsJr66bAM/o27tcpMuXlwlQqmNxDSP7pKPLsFrUuFsr9qk0DiPCcuI8HYwjuG51
1vE2G4rFsGhln2nt0bVft8VZj0Sty7EiPpV6Mx6xkfZJrHkGIWdesfNDyLLmNEahbrEd/nFzml3K
il8Rui32bKo8pTWtaAZKo8Io0D+e87CRXpUemJwORVVca7nF9tBhVsTnnUUVSf+Y+VnTKfoLllx+
4cPikwNh4OVZ+P5/r4eYV/7ypMYb3UQIHzV5aC6Ih4CzoobfRyLWI7ZPztuHZpPesKvm/Qw1WDZs
RqTFfijKH1CNg+8PDAML0JUOxenHrrN6EJSXFZJeOXlVgqIKFyd3gHLbyIMAqEfI5J+ERr8Afi5i
6TTJw0Z+FJ0fg2hE6iiWB5zAcEtbd5gc/kaNg+N7jgwOohj0jtI27PnQIiJrhg8sIUEFZzX/kjmH
K/009dJrSTR6WF6molgDkjvzkGqs4RU1ELaf9Chu4zn6L7gy5GckSZf7lllXInquGKBIzakfpAWz
L0ff7MgcQ87phhr9bE+NKrV8fncZoaStfPcEWGXlr2qHkA5yGevlZfdtAWOkINFy7Vp0aIzd6CM5
JsRs2Gik7d56kOxNjWYxpoDVFh2P1uz14GDpFJVQkU3PifSyr7PCNXERbd1pmsjzQmN1u71muklK
2lyqnjYfw9Eb7t2vIVd2R3hrnX9JuNeYRmDHwzeFIrX8SFyIyE7XOx9YneiAxR2j+S3HBQPiJCjo
exvo65FIcKa5h5UbRi7uwGM++4zk8O6KC1GaDhnZCXk0H0Em4z++DSrTKdYOqK1SXafbWlWBlVps
iCjznwx1zHmmdZVhSnqU8l8nkf+giv1K22a5cJU7VsrPFss3kGb7r4vtQouMqikelhmPQdU4xdGX
ly8yxYP1oEA26PeTugdYVqTjMPwzlL9F/JJgiIXgf69QTgb2RLKxXFRxgg2FJpqrlg7r7/FBk7F3
UeAPSjjwaZ4hAo8sMs2CfIvlHpFPCfAhv5A30RA+bHKIBA/Bd4hOn0Ei4Id1vUeyutSGZ+3wwRfa
yamsKi94ELQlK0g4ZjwYM0Ld7QbNfjh6qX/GQpUedp/4YLft6FBsiT/CFydlYRyTNUy2CIgEtCb7
mFn1kva9Mnj8B7P9XS8/4X+7nuBTDX2fSO5VMXKuHeLzTh6qDwERvKCJyfTfWVWV2oHw8YZ9R4R7
Af9c67ziwfNvhCVWuHTP+4vM8VEnk4t7xvHbzhPyZLUeswOPvRLS4sRyVIozCMrfnHEcEJDKlbFi
TAbnNZH7SL5FVnfxCGFZxCllKxzV/eYvR6zL6dFAgQ+Qrxk0UOtpAjs0GWhc7s/5y6FiZfdccd02
xpPrhkuK6Dm6+4SU42uh1FNs92caozGrzxBHUnNYPDxuj2JhXgTjxrth8T21aNEjjrypeGbUunIu
ImUuQlcjIdx31r5GVCvTM2g95eq+LhmGUKdtRdLa4/rRGvYBNhjJJdR2ONqWYbzl0IiqQKMx6+Ir
XqYgHuVSfV7GFbRR2H6ObrZCfbuLeEpxCLWKQ7yxxoyY+B279WIfjt3dW8bqPGI1GrftrHm6L9hW
hmMtKLweaFIV8ZR2k1MeN/2QwhP4YefwAE879ADk5uKUJG16Ov7byuPw5cfJJctujHrD01aRg8iQ
PuVi7MouM2asHnBJTrfeac8wugj7yQWaOhB210uIly+dyj/FD3gnmg0Y4cDwfpSFcRySmoC0zpqx
kO870GBaoLoq6eRMM5KqhOcm0mdTfvUWOx0GbblhmlEh7r9EovNL7i706M0UGLStT951eXTHQ9Ak
FXwEI/dftrlwHSrhYMuzkuAVqpamfP5xP15kaw1vveavuZ4ljazSSRbTa7tTouzMIpYYwgVBJkLu
A9T0A43CwK7VK7+hFKozoT1CfBQVMfCZo/kJBCvugvErlAJAnkKLCmSN6Mfjk6kW1DS4d/my9Vm6
vjKTeIdfhl6U21hJ7fescdXusp31OpVays62ljJK62YrBwtWF99XGoTrIY+nwvDUbp6p2LNVzWAE
3dEgWehHM1EAI4v3txAbXpUrl8sjJsLA82QepxNmrtdlnXdWUFoO4HgvCG3U4oc7F8XW6rw1k7bB
Wuen3ZYzjhkgOLfi34rQu5NY/LqLSLMOysanr3eXGgEUpoCQxOFNNFCrqSgrjnL+QSbRiVJtdI+G
KpqZ8cEsnFY0nozcUFPtTIah1ftdaFaBi9R3QBOYMDfzbQk/nPJMWYy+VfaI1wkDJHc9G40/L8DB
5190sW90eYItuCXUdZWNVOV055YQN642kanY5qzHFFTOFoTuaceBmm+TNXzreZSUUhfMGSjG0jKp
jiwg1EydC7b5QoeVQcTzMkpmIts37EEWeVo34Ulb8tVpWWa8uM+xFveJmIYb0WUjgOtY1Amjviot
yeZu9xv0OE0Hj4biT5goZi/sn8Dv27Dxb24xpmWLNsQx76q/FW0/LRIpNVZLsSYxrB5mxMd9/Lo1
KuBmbnw2PtdcIxC9Qs2Q1827O6PjhrCQrzZAMif/Iv8yR7Y4j/UaJP++lGU6G26J9zEvecMjr2E5
FbDrTlQpHJ2VYDNuaBBcaA4oILoRGUwJwlf6XP/mWEucysUkL+5pMFE7/uYsqsLyRMf7GDTT2Siq
YkJUsPQixLr8D9obCd7EJB7p0QAAgsiT+gJ5SE1BeNno40m12S2DxXFl0MrRag11TNkjU1+bK9Ut
SLhO6Bf1IpNo7C4YW7u75CBnPdpeJOBNsd9BON5JiGTUy+uo2Bky1/oRrDCyXx5dzGbiVuVrNtXQ
SVSTZV1T0geXw1yGYtzM0XERE+G6xgFHtxpnXFXJsSVM/Sm4yRVv102dGR59/uGKJ1VpMhHZdeqp
nmRrVwYAraQY7UaPuVZiR4suHjzwXbYeADGTGOClM1J3MnLdbJMGlxB6cW2HP8QMuyPnLRZ4NX9t
f0kNCx01Ef1ac4TR/iaGDqIn10BIVUj0Wp6/LBMv1w1p4VTrnTm/ZBJBe507zHaS2OWFoOrCFaf3
IspzyAFlOM4DZOAb3YYSB0KV+i7n0s8ZH1RLlB1dJF2uJNM6jurCee1+KC6zvXbtNsZ7CAuSfIiR
czmeMpyh7n7AHMc9tqy4Cy2WTQBeg89gvcsyRtppF/GTZKiN00S/yxpr4iaX4iP4uFmJqfQqhW3v
J8Z7l3KFdO3XltLc4fmjuX10EppFFJym0o3FZEdwq87/Q03QWAn6+wmzsnrWk3rJtxL2rAOiE/FY
MloeKQLpTf1bvofGOPnhv1Ma/23oNiJF+88xXjjtxMuBkZRbqFJI32kbTNbdZztypAb1FYgno4XY
Cy13QJWl5M/NGufiCPtn6PlaF7VNZL9QO4K9DOjxJdlUxfVYvACzXahjqEwXLft/v4FdlEasUjjq
YyKSaRvnafvvrvCm4sFDHc/IxgFnyeJpEJQNIeFaIPIIhZRcqDmBnXICqLBqKGZ/VVL19wpAdfBM
B9NmpgEUQEBeOmUZlRkie9MkyzpgobnP710G6Ro8wSiFNOZ1+YbSva9Jnv1HTnpiskhgDH8PQFNX
fpP0bLspbZsAmYIr/dP7/3OCgYemP2ezqvx9mCWCH0fjSZC5j8M3UEvJnejKaX5JEAlFa6vKniHa
mUwPowskyXNv18Q7cF3bvz+XdD4ONc+DIAB9GCNnMZ+bQoVa3tOGSf8JsTSf7t3ilidrQ1c0YUQy
PtX5n03JfTFnZUbbHkTzpZeH8JgOiLFBUWBZxQrck/PZ1ro1owVuR+4qy22+0cNHKF5/FiP+68jb
qaYqXGBUNR2LTLRWJKGc9z0UYgwfoZrem9KdrOW3LArAfoUdsJgtW7xqLEB7CipFYWGN+7f/6FcA
L4jd74IaBN3ty5wVUkIK3VJG5lKEAw18UaYANcFztI+IrzgQQ4xq1YuUh2fAV1c7db6T9d2sdcMU
3P7C9ngC1cCyxjEQvg3+WGCI1AP0GLsS966fFylPHYYv1lM4dRkEiRozEsCtmUGo6xbfKLG9ifLy
hzPP7z3/FTu8aeUQR3YRba2al4a8zVWutlRzwA73womdKwJLw3ijFCX8/x47TGbNW2QDE8QXwP0K
B80KtE050oShcEKWNt4hLeXELzHJC7dWA/vhSYKLsDFUSi5hKFiewvYZGWrljtmSq9vorPI43Lwb
J6qprhQtbQdqUySheIlKSHphxRfeddaU/erLSx/oCdSeLdHxQnMKr4lviHlyvVFO6MmUbKe7P4qG
t5xZQOAAMuUlWTj9ThoK2vIXc5Xli6aIiO0OMCWIq4fWL8FCW/g6Xb1Jd6Hj/UN2VBzKLbNDIMZS
2YKNscVuAG5h4nkNwW2hmXEX7HgasllOCk5mZAEWrWmQ+pnp/0tJxJDC4rekzBXHBZPsJGMNMjIE
XaeJjUNJf5kWCnFDQt/CNAx5v5S++DxVrYSFZ9eGNQqglAEAjC+xmr3VqAdgi5W3Xw2AW3ZwOVv2
sVNcjqroVQK0FLqyZuqjt6mTrcIKTsyrbehkD311bDBvjWSwexM7meaUBtU8pYRcBhpkTL9vwnZA
R/TI5x7ieRLaL3XEFUBwbmLQE+WNVGiLy//6tt4e6z3P11t+DCeivlKyOBfzTBR2+BcDywB7jiks
rzZnP3pM3hgb4M3ivUCuE1n28xdvNkStgmoAAcKsGKEfDcOkPMpnI/cAt/XUaU2FFKU7qwIhKcg1
u7pMOdgcyukMj/r2hMdVmvxjL/pAQYebjmwvsTilhvfNOZ6n4JFLa9f6BaeviD4ezjTA3kVI1KUa
nXBcpvcAw2Xg5oIHfWG/VQ7UJIw7VE7KerV7NzAgPmA0PfwASnYA6j0ZWK7pG2JaVkqSR5a68RM3
rEH5DBeUMXkiWi5qwHfjArS0w4mLUzcoL3D+vyHLvjyrMDZi1oqvvHDZsSJGg133IP/DcRVUNuUU
7A+RzQ6+UPW453KJndj6Z+RyvMk2vX3VuK6v7unw05zDv9j+/8bSXNVGjyATuRQGwMajwetYVmhB
BBT+Svzub9cIwbWPaLDSEqNn7hqOhZ++B3tOj5XXXL1imTSvDmyJ/k66vErbEKxRVFBtYm/0D2HQ
V9eIoLjuaV52zmg9igM1z4kNuFqRKmji2wOZYtdVs45x71gHlyqrjcFlwG8vi7uh+BmsNCwzniAG
eWxAAoSGDYcvf3l7uZSIQ7LNFgxIzA9SUIzim/N66cGvW3vN6VHNT4AXwqUJHK8ZVdeg19wjimnU
BY8qxmVRxaH3t2XBwOdd5BzRez33Q7tRjhNRn0a1Ql5hgsvnanB4vZwxbAFZLx8Z3NVdTvyks5JK
asH1LHGr/7B4KX3Ur33VA1jZxnKf8WGkpK8vd1uMRrRAwxVxLwFlqXsW6LoNRgEL+ZcdufEeBvZn
oqXjpcwty7X5yC9Lnn0sG+OtiewFjtQkU+KCENOSAMhT11jQJMV41Yyfz5UBLCVMR6k4PRVXsNC5
l0X/G/K+MW5svhWDv5N7v9ua2S2K0J3FWJhJWHYYn8SfMA1miKDxgLp9QYdi9ABdBRpkJwrfgfFJ
CvtVjJhI0BlObKbrynwETtT4jJnXIAzkLCzPx+9khsVToSg1mbb0KeuUZNtRfsTQFlIBJX0n8Rkl
6wEUhqyMwb4qNNil2h/sPcijKdYGxOtsBTFzGNS5sM8PHPxWy6+obYA2tMU0/bJpSJGkJEC4LopQ
pLxJC1OY7PI9ZpezYAL6zzenxd7xQM40Y6jcycmp5VtbwoGQ+chYhIwQGlH3yYXi/vG3sWOBoaKf
81sdzNp9tXVl4r0NY3exmwj3QQUoGTPzxhjFv5KYnqmiV0Dy2qP1QZbOBU77/8AODbteOEyGSY3f
M5+AcwAEMmAlsYD274wMZUhJ3XrjjL4QA/IQI9g77nQyBLcnt9yl8NqUwzk8o64lMWrImC/Vw5hu
YjOvneX/ZD/VkH9hmIM59M8Z3sYKRGc31rG9Grx3uK4rZj+I4up1OKl9F+UoXmGho8n9lXxom1tt
5xBx5NmT2xSCB+k8Z8thXOpTbRICbuSGOBg92eIe/QkDx+7rIeljsJGkMNFjOV01JeVWJn1raL2I
KvDr1yyp8tzPMTwHkKSIxUwJORK3+rk/e3i0jMnAayRZxYk3esf7j8pcNQlDTQ04kN8ZBZH9Fm+y
0ZfCrdsWLPTurZjAKOkhPhk8+m3hDj5vxxP8eRwuYRCBBe7jqRycBm60ymV8SG4IUMcdKW3NYBrq
Fo+CgzoUB55PbeGjYOrB+dB72AlWi/bYvL2bZgdZw+J1movyE3wgfYHrnv9eAaT08SzbGB2U8eYH
W1ehRE9VsE6+byZ4o8/3nGKNZys7wlQknHwazMOfLB8wpiEEAzKRKiCSVZ4YvGzrWps74ZIhT8e1
1VNLPZmTlEq2Yt00gCTK1YaACrfZE9hmQ95FxsHD0rVStl5AZqYpPehEyXknd3U0wq11J6UiiqZd
vyVTx+8I4t3sC5IOm60kejy0j8gny2Cr0jIQlhq3SxqL38MrpUBul142rXNW/b4HmJpKdWS1Bi3f
cziVrBUMy22LDW+kEPGmm0STY0qDBVwK7zwSmqgU7EmZGBeGYZSjljBYGvWkld962ZI2TVrSnmiv
aBodhioS4ACvzVFEzVpQRmbkTgHzLd0cuR4o2OrW0DftqGKJXFiMeIsL+1CVLyCczuNVP9C9Ngm5
G+wQ5Rnu3UmnIiCWl8ZYudt+EE4tjuLKhcNh6MFlDt9iucmhCRDLuVkXRucJ5pE8jg0XLEJL7aEa
P4XBIQe4QYJBKXL708D8udcAXKXX6H3Si8R8b8XZ8iR6AogtpnjLKCItQ4sCa4EjYFFjINuAPgQi
bRW8Xz8fr+3V3NvLOBXfTJHcZQS/j8ck5kaOzoucN2K9yhtCGb/V7hLNjlDzcHvGdzeBgsKhV7ib
OC1UhjNKrFSkO9m9I7A8Vi17Sud8xEZV11OsiT3q2F6pzavhbkwXAwIa5+3KxH0V1CwO1zZGLwJx
OYmWuJw01Ki7XoHmssCLeL8JIzk6gzIo0CDf9GLLsXxqzaLpdLAlskLE2qxOgt08+wUNFrPYuIy7
fbKFGHNlH35wsRURruszTquxXSIKilToGjYU3PTn1/kcSK7YSd/X4oEbGYMAp1QuCSQ5vYVTCNPB
yPmSFiO49YV8qgo+6dtU0g3oeb1MtmuPqke+uriYmfd1frgRg21CF/KcOjmYXhmVn6kNw4D5YoDf
SNbuwaUbXn1L2yuQK906OoNVRiYI9+OcaaGzeSP/1ffIQEVQlvSZ2G8RC3QbAFuraWoGI4x8AqI/
Ve1zIpjsi/KbBA+SypCkyXEwGCshRSQkwzU8YtpFzCK5SgyrcoDEEjgoR+UAT9xKrnTuh4TVhYdp
75+d5qsrlh8XurTsIo6YkdZazGpTPo3Bs/tNwd1f3yz6iUPrL7sO8An60NS13PJGCKUXPmDJ4i4y
J5GNrL9F376tYdk06rguYhcjDK3ILYZXqSSO40ZM4fmSXWYU6kB126v76LRJRJW4RDMhukPBDtHv
TD720vE6pF0+l1X6XZv1ewqFkXVQL/rzAvTk9jc+jct0XWikKk360VUrBHpzGuhvwAZGjSCwo7GX
9rySPOmfSzT1YdGR5blTmeAevnC5WecvaXv3iwyFHpIKG15qmwOjQGz6udQ1wwh+pm3euOy0Q5OE
1gBnxoZ5BXwluUjhKBisbX+hk4oJNAusgeYLQguW1YQWKwY9VEQlir76fmukiKmBUqLDRSEXGx3m
sBlYP/7epvM73D3TMWdBnzRBXq2JkYo2W1QrZTH2tj3fPtsrUhEdZ9TtcEJUB6hxWpvsPVwFthSP
eIFlepscc71B0lBRZXD+Imtv0uQ5htbVsn9bT3MtKO2ENvNa7p1ocAmxtXtj6bwdRXhSDBYhCn69
nuFJpyDINAkqioyBRy1CBvSer3FtVL6louGof/uG3tzssLPpiXfJ3LeTJlaJO3eIn5WpxtkYQ5Dd
Romr0Kku9g3bxz4hMvmEoidAKvA3lvK5ZqpQTp7PMg2mELyci6SlyIi3qex2ascsRC9KUTV7s0W9
u9cRKWCT2PhGL2mDZ4zFzzy4OgiFSEptZWQKOm61O9gEtBVzZTrLtUJZ2723ZXyexMLE/Ogf4A+c
70XpuExM4S2SqPna++F6jmtWguyZw8J7hkYOlVdfHjfmlQZeU8oAc2wiGuU3pMUYMhtQuoDSyFP1
dtcMUfiBkCIbmyhTVIj3jvSLcqnWBtBNJVXA1SMBsL8wZ6iTBOuhKssNls8t9/IjFbYKNnSDPlx4
IvJ09TiI5Cr+J8UnKOJfSAYWhSbxud0ZAJkcU3cX98bGZoTYiSn6/9YoEJ8gWpq9MYk1j7reSEJ/
kyB3MfCfYq+cgL37If5I8IViZgV5ce14WCDuExRNS/Ww7mfTwJHGvFMQKLn4HUcfuh0ApBf6oXld
m+qDrag+0P8IeyalOoibpxoM363ZV/mPqrjrNR8Q/LuSEKzeu2HFHaY/Jj1fWrddNoFCe4lUkLPH
AV0GLKjKxVGXnDt4B+2KjutlsE3HSEhPhdS8y0cGm5Il4pyHyYPTieJpW8ExNrejRKyCLBJwN2Hn
n4Zp6IWFRzCESK/BjEJeEdJKIh7AsnIJXb9iLqUnyJ9cU53RdJb7UadNtR+ip1SxN8ZEJbrcjAqL
xd8J7yvpbf50eh+nSmGFWIswnhV/HRY5LQHQLHshFIWR8mp1lUkXBWi8/4lGzWRRWkgrAX+B0wru
FcLD1lO6cPvz7tyQPzwvODQn899IGF7Ne4vQMvmcmS+DuzbPDgyEQhXfcjzLhQDzCypnL9fKy6jk
Q7KRdsclE/2y2C6PkXfuwJk+hqyePkZCnBxrRIPKMilfXKu7ukxvJppxNkFB2dg+ZK/8iFSOG164
iO/4ZG5wLWOiZdCnI/a1EabtiWgcL6GYGzbLubUkCtARyeUllBpphRQu0LmazZ20dxaFaiStXAVY
/WU65xU2DLyiY0rTwKaXq3qCM9Jn/rpOWZALQacIKFHsOu0fCAJh10CRe4xIpUdc3ZgiuLdMVy58
OsV/fWXUCUwjDJNA2VL0AduSED16MvDCHKcctY28FM+AvcqyrrrIWaJrIgaFUyFSjbdH0IRwgATc
ojBlGM4iR3h7nmdRHfLf68IlbqjjLvcXIpYlLwb5FmTC/j+8p/mYrVZv7edjBOzsIYDTGRL7arkC
Y27VgZWTi4RCUfCevwI261fHv7OO3SLYMM3owSczgL7flREL7wVuKqzi1O5FpoRSIxckiFnUdEap
UD5SFA5iTgNuc71QMZd9ufBX5DGAdYAyC/nfRrJkFINL+jZp7EYeJ1EXzjd+XoBVDM4GbyETuWPc
zMiPDEt28GfN+Wf5Jr748o9q+1p6H+K2lMSu7gdLlRifa/OjImcrAfUOdTpCeI0E+bcHQOK0hvGZ
hckG/wrohoBUb63H6LfqoUqD+ZQ/MxQooBry+lXuzw6+WZ7rIPh4UpdDhuM3dugemuHGK/a+g7yZ
7dOqeioTE3WVyslbd4RrFPlqCNS1lVgZK7XOqqvssT0CvSAiygk2q1U47FNwyIYmiGafDy5d+M/6
/TKa0tJCU4R4HqV5yUE0IToIUdY+Ad7Yieg5WtyElfClwMPmvXJTRcAuiDp3qJ224Y8AoEIbjs9r
A4B7+WIpZg6xV+IgfDEG1rnFdh/0kOqJ5CZxQl6WFpSgJQSODkhsb3sAdbDVUosYmGl6Wf8iVVhT
WkuwBAd8jCvHIHDwXuV47PR6mVrBrIn7vMKPYiDh/A8KDWGPFJmlS7b7PU2n54unHSsMW04NPMEY
k3+kMQcXiJVq5tBbNZo3Dkxm0cozwLcCCAhrz0gz9Dtfn0NjFxD1kYsEFim9ZSeBWzeaI2m+Wod8
IvxgtLFpm438pp6ij/carHu4B8i1oPke3YivZMz2yfcbBmqUIdmWVTjk/YVxWWq0322eDHi/ZMrh
wrk5VuAqYnf1Hv9Rp1zX0bsV1/4HahSOzXye8tkf4HPaebutBF9sNB1D8FvDnmMkWL3c8mO66UV2
KEvWgCzJESFV+QkH0bzKj8adIbhpL6CbTNDPz13AW9rXCuykMYjKGx9lHOfDdqE3/NnI1uH27BDf
Zf+lN2/bpyzygQpqviUMipyfr6A6mkyjr0syEoynQfuzv9Wx8ky237OquktZy1L4ehgHlTTZwoZP
AKWvL1SS9LqQR+5OvAY4nTcIisgY7l6a7Bquh+m+fahHj5N2gFcQRnyoveeu+g22VjVpeRwcq/bg
5jgLAuUNLnuOvpLhRQyQ/wKN0M4uVqjc7r1HF5VTLcZIyzt+hPgmI8G95KB0LFT0F6t2k1cc6Mu8
Dj0nhOwk2+eTq+2mbyqWAian0cM00lpXnRq2SvMpZgSVTi2Pr/fmVimRcjSfK+VIyGjDuszEc5mH
O1N2Adn7k057eDkQWQ1i90pGwqsp4QiVSclxaLmieW7U3YpiK/8qNdvAEwTt25ruxEDzZzHR8rEC
Zm5PwOpR7ULbIFl0RAnx3wEghZYFP8NkFmQm9q3zfaNCnfjKwqxqd1NtKPBqE2iZSYG9lUOKHkxj
CZzq4i23PTnJPjarPxU2pbQIOjJi1sF7wNMOVxhtTouY9Atp3pbplBAh24kzmDtzvpqWtFSb06GD
qGYmhwz1npgpC/YK16U/v5Vsb52pM5dnM3SkZk+LZ9uU6ZJsSWaylNQ9fbwvcvIWrzKbwU278iTV
eUSDC16D231+O5bTBdPpFDuFt/+Gg4cPiTTs/cUjhofKybe6IKhiDFwaesXlepsznQyypT3izaix
gjXB4UbHgC0H3KUKOyx2rjr6KPRDNgcSl1pjiEJ9/DX60BP+3dmvbqGO5yW90NAABpODmE0ykhgp
i4jO9TdnZ5pTyCn5Mb+tlqJ91wkkzJ3UNMLE9oo7ksmFTi8Kvfdyr0Rhza1TiPeKF6fd8U12rURD
gsz8JHjoZIs/o0tpHTd6+D5IpT3tyM9Jxstt+6w/P6R83ML4Sc4sKiISyG/ntMkJj1BsSQ3zokgP
dOamSQVYEp1Zn0Gj1yo+uWjLLnu69sKjKtow0uwED6ToKk5d9bAG+FA995vFhT7fZr6w5H5c4pdV
UPeYiW/ztcMMM1OITyf9wlo6RLwX1qE0VYmh0mo5Mch6AN2xCwgfxxjgMUexHMtkJ/v2iSZfh3cY
YEAg4h/E/zKnS55KNJ/Q0QpjB+slsusAsN6qBSrjCXDxV3HRbCtcWjN3fAKn2ojmzYTsoE2XgpoJ
IS5imrd6dsO7LkPlFmwIumi2mXXu+uzjjrKCEXiSUkQgI+5Nequ8W07ONnrpgTckvwyZBvmDEfrt
aV+y6Bfs78bvo3jPe4zdS8o6F9MQ6AT2kqffOksYKEuS7fE8jCoUTXF8bSLgmbMRRnuu9oXKZOVn
4O6ieGyVe8VRfa3CgKmdy5LHp1BmvBrT08pM2nZ6fsenka9/o2S+0k6AhManvELMlOhh+GaqzPWY
eWqmhQsyKXXMQN2VKWzTCqQqOBgvMmd8N70QxRulzdHQKYN8rGek7dHI+VgU+ReXqOq5NLGPuk/b
jIZqO+XiIMi0lQCozAJMTi12gZaFdiBb4p3dV/idI12ZsL/n1hqRDTM5XeINDHNmSjfysNLe5/yS
qnEoRo3q6Z0t0tuGu+eWuTT6uIMsHg9fC3/u03u5QMH/6Ix1bfOzptKK3sN+NK7F3Wcemr9iioeP
taPbzXvbcIt4zjNeJp6TdL45sld2SdN6xUNOtcZ0O0spDClswJwM4Cn89Ysk8VScusIt5lte0UWE
PxA30Ic5BOxwQg/qJsGWu6kxKaiMhp5HQbRI+MMKn1mc/Z6Orpox+pyCfBM2OaKxpsXFRdrebkI5
u1COMzpxGx1HgYyO/qgaZr0tinL9fQmy2W8JwSMrtxyshvLJkJDC3m92/ZeC45JLnrd4aTYgPFRz
G0Ay2qZa4toF1ydU3b0SZelyoo86eGqoBcVR4SAkqKM4FacoJJx7goLzeLpEYYlamL4fd7x7uQmO
S5oJUROHT1D8Dfx8v4LXJCBCH1uFTZBibHrghgxqx70xYV1CwJDmW0RRjTkaq94yEvrSJYvbs3sU
bbJM56cHXRMBmd4j7HRNNBC1832b4grA3IqNcvxl/wNTg+9JY/XYtbuq8cxstrs/2dhjx81CrRM2
BRTu8aOpLeSGwznudhvn5PDosocdSjhbq67PbBssx0aAQj5Hier4LbD4R8pOaG+Z/mIx5Jk7c/aT
WGoron069V2DySu9Zhan1Pkr0UvEzUsEBkaXuBkdaRMnIRBhb1iSKPtOSCIcl9v4+1Gj9FDuBtd+
Ymt8sQ/3NBYo+bNmEf5RxByjeqyBsyK2K7BqjhbvcgOl9sswT0wk2e/PD5FG6YiOCh0YvGSakSRm
KrQ6uMioDa0kgbbs4mejTa4NoZg1zpTkxzs5rf7XcintDNLiDQywO6vDd7xFi01En6PAr6ChDzIk
jCsgtIVI+9k+dHGG3z/1yqBHp0UE5EIvHZU9A19VU6chDUoKjP3lWbnSWW2W2PXhRClkDCfJ235w
iPP0lHo7wlpy5qnjHikXxXe7xqMWlas0BIUrNLyn1tr+zAmICh4nEpzEJAuO4Oq1huZDGnLRv38/
344+9Z7QX2U7YKvSvkfif73ZcCAW9aO8K1+7ZoWKBEBP2hsSXi7/hx//eY+M6c1Hu8GvcR2LwmyG
aLtE0U9uF7D5cL6oETIa0VRklRD5xWJ+Vwa0Lw5xvxDMc5ahmvenC6ynxN+t81/mFSNxav2zBHzn
4tf04WPQAUWmwyXDBq0a4ATMBG4+zpaJkEyTGGtOALyIgdMLaM4VMTAu15sIS/oyq69V3fqd7o1a
tpeEUWe5ZOtj7dqLElVzZCzBid0brkUW69qk/vBfZz0jv325RyCT4lfuGB3nOozUyeC6zxEEx13F
aTb+cc//tb1oKhsWt+5m4b7hXNuRODVNpUl7ELKBwUVGG/5Zm6TLEvhUk6SuU6wWj0BDuWP/8+Xx
PmC5gIhpmRkj3U9JcORlgZhBrzc/HHErIPnl1AQ8PDSB+5++hiFTOsXcx4JNCMlKotpzeOG4sLwz
IllBK4kIr0ELMOnEhzFUT3Wq921hTUU7w5gxprXRPnyKp5qTwxk9ddB8dDHBuc7iPPOD/G8Xl9Ur
UKR7OdG+AOYcb+JW7w4Lg0iTXFz0dDWNvEttEBfwrpoD2ZgwTvDHNUZ+AInpHS5PxNDelJjGYd3O
T9Di2VVFKMo74c8F9zZpZxgn3nDCdcnaQIcrmSJDMJD7sYzFYmAE7OPmuy2U/02lV3hHNIHtm3SL
m/aahBkVic6bLGOVnsAitZ8SebkW9u5+UXRV+C9PHpUHSI0QAEYZKYaYYvLA4WHCHC98pJiDLdal
O6gKce9S2lQssfZk3aiGXd7b9eLAhGbftUH8UCNnkezLvaFtc5LjGCzHo8bZn5DQKzODxORlbue0
UPGiU6tKzJVjG9gRPLrRAFaUmnpsdf4hLgR/AUFPYImT9vgoYvj+opTDFztjioaOjENNm3FHL4UB
2FTvDFG5mBBFmHclce0nEyghvYG4HVd6nbk2eIJALIPDxM94w3xuMgsO5GuKtww3GqyIe9ujMHT3
1XV7W+D85oOGJ/dI8Xq9nULrFnkEUtaS0mqxGdpynoP+w7gUEWrMaeuZMjDjoNx5CX0ierDRVCPa
oKnYhwhqFnCri9i+UN9TD4VPMuN5OSKOIQwdIvKyUsJ8dtEW68tkMnsCTt3GBK7ZKR5n7XGyVLr0
6961ml1bmaAqQLz5xcOU3z0yj1aFUETotStTTJhGqfc+qAGBL3afqIvlQIw6ihoMFGI8uFsOtrLO
s00VE53BW4BcGcV6o4J8RQhywZZvbtkS1S557c44sgsLz2I+ThjqMYiG4MipiSkVvvw0MNyDiELo
nRwtwFiqmwS/aR6FZSAbex8VMz9pYiE2NbQrjgoI7wByfQvcF1xAVJ8N2lJY76q0LIqZYrnCtTrh
+K+O3E1i5SK+BFs99EkF8UCTDlqyt+GP18E3r1IU1DIwqztbnlcyf3fxoB/0NoNxc1+ZoRq5bVLT
xIqF8LBmBETdcoKaD5bqJvheo3LsvLUTpxs6E0ymOtpEVEYo7T/37FSlE1W56QevCmE5ivelSktk
zadCoX6PJvuM5qoy68OERCoWp5Gnx9J5vbEhVowWIA0qRHkOouCHnCUQ4xpTczn07pKKXrWG1706
4Eem6d/6jfJPBc2Y3wKany7NDbT0F87/cu8IniyT8FwjcZ5MRSBS332FY7Y12vW9u25k57m4Vp14
atBpZUDNFLhk2V/8fqhu8ajckAlZm9tjOx7LG0Gva6mOosrgjbSli89EEGTJGsy0xhgun7NXSBTG
CuAtZZCpEmz0exUpyQ5XG3Ge/sq7RwXdhTjfz8pihdiRlvKVB19IaBCVt/najHjRACySgnWwkecv
zmYUSFneieUXvqB2uLfFhCIxs1qkT/wRJd719GB3Vr5fAYuBZkMzqFPywSzlQbxsdzuNzWIPIgbG
K9FfZaM2jqELvVXFbpQZ1GDu1ymVs1thNh8iNxxeys31mCesoPdA/dZDrNcXsLsUB2DX6gc1Y3vq
MGreYkuKnVXIS37Q/a//bdjgkNFgQLZOS0dzUDHknlSwcAQBu+A53N+RTkDjEkPzOyoRL5haQASW
qhCrP+b5dqGPXjiaC4dhKeJHDS8SuOx5WUeMiaZuWzhN/9rCX4loqqzhvBTovDNWfANSoAC3VTM1
WPOXaG6XFOeX8Juz+vAtquXWTuaG2cdTYgaprEayconUcf4ZPhUK1csbU2q17AianQ4Ln9AEbXQ1
d7gSCFxRgAM8zP224YTR5Pp/xG2MDmhg6PPP0bF5Kg7B0JIk/577XevjG6KuWSRRfGj2IEjP9IUW
ksI12ViAAwzilhrVvygBO6lG9arUyuvsNAyktlpMFfvxEyuM7tJWH0CtbtgEPz5bJoEzBFbu161I
6pUKAeyTAB28+W/3hrst38WjxNRoRwbS4OLIdTFiKa9Au8qZn9EbGTpNQg+j8Zx363wbMr3nzc7j
MqFi36I9QjqJwZoOA0KrC8aUa7lyneweT5CgzpKaxnFOftPsb1C9zPVUcdNz42MJ7PWlEmTaH2/o
VQvDnyP0Od+QTMt8pcKpdgWCbWB5/Ejrzx3GUJWNPoQUqnqlXB4OaUqZtnGa4X62imzblEljwKmf
fAwwiUecyzYuDhB9jjFFuDdynkZaycyP3Lbyn7jSSBlL0wDt2alqJtK375zIBKwe1WAYXYBhl29F
LpXW+ua/VZg9qQUPBarey+/GITmBohnmakMGWx/nw+fvohbYcytj/+tJA4OujH5phkjLIB0lyGtY
3GjUApmevtO9qBdGHOMpV8mEenR80T8GatRBrsybY97e22pM1bmO/bFehPDRi1VAesUFoAa3E8es
V1T6nl7bkmYnV9Ro1LguGWHIBMNUhVrsXb5yNVc8jOposJKWxT7Ljrd1+MU6xuC42S3rvK2oXJ+w
+m88f1C5M7pOJORoFfvzP+gaDdvznCxpVdb7+jkvhIIwa/VVJiLuyLur4muleq7d58jfne8jbF2I
01nrOUNCHnqOuCZZJ3R+c58YGaod8k/q5MA3H/Ol61IT8iLSL7bXyZUHMvrGIIBA6sR9aQb4gYde
4ny1A/Kosp6hluG2/+DXWBrex4f8Q102D2LhfZSmjxeX+LUtDT31JOF0fqC8fkJm9GmW/0fL4wI6
OO1rr0UuaywJicUtyKT2O9AfaFlMUU+izYgiuOJm5kX2M2NCUTEKYuTjALipV1q58pOHPEB6uAPR
DCDdSl0oTB1kCBmZ6HO4gTLyfx5Qz18H72HTCiVJOIbYpSCgY5AlMQLGUu3c9BRgymNK9iJu6KOD
f17U0N9y6SKijhUppTm5kXY/p8BLQGAv+dwQUZNNREbUuhNgvBc0mbqaSHJpHEV5QgjAuiHqYxIs
9gFQ/mtgIHOuC5hwPKynL7oFki0g1S/P8oUhikKBGFMUqUQXgBUpzWtboNc6J9BlEV7OxiEklnr2
3tQiXVpn6cIOWv8TFwb6Za0EOklxZRsUb/SXCX+IFOgwi9kPE6UnX7kIWPu8YCwTwkKol+sCSVra
77cybGndKV1dKKIFwwa+99Y2VQwoGRJJaecQ09JRevVcF7xawshoqgupqYj+2ygcG+65+vOB9Hjk
d5WKs+PIZp+AClvhE86/EHbcbfpKhnyw0EFmqe+vQdXisIFiK0xrW2JsC467LFd/HmQMLRwL8qML
ndHVH341iN2umZ3GqR7tgBLKqs4Ldc/fXcFpnzKnawbThhJWQW8j+zYozYnYuotyUal01ZDj/jc5
6L9awLRTP5lPfFDqftqSEGbuIQwPzGp/Q37s8FU1k4SUeh6Q9j5Zurp4s5aC2eQ6l4jp9bbQqRzM
LUcvq/h/FwzHg7f+Ri7bigQnFYgonTHO5WKVmJoE98QWjky6kGTMm4pEBn+Y08EU6jmjAydrqnCD
BUqKKlHHp0A5SgERWOvuaCQ2PF98zwnaQFOlh6w9mlTR3VSDP9CM8avrs2gAHIyDOEjbqhMrV1Bf
qwTYa5muDhYp+Y7Ztcsx8DcG0x5/x2+sVKampye1tsebpIkzSzO6oUeArBfwvtAizB0S8pYd7x09
D5GhPkJNJD7CGw7QY97g4Wme+FrrbC6MKkNP/8BVRb0hoGx+iCQPsZ1OHfCGEti1RQk0MhLnne5a
21gnTO71QcU/iHiBUCOOyMLXf+it7XEMrYM5BXcPNVLyNgEeLoG4y9HbO9ve5qrIJVJ7302fhso1
NgHQRAFBTC3hWzTpRDlyn8chLWRlFShQQtxX3NIxF2fPdZRgZZ6hVO16Abq76cbuUlceOQti/5PR
/syzPDYUg/lIUc7IPAkBo/FFUil8+8Q1gjcwsGjRHT9rkdbUDOELSf98UoB0KtlHWE1+gYlRkeYQ
OX1aLWUaWZks46iS/wSFLvL1lgjmVSENEnKMNXXfMMxGSvIkRVjNnNU3VbLOsbZwYeDf5wToa4sr
35zu2wpyB7cX0LUzDz/uYyKs+dURyFO7gtdUiMje2nldLleQeK7F5/a8Bivj45BRLdOdfiG7ln32
vqqFYqCRmqMDJzia5p8xPgSbeLY/sKKdejecA4fhZzTANXoVSISBi4jWonzcS3tXwyaSRxBhfWit
Wb/bws9Wd093gI6v1mfzxQ1rLlWlirMN3X7XBXlEBRUPFd8FwU5nBvBq8eW6dRwWANEr2TiXvxxr
qTxeqWenIavoxvZLj3Ri76xCW1+DUWLrJBWMHGZDQibQNSTiNMIMAvSZoVPna5KXEmbpK+DH9s5r
fQOeF2PxFMlBZayNrmAJTRejVy5kLAfVljNui4VWmhA8fnuDZFSCkaeWxPm72G30kIet/HXJ9XLt
HFisMn0X1mY2v1Res3gnJSIrdkRfwXVOJ6tIPm/nnxzzZvvS16Ykyjb67Tu6N8EY92ev0mn/WmH3
/EPoU3iZQLxu9sHZfKCGAMwCPq9YE9AmP7B5BuQegcqKUWwX5X76U8Rpk6f70cxZtDgdUvvw5Cr5
mod7V0Akcu7Ia/PNy6+IG8IawJoFXx1sKYSsG0ET4TrK8GHVaSu98NumfvI9EJVJ6N6p93OWefHw
gF7dlA/NZwX8ilxU4xLv8M5owJuyLTYIwAeWcndb++UyIaaY2sncn5HmLfXUiGijJDmX+5Wnrwhs
JLD65d5IEyoiuOQYz1wjyxFaBHFPwa8qnlV0V5CBd6We5Ne5HhAFn1hRHkcWmveU/oMsiPMv66Im
UhpE/CrDVv5XK97abeucsBYWjfLXgP0P+VfQiM0KNaaVQ3UDhweKb6/SVdvjAnojEKCA7pjCD71g
gV7WsJYnKoxBf8RkJtNCBCmdbtOqdYAKv2KWsjUfFNxaioWygMgBZ04PL2oekb/jcr27HKKOL0oz
ouD6vNoQq6k/mLu11xFLHUhP6+CO1G6YdOrciKUqdH13+XjKHk4N5/Zx74wjNdzvXdlFdsacycgd
HGkw2mkIg5PcqnkLhXZ2JebGCDxUNQQTwnof+DNcCuBUw24pQRBEEtpnl2m5CFzEhUXkPIMIbc9r
v9REuzr3qX0enRlntYD/1LK6Lnt/9CBXGjYcFpl2AkmCG5B2gePH7NKxqqrdBixfATQ0Ujg118yC
cjk4q9C4wKPKMxAxaFJeJgXzuQ7cjq42CybyRcoyrR+x9hjCeLGHe6yERQ/RbymliJqomjxDDEnm
IcE6qOd50xWDnI/fiIRf7+68E6UKTWuoF4soAbCQ9ETwoN1FnUhxfuMEh07DWxdU+XP3F3yn6IUF
ElptEyetitWoACVlHGxpuyAquhflUx1GUj1swZX/q3gy2QBbLJ/fCpS/zg7gYwL4tQOa3LjSdRZ0
voO1kLGPIFvaF6w1QH9m1UdEBRCdu3UyT78zXCS+RjMlYcanuDU4+Z1xH9n7oA+v7VZZYe0Mo4pB
wxdsPSkzSurzzIuyeQHKF29pwNW87cz+ZuR9A4aeSZ2sdVjMU/8h7LI496c5PS59SSCSepGxS765
qWA/8WgXddmOFUiO3X+2+Z7Nn+Cb2SOnmftJ1Ns6SOjYOXAHkVkci1F9KSGw/hGpGia07KUvHk2O
+W9WeXhoCG+dLPwsX//nvDFUPw7l8LGp6c7nVlL31OJ0aJ3LJs0igNKsfZ7cBJ1xDr1+sjNx+dnd
gxVPOCLRjRq1jIrQXrNWWXLJNLBikGD7nhBi+JajoeEZX9+XuUDH8sOJPVN+nxtYtSnaDuf/U0s6
MYMov0lyO+H96jqQk83xm15f8GbLeV7cquTxb6xYiXvTC2xBobXO4v6yXzzaRjNzWEee/8XnoMTR
QR3IVzUON0YS5kXP3pRNVGKENFaUeO2Bt07UKK5kJbTJ6wKTYTcRj8lA2sLFvFSE2x7qnxkI0c1D
euHKHS5TfYrk72Tpg3OV4YLsxYX8YsZC7rmTz+EO1pFKyzqMktD1H1+YQ+96Rp5mZJ8IkOC7ht9r
fEpMeR4abJ3a0H9S5nXZqi+c8eUdlXWnOL+Ch7TqatPBoo1Jr4UytlcY35KYw+dzdx/SR+X0iKlI
uSFKyQvIj9IWBMkSry30wWSMOi15Ia35mRvFLi9e5tn1PbebNL9I75K+iyB8r8pG2cWusMn5Ah6n
sZT/Ku/T5ZsyNHuOtzxsJ5TtU5fTSNZEw77QKaW+is1CBOvsOpcT9j3DwPPa6xvCchgeOQi51tMV
iY4j5EHZ4Z7hmChPWR5kJSdWBM6wOKu/1iHOhT1wPcTzT1/ZAsih0U3TFWHpDrUcMt+UZ9ypmrVO
XUvTqB1NbP92LFqxHiPcJT1iTaLHLdPuw6WtV+p+n+bkwa5onHv+UrpF3tK8PgtR8hdGCXHF8pBh
inOCoKMxza9cni8I+yAahmreUBp1bxJozlSL5BnMo8iHeD0Fx3t7sCaekwvDRFcu71GrI3qwfpoQ
n4GSQY/80u+VvxMruQb/qbEk+DXe+ibZB7pn/c3mA2QjY+cAUBQzSVUW2GVGRXtrM9go9QZRsGDl
7HchEeKH+ZS6nA+iRxDCGLSuYnLm9bd2yT7v9EgGMVjq669kR/LaQORMDQP4JgaKI7FO/DSD7J6R
PYQNC+JfwwmapTc1dSBF/6n+ULiOD8onJAk5A8oOLqH25r9ZhEDZpC/N2anpI60l6R5Gmr08rKOb
KbSXYp0eukv3Y4hsezU8Zml7XGCR4NekFzW4RuOz12+ZZFTI5CQ6QZ+g0xsGFAQfY7FKJH8h77+3
iNKJZPyg96Uc9nYE3t9tlC7yVzxiqTMDKL1/wwzxS/GMvx3l1gom8tlThQNUr3XT1z4J7PXB1AhP
rx13zxxWUjGstgN/VDQn5nH86zTY4B56YNH2Bh5jkbvn9RlnzziyK9LxC3UJnjnWTk3D/qDh4W+b
FEXawSy1/gbpzP9SPAEm0DLF3bRfxIm2Fo59Hbg/rdvmhLmOKdQbhaFeXZFMyiP9CWP1GpD+YWJ1
NJOeejN+UMViyyK1mj/OwzIQlXmwdWjvP6/dsl6jwl+Eg8if5ZJ6N+9USbg6b4XEb1xSIDkITzHv
EGXCQcAq+/1l8eqQ+l6AqNUg76y07cZeZbEEB4dfhAkejGdPYC2XJvf68JIN7xJjwL+9CppP2QHB
tgddnjG1NcA4r0OOZy5J7Mjvf2rJPk0b7lzpt0jJHBvD5ZHDoTIxbGh2i0ZHGD8gSAm2vxnh8Ehe
/HyA/ky/l1HwwMC7rHOjiPy9o2qr/b6Wzi4KLH2hAnlXYwWw1T9XSCv+xgK7IeMAdT2noNLgN4ya
VG/sr+7N0fFjH78R4UA0e0yDRZMc2ZqZESi0WcgfDdfxKnwma5Qo+cgcZwfNC23OWlASeevqrRFk
6h4x2LF6g818oYU7RzjzmxP0qYewGDNXn5xiGr3/PpE1krR5O4V60Uorn7XGAKXzZps5AQsXmfES
fjvouPoA/vQXQJLtooQbxsto6y9gmAvKL3/z7d2ljK1e5KDs8PHpLgCO/h+Ft4+huuG+Mz0dAy1u
C5Xu0lTVtYatrhEgC8ReQ+5MVKRhP/WGZlWzbXH43+Ok4MZndP3c1ZaSeHEFyDrE0jfddZvVHDiw
gND9URAKoprnZznG045AK2ZfocMbJQ1OrqZSeGSjrTQWX3XXNj/MYfYMXQpgs3bXqZKsP2XZ18Ao
IYgfUBN30Cd5GXTrtRT6Yh/iw92w7lfLJLx0LK7O4x3CcSu35yQlDskWFMuSdWxTn+MN0EUlqM+y
YjfkllVxvF5fnMc03bnLM35DQbj+XHaGb5VlC2NcGUvfkqhLrcXO/+4E5bze2j8vnLtHCBodvqC+
WF86DtN0W9IpurvnpiSkNQrzyGQEgc+tciaGBPGDg9S+flxE3lPNmZFTJodVTbFlwi1/4SVlX0/l
Fvw9lkD9Luink+QcKQ7fxf5sBXmIuPjK5r3/3DRGhbu+SAN1WbN3kHqzaSG1Lk3qH81DhfkKBo7A
SQyGOjL48/UGXINX1RlC+T+ZaKimJSGBtoMsWlqTJV3WKSr9Fu2786wO1cBPO02XC8Ol4MWiiG7Y
d+EN8oONhk+IMtmtW+RBzoizRXqqtcF2xkFAcwdEwAnIr6pm0UPdjmTIQkbFr7r74BV6JZt6SukB
8tMd79VLcFygVrmmJm1pvmDoU5PizdFN77CDfb4OdZ36ev8LHVQ4hpT5AofSwh3/i20wwHM7ja0l
ffgkOa+ROEbszhHzcmNrFkk23LZoA64qpUvaM2xgAUd1SrQuKVVqflMTA8RVWtwTkmQxOQucYWg8
c2uP2dVK8DpgKpw2Q/f7hUeCjXRxVLMKeXufu1LyDhUeUZKXyCYTmhGFYad6O5U886iCFBFXAucP
QJ6D1l7/3uoG8Qx0xsEDdrN30AirKiJgvA2JgmzZqHiLD8ILQ0qp3m97poZzuGDLLUf6FQfGYtAj
kwrTN5o4zM5sZ47se4Ell3lxDDoOD+0+3jo4jgTjcycGRjcHvpm9o9n7ollHGIlJ3Jz6/6ze0k3a
m5CBNydzbZ2XTDvdZFuOmDn2wb3hZwMqyb5o6Zh9uBLYwuTJi9BbAvgwFvhAohWbIePbv29FQzvt
VD89DRe61nQwej79xfZZHz45Oyx6+DuC3SAH/sYryBTf+lyadTto6IJsEKEmkMJ7vGyghU9Qb0V5
Q95Lbpa9KLV4TJuXaSjcjgRIqrJYbMMyVxhfOb7DIP5Y8WfJZHIkIszcZe73yBUN/gzPj2UJkmOr
6Sy5l0okHAb4C0yRooP50ZYwt4B64CEOOe+5XTjrAHKO9mRTmW31C0Ylc210ug4niNA/aO3Wo14K
XNxc7S6y7QLC2nbQq6alddxA8WYFWPDtn5MgEbUaGzdCrDGGkpDqqn9nUq2l1AcrQuf9MXeZWsgn
f2jaS0TbmOBQmxFGp4WeRvB6tGwmtXLp/WaoC09f9tuwqOdp3U+g3ivc9xawY6ZbdzVCLf1WIxbp
4WQAHUDwPaburIdwDn63QpRrPD+GdKpUQ9OMy5VRHDX5HttXFg4SCvkYgyGsOPtl06KQheNkKGVy
prw5rWlaNnSQYp6sfdJ47lM7J5t7ttIobR/5uOnK6bcYeltvCzKMy62H1NqTB9wChs1OyeISYQ6e
HzSLfbavNXFpX2wB9R2qqjwAx9Ie6g2Gg1K8HbiZTf36BuQfUdZgHQakH5gybOjfOgL1/MjPuN3/
2UDkGvzHuz4su1qfU0aMQlckEvjRISIH6L60yCWDehtIU+8sUPqQ3mkojMkbxzuOeOhsYQ/PQgIW
lw70TuCw0ZNOLQ5zH1/HhPYE0feX/fyLehUmenqDxFPdVliJT8f2hvdlqPq44W1aJEBnLP1EDDe0
7POqKNL0tfPycmksNkDKRD7md6YS7OH6KxQr/q/CcnnsgStmERxVnlAkT4nPisQAoPNe9zURcaBW
qNDCY1WlK+h19Ui/VdR7Ll17vkrFRI+LNABmXpcX3OaMjjTYIhtnXtlqZUdxCRBTppy2Zz1/Wt55
p6pSfq1u59vlH1vFdMbJrok3yCaPFuh3iTOyqr1AHHwgzqHCDsslw49QNAu+M3Q0nHvncHZ0gKDG
VZXwz6e4EMSbwqKKKxGdNtvYTVoPOm/jhh3MSZVmKobesuLUE/URJ3NhZP94PzCN53/vAq3IXhpg
N0czKNys10+Hu47JEfBsmtqqR5ITiWkQduXB44b0m8yg39fPtZRLVnPeNuUHvrGAzwrBlqI89t3O
iAOj2lDhoJ1TqQTepdJ7O7N1Y7B9Vnh6Fv20RNAfYz4ureZMS9+KIFYeeVrQ9CutMD5uMhwFyqCb
LPu7V2vAIuVhGjNGF/Bs3q096QPbsujtZz7k3qYfKjFsIztsvJ7dYg4gHG2XsxpihhQgD+ku4SFv
8okCGlmGD9nAOgLAXp5Je6hoeXNpiJOaKdOqpGguwMUBFI67jWhP/kfL3OZYI0J94ZzEWOYQm/DC
kk8fcytrxwk7Y+6rynWJNpbsjSy8ZXz2KAWST+vEur7N1dFoW3RKVX/Gw8doFOuYYx2oavkcs+fd
6uTgYfJwORiybVujSjk5gWVQpdhnihOMRO/IKr56/11n9A5a6rrlEbOdszm2WRLScWzwg0r0UTTr
n28F/iSEaRXSPD9SsvxdyjxwtXmv31mzSG+e/6QpVRDrafJ8VFDlokNgWnzzW631BYqFDm9ZzDJy
RPGJHceBF4oivg0UAnDC6QMsXFxI5LF91cYboRSNKfF6GkI59XsalktacdOAsIykJKmUsEIIKgew
Q6YZpaxdbW2TrP3qSRiObB8/PzTkATEEudwzoVI4RQn2F7leZxqVvZmlGovRSl2+ebHw7/p9XxnM
HVJPV2XkkGfg8z/FhJd8dtG7iifrWX2im0zZyQHVyQR5BjcWKL6c2fSVvMqebZtt4Kv66pwuZpkI
K6d7N/SJECcZsEG5nYDfGTlgYQ8z+vDOYGQbvQv8UGTaFdv+8rC/H81+PNX2bOW1jXlzbDVROe+u
AnwyAjR3TI2BNtUddbmLZRxwp6qh+Kz3EcDZX8mCKTW7aF23puft9UjFoAXOVGeRNq9XrtGUk2w2
eiffR63v3cAIP6Z5cwjCuCNNSGBW3zy6Z35+XednpXOio3xm7acOb4jOP4nBHV84+wdh1osebJMe
mzDKgyW99P9zgs9Ejl80E2nKF7ONRk32fDyDHBtNogsvJuCqwqBnWx6EyzyD3HVNM5i105Fv9IK9
b8M7KIfhxsBlYJA4f8NSyJgs4jOKA6PNii04zcB4nkY68wg0gboD6dyoZN4QqPqVtS2IYj9DBP2e
8bEOdXSBukk9w2t6kBbx4etUHQdWg1KQIYeBJSdwS1Mss8h7QLJGQM9Gao+eExug6Aq06gEzOUwX
th2K4ntRb3eWQ25HfUcniOQ8Ft3LzqjW9x65R/PJD26VSyk+Vm8MG6DSs0PbbK6eQxlrEQRZcrfX
+Pf4sUFpWNClFe6ldfz0vKlLpjtkjpUt4yhnZFiS53ZT4z/lxpUCwgcc3gqPtlqC9SiTeZYC6KOU
c8UK8DdEoZN2XK/+h+kexzNpG77zXanrkj6Wski0RlB07gn2adAy+SieHVeVCgtEGxDPl99NdVVw
67+H9an55pTq4YsiVv5FkPHqHSOxslqjrk9iyNAUjvHPelwHwBMGPFBchUxC+dfqvcv+OWnFjLQ5
NHvuj0DuvUNu9wYjIu/HuXpLMNVuOQQWbX1oUGOPk5H1So90aEOoTGqID7BKoyj55paU0ElKCfjJ
0WjFRFyaJB9FgMuSJETpNNzNPeeJUmCsD/ck747w1MksLVONJZ5FhQFmON+/OnW/WPEIyFrrK1c+
8o5yjQQNH2R9cfhCXC5ofeAH4Wb7B3p8p5KWn969tV+si+CoxIzlbr03uO7kVFddtiIBpAirbAxG
B7B2LjV3zNwdqJVnjfsFHiTxugCoNUhAkQv/ouAScF1o7cYm7Ty+fMQnIXYVlqT08KQT8RleLeTI
5x0LzQ0EB4DO3m3KJpqd26K6ElVaO4yaK6i2z8U/4j2rQK6LXcgwDMiX8SthOTeMNMiv7dpKwPeW
z2YmAWi+RB+wlYkVjeFz38dqHofFWoikLu4jsEpTZ0js7Y+I1ePeEnz8WK1JIKfgKlKfwoQfyczK
xZiZ2XjYKUYW5B7hwguSLuVCMTkQPr0GvQwjsQ+tqyS6vSlWr/MupLhOTr1RX43z/S+Hyqa6oTAs
pmBH96SvnNnIaF9F+dBuWQsVM53Fu5O2R3iJ2h1l2RdvIiJ3KA67VWm6N98eburfzrE5SzQ+zS4H
UipewipbDnNBJV1IgOgSYZUh/VJfJh6AM/hBVKTbV6P9BUAkCB9HYO+isO4Gz+i0rBvnUmyjQMAa
LWkb+r3teiToEY8PyM7XWc/u7h8c+z4grZDsUu8wswqXM4dmsLfYT7W4rTJ7v8/Z7CYYouiv+++R
mpM9MKxHvtHLdFBX7/bMzOzUoLzlgsV6FRs/SKTn/qS2hUGU+cHIXtuIGbWEaLQZpAqivVmSNMBf
P+h/KAFJKguYrPHnSy/folMZSHlcHAgfN9VUYYc/GaX8uUV3RztjqszrWjgPHKufHxbXhtP9dQtA
WUPgBNk3BfWhsG6EZtv6OvY1gZin0vu6KgIq2yiB37/H8/65euiK+/UNSOEVO66ufJWgrExS9UOQ
GmRhBItggFZy4vjAmStIKgbDYoANO3OQJiJsU5QGcy5G/Le6ZxohAgnAwEC3Avzwh1Ey1Liuflm9
2PurZu0uDcOaSTf88Vr2Wok0FDJP2bEy9YdvcDm0rca0r8tsnLT09Ksr1SrsqciMTVP9BLARxCcM
lkDTMl+TIShWajzyDJdPj4zoDsR2Tt/NTjcj94u8mc7siTuofNOkqSkPSiT6wHheKRYVfK9Sj9vm
7uYvwEcBAX5owiYJPbXE8AWTLYs8gH6zvRqG6EMfmzHBn0dhaspZcfZlqjGLxbDwCP77BUchkdFy
aKtG6iRTLgZL+JNwyzF4d26lNw2Z+E69TrImLWuxsp4APT77TjY0Fdx20B6vVzIQv7pSPSwojrKN
7YN7DzAj016oxFXrOPYMho/Mbq8CBq+Bznug8NfrtIxMHh1Bb10OeuCkxXwzEVV5DOBFUdV+hwqt
d19Ju1jsoEOhZtDtre2dOLMqUpM6gQnFcimiVi4G95YzUg9l3G/COrWAqh+qGFOL+jOsG+HeinFu
KxBJOFWRMP84FEOdAaYuM+KdvAt+2I6HwO0ndSo7G9zaswSBGNGHS2peEB8zFFwjeAePsNGBKJMk
pCiKF4uYB6Ws87bVvR7JPyILAvM8qSNhl8kLdbFh7ycnN+V2iWyDc3HlmQBDmoUSIAzOAnUQIUPo
nT4BWrr/zRQV0727N0JqL2MH67Ub7vB2fBhJBTD88f9McAAcSaDxPFDDaz94esbKgMlolfLn3qz0
UkMq9lVcrwjJFdVu6+ZpjVmOw8ElNz/B8GmEvdOpYs6BKSzA7xc4SZPJY0uAZ14n7TiE/PqJTe61
w5W5RvNgfKtquvFxrmEW+RZ2XIHUrDN41Lkmlwb0bE2zRogAEMDClYZuZMbBn6lXIy5FRSYKGMnF
HExaURvLzeoweKiUHkl12fl14mZtiv+IqaEJe61G9JSyHRun1A1c4/+Mk1234qYzRIhT1XikOeV7
Vfk1EXgvCZ6ZspQDUb9Zc6oNJto0OFDyK9lhvc/hCTL2RxMufNCi8SEu4M6D05DjpPLubf/rBYra
ww5OayQCAjOlTWYVungFVdRNDs4Fq1TWb5ldtd3bFbf2EaeJtR6PV/HWyYMO0Hfb/6Vtcg25IKTz
y/+6gGa2Djjy+o5N/X56ilwfIbMBbL4k24H6HeJf3JfbCnLOwNko5AoTAGtF+KB0ZFyZFh9ObfmC
i9JgG4EWLF+EYlNcDo5AmKKk+5JMemhoR2MJSYdcafBQbX/MPRoV094k6cODTuwMew8OTuraWJiQ
325qGq93kqUiuMBs5cBb97fZtjXQqomae1CVpjyI3tNYH8loCSGY/Th90CSTe/VD2SJvW5ArdIdV
48vXauVo35YNEJ+XdK5ZHHZHws1ba+UCZpf6Q01c+QWnG6j46vcjLDWq+OrZy7WOfo9d46Mkqrrj
FhQVHK1YgbrhsSCWn/e+T54Vui0BIlmd47j830FfTb/qbaEXCeJbEOwuLJ0DiHV15Gk/rY871v9T
RgUlnUd+W4Ym9f2XnB0G6Bs//YPpX0e68muolRUYTaQkxblOZQFehTLu++HZh93ivOOBuuJLerQM
o+WNaRmCUxqHnp4WGTzKraNrRpLcS0iDshepF3O4jc79gIjK/AXECp8hil45590q/G8lBznBDUL3
hKx9FUvXGjiGyY5EJ/nKBqWOHKF0HyeOHirmQPTv1+oZQ8blFUA4k6PhJfuyx8ASTvBS1Zao0GsW
6oL2O+fNiizrpiB1VEdTcsZiZ66tmpopUeizOZZ+ozKxonOnP+DFbppGlMjnZHW4ms5w68zw8zLP
wxLEP8Kr9QDA/8efTit8/69A6UyQ9Iz9EMVzKTJ2xiiarw3SRNkpn1iJF6BZOgsg2P0Cs6QOMm94
rD2ZT2nLBGH4UD5fIRGSe9UaJ8wyKo5ATIKC6oAz3xdKBRVqI4dAm+6fCrwI7ayNEwbXv2sBBwqo
hZ2h/dPSZ9yZPOlAoVsY2nrki/L+ijfabHZNCR0afbJWk++PY/+F3sT08JglOHD40UxqkTWE0U54
cy2964jeBp/Ildbdk+HdR/jvUBIIm+FJA25+XVH9DCkXLSEn7sRHe/owBXdwWWde6CTzvT9MP+3C
flHDSeFFfyrXZu4JzuIplFulFHdPcZkEBvwNhrJ5GYeREL4g1ruDPlADB89xtPFuZztCLZLs9ejx
v8m0pkqIMq+1IVGh9RaPa3tZNJ8Oi7kkJpQ+cxNyu9Ch00PjnX+pMqlWeavXhql5XLHTA1nvpVXP
m+SeGstlFZIa3njpbxFbKzjrs0+MrtKR+q2Y8J62GOp/pq0Xxp8jQNc12jSLZqic5zzM8mYjSpJK
3oCgy65QCp2TmhAzL4nmGzdjqCmbQcMoD1+HqOR6kh1sctGb5JT7rFKXIIs0KWmVXQ9Y2+uli2CH
LIAFAOfA6eLvTpoT0eA3wBaK6R9yW2wjViZm7PXCptW0sK64uVKD5/+3R5BJoI5MGJxGwPPsUB9Z
eq4M5LfCXJMNrUlcrADlWSjgH/9BwrJ6rPHLh3zSvKW3fwuBRq6QGUUKrbYk4FXivvt+aMs6oQG7
Si31Gx/lloTS8MOJaJByqYV4s91rmXFWEyhnLsxEpsrNQptPKQ/BoImx/APqw4CKR9KkKikt+vEC
CscrlmkcPVzYpz8Ng0X6O//1MFitX4FMkBFgWWyPJ1cJle05f+331ScL6548A0Qc/8d0mCp6DYiv
feKP/q7LlhCmF/HPvuCgSk2EYjYxwv/T78ZAV+ZD3a25r0kk44RyTDuQdlEP04RE4mCGI67oCwCW
7tAk1mV8n+p4iFEtJsX97SSFB0O6qve2ccm4HRjMjIDZjYNfKLObR9Qz1T7iIHUvtXRH/l4m90Gq
x2P7nbE7T0LRWkpN5LNK/GFYj+YSfFvZ82Y16pc7PH3A5RxpSWtBEybnnLlD5JSsBZlosmC1tqHx
V8iUgDa/k87WChcwLQJhyYuRsBtt7w7N67F7yrdPLq1eyXbybKAOcONxFOhqGB+1G0B8dvZQy9RG
HrSdERXMJfcE/BfPuC5txWcd74MjgQAQ6FhMXGp8S5M1gPbNOWniFbArcG9Blt5iriqNIrGlHf1V
65AMVPqcC9C6QRwriBTaJC760kAxOu2sCl3Co5P6uZKkaQY+kfUWLDC4IfSFde4W5byf+qkr/Wb/
5hO4POWtIa4VJveGc536+nswfXEU1yzdtXW17cvg7m99vDZtD+hiJ1I973SXHzpn3Ouipge7WkTD
HOdQlDBmS9Wowqh/1pHVzKMz4dBf6qip4lX0YqEffx7bantcvpCldWp7grKAXiRdJKwok7fVXTmd
wE9boedbS6axJBhXe4p9PPc+RPLVBHH27S8nVnBhWKCFcD9eRlD79f71V7KnDBqEPo/wJDKHJoIb
cvJJ7ubwoNLS0irH785/EpQRxHOmQSIJxj66aEd36McpCK8RIBA+edH5CfVwrG9BuqlmZOirLMsG
/F2Zqkirr9YjGl++PMc92XfsjL65m85plRpVKUVtIMjCcne/sJ+VlqPU0l7pMB+uW+Yh9fkE8rSu
k+dq4BryT0KsSPAezrs0YvfGjlwpI/qQawJRxr4vZiZzTXZu69VenhfuCuK5WkNzG6RxWJDGs+7G
uE1LCOCBFEstweyMRmoOwIzaQo6lyc4E3D9uLjjTRMy/YAeue3rlr6vYsDBRrN45Fj6zYCWCrv84
uMl41ezNvMxNd1doQjYjvSmSOIj+yKWAdLADnPaB0Vm3fK/i7SY2Ej603eMtl1zu5gI5cvzqjEY7
Tzz38Fnxdr5/JXq1WAlTOwQgBhbt3SvNduqRGp15IVMSn7lmW1so7LGkx2hhEpZZ0o78AZMD+jxb
SjHDHRLBs1QC0xEL7t+vd1kSbQs/b1SknJnJnPEOIuGf4Xw/KzXQBXTvi74YqggXtLwL5Vfcle5G
QdquefpXPyQmnMKvOqbXNsIasAuS2HhpnElApUmdpddDGsCzWFsZ2Y/OVCoqEI88fvsQe8MSTmji
yKHB3JqZSq6aCH8xMj1Bx6EwQt/Axh41RiOF1TOlCdNuXzJRpDCzXauPqkwHWo7cCyI1P/yTbt+5
n13eC2dxgr3mcF+lLdieZ2iWnzsOYm0UQHNo4v+KRLelXHGq3Oky8bhQG1DiJFmQQGetCSwn8qji
c5rYoruTE/lJ+gesR4VxtZ9cgZ8CG5oNe8gOt3AwiApRNT57Momgi0C3NDyigwHM//TaNm9SFod2
Bxg/9+2ied7iv9oTkiF00B2+gkeRlS5EpYgCKLNgaYMa9UREmzboH7f+KRRnSxwWOzPPWcr0i0kO
vH0omQh6G3fqgcaefdaMEaQLm25gWEormpDwqCAZNEQpHQRip1nilpAQD6+Pojyf9ffMnmlpaSPx
iT3dS7BQRA4ojx776tSx4Z5Eiym1x4eo5rFMq4/vKndAf0DI3EDHSEztodcLhNO8gGefT4rZa1I1
a5XhWvllsYs1YNLlJZoqvWkmrQWa4FgFY6m+adFHWtqE1lWmshLigu9DpfZE9rRYx5UOMGxtxwUp
Vmp8oLgl3bXtu+Ou1z2IOENcWPqIs/3X9fxqj7/TI3tSywVJcZ0/6HRt34Q8ipdnzFDJ11fWfmJA
ViHmbe5xXodB98ziYJQyLPvGRCsI4L2h5sSGVa9e39xRfenRHO0PA4GhDEL86j8j2NmIMiSZdZQU
adiYt3wYK3FM1fvNSucVSymN6lK+tozarplyBQiVkGGrBYUklNz7X6JrDIhRnXWpzkkKsU1blwdb
2Hcnrgq9nC7/Y036g44660uc3qIFFsKCvXRBPzWzh2obLJVe+Mhs1vFZiMItjTBvHosIorTU6Qa8
rA/wuaTZuvJjMOubj2hmslKDMLgClHgCDExcVGVpMhXn/+uuRTX9ZDqCcZMoD6crFbAOTLiN1YU1
BYoRXTJR/ubHnGLkvMWLMjG0DXeaFEcELm0uDaMW8Kk7NVXuX13i4ie4B69hqzNreZPRq3PZHYBw
wMwgPFjlLQ2wBDnBm6PN5ly7MLOOR8zgmdzNfAamK5K0C4Irq6FP4qTtq2lBWTadIj4TzpJkD5jf
TV6XKjJwQf/vWn1Bk1vPti85jLM249179vBe8h74ZiLip7x0GndHxe968HqD6mL+RX/N8RzwP6J/
WWS8n6MU6cUqz9kcNfRvh/MiWb9VXrTa4m66yzRAmUbFglDFecHNHjf9UgVLRCKRi/9chZsbe+R4
SckYHdjz6NPNKBnpFCvibt5RA6asmtAezdCd484fj7GGiV9L5Y/iOfCqAZvXqYi4FTQRagSIO0R4
mZ3uJvUbN+wN/D70moGYVjewE2tJ32IZ4d2XfQndLOVvPB2oO6aoxOBzZmHovZd0+FS5KFfS+EWx
oBiWXZi1hwl8yHZiyfn3sZDQyVVJ/zy5l3GSPv7YGm4k03Ff5Di2kWjYnDT35LJMkGNT3fNRsiRo
VSPRtNt4JKZPXdhBGm7u85JZyqCEfVsRaDToAezxfD4BmAqZD7uaZVH4ZhafbNumT+WraouzAK7N
NoHWqvwoAL9tE/240JpnbSnhc0oRMWtJxDYfLcHaoyrgc61A2yPxfPGWicvrVLYV2hLNcLOGS2nR
w1H0ZaSdpfIaVoJlufwJ50M4wlKJIsNCkgB1LIwWwjBgfQ9cCJtgBCDBDRksizMvB9D94A2K9ZOS
pXLcrs5fL0FM5Wl1FX2EaHwwgZOGdsKzKP7X6auO4yP7vMpvn/ZIYWAKdrl0JU+JM9ylv9cS8NB3
a5or2pkjpKzfq6+/PMd5T+n6DMlL8rUHuQOj86w37l3rOqLZ3aGATCafAJC8Kvb7Z6qwPhbkeXNV
McPhd/PbkwdmoDRjH9mjaKm5t8b8cQdHr+FMYkKST3cTfGYHyVv2k4zyk3ZZL2fh2vpayLZd+olS
aFRC/YykVk3Df8Jghi0K8kWoN54cwuNzk9tzv0mmt8ghPK2R6jvliwlIUdYjC2gycnvNE3XrKuCK
0WLiuOyjhZYsCdgfkT1kn0+I9V2gtB2Q0TC2qAenI1zf3MxZk6D57q5mJ1Gd+gGX+kxyTYWVbbj1
SHbWWV2+Vsck7IhPTL9OYTUEnj0+Yhy6nvF/+af6gwB+sUdRtyuLq5mFrEeCi52XLGeuRUThgFN0
pLLfqIk8kKvxts2VOHMy0yuvJiU8w+PwEUJQ7Ib8a9HyF+nLlul/5FF+xKJefik59cI/hot2P197
wCS6VyII/IlPOfxRVZEfZoPQ2v0/ACTyqojzVI9ri1Nj8V79gvY9hFLs+Ccn1TQEv2MJ+SyqcYP7
TbyXPYPk78yM+JSVe7UwZ036mCq1ibijXzO6MB/6YcQBnstNc8TwmIU6G2oaN4kvK6/ETaZQTvS+
rlzEMQzqU5Dsx+mSJ+mdlRIe53gbOuiqRPneNOOjI/XfsvLdMegBGYQjjtTkSGBReSdZMCndzDtu
Suyq+MZghWQ+3NDzEek2243rGGb1jpfHjXJ0Vh/rFwDvbj0PylKatOl0RPHFJ5hY7Tp6VkR2ylhr
wENIEvmrAnVW5QfwQQSYEwPfqIoc68uSEbb4qxZK9J1Vpx7uGyKxIotUa6Gccku2ACYE8JjKo0mh
7WepnRD8xLmzQO8pnytb8HBqXY2EYWoMjAcqo7faBgh7lgKXSRETdNDkzGklgScpkHZsSVy1KDHO
c6EM+vvY3jp7l1/TpEZP6dWI64Tk88bMiUPZRxWVo7lHbr0oKVbEtqeb1CsNq8NOjPBQCP4Z5J3t
BrpQZFaiKbfDopjRnyYBKfDcZY4i5ACNHLP+fGE3tj/bKOpiT6dlfNmg2Gl1ZsRmc439HAwnLo+u
DCIExCyS0LoMLfF5BW3WYXmo3a9Du+zou7cFazugbRi9hRWUcF2Fw/29fxwQdZ96UAdzgOmQvbaH
1B+eKOCBJITnQysE5JD0vnrr06K3Gyicw4/1fkmWmylNAZrG85+vmdU+cmbxTZ2TRi4DzU5w+BdV
J4M+6ibfQrxL1wlfpRBCJrZEvVchNSZkCEQUZUvhPiftUKANH9DxCnrE/cpYv55hwgvE56zr/aE5
GQYFrgWBtZoYD4cBjR/GIRoUwBpsRcOTzW9EkQQsvSLZcBYqBQVdlHLRVEr6zAbuBV9xIq2oCpu8
W/4Nd51sAVQLLZcmAOGjDyKSeRr3mmEou+/D2B8fMDazeuuNq5NGQIWWaZqUkd7zGSIXQczeeWV7
CqVdpsMEdjvAab0OLml9//PLXuKWUhpifLjve0rYJyB8YZEOK1x6KcxCmE6BcUCR7tb47Hmk6how
cx3ek2Y3Mi2r5Z2zY8cR7m9hQu5QfxzGszd+v85zF9l+VCUEBEDiKlgcob4MDWGpoXoEpBqEi99k
DWxkjFEf8RdIaa4vyis8qR9vOtdaFQRza1wfCRjxWa/UILtiCL6wIhH+bjlyESoJx6TGTDrcnljA
qdRZ5/ThGgdIL3VBrOO1JsL3HHPHnKLEMg2pkFLXDSX/eeWCwXy6RKbfy637ulZykA51zdfI1dXP
guX8fWi4+WLj5yXhvjEx3hwAX2YrwH0IHLsZ5Qr2fLs4wkIUsNsIVCwWBDNzQ3Slu9HGfnDZdVKi
RprG/KJ4zAJTSfF9uv+FaTO8onuKjHqDcCOIocIR8ECOe6u/IMcCPvaoQZwA5z09gDqpag1xtEpX
0AB2b5AXQrzGYdXsrwPClLpZKcGmrShk9HeeaQSZqofHDoa/c2svVGy+m2zXSUPHVZ8+ZW/oRSbT
Y/yGxL1GFirP425x5Rg53YGFvsFR2ctTRY8cMnZBNM6QIDVwJTXsZkgHyMFVMFpO+t3TjM6j+32n
nq5+D8jnn5R4y9YwBOitsFE6rJHlO91wm4U8j5/lYOsL7HXEFrbYjxaiCWShEWdNWInyiQiJEdST
EiC3A8mH9R67S8fcgME3NLCQv9PK6+A06reIA9X3HAZHfWKfNkyDHM3oKN2qCDbRsUee4U499jF4
B5IrsbZ+6KxYzqhoxcl5JySr/8p1LBRxceAq1oCf3IgDORUqbkn5efu0v0TKIa5dqSY2uSZTetr2
bliRkUdaMqjH78YPDbzyYwBRnavCUF7Ak4zcaNPTEMeR0OlShSAyIJrwS4hRZulLGKRPoR7rO3Zr
+qJ0TeK/vJ7Wfqg/Lv5aS32P6K5v+NlN01pArH6H2iC2qaDb7fBk06iu+tFRl3kdmMZc4K4Z8tgO
Qt54BSySFE5RwxJwBusGv9GmSuXQTp/x01F/E/cPqCapuVwr2Gy19VNMMj9jRTeLNKdeRKYIhET0
qtycKtNjBdYS+hSJmYT/ofHDjZJiEYrdF9ehckgpqvx0OdEE25opmFE2tg8lF729y1DlrUZUPIW/
TKKR28lTK29TdFZQk5SDdf1Au1UxRAId6sBRfJAUc6yC51qFEfvXKl8hZDKH8Ufsqv9x9pPIb6XY
yFUrcUd3Ephw/vXjdFlcVvpCY4EcyoA5YeJah1GiLevcDIzeiQA0zz5YBzMK6duG55514iAMhayc
ZwhpOLRI9uc4kuEv94ZTZjqRhU84MBq50U+7UjIgfaYlnsyZ79Gntu/tp5BPb8zzwIzCOlEc3TqL
/2cDRoZ1RBSQvjftS3AMusSjP+pfO/z2TIwDPQhbN9yTYKYW75mPe9SSrALDnQqqrD2LFXTbMtHj
bkqW+vcKuKNzlK2i2Zstb4uo3z79Eh56Tn1CebV+zA8BLIdB7wFH1Yk6PzKYe2ColoC6Np8z+dBe
aMyK6JwpeK9l8xZ2qSz6pd8IesHZGpXmzTaMHfwJ4r5EDOBFl3Qdn1YsYj3MhUP88HHbVUFqhN92
lLYJSSCjBPG0o+k2GnK9lbsYopgDVRNpVaV1zXTpWVlUHqAa0XOK/Skb9O8sTV1OLHIXCHs2b5ij
ZBIvcxvH/Dgvf+x5ZfENQu9UpCNMSBeybLGiOUoABCon78TpVgdFzLQgSJHZ7FOJLaXEsqtBFPXn
oPhxrTSHUm+4OLYvynq5RQI8J/w37XYMLjmz1sRrWcHWxVhXx0hOgFsgAW4RTUMNWQ2MVd3KgSZa
/MJCZbyc+izwZaZKufu981tqOyBFbMNn1Ax0BhXXRVzZ56GT9qTPPo+g2c64x5h6F5K1YQiBYA6y
rZha6SBpX6tNVWif5CL500VKbPYVAQzUVzbfnwyRrwwHJWCnNLT745xA7XVIxpdoFL8gA+NtmUiy
2ZIsB3tSQ+qQeoi3OB+tYur4mXGJbLrBv/il+KzLYAlDj5As6wZ3gkTID9TOpPjxV7DDxyxVJrXb
ugB+0uB3hvqX3MtQTOiufZ6a6AjTNnpEegIkqDPaH1Fd/SsMwvZeQyywRzmYrn+YqVuxpQWrBgZ6
xiKvTRw8kbiSQ4ysgybFwnX6t6wGyHvEbZKqxpiBftzhyXBYD9kf2EzRQFedXK/fj7piDmNcYSjV
91P72xd7aoatpLLSUax/pIeHnNw1XoEs/DIrwahy/8P7e4Crl60CwvDI+YvU2NfcZkpjeuxnr6sZ
IyQ2gw4cywgW5GWMsyogyNJxf3O8Q8Wn5dA+gBUf57QXysrHRhVD1cdeujZ9XtxvlsR6664xMakQ
qehhy5wafuPXht7p8aWT9XocPhXMv7t+ScCFXDADBfXf5PicsSi3h5rQVU4TWkhms0v/78LxFGTz
IY/D4uHj2H0h3svmY/IJmGZYctsEyvAR+wV2P5KBrF3PtebrQGuco+dhoSccsNGBU6lc5G6SNQaY
emGAHzYFCptYtf4i8KnaS05bXRYKoPa5ZJzd1rcdKMO+rLT7vVnrQQ74HyWkGn1aRdXwkK5KYeI1
q8sHF/9NRrAaveboE1bcAXwUgQCP6Gh20W7nrR9h2rbORCN6623rq4zuLJ0laIBrP7BDXFR541bc
oK3odZ6Cg1y8my1egTAC0t4M9WrZnq1SHz8tmOktyEXxtGA6AaFLzKc8Lbz0fp928ytVnVD6eI0M
7CVOg52LLc3iH+Z5gBqD5E9RuwWCcJfpWhTunBOuTuVXJJt0Y3PylBKjdtk/byL7DTmofsgPLRmw
sRn/7HtzbF1W41TWh3DobUKtpXI//ksU/vJcgPOwsd+vJ4ksvnNxLHb1BNdXSm9TbojlTjaAH9Wg
IOCD7RSlNtp4aKBxeUwvcs86wDGT0kJlY/84qbmOVzGTsRwVhui5GZTrzugAd7YwRW5nVpshMtFZ
AScGdY2jMYXV1ahaVd6NdnfHoaaGtin9C6g6jQDOkCGemZbHflq48u1X1btfScYoQNcOXovqHm+h
2rJkG/w0MltwCxmmjXFqd0/3vmR1+fuDpl8ewrCV3fOwuifgKxOjJfFV2CUMwfBojzL1NTB80QBL
OVlwHdhFFbyKoOImC8aa+BCnR5kEVZ65HHeqHwnRfO1qc2svnHX0ZAHuSDbJStLdJYOcPEwt+2x5
ow41xYnE33mDeyiWz9N9A5muD/5+GzmwFKCuDdEAo3RfHYLH1dcWMFmYU0EX95kWxP3mxEYvEDiH
eE1XZ5fDlWNTovz8VJJi+Amk+RfhMCwMxkKXya02an6nzEoKV7tXXwIOO/fLdon8ww57OaGrb9QJ
8JyHTtgzIzQB+hUShjTcRocjOZihbl/YXvI5hxZllUVeTYvPg2MMcxMyJKdDnRayiJS2du+5gLkM
Tmp2vAUR8vK+Zm58aCj0kspSCobvUSH+dJeqp6UBM+BkMGaVe8+dQJYrF582wR6D1oPJL/9ZEqUv
TspaJpoS5O50iCUG+mrydmo7tLALHGXKrN7z+gd92OLoxs5zHbtmNSWjppf5JEXH9vv7tsKl/FfW
sfeDDt0yCNSCSGYO38T3eBcPtjkN25TDECzKFsHvxkZ8DT/epAWkGGtqh3qTMQ/mCvIUyv5hK35E
l0VW2r711g8E1WspSFoM4tzUNoAXlHDhsTtMX5YRXBQL8oL0o5rcjmRCDFFyHl+1m+1MSZBUyMCV
LUel4yieCnotTGk1DrT40/R11kJmoPGo1NtWcLVQAvKGdBNxrVu3LdMZfJScQcYrDzZSNd4RuCNI
YLQHKHEGccWfUPmqESWJkPCdE4QHHT/6oXJSXrq4ywVQ1HMUCIlkvkrgszruuL9kyzmtPhcsGoVj
OSfxMiJu+9PLkFYJ1LREiQ78kqqqGedHnh7lBF8kDLqRIwd6lkysz4l7hxOPua2B7s7xGWMCL439
0ocKu1slR4kwCrScgZpWJIf1ue7no4c1JD0k/JwfgwKOMi2sZyAVJWm43MmodlTzg/U069sCAuu3
viBEZdUakwG9zsC1+Gm2Jrd2WsXCtzuYbN5n8tQHkhMVtCF4vc1ajMAf8JxW+9CLw1HhYjKOVAoW
YD0/LltSUiflvC+cl7492TeFj1jWeiNHSROzXgDTVERLelDv3JZslmGdAetWJMspj3OwtR4Ed9yt
Bl0qWvbo8BwKEWsZjl8ngsV0eyUu2ESHEBh8mIuGkq9mQLNzfG8AVs+3uhBJBa32r5BWyyyFlg3D
H+aMr/LFRJulM0P3q6FaPf3B7FegltPVDUtQGuhXn1+5xXBGAZdRG0q+bN7Dsi9qXcLQabJY9Gog
yG9P/78x3Oy5D6z7zgj+D6nvMFo2zEfbpHJlMOe4JNRZbeebt3AIrxg/LE1pSo0bcUUzreivIQKr
Obbr0oqaaMX/tKP4wRaCSNzuHOyBLU96hmyJamQHhGij0+Tq1zNOq00IEXp1LcvT8fjqVbWgTlUM
ipr8jOE2d0kl4V3ag4dw+G4//imo9WMT6z8YV3YsMUxh8+HOAOfuqmx9fRjtXeRZO2rmt2MHyvtw
SiL+Cre/F6lY4EIiAFVY3y3hfzykD9h3Z11M32ZY91u9UkM4uxgUWVRwnf1m9+aaKpgAlNoeEVgJ
9Uwasx6Ht+TAEUbl3pwcmyauc68vTV3JCNI90ywmgDm+ubUz2jQg6Jffa+bIuB08NsPCeWnwrGXu
O8PM9Hi1hl3DDepgHSN2tM+ZOFt2oGA+qJqYezf5opDgIyEMUbxEKN3hvHDL/3PhotaUBaziFemL
kMaQEC8GUvlXua7JsRakcH0Eb2RdqOEIDS8y4zp+J8dztRYqdTz3+jlai8sR5HAud7kSsR231wDo
xcU0KNoitSSUMiVp7UNGKiHQyU3SfbQlh85TRIgathU2K/ZcMW0nMURIVcgWUPMR4iIudqfDK6NK
u3Qqb97Y16TqNUhh+5r7uHRzpFpSmT1hk29KZafqHI75bo6Cf1m3xKD87ENWkNlJZqv5cbx70skI
eu8ZmPvYXsIY1GXFrQa65dP9ndzeEBlcQnX+w713G67dsGFiyhHtv5+hpQ0KK1SyYFwO0A7ZohgN
zRPwTkpMUWJTRITC8v2RWokvX1d4HphuWVwcl+Xo39T+tC9O2n8/l2qzhNJbMvn8L3nfzweTkdbu
/lvrx/H3Dqj9MHhkFbzejbBhojbC19N+l5E1onhF/7EiHEGHsGoJv1mM1qDW9/tXADFRcoIfPFyx
QP8J5epJz5Wa6HDqB369koa9drUgqo8FNuZLb9nUigK2UUbrdC2nucHaqI9WGTauH4ByyKScOogG
8yzfMVZIoqGPRhzj3/csyM3vAMuadnYBbaWfN2BljmjgdcgLRpZmshA6fNrhC+JfVN955AZA0CC7
oaam+pse39hmvnVSX2C2crLZIwPFojEsvZO/LFQ6tmTDYErOrCHYFdG9mI1n03NOBYJjNoLiFbsh
tR4SzqtvrDqWQOKPn4m17Azs9d28mjluFjadnKhZn94X6J/Pqo8JI2dZ20PNB70jST+V89LlviJS
uuX+6osjoDg7g4RERfh9a6W3qQRWusPiTaNS5iRUi5hSz1gTCN8fgtfcYsZavMxEeC70RUSy28aD
r2PRAQoPfeA8YgUf0qLtDDkdqoVaJDwRnc9Aaj2veyWgAOSD5rYTYA4Y1JwiI/G3GBTTWYjBaSku
U7lUh+Ud8QznkePnTp0lyqMfeDG7Be2/pRaocvKxAQKy/34yqeK+lEFkIytRkE9TS/GuvrBXtkQz
85lhukZCdxeT8kxxCSmZ5eIDo7aqWg1UyW4I13Q8NqZWtjuwQG6yjuAOd3J02QyaXiIO53as9AK1
Z3Ld+5hzy2H1K3/U5DGdalX+8HRv1MHGA16bZAQs/90zmiSVniMNdXy+I8Yz4vly+QgC5GKAh6XA
TJtiCbCb3iHr/FmDQvLxKGSst7+Vvdq0jXTygbtgCDM5Q7LqSGUEKnFbwb6Ob+3dPiB2cWrP+SNi
w8suTeTv/tfOAEtJq+L2VOeOpOBFVporRQMjGBiAt1fKVI5jo2EMmzgJCGxjqaDwUeJfVmB5gzf6
+ASi+TBJGa8NMCTbZfahMuHrJCa8tw+5FdnurSuEp+t/vdSaJR8BSkIRwOsS6TAs7NIoAzxcGOsT
rv8xpP095GXANcRSUZPVlAEMRw2lIBXFiSknrY1b/NMCUlkG83bdzepCuPs66bCRsQ3sjPgSS0jU
neCqtjsP6ie9fdqhlhCZ3tSLCprZFM3fMfn0jwq0Nw7MWGqamGA8gZr6j2cDNw8G5Qw3hr6QkO2s
tWgmSIwejdaoj4EwvCN1jVjYwci+T4N9DX5InnlxM3VRKJgkor6mc1SPT5D4KIoFBR4LEI7bIoPl
Pj0CoAoA/MxTUiByHdeFj6sUCnSbjYYGzral21MBANdinJd+K7Jw07hjzcVFEzWT+p5L6YXybjP2
HlvPHtvWhAwsZ9ZaeIQTQot6nXDFgYvz1J7kYnTUXr2+qmp94hz4k9QfnPb1Tkzv6ODCMwtDpYqk
12qTESUtmCIRwoAyrvy8yP7n2zf3OTp8qhvKiO7JgLQsWobWofKDsX59X0JuvK8P+nZuTHJ8hWcz
iqIAYaotb+iukxLq47ylMNN/eJ0lVTlI3xcI7MxDAmY3PjymnpNzUMtwf13AmPwHH/VfzxdbCGTl
/oF47gRvFRVngrjv3XKAVJ576NuFJEfYslySjzTJHCxs6nUGeMXIj7y4xKbvArAyyQgzyUwgY1do
6B4cGWnetu5Zsy/y2ktW1uI7He5UDr3BRnePlHltXYNtIomeuiVzBOOw1kv55a+jw73bxi1uDXW6
hQiISaQKkLkknI2zgp9zdSuDqy8tDLp+zN/7Wvn2ildBys0ZWGalcYdE4lL9XjMsa7uNftWWQIr8
c3Q5fU+1PN5ZxuPpV8vf0I+BlH1YVujhqzHGYY4pHxhiTVcoULWzXcpV5daQNrvL//OQ8ivMocKS
vwEllPrpiPTeYqAevjXVn6HXzOO5sSkURJYJqZ9pQFVV2L/oivGQvG5YqF2H2nPXbjfvyehLrBog
TZUpy5Hraq3EzKji5p5Qn1LC8JycWH8zyFHgVuoJ+PXD1XYgoir4cL3kMP1n9FkNKtydcI4ndInF
eP57mnTE3aOhDKaiqvhASbdqxohp0oOrPJanFbNv4PjYx3gE6DoC+UENOU/R3mtmMICm4iSL7PDV
X6/1AAjdgkExg1qdhQI9jPY70YmwHPhnwPNTwbPX0HAN/X5o2yYf/IQDjeyevvwS6Yxeu7it0MPj
ZvbLHy5737TOEtTNgmUCUNrEvzm8kj4sxG3huLE2WFSco5jXEZpzHqgjoLar8zucN/2pVcdQqJBZ
8fqLLK3DgX8EEnzz+RIdqVtN+iXarSY3mbDrzU2cVF2//5G/VXpxzZ80Bwf9t0yZNXoM1o8Rz21c
jOqgbCGq31sQOrz5diBxXvYp6JlRcymSPJgbnzpF+TtrY73oOMMIIcOIdN0z1+oOonQxMf0w+XOm
uOBVZbDNCIhEZR4fz5u7ecO/ivaxqXnDi5+f8X2Zp6e0wEudX/EqbHC7TuYmhy37OYas2mmijCYh
DQYnjzKNI32DYAHOTc7D0EHg+cRuLfzY2Dbvel4IXEotpK0lyU6huQrb1giLgeG/ctTlj7etODth
CKDKr0qqT6tpD6dEULxOFlqM04O3mzxvM5q3vR5x/eFRf/1+i/lDMG12eHMuw094WB6AUYZr0K5n
mczE4Yj99qg5wiyQ3MFgp3lVegfvKl0NcTgDGTlGPsNIPUHffGCoo1gOaPwJTv+oNYg6O0NUoodk
vYAY9OySq5ds6HBmdMLp1uf+cKXh9NXnOBATdXfV/ij5k0zOaMSAB9A2ope8g6XbnPW2QcEMi8Vq
b2LLU2ADl/cKGtDo3eAEJ6TpcNCo4sQbJ3WfA+gYquvpO6IYST4fxcY3D3imaiFtpDknSCFb1Xgf
hddNUwpdVkLBp+fXRsUl0WrZXB33rpKnekPlH8tKxIKLsPZndmXOdo7emygxBiIc6TjcfmnWVMlI
hlk1jwRSC4IQ8pywMDsY8VG+UT+Fz9bG/SRF7XsaCGI+2rkLxDjGBbvz2uRNR/IvutLXZ8F3M5dW
y0ud5hcUCknlr4CsMlio6mjm7axFV32smvOK547cFns1kuMACGx/ZFNjwru80RA4n1h1Q4TtDniU
vMYpZY4VlyYBZO1aNUlW1NkaWEh0EBt9ttqsvvnpZiql+BAi4IxZQQnqlKxMWZK/Rq8xRH4n4ZPR
DlDS6iDvlHeNotj/IQIcw8UFGVva8mWkPqX14Na/h3YE1PJ/Wq7TOYOjYjiZ9E4+nFobz4KLT2aB
T/OSvN3Zf9vcDOADlDJRi1NgdreAS/sY2EXmoUbAPMUixkJbInCLPBrcjT/qAj90a4h2g5923zWW
K9nXy7M2ENgiNvvuFedIilamNQN7RpX9fJwvXzriAATqc4hbqiNU86xDVGpWAW0s/c6DWysiLCMx
iuXTKm5ZxuisLD1BGm1ujp+E6EW+FwXutuzowucHO+f09v9oR75A4OFgawTopmIRp+AGHqXrt/VE
ydXnooa3mbcQ5oj9NTbQblZ0COVcvHPVlcp7FigoUPBxlVyc3QvmjNr3um5HkFfx3XBii93r52g4
m86aOArx5XhlgAeSGi8qKN8L/5ar/9FkqQrwcGm/efo6V2VYjdVajo6IbgtrdaxUf4bZrV6SJBwV
SBX2LNDhNiOWlexBUyVqbUj3AfygiUjDu1sTvX0+cQh+wKaOtD6WIHyAuNb5hLLA4VKOvkWjtz3c
q0SruBCKOlU2/OtM1UO5HmlgLbVPZoR+QRNlU4xnFJBw5ZTwEynd06qg7ahoMPtwx/J6hrABiAmg
xneE+gGUP+FAJuOOIbxqyBSgWQ4yCi8W6Ixoc0uiz+NJa8cT3Zsw1EvJAkTBeJwfYUDbsNAkL/IY
8osFGfDLM77P7lChL8/m+rp+stKZr13ip/y+yuZXJCQoXWCICboQBENQa/usnLeSJZDgxezGNZ81
grsMPe4ITluSYzy7pmKX9o8GtCP970m5XpVmoP+YPp/pRj2TzokzreTGfMKA5+FpQDz/NWHZyEbe
3yf2roUANpmMq/fcBDesNtUAwxSoCdSUSQoUAX2LXo6bFMlnka2s8/UaFM4aqn2X2SI8KfhbreSB
Vqe5dkKmP06O8EitWMh6Elp7fJDh7kVBALiinKADGPGjhZEnPvOEo5gmILncSo93/UY3xAIu3H6Y
2ePSSBjkEmTAD3p0gRf0yb0YE/Q7AF3PdkuoWlR7Zw2TVRFedUwz6ZUaQvOa3mygVIPkSs21FYhp
41Oz5jPGXOSpENQFel+JWSALH4aKrJ/bR3OxieUMTWmozRdVSVeR6uN74IMHWHzJHfGAmg7jL+GE
sJjptgpjq9ELeWR+gzYGfVFZu8WWJnrBRfFtBLa6IuMqDCiw1q4x2L0hJPl+AnqfhTDSizd9SOFt
o6uahlnJ4bf/+rRg3NASMadgkSK39fMPnLc+9CtzPJ1kc9Edfmd/s7+j3HaLzkoqDIdhUF0j4K5E
7tjj4cGmcv+gb9eoh9k+0vPHZSElhhJfh3nIxHHJTIFDDBB5jpcn8LTaVcT6uZUktw3fudi5AYlW
VAxA0TudczHypFDClp06w+FmUX945pz3BNPyg+GP44+iasI96Sp1xn1zR4l3uHk1yJSLTvZ41aGb
JuZxRiu0EiZamd4nWGVPJrBR2roMh1aP8XwPaXKD8078zrcNBn6UiRFCL0m3fibTmEcb1/E62vpC
35bBT6hTYxUDYdf8YTPBvNsqZ/F04CuEiRbVjO/N4U/Ox/InoDqYIgNFiWu8z8tjPoJyIZVZTGvR
WqntRU0nDUKIz5Lo1Y40KZ6doxZhFxW4rPlLh7ted4qvFptfnTjpPtE0wE98GA4PWYaFvnnP0TdO
yTbbEnKY6fudDhNwkQQhZ+PX2Yn2yKO6HbQNEOckhrA2z+qcxoVHwn7FlzAKfINd7ZCI7UfW+h19
wQ8FDtEN61tP+ba94NQ1H3wu1sG2ACZ1HPPodt8FtGDwAp8++orb/rIXVYgymCahuXFO2fa0rUDz
KmJGg3qURF7vq+Docz3ywxMQv4OjmJgzr8oG+jBB90CZcjy0Y8sAYeBVX67mx1G1W9+1ZqRKrPWC
upMXYTUoPHSblXs4DHNXu1yyi5id1ADn1SG/ERkaFby+ppxWZIQBIF2hkUNFckmBXC4GelL4niaD
zpKLnSQrvWh/Qg1GGcV2dOEyTAfrrxiR5vLIopkDzsQH4Dd31JLESFb7IkGVFk2RGDD/3XE25YfX
8xaK5BTVxaVd4DIhrZO+QELvSsxn8uBD/bvp8Jr9uB515PwAgiEvxphwsgtyfIDmuxoQRxDNye8R
uS+N4qkMdTataf92GKsTN6VHPwRyyLs4LNSdCLtkJBmH1Y7MLixeVTOcc0B/y2Op3XlBFEMklI7W
pi971iyy8yhmQll+UQmjlCDqaCr8FGUnHssdXNVeCNEWUKZmgZT7A7qiXZjjdPE4sssY9qMtlkt0
KGZ5z3KAo6Iy2hc/FzsXMzN612Gq7aptSsTxuWdf6+x+zyp79M7l3JrWDPsTnmij1bm4C+t7qq1u
TbRPG41SaR33tR2DZ/RTNQEQAhCdS+5heKiXYqAW6bOLfsz4WW27E0/nOowKDg8kmqDMuPTv/ysb
QnGtPtblYJbKljn56Mmacg2pqQfLulfrmLIDGK2elviB5PTBHmhRSJ37kAG41rwnHg1aJ0j4Iccl
IpG0/rjBd6AJ0FizBCtl6TH3bivP5UlY1OUr5uwM+lIGcrFPqZ1DchkRVb454tbcB+nQKNdtgwPr
qXUlcF7s+W5RTL0jWQ7U3T3VtupQQBCC3SRbFik4o/qa6cZR5dPjaY0LsNy6uaSe89zrdPLF7CLN
GuAgHnPIDGiYCNYhZWMo6A9qPcD3n2keV8l7TUNVAfSXSte7sJ9dlNqwXtvClGwDrXQyhIGFp3w3
+BAweB4OSyjv3Zgz4nCUxvfzHv0VroL22DnEPXcJW/yV8taOTcLpCiEylHsj4v84xbarP8KOrXsf
/B4xFg/jC/oTsGBai4WeF5wE5mve1A6xphLSs1sV16UngupykgxtaPIIVyJ13AjEiWRSQumzH7P8
5hfMbERr+xd2dOXlKAKjos2yWzhDQvQorKs2uU9QjzEQSnQwCDTXXtPhvMmSHUYtcADb2B6fnumg
47JrGp/wsPrGQ8DcuxEdgBs+o9G83Hpeb6FX2v/gXSR/SbthDpJ7QINf9XE8zrwD9HF7RvBLW3A3
TDrYG/FkuZ+D2b5Wiu1tavZhQ06vt/6ay9QGaJqb90cDevH6RKL3FYrQIxDttfhXKuwzMKqVGmrg
WrBRD5yDnQKzgwGcw3S3iOQUi0KHKMX7pbb+rompx7kZhq4kgS1K8yT1UH/OwISw2eLcMk+wCOu0
ZRQvGeXQAdDT9QbALP2O6NE7nTegjnrmyghuzW2QjxLYFG9davObRaSXWf2R9bYDkiFXPke28y23
IYCimgr0YwnD1wItttjQIpyuOTJ8OBLldHKF6vfWSX4oqfIGQAOlHdwmPzfVm5snKo5zixEafZTF
yE6mhxq33/XxH4dmzMCeOW3LknPK4c0hgOP1xDk5yWz+iXpxYhcV6dyiSOmi7MkPdWBLDraZumGd
Tj0WnsDuoxuX7kxGShCnmq32+rbUkOZIqQ9XGHDme00tA6FNZC8WeMVaN4cQ2A1aGYEBhK/ucxRR
vCgYrGe7YEOGc7fDv7nEqjfVKAxda+KUfToaqY5NNHA25/3NJFYhmUC/QdvYlLDGYWSOKqXSvy44
2YcgOP6X9WnFm2TTXDmlrxdS/vlLA3sz/0+RoiVY38QLrMKQ/iynoDuhYF7B9n7N4SdYrofQsnux
RpF++LGnaXt27y5LiRJOszEMZUMSnW6fvCE+36w+Pu7Bh471st/ucKQU8Spe071dqHFy5KkZxbwf
jk3Jzt4q25BIjYvY9QYVWlxIEK4COARaaG4b1CLrhYXQQ9YZZA1wDMM86Dw/xO+yKEc/F+alBevM
KIpgLP6BAeJyUrM+ZmIJK1GTYHpJlxbhHw45uIk7FkHyLcqjxvN/2o5j22uQX1IDpfP56EM+Aq5/
D+h7bcQ745SZuJS8CwcZNiXRnROB3epCt+1o15ovqZ77uZddSG15r9M5RcRrL5e+qy6jVOg8lkeC
LIjN7pqvGY+ySSJsCgD0HPM6AfslFdVyQi4V2GZ7N9lVlMsDPfxGjhfTD4rjOwztMxNKk2F4UMUG
iE3p0wA3W5qCsRPKmv+DVrW26YxH7Fwhiz1X2uJuLw+0ApBGjGU1XtgpjSY1Gse7I4yP49/PLWYq
HCMfvgpipGAyiFV9Zy5AsUp8HAJF9WTqNr4tlVnIBttwZP0XZyETwRlKqtF3bJUc12f7F62aDJIa
V/Lawlyf0VFB3afpxwLl82bBgztxm4Opltc6KjvoDx6ciP4jZNqSf3zax89kjmugHTipuP78XAlA
0uIKkfzNAajKhJI6ZShAN0D/BmIq3YttaXRZ1IenuzSXH/zSLrLtbCk4hrrUrFkXPmTltjA5zDjm
iB6d6ju6EvMKPdYGFCoIKnLcEQK1k9NsZV0+yy84cmyrYwGkszcFoxRKqOCnE3GtS/wYnFzaGhE+
OSr8LsvtYEXbwWGU9rnNxmCT2uoL/UfyKY88z6w/uiZleeU0O5ratwr8s5nDv3O0snQPMRB+NFtE
rOgdBiLgVI9JRuTz6muxw20F1Oyc/6IIpDkDRsN1RV+ChAtEptWbwK0cnaEaTg2rT8r8QDBXcpKj
WGXdV2+QUvFVm06s1E6wfGrX0v4+scvbA4hqa0oGdEkgXrd5d12ZWxRDJWi8/lZqPptR9MHLHVdg
oVN0mKRkxGYzH2pBN5fhPKg5MX2E6Bz1w50XcyMjrUUOzdsZW9MCpMx+oYQ3bt0fxHOZBZ4OH+Ae
tR7a0YUCcoZZdq3pTREYgBOLjvBdOM3RAW5JO89IlKYMVZTOVBUa0huy9YKa2Win+eEiFNMf4RFT
kr/3XvShq5Q1RgnqY9berDm5DJxOfJ+MoLAauRQ0Uinx4tfWNRCYcI80AXgsPT53UESE24aE8dbV
I1Ax6uKvQcuTt/siFVC7B4M83n9Q4hFh6aqW+n9aFoAuXSCUGOrsarPSVI4vKgfr4LSM2/Trv4q9
j3Nlyd+eEbnArx3dWY3yydBYZ7o6j4sLf1ZSk7cXIrPblI+9tkHDix7gKg9eL3wsPxKc7zyUrDoY
aYWeluinlBe+iCjx9pcqewCXzxIeYlW/qP7RBmCHEgrgmYiba8fUUZcVYvnJdOEC4uaireOuYstL
FlHdr7HBmK8nbUHGjGCDBChwWJoXBPQFbKe3gGjDzhLI4mXBC+FqtoUrYqBQeCA4fbl6ctcVYBHi
/qM4Q4bSPIWK9jTkfQfHq9Q1rg4m24saXKc9oKMx/1uOAlxQ6KPK8tdYb2JOyTIW7okny7hrYyoU
thkBUQTOmy6ifEB9VjR7v37MdUWmfqyd3XKatOmPOREZcc/YpUtvT3A+z4k0ltrJbR1KxdRoWNvI
gkB0RyFE33eq5z1D85SCMSJt18RoWoDY2XxR3U/6HpuChBe1uPueauqcivcIAYL47x/8oWQHtO5T
vxa0X2EA8K11c7ONQMvKEVqLLxyDMwW4ZT0esU62IB6Ob5glciCz/odvklG/HLoWkmm34ARLI6Rj
1Vc0NQQdNWt6JGlxbQ5fx1JD8IXsH2bszL3i3fmNcmt/vmpdb6D/NU5K3qAIBBlxYT/Tnl6hVgXu
6OLAOQRHvPrjXuDBpGprkwsHUskVTo3BrNmfR+Mkkrf3IOZaT3KX/8h9KpO5tNoJXaf8G1UgKfmA
tm67MlCoMoDCi/2yRawZoivb75MDmkwr7VDhG4eUmHitBIrwyW7kPIrmKk1TzLtbTEaOF6/gUt4Y
mRUdS45uaA0Ac1YhQmUTA7eb2JdVHP29ovErSUAnnlcxHURTX12vY6ogsTLOJIT5x4z2g08GRdAe
Hk8vP+qF6XWYQxV+h1VCYkecBnzWFQ5NLXkwnkskN28z+85EiziOo6kCtLKLD1eTKjqoTVDAzhe6
BdRtkjkFhFphq3jcEleDNUGCWfaNuA0OvnVZaGs32Jax7evldZTBDtUtxatumB1H8p/ew/qHgDJU
g4/SXYWvODEwmn0D7C4/VvW+/I39+crLP3HvlXKj2y1HG7an7iufFM/aLdKyf3KS9q2eYWLJcyHQ
FJp4apWub60tEyzvRPtWsPn9ziRsWf7IqvV9hoXy4gZQUYwOWHLcgtNv8B4xRtsu8pVI/NYHDGt4
IMpYUef0XdPpjIf+EY33K/k1E4TR8RjpwLMXXa6iqJISghVFX34BzZYshwo3eX3hgTKFm5A9H21+
ZE85MZCuDuHyZ2I3zlsKu/rrbc1FOjjkFyX5CSgRT/VrxrOdE9RenoOaflYdv6clLc4FlAsqLCg8
wvJWUahFg7UEWiPg5N1kJR5lLBq7Evv0L8rGgNsI+RlTAfmw0mEPoKgDcrw/GDankkorkxsiP3QH
GmChGU6ooXKzvPFbYjbl4a3k6DS7Fu7C0a4sySWt8wlVHqjf/sUKgKtW3DxNEJZ3gTiGf7I21b4p
KMjzt897z4zXu9dQzgY7+jfwj2Gd7CcwA275qkFV/GXxLhzSevYNunTB/ax7WPxyfsSxlPudFXQe
z9NCP0wy7E0t7PrugKhSrJtk0xqhSWF/oc1OFYbqjzneY+Pw8Lin/RlikpAeeXB0SAdsRszCZZg6
XW5v4p1N8c5CnEUrECoSaoJmYxMccw4yqdHmc2j59AKbemX0bZPsAIWqXAWm3rH8xc7gZnnm+/mR
uhx7VGaDTS021pRoYMVzuzvk0/zyJ2se1IVmnOY1E1731ljvmURQ6GZFrPY8sntZzjsuAHrMxhxz
+fXvMR41WEDf4Ptvdtuvy0pivcKJt++yETsmXyRxUj+/dA6okKomNxQVCf1Crnl4ojbJrm/JmNbs
a+Mvgv1xzwviu0vtE+V8jWPQYE5xehpy+3euh7+Je8QKmyocxcUJk1KeyC4n3Aok/FCiumNZuQ4T
JrHBl+5OLovT8sV8kVlb8aQBhdhCqbJZF0++dLV6Mj8ry976WRJcU5Ib1nSoHl+m+YWGyIwlR2q3
ugkL13jSwd4ETCVLKXPJwKlRY+WX0XnOKcSWTNGT3Eg2vNIqfv1RCw7cH2lTthJbM5Rzfww3KYKV
XHLVkOeEupOp7nnrH+BZcVhZ31gmZWKl8LEyPWF8teWjsVf3HhpymT+UASc0d4qEFbr1v6+Bc2+V
Rzy0M5QL+Sbgpwct3vFyV8GSW5GdtB49Qswg50fjI4PRnBZC05cbj0vhLaz7yuTp/Y7pnhGUXj85
cK3HGTe3dRjTas8qR2fNu1r81fEb8ShzEVMSS3jYqvhZfbzCjmvh6k2L/oaJ8Pz7I0fPHICveruw
2XDasiPWiNj+23OvCmfTfO7rzxop5h62ge4JBia2Gb89bL0DxJMT+2ajLyfy5iJ3K26R+y7iprYq
VQtIz6Wp6Fgmu/u1ZcqhQO9qh4PS+0gd7JOqhxSwsHQycd6F6BNuqqFxhZD082Cze4d1FdiTGcPx
IWp3mpR/FBeDsCjBVXNVU6ScNW1ey0BA1ndoPUyghTQOb5vwXrRBYtuyAm59gUWIHBc8B4oP2m6Y
zzPxDWjvJr6cRRbjnaOMB7voWvWhk7M9g8CnHEXjcycLkvi9ZM2p3bh3kAssSfGv3y/30Aidgtk6
c5zz3TxLd+JLn8flcjcKYtfZxA8/OvMTeb7k9mMZdlmQ7GTf4qKgzpb0uukcUilRnKn8u98KWGRo
5uvzXVj2CPolacC8neXd33qXUKalFUwZVaE5z6oGGgvKubfFSqDzUeXFBznN2JIkKWfrPQ1RKWtM
DfZF8q9O8oeDv4fDG3yXk8rLl1xWQuXgMFmsikVp8Iyh6r/Ln0MlmC6XDgPGfh59ELzVwjC1BL4E
bwOeB8uJEmImsDOytLe0lpEyMCwPUVjr/+euPud4VsJHHpbQEmEEpARHqMmdP8AcJmd/YdZnqkDg
JAHIZwPlXNP/v8nI5VPGEYmBbap0Oh4sgtQorWdGrcDtYv1gLS6xjZR01bdhC4pj5i1W+4y0x5kc
1Xa6PvMo7Yze345FTE12wMJI79IKpRwpEufaVT1Dlg/Nb0obr+q6ZI7ISLubdWGC2Fel1WDBqy+o
osjQ9OGnYfwkJPly7BhzWEYvIOw7HeixNFrki3vQs4+0YrS0J+EPGJlb1mEIgXwV0ckL0MM11mHD
T39UCSVn4f13SuQITEMeixCtNoqGppL4nrkSh17v7BesVYG7XBBPyGVlP0kkYcttVyRutQ9k/fLc
mO/H5h05sr6JYifUxw6fnoFTPUol5XLyWc+yoVYPFXTLldKkKagswoKKwxbkY1RlXVoQR2sjwVRz
RYaBLMAPjRZwLVpkikCXN8StwJ1pePv9NXSeBpk6g+ejcn80HIJZ6aiIQj5WAc9GoqZ38VXoN7SL
e5u6ijYCYAWqYkcrjJnydWHsduknYhUCeZlp4tgKpGhGkcbcPcnnjb/0PNIR4/juQMwJIDQx2sx+
aB/g2Ph0GUyNOADiNgYFIuAR44IZhBoTz7Xu9OWgucWoY/zOz+sim8+yuc1cqWfsWLHwFXZx4p26
B6WVjb8SzOLGzJkF9eT7WeoBGPP79hbRlpGbPl0Gb5GXOirINspcK722MYb/zRTNIfsAL4tFdZGo
PBl/mY4V7TXZamNcbcJMqdX/s5O5DJA94yTANQ/r7Fig9e6S8ojBhz+gHTn94+MmrCd2hZ1sfRiH
zsKgW0q4WLDv4s4E/FPfvVXNykALsMz84S2F30oAbKgSHfxsoVm4W0z7gZqrmtMmW00V7lqTVQFz
nFflxVgoyW/l2yq9GoJRRFvW0XVlRNVh/r1RVYPIncMqg0K9pjExGMTtxxuThHwpGoYNVzIQyVGC
VPeSuJrKmDMq4/Ba2Y3G0YERNY/SyNUr3kPGbA1jOLJWR6c/4kKIJOxjy6micsYkwxqh9wUc26Mv
WqtxVElhWahtvM2Brl9KC950YyCNHo9raHBWc3ATzwD4Uq3ZrnFXOHyk0M5XiMLYz2+TVkFxm4Vn
xg1MOWOGZ90i51IuH4QrF7nAIBMEdHDrixCsHrX1jK4lZrIBB1C+nJScxWFmJ5posUHcnd78Pxud
P5nVGKypkd2aN7Owa2KBoAzCn0J58OhKZ9pagxxMOYLmAFGwTsHZcg7l82T0rypQ9SRgaBHzGZkZ
iLsb6+xzKv3UDQ0qYC3ey46ffIOURuHcAmRU2gauoOaH6/caA4OW9KPvUvQXL9TcRzoHuXoatIX+
L91P2vIj8Xguy594Ozg9INU/Yri9buDGqseZMj/GzHxW/lD4raonVx2ACgu5sTdQ+GKdr4zy6e0v
7FXWRHOxbcgw1I9Sf/O47CT6gmnKNZZ4sPi+jZbwvuzPoSIIa5fi8RflGOvaF9zgn/dm+yyT2r0h
E0m4arZwofmy7Z8y3C5donTni0BJStZSniw6A4z/Jd9lLptINXmrfUKA4JYcxeilaiksm+XRMlMZ
bdYpPC65zzb/j19XDzwf7+lb/2CCqkQDLqLXaGdHyRU/MB7rGyvbD+hn3JRcQ8+6NQWnVKLOKWKM
HTxTq+Sc3cc50DUU9ECqd6C0otbr6SDR4GN7DPCmMD4C7jezddykgdu+l3x/TW4ruCmCz7OaBafe
/0Ctt2C/XtD3ezxpj0lm7FSzQFO0M22SH339rVUSlvJWbme4+y9gdUFpXye+7V94Qph47rVlB/zc
pR/ay2X9fnRg2fIaetxpWo5yKGkCJGPWedaHeRSGE5h6UM1vkINCvYBxCo+luMNLnfNvx2ppTZzo
5egJkPnUWPkf8qDl6AGm7PHxyCCr1RhVlcSy+Kqds/M5Qmr+MHfW4R60wfdcUalNUqmln1ExU3c7
xSTGgqzE8ryurqfPAMSA0yux2RlW41M5wSFiJG8jLZI3rnSkSTpQtZHi8jP5bzfgukLqAPM3xVd4
tmOy832At/rHMgNncFg9j+o/CE8RFm6yqC+utTZ5MxKbEzmDC6IWAU9eL2y9vTsdQrp7AmCBv+6k
D1OQI8H9x1wFW+UHuCL7xZz/tDxv32INxuIWYLWNCl/KZPTbQdoMfkhQGO3lUP6ggfWNxxw+vP3j
2owq9AhV5IrNzvAZ6oGkoNFZXi3X/8oC/sJKBn58dGRz76m3v5TzQBUBtSoInCIUdSX3Eo1CLucF
OlO/40i9ur8NzORYqLYw8hDPIfoyXTXIwOqbma+FKK1Q6o24yJqQuvYWqiHtacaGbeH0upKHxRZv
quTWXov+oA8YSclCcl4i5nMANRtpCzeFKtGvT//JJu3c7d5dGrnoYGYylToU468jTiWYKoyPYlIg
3GNnBKW9TIk2IAtnJJnyduxDnLL/jDMs7vtWmihV6PW2ZOiDXJ1dNxLNeXO/Pfbr11JcMc9vYs8P
lFgw5SmLiab9l1vSRsSlEvG2lCUtYdodAVR2HoKlLlitIYWJG8xdppUbaAorie/r/axkAfbJCImP
X86bhZZtbjGQwwv/rQ36qUD3i3mGc0aJS76vfKZJo/7wwuHl6DKNctdYK8QQHTT5Dr3jf9Zu1d9C
yjCig3X9iOtoCbokiZnLwASVJ1ZKq/yT1N1p9Q6zeaoTW8cBJ0KXY1R759JyZFTNjTJc3xGcs2sr
WdmTGnwzjrY0SXlHVVAnRLAr1dv/mXxhh6v3gsTXtEGzU1ipMVekqcvOdzslhQgiyfTUFcv3ceAH
B8DZddKw3h39WVggsA3zKk2mIFL77jV6lv6mEYFfoFB+/MN8of0ozFF3p1ELutVQYMLwxRTeAhlB
08XDicLsmeF75oSUfi9pbiAZKURAQRHa4kph5FJBQBEf2ykqLgldesekYmybiXcBJgc6BCgDAnT7
j2uQMe7LHFrz8arxpT4rSzvK5CRg7WwuGA/PeFV59coEppqUOfR/tnIGpV48S9DMKWypU3aR0104
YIjC54mm3H716iwv40J4YVp7CB431eS++YF94S34vqWiIK4UFcVXrCpNfhfpJWvl8hyZPjWiyqaz
aF6uKFFEZToyEW9jh2Z50j7laf7TVEYPyXANOK/BAI9POrAGx0BbHYfZaVtuNdIt/x9TzPsD1kAQ
2c1ZJ2N0YQxQPtATppOTAfSlbXMuGbNCjhsQpoBFVOKLXfqHyeEZ4YFJ8HBwxZHIJXmJAE6RvppH
fv0zSjwUL8lJWhHBlojNBGdTmAb5xvXQa1Ij86ZOizkF58ZJyhyh/ykwCd7V5SHoBE/WQso7F/Ix
iyBBMWOev6qEW1tkvhBC2G9vcCD+tFnVHnhsUQ/oIsWrEstzhf1X/Al6OITDXm8yrbnvYtLqtChk
toljwXBiha2QSzqRd/Z3igWvgsksuP/iW79//ZJuRyEToY9F6yfB9ce2xr6tfzlR3wbCNXby1nxo
zPxadGJ+cxJrIBEeqF6X62T+PgSokpUoO2dPoQCIHSYz6m0Wd5emWNpdZ55R/ezh8avzIScznPVy
9IiKeUtvTyYohycMe51Kj/j+q4zidnmk02WohrfUIPMlZvCVQOjvOACi19lS5VxyJGarqc7DU5gB
ld+GPGeyDVSIlyNl+z3JVSFgObS5SrtgoBaV1RkbPtjqZc9JgWx/8y5kptQswRNtT1fSNBs/ez6O
aDOW3YWUqL3DIaVfNcwBYXU0eH+KtoEerRuhAj8TEzvMMx93t54B0vSUzGT0Nn7qeaXCjzCwvVwU
uatUpvESMMn41GkPkJJUVFSqADEq8RR94VfKJyLzZxPB0dKX3Zwj6QFJY1ccrpoyHukz+Fuhlmx8
Q/ZlIhmCOlLto6dQdVWDqxTigqVbTgaEZJYXX8+s8kPCkBO79fPVZBVVpLXm40tZzv/EWzpRr682
UVWt/7vWRlbezrqYUsyl6cMQw5oatDrt+lM19cjS/+2+MlZWlpAsS8Ry78Ohh2XOdFsmdg+wZr9B
vPWyLgcQyIh71Ln09Wx9qzR5IcopxhFROUkPbX4xPvcxIZQYWZ3Z/xsKzxk5taJ9NAdmsqIF9oHj
UP8KRwa7SAdWts/mhmVWrOC+IhVES/mgg5GcCBUgcNvyPxp69gLGxWnYG16JZlk0E4vLB7dN6BvX
MJ77wxD7YT5MyI00NrwwGTuz2jkOE0ddpUa4YCuhI660yT3Qy457MJYOtXHSHiNJMs8hTKpoK+JH
Qqd9w8UjshyWI9Us060tWTiWtwq5WtFvRrJkEQCdV7HAZn4Hd98BCiyzLxbIX+l2anS8vmg0dZku
W/cEOLpiy5q26l11YrwkWYROCeJa92GlEryxHqruckIuHFXwLxGWgGr71Ci7y5o3jkv1TkuLuTQ3
pyx/L7KSXZekZLpyC9pAM9h+FTzHh3Qrn3k3Al7nqz5EH7L6DX3xyZhMrBPZzm0+IOB+U7GWWutF
hYELXkAISs6sPF+zp3xxwuNT9dzgkv/BBg4/MR0OCHgImFgy6snmqfyIMAVdj47Hkmi53jYNI/0q
c4HPSi9R09Xqj1Kb1X8RN4x+G+krHtrhtIqUTM9Q8Y0k27zA7od6HmtVoAB+G0HGtSqkteOVnq0T
KTpCLE9DUOtKO+H5w14K9L4mnkAMdVGdgd4bHZpY+O7NRBkf1/XrBkVKYCT7wAPvBIbHDgaKXdPe
lawZpGvOL5zdA/8aiNMsRmalMMlOjBd+vZOBaaiZyEecCCTATViUDOT/TDWL8Z/fNkK1BjE2sml5
hSioSXts/0Qc/u4kM/FKBw4Olh/UHknLxS0rsX1ctDid6JENMk810b9n5FJD7brJs5QaM6d2Huo0
WLENnB6+QulH047SU5Noyc6a8y0AoKL2dvnBhwG4L8qItp41TVFId0567XdxaDd6i5gZs7mQ1WHV
wzZxWsrpOf42ZLDqcsJ8Rnap10AoXTesBZZndmoDhPM5Sm/m0g06b9DOe9Fz7GmELQ2n+PNMZbFo
WcPIT5QFn7n5UmYgqrKt0+vg/Qolxaiqvp1wkrmbCn3Q9s9fI2TztR/aFYUiIx/A9BTm+FAx+knn
gbUwYoGDcPpZ6RBhktFmSrjQwslEz8q2plaAnpjAuFjWlmeBiX12AbQxDZ9Wt8Yhx5fb0/t7N83L
fQ3VDSbb37lLRSgZbt8KTYGs2lnIz04Rsyet6R1Cttc4D549/GV9fM3Jr3Qxqy9pPM9VmOswXgAh
KA3lq/Bz4IJPwv+20ib7EyuVqkfDG2xBlWoxoGVbl0r7IZ2UyOwHr4BU1TIMaCoTClTd2BOpsz/l
j3PsANcd9oTEI5asIRp4zzTpOFWEk9j5sfBm+hKIiCQ/auVJbPs85tFxpmxOqf95Op0xdvXKHdCi
O0f91+ZnWcpbnYpkbi5QF+BphTC1diwHYTQ3yiYFgMuXw9jB6PHI40wWAh4bTsZhescD1zOY083i
k2tmNMX7nQ762TQ0J6x7lrIvm81m2jEYf37JuxXA0MdvqJsvnLoBH5G+UhQ9gY2j+c1e56KV+LBz
UBDlSvM91sAjijGniQNnnxbWUU27pBg51HyOWXwPnzbtTJaYDLsOZncSqniNhIgrbqFUqms052B3
bnU3uhkDl/3SXvQSbnpPrN21Inq5RzSCphEDDAU92E+xW26d9w17aZWm5k0YPNCOa3Fv+1MYwBiW
i9AkCJfZNWCmmfNJ6BtneK/yucMBpKujvj19QAjQCZKvrGvOW3eSvX67FJdqp5TipFhwXnvyDfeR
Au37D+6OW23CvuIHfkHe1JZof859jYuO8VgYIljqhEz6CqCYvKS4JNTJH2l9PptttDa/he2csG7v
WwSedcmvsJ1TquXwn7DXZ4zeA4CYUJkYcb0ZHuZXaa9tOXTxk0BXLk1mLhP21qL2WSLJr+iC1/r1
uAupvfZr4PthN/StumhaqYIOak8GSDAXaQmmc9IbJVHosgOEw9AxTChd0GP4VPw0/5v2SIxhF+vT
R4HDKX6aZfq6rY0F+2oY4l+HkhZIwHe0zQvqBwKp8XcupoeH+yMlRgrXelUQnTj93cbUezK4OERE
xDhAPi+NN2fDjPCccsUGZUfMzfGTXB364KuNHylCgcdTgRGVKbjAgDdUNT0MbfBzSe/hTkC2io+D
itJxr8oC29Ya5ZhJaYk+1g8graCEduLeLo30L52jn0nB3frX0N9+CiFYMo6AzOG3l7aaonq9Iwr7
Gl7jxTxrljamhAj9nmy5qYJv5LdmEH+Ui3i9XipPgV1zn7yXOZ/UX67R55iZRFGoVpMsq0pseKCG
4HXmGfcv70gn6p/xpLNDqGhXhcItUNRVgr2Aabp74hNbAxzyXT4cBdQDxm9WvcfOPMvucMpLs2a0
KJX5iMJ8Di2BGORTBrVZtSh/s/qrCdcnoylx6UHPtVe0LU8xlSmaVxT6++RzsT6+tdbZY3NR+jxX
ALLc7DXJ7ENUZqShvM0sOeEDAh7of+9da5S0o+UKIQBiZJ3gs0N0Nu3XdzS5mQz/7zQctsJbm+1Y
dpZialHnk0fvITYTOrfJuIIgMmX/9IagKrHeTnDxBPbcQJR+jvSrzrJYttxmjmfyjtf59JlOHYaO
/IYVv2iZM4ag9FpySG8IWzAHMUOlCUj7eD74QrcFot6o8ncsP7+VGC4xa6AV+uenS5MZ9EZh+n94
RctgyxngX+svBaQh95Vw09RcIs+i4+0wjP+XYeMCkBdKQusnC3yvy40kU2XTT2VZDRz2XMEV+CIM
vEFhP+I67bCfngAx/4hzB3Mj3/4BGzJG5D6hjvKlNQbOm91XbxAuqJ4ItLv+ICha6aXvejG2bgiR
Ph7khiN1FFEmWUD7NJB55fBJAfv7stf02lnoFX4EiddGbL/m8PLU7bxoM0FOvPE2qKzAvoHW7uWI
tHP1V3bv8IcZnVxiD1d80dotVhi5lSo+FCdel5SpifawlUqob/eLFVGMhcwjIDoXmp/MyzYPRyv8
PqIbQMyTxzUTOGqhO8ICOTxbNa8L9SL/iVLCtzPp1K8Oesz6GCNEMV2lJ9uCVM0en+up0k+L7Q9T
aySaoqhUUgKQiHhN1Qs0uN96Da/cMfUmikmvMzwCrpzzZtavdoOG2gEmd5Y8Fz900molXKKob/w8
BRrYiQAQ/YLgYHzOo916EyckBMm+hApgi/BxQmdO78yKW5d2OmNDdcEmAKKaH3lmGxBFYCToE+Di
n0eXS6RCn5OawD6DC1ppZ3zHGqSDEoLJu1E7MM5ltSMfaGEq6OYLKZm+AaaedW4S3R2UMXc3XAR3
sHbfpruxpLGUgrK/J7d1Se1Mi8yrIwb4GgIFStSsk///GHOf/i8/nOHE4uAvp8wGkfmtk4nDPggb
AX3np0PAZcFPLKC0pvvgQ6PEHs5g82hbJdozhxhQvDO6RH771dO9NhqSAzF7WXZyLu+BBmE41DPb
7Oz0zLfh5ZZ/SGCX+PdTX9smZdHZfafqMsVytSrp5GjJ1OrJH85YqkqLgjcUVVY1zUS+biSZGoRO
kbEOUmDAg5fCmilFpIoYsVZQpwvbtNL9fZsa3TTzVAzhVlCbESYalZFLebESrKjOI+QrC+7t0Bfp
rqMvfeGtCAlAcwJq3aP4AFhUQ/FnR190pIFGUJKWeCyHZyjvwkEpa7QHyOiae8vJ5hprgEnoynhy
aKCwiqEjy2p3D2e506PQcNInnyZyH14WqCEHh1ZtgDSpNbPSP+8zXkvVcswOjcyKFynvzN29D0Xv
ABpV4ImvxcNS9KBOoaZs/MW5iFRWnxDE3s5z+BmM2Y9J7FSu8YDW6bX2ef/zngwv9iEVFL1GdOrC
5o8ss1zhkqpJC/cB0ox9XnBcnoH/eN20MqSrAPwLJcMDfzW2ZbktRBwxlE+I5E668vG9tZKgG//z
3C3lWVclmhH3TF8RrwFkKvCpAgOuot48QLaBpmGUkAhEBlcOuJzKNy/w8QSh7mXrlAXvgy1Ug8gl
RdXMlP/tzAW2Yoi1Ukwa/j7pfN3C63UGW2xAXr7lgi64PKqTvG03ceuZ/aHU22Y2LJEJ6poqGJzH
2Flpuq3/yyWUs5OuHCw/vkm5EJOTbBuMS+3xUIf0cIiB6uO0oUih27ntKe8KHyhDqOKme+mu+73n
MyFb1AKi1YwfGspQb2vN9jwRJ6uMt30J+L5+Fi1sEOeXWUaJJZb1MehvaxHEHlX0WQTK71l9AB5j
rJ5EAYiMq+zQIm6s3tdphTJ0UYU2FzBke5DevL0+A0CKSueJp7Ba1FiUT8E8icNrX8sk8uYmbMX0
1bPqgNvkFXMCbPpWz5fHYz5RXarbS1o7KZ5WSU12CKUZc7r6BLDM3gRC4O62JwRG/iEzGqrMn9Ag
tH/sLcIK3csriAouqLbGmzqMhyMUrPTuOPDWVRxP0HR02zOZmkbjxdZMml61vaFQi3lRzBXjn5NJ
XCfUw5bSUU9JseqAyEyAlslmG33WUbM8+P+QLeHWTbT7vGOOiWgkMAmg5CSqPGWc3HoOgk0SsG1k
CuANWufH8PPQ1MEFppS3L7NzKvnIOklqNxdFphV8xER3cvTzDQKCyR5r5Xc0B8LfvlPUyx4RtG7Z
Ut0JEuz6i28LjiJOZwo/Zmnt6jCufmGKaea7dAV0QpCbV76JBa4KNFy6kiE5ku480A6hYcVfm0Ht
ZloLh6xf/HlTZIg6fLDi3AA3MZytqSN2Xk7F0j+S6Mo1khQen96+/O6ZFf8y/KcXlq6U2fGQBQVr
ZklLx7TPcACJuHqcUM7IHdHCvmNQGwCbsEQNXnde0/4NaCZzIQuJHHr+Kpbwxnmp2abd2T4c/+/r
K8LDqbtPf2OzTiu8ZEYLJapxZDo78ODsd9yAhoeJC+TgSPHk96sDe5IOgKumla15lv9Gmi6p20D0
YUL6W9yaUz+G3Owlf/rk2Qgyij7BaP3SmNQ2zc2lta2P6/40GkBE2ST7L4AV6gCLC+vciY5CdNVu
vv1t2vGk/qxCIKzKCzgoQzEYmW/oxFyQnk0HhO2scujamrJD3OljdaLR+rOwKAI8cuRTtyfnsdQD
8MVDc5CakvVLX7K2Ap3dL4MVY5Q41SEn8cNwng9YvIs8b4rFiqwlLhCJvRK6nXZNL+kH1t/2hnq/
oWZLq8nRsWh8En41ZFcj+fDn6f3RdDioCohxsafRSa2XfiQkyGrn/DzdvAPTam4Y3gF/Hz86xdJW
85oRetFN+G50gl/lP0ibX+px2nFfeD2Y6mhh51pSfpNUAGG9VjNqlBu5rUeYdeYrnovWxNC0wmiS
10yd/EO6xkjJ/rl/GmVb3iohmBvkiiyOcuOo9OD+ajRTqLlIcEtRBfLvCleE9UjaX1WYIdy/T4B6
hHPoGaYAbn30o9dDuLYJPMxxJLiyBMHlNYhvxWgjD/VSD7evO/GMOL+rm35u5dUIH3shm+HZHB40
WonWVU+MbyKkjz92wLtWlsLw38x5dPrO9gt4YJ9y5Zbw9EZHK7qF0l43OtcIItj8fQ9WqomEQcWV
P7Zhm11F7VdSqIoCZkxgBthYk1uAZBd6ppn+j0EyaYNs7wCxIIbPypZycZJdAYMYItKD80IMEG5m
l9YNew1Qq+ICBPwWo8HaTetTDwRIdYj66IIfDYspV23Nz/bTIGF06y4+1AOsGlKxFj1uVbUc8FzE
HUdAa2wrd7d3IfO1xeCFPr870CBCyjhAXsp7F2LI1oxlrmiNkTk6bxrNgMbvWTa0vXrrjf0/JWZv
nXhY7/WsKo+aPdcdpDiTv54SBE6hnmaeOWyBRrs+wdIAC+hbzTmDGlEbstNK3B2WjZmiai+Nk7Uq
T9GjLJFJ9jQTawkhWkLj8e5ROyta85h3mCUzVSaFyWEBgBHWLPbFLG5N3/oYpBDVDqNG94T9Zlu/
JtQ3B8Tu4gSwfAObU/FF5INOnxCrFKhmQpm6KVifhhvZIYIcExjK9mJ8eKYmC6Us2xslZnYHyeQA
/MzjGh6WeV02KiAk6hUBrgldt5cObIZrGykrjRCYTmGsRvTzkkr1oaAUSda3cRxVWHzXmpSj/k3A
5vko4yT1feJjyjYCnCPReQG+vhZg5imht2xdjfYbvCc9AlsnUyIrLSA7bGCL9gbLgkg5nFDduXMV
pj2kU7XjG3oQ4nxYi9PZ3BzgBsxTxGDnxP1XCrCquY1N46DQ5p1JoUXFqWCu8mV8krsZ+PvyqfFR
VRU9OAoY4xLMyDvPNHeezG/Zef/ZuElQHbU1cM4RZfQ3bmZwdb9tBkASam3krE5zWz91ciG++kDE
Dbb+iChtMHfLRkWcgquk6ATLe+Z+yqOGXANdX+1Rb/m4ipcUgJX5dzZoYjbSBf+XqUpzqFXAff5x
kysEQ6D4reCvH8xQbv2oDxza2tF+wc/uqMc8lLoodV1lY71vCOHncIy6Rfv5ZILv5fbJvmqj3nes
apz19DPEWZifGwPd7hS66tbbTS8Ieq8TCyl65glCcCHe646TOh2UdfmTAXWYAWagEpRf0z+196Yj
Q08OZNPMl7KG/c5FI7X2xOjqsWmpa/MwTDvovaIooADmmO1csNaGC4kq6GNyuVORdoiQa7Y9Z1br
O0aFJDxLHf+WGQ91r8zh2u6ON17v0I96L2LJEm4SoZwSeKD1TVxQMmJ9Qt+9DDwoQjhr25zKpj08
brPxjGtDOyPWz0EufIXMgdoxsmexvuzxjEXYrZbcXgDpyxM0a1mpI42FNJXlMGkGsKq6AZwAdFqM
XPY4zha54sK5MzQwdUwIhhyvv8V7lrBgBvf0NGPOCgQs4mtQ5+L0q1Zjy34X7wTPEeDOcQ+pWsQk
AhWo8qySMx5LDRX6zcNtBait+TBzvNB4HWOxYxtC0iyeyWf9No6ea8io2zbCygfg2k2qeDQq77+1
TqgDxB3ldOa5A5Y+qOzmOdcbljvYMZ6EkvbOz6IBiALdoPdJm6sTLU4z+B5jpFddznytMFh4b3V9
eBQh+Mo6ixT2DysUADR6JxGpmF8PmAcviAtbBz67E5sO23iunYMliIeTv5wrJRz8nTVnm6kNGDeG
+hT3toXWDFe1aZZPIFO6K2YBKeD+BXPNKtfe5q65lCqykP0KsHhBgeTi/0rGDOHHdXgVD63tsWl0
BDsEZM+tWfHhJ0h6Y/YOol1hXwIUAc7c+dLBiIOx0d7bNZYOhQH3Sp5bipxryVFh31mjt/2lW8kX
gvXtBbUP7rU+NMsvkWLu2LaZSqWdgfQ1Wy7WyzMb5MjO4RJGiC8NBP+FCEsmHuGB0c7jV8XJQdK3
x6CkcBSqDiMkHM2Va1vElnQSeJ1vurzdN3IMKQLDdF86NzPYjkUbnY2B2L7ygfM4HfULWOAb5cit
Uu1Up4iN59dNM3RT7d7UvLYoUwF+M/75FaHVcnDqdCedNLyMPV/GIgDozHlwjWX1XwtdyZ0DJjT/
k0ej2ePEyFjK+goY9OI87WkRUNprE0xJ3+3tX3oQId+TGhnPA9SP3x0UNVwjZk2tRQdSBYGBL6lq
XOyPHjvwms+bgXNwKwrVMbyhFFpJ2t8GnLcdKM/DJotCwshA2jQuzevNmAxIu1PysooTW0RPjhll
vhDlNoJtCBcnnEdBdq4ncnpBNeOWO+WVnFL9oUNJV1He1QWcZ6709OeqDdfq0BP1vJgye0w7ERuQ
5lvPzX4GcgiOCFSaYvKSRC+bB4icLXxPb7IFXtd64bbZRhN7BnWXpyUFleYMzjF47SFa7mF7/ZS8
NpiZdQA59nmq+J/Sm25gXrYyZz10N1PnF5IpLKW3kmCNcIiKHJjVJV9IFKkgrE17RhfcOvQgHC2c
qd+KLyM9ilMhO1GSvRjDgFcI6kFqHVpmMYZUVUsPNmCwbTDN4LQfYtVXb3Z9TQtgek1+otwWqtrq
YxXdSQbtraFcCaSTr2l7CEpv7yFZK19zWSz5HMimHSquWR+cGSx0AIy2EhuLIkM7vGeadFx5ozO0
LQcN3chONfJgArCUuUJEH2mOD0v2sk3353p6TMwutaH5DVVcghbNkeeyFUO1ZQqFReIjWBZBYfNR
/WBxXiQBEVfH1yCkQ3yWwSGLYzE24fix34dF/rE9obRLl+/1qzGmRZpeVmaJgvUS1QyHYh2J5HiG
P8oYSPuBGykxwIjLzyCMih0ovl9bCsEBX8imA6UXRB+klIbRn/nqgvAs5Bj4wuSiYPysZW9nlg0U
GaNWp6j5ptOJHtWjj1gVvtDI4Y3Jo8bTDfH/mhHSuXbSxoimi0S98ZrGmcpJp30d3mM1E0nCeEwz
xvFpjuhzyYDu8aeuK7QcdvMlQeSB45qvVIgKHBUbylUmgtibsk6a1MYl2GvVCkIWzTW6XFObnNrq
gzLtvDa9/eWlCNp5kOuA8DHchWoeScfFoKfbnhbTuJlA13O4vuRqsz1WSCCfFUsSWt/ig8t3T9dS
ZlKwxOFa3fBzEzlZg0Cbusip+hZBFIluihZ7Rtpml9ssqpkGEEc0n+6zAqoa8S5hjpx4is+TpCmT
/CozeW9qJUxKUBUJ/V4Mc3RGvMEAmWEV6NXCGhTbMlnj79yQVkDkxdbmLIWPKAxuecX3a/0XaXLP
IQkdIET9PolP5h4R2QpDtF6PWzipwecYKnX41DzJkamQ5z3trFfX5DoW+iQncYq4DBsl/SdgF92L
xb5pPunbf5PUeLqLmmHBIpI8ZWxKeGfPC/IQrfuuALSyxt1G9GYKQe0cROsqAj6VBfaW0feMz0LE
C1TtqgXDbl7ytDx51+MRdcUBQCXRpY7ugpXosmWr89G6teo1DK+rZATD4ypI80jXQdZA0i3JwjsF
zLDFsOHy6gfawl+OT4BZS4m9BXGtPEP2EpdrsWpZvefTUcdgXF98+tBvhThwT6NVFE5GKy2Yzt0n
Gw9k5J7s378XiRjEkEItyUSfBCQHOKCdHX2A5md1HRmME9yr3qiZvNnxvdbmyBi9JMyWohHr/+0F
Y8ewKreu4Xdy5f7jSBOQFoy++CBxPMdulGSsWvZJZG7Z0dY4SaSHR6WwDP6OkjYEwqtxDRWY0/Ce
IcQbuCEjYtZt+0IiVQMu/dlsgedo3wkQ5BjbzPQRrUPhlwLi75KCZHgKr84ae5ACgPj1evn5b+Uk
mAPdtkr/0Ow9Z/SDiCe65HRU/Cf1L/O2o7CB+d5xsW0w30mIU5gFYzlrA4tpEG+QJiA5C1mBcq8u
qasX+ot6Y56fo0YPnlIhvtG2qW2Hq/nSQ0dQ3UepDOwuUiVpAEvUUfIfhABJbTmCbh/zseYfoF0s
jBolZ/CSXZISzmxZbtqfsVRXgAGJzxYYMS8DFNs8cejj+NrK46GBnv5mCuzzsMoTst+3r5yhF1kn
CPh49tZfbfwYvd/bixDg/f6t2BxmsqlaOYW1DTGdsfPmRLO03LlxOO5g4oxOQA4OMlDNhTkIxdvr
PH1R/rZNHTCCxNx1SUuC/J0Uhuup4fQaGQJA0NXw4V6FD+C9/jld5PsUA49qbAEBQWRxmiOurUpC
XVl1rQaxStiCxP2/aiO6jEZZSdaT00QEQEHczk9AoQQprT7wvVEGlQE7TBDjenoI30Za285drvPI
0bzoM2eQhl98Xb1te90D9HQcYSQZDLKLBfTaFXV911qi0b1nKCLZhr3jF7fFqPlUdBh1/HWIe1AZ
6KvG/H7zq8ZzUsmzco1ug8JaweX6RsWlhZpKUa5WyoHUH6qSIXrnxS+2y62jntVo7entY86lGhM/
jnZopg5FIsbAyQD7Y3khZ66gB8aHF+HqhkuCS2kqg3AmcK/1z672ELD610jN8QOqEdyE/yEnHmor
N4I09Sp6y1sF5F//3x5jNb7/rxSoYP3f67etsb3qw1a8cyDuE2YahL7871nAxkZ3dVt83MYin7K+
E9J6Pwz89uwCOyX/Gum2wCASlm6UjMrwxYMalqqNxsy5oLWEelj5v2rmNqIrL/8CIHz8ra6hlhtn
dQFIcg8XOp0hR8IYWeYUModEaUBYxpqRlh/XVFrcOQn8XEsihClGG1CHbFb+Y6d8LfG3LpsOAewA
PVM7r3oA1a1KpucrA1UObzrjfMTIqKbHL+HmEa7lDv3qbQ9/1wxFExK3aBZHyJgXcmckLhN7/ijb
HsZ9Er+y0qd/TdSfQXeQ1quKRU8IbolE9OEsoTvxLmaaovPkbhj3fs2DNVNZkKJefC3JS9KTrRsY
O2+JZJf+oo/Sgx9HKFZXPbUBSgPI5tAFAi8hm943BDjhjdJWxka0xiBCqOYbowKewCaKBXj5ferN
ZT0m8Efdq/3mc6rPjhHupfmPxRK3Bwm5xJseqyIC/DKVd6owAp7yhv6tq/KO9MFtvpyABojSzImD
1VMG3Snb4BpnCagiQHO7vz20t5BHftECv4ClOp4QsFE/C3jsC2p2eUYLNmI9rfqPesqGWmA7m1bi
4ZThS6MeYIT0VotPv7Hb0xpusy5xqqDxhAQCEdxjJ7QCRDWS7xMdHbcn25IGfrMPdYGfYsFuJpYw
POwhXd8mZJWzif93TksoTNw2MZ8XhEcYdAJrEcsUdDppNlrBSzdm071oCB0bm7C2LK+VPaFlOrkq
ovOAMu+pQLYbC1VUs7nuUaArnD+q0cNL+BqmLlMQq/vmwBuiaDQl06uTZ+OpBCBj4rXBAvN8utJw
u6jxOm9VmBLjVLT1x694rW+GFBfnX5MWlfXU0SMRZDI1TdIjnrksnjNf98jOey7bV46rpjntowyC
TjkGY0ex9iPNYlZ23UMagG3snK07ACMTSkOH3JhAC3xBKyy1L9/cDUntBab9xAnMGm/rX3QuA3ii
WV+UzLt2ZqrE5PZR0H+xA10HkQKPbIwNUJIJtmfNOl5qXlZFDB5POKnlCimzIQWd91r9r8Y+BzrL
7SkKjPy+EPTX+HlprJigHmTXP+GvrGmfeLgbfskI7jdnBTC6FgWk9g8I0pyTLnEfAbHmnpFQlMPy
6zeTsyFNlTJS/4/yXXr5ExajDWeraSWQkM8aSdWjopSzFOtLbM+IKGi0FcQglQlth4Ejiz+HTvyt
1ULkjIvCA3IFzOQZTKo47e0IofXo3vvDUL5WgLcVziU8rv1WNi3AmBtoFF5Q0DAi32XTkWLBFobj
0kAeglithFRRYUC5zKU/GeJf7pru/AgdjCLZCPr1fX698Cl2iEncAmNBkSTGYK2yeQopWV0Cp71R
UP/6pUHiUmB4llhdFHkLbKzHvwail5IRoB5Ev1+M8+H+ZaHF/b4x+ZecuZjHfWO8PumXkoiJqqvO
uzuWYI1q8iST0yBVdWBjtAIufa9RE0PwXOGFhjKM7bbRvOSo+3aMP7edu1g45y8EL+ScoP7Fm93w
MIvCEeT5AIKF41YZi5rNSQZ1vJrchZIQkjI2PkvZZfoRrgupXdS4gohxa8ckwhwiTLjgTwtntPxu
TIIgnRwRD+HNc60PTwHK3eY4TZxV8MlypiNqX3W95hnSTFgkuByfwv0Uwbi0/N0U8sMJkVf4c7sl
wWjR2UHpipxckuc7NZU6sCStIsdWlEaf9DIXlPb+M/M5J/aLr1O+sJ4fLSl8Ggyz5F79oJtdlA8X
55MIs9J3WSerCCLQ+eYy8AqQkmIDZGMZ3S8cS6R54iVv6+QYeOUbkSc56MKGLi9GEfePZLoI5Sxn
iaQHvl61CsBp0OhJhMh5LsDi2RxRe7/NIOQg3qvfwKqUDWmPgOj28ILUHiz3IXVlQlXtFGjtB2oP
+KkrpbzOyoUZeoS6dz//MHkPxb/UNcYNrLUFVJqfiQAGXItZ0cU3ms+vAbIsrTJV0jBk6dOGYHRM
YIePXQrU730FjA7S/5yo+PzEprfbwcGz5GtLXJAyTdvaJL1+d3w+KRI8S0oZqtxuATz59oafN9zk
PMlTLbjlZkggYFivmo9x0R2d+2abyFyDUqJWb4ase16g23NpfIb0ZgBuF0XkCKSjzamEKnwFeiZf
ELTi49AVZug17Bk5gDtjhG5DmKo0mBeIgaFI01xCDcZy3iZbxK4K1Oz4mEZsA7wIzpvHpGeUkQOy
AGZInh+5SUm9X7NGnurwsYr8SYnMxXF51eBelaggH81OEhqgpKzLZb9b5qOLw8ehKeP9szHj+Iay
+YVOShOs/tX+0JIMrj9K6elRcCmU5Mlo+fK6ww6guD7RrCPUEk+rQULYOSO5A/XlMbhDipiQPora
dhnTF4qQADPh2Q0VCkkerujnizw2mwQlLMOEEAUAa/qOr4VDKkmQxnKFVhpMC4GvPNmOHI1UAgnj
G4y90UZ2Sf7NwgXN4FGwpbT5ONu5CIIS/yA24CVWbSe8NjCXJ5DY9MFPbCcO2F7rg3rKbqyGXwy+
QzoDwtAAzT1N9Sbf0puaVLWiagRqIJmCETACZci9z6UOaZ3lVrLMNJzRqXWWy0ksSD/ORtK/j+e1
kA4fy3UdUN/z8ibDG92UzVKwCzlGiTVVOSsfD4K2CHA3eK/tff7jhXY2++KBZ+e/jCw160XFPViZ
OzS1xcKydncIAq32OdEd6IajJcDLSiPoz05k1/uGelBAjG4QHCp7ZPCSqG9Ohum8V5tfz6SzrSVJ
IAYL/JiQrrVXBFipufL26yN3igVfpNYiSatoFAWTBrnGVeFgDugQkTwfxnmsXrlaqglGdscyXlsB
AgSiaW8hAjooDPhLs08UIOo3OvEZRJpIhlEDlJm6RSi1lFCQCZtYhprBMPrzp3swaC0PY8XIuIpu
+bmldjGOF4nP5hAZ2bCRO6KKcRgsEStE+LfKVFHhY+7Zq1HbIHmgoKRyD00fT/RWa2M9pSIBhuyN
Pjy9OafkmSCJvJ4YuY6D2qOw1QwMmx4//82S/ku6fwPboS1LOhHTAdZRd8hf9KcJwsfkdByJ7dmS
aCYWx94AHZTpCz2JRU+v72Ig3mw1g8jbugCGR2ILixg10kThHMz98Z7KvIaeZ9FwoR3ytGkuP+Uu
z8FLYi9x8/JJF5VPgq8rX/wnqlwbg0dZpIEPNsT87mJQTBZHF8JZWzeq3F+NY91eerMsJsc4iph3
eUfsLIdLDe36boYz/4HBhp8+4VW//B4906MTbCqgzNOpOPsDxQhGcbS4g3tFGE38BVo9B4lj+6c9
73lnD/2G2G78+VQb4oI+IKpgGTLpcLfjVxtLnSkowlbp/cj9vICXpG4FfiP0rRJAL978qW46gZxm
RsD+aCTm2OrKg4lPsBLTCYcTViLctHd13bkIWbfWViFje98yUiLMCV4Oilgc5xy/9xkDR66CYinF
6ib0LkdM8rJDEWf7npJ10eU+VgmzjVdNAdKWIxXDSQ8vPRFjrQh7BW6xbRVmNwU1+/4x98oOdBgf
Mj4g7B0mYbcVuJtR93oIYVpi5YDqkKbH+2YGtJyUGOKzRkZ0BMg/cpB1CCC3Kt0bYE4CVD413sx3
Y8LJFqaURI20F6Ojt38iatdMbnnDiq3OBHsT7KWQG6IzQLGXhyW39XmctWXULrf0GWie/KGZyB2K
lUsI4+/paAjU8MdWYymDyxWZr1PmMrNsMzp/ev7rXRPOrC5QnImDuN9OJN39v9MOnljCSh6lbeS9
xKqZHDwF1f7X1BFW5CqNVyUXI/qfaFmpsv669QTerZ65yZ8FyguF9t23jHQpkQUsItWyvvpF90Ck
iJG832/99rHmpdvuEG4D2BloU2Pzf5vsbX4IUMBfRb6xPrujYJc65w4bOWkQXG8D9LDZFVECmaaE
FuB/IwG3iCN4N6MZrD5bGws3/TMkIYChukX9sWEDRzF2QqQgpXRhHNLCgwHkSsgndcctScGZckHf
5tBiNpJzhyHjL6g104KE8rk3UR4JHBCuVa0tybln96Y0ROhQ6waBbU8/eRKZvTj5pETiX0D/ENdi
TeJsfGBzsBN67wOUAIwY1GRKp6o0xPgEGCRSdsryVf40alL59fBqO04m8oFlz3qhFQLYN1ByPFlB
VSk7aqrG+MoMtnHWTNYF5yikcis5g+3Ctbgo4DFprgburmZyFwzUz/syp8TwbYEoZFPdnKjuvO7y
qzsI3AwHPvkDsTKT7maqyRN0hr/Ux6z9iBE5QamMGSHfZFcEymBmgxB1JA/OS/ec2XePQAwUV4pP
Aj0IzQeFoBbt6QDIGV6c1J7L3XsrodG20OxaDTEP9IZUcbHpY+RwFRZMO/Z8qBvtaDtsp1ycvEbE
29ZrAM/p5GeyOxZuIJXc513IEnm7G9VjluzjmfxedSdTln07bz+JfXKvb7KeIC+2c228ufS83KlN
/CBPYsT1hTsZmsxfCUhml8h0PsdphnFzSrD/e1yxTXQJBGDC7KMM0Vja/6RYJQfolzeuu+rcl4Lx
qcV7LQ4DRpCu9FKtAiEgXJGRJF4Ug8PhIS8yhepVxBnxsHAHgg5bmwEhO7DZ9edyJTSDXLnh++lb
Tnaj2PRURqVR9srEUfz6c0MrHczsj7pdhYaRCielUAk01BnxYz8gua3WqtYfQHeJ1fn9yE7hOLTm
nLmMEFuKx9W0Lgo+jkU1f7cl2IkdHIXpu926VRLt78Xc0IKE8eK9oi7Cq2pWv4n34xQ1vC83XR0O
Sl0rLjxDAt+nCpFtIk0CzYxAQt9xrQR3UN7H3wyExHSvUw7Lr3FOU3GL7XLiJYF94rFz+VEapz2+
KJeCvm0B9lOtvHgITjHja7MrqihffkIbzucgzel0DVAIpeHt9Umpq+z68E9xPXzx6twsoVB8bIaH
WSUnNXJeU+5gDsvlsqvHclUOc99f5vMkHanOA3VGH7ULGj/RIpoB+vzygX4fJSMkAB+3qAj0OohB
6G195eBMQDQD9xo9W5BKhr3yPTBKF28Bdl8H/8BUQ1gfTFPY4FQqaxbOdVvduzML92cScoh5CoGR
wrQNxnBkLA6t/AhqKPu3FR0f1WUBl+9xE6LAzOrj+tFJt0ids0B3SWAS8fH4+DKvOn6oMMArxzLs
5cOfMkh7McC9VMSVOwq80+RPGVGkVlzXoLH93k5Im4Ehi4XVwqGCKk32WKzXq/b7kDJr8u3G2AT/
jCu0QwNfR/ZCHjEqtVKk4I8RqSkqBBT2XJJz1tXvtlEmYmiJOD8ZVT/FLfZioq8E6BqgEya8IotU
hhGC1+7iQo5fa05Otwcs/ZWybpe3c4m2mybP2vDK1zGAy72g8AkjvlTPmpkJdeUl+ZbkIJQm0FD5
YC6hoA0MrB64h/TiTBTnLnbWPFohsyUYCuH5oJWHqq1eosEoOfdeKBq6DHoGtd4MkG0vYojV1liD
BI9fqI1ee9TcHjgV89/PJoaI7oZQekyAK4h+lF8yg3O2VWv9pTiZmpax/WKW7FRbqdHdxgt/r3B3
BD2P9Hm6mObHS6boz6ub/Bb8GMJZKIDuarNDS4BeLFyffuyAVdxhZWcY3WHIG1dA+R/3a4EfiUQH
n7OR50mo72XCp0OONt4InayySkN13gcR97fO5PJAWXguOR9EuQ3ZOAa2T23xSv+Tiu539yAMjxXn
Hw2tKWOWbP5ZbT5BtEYxiYjNzochll746HKcECPPUKAZmlk1N4CeENQsyvP/VjsCXDpQGA6stllv
8Z3yIDWitJDhugoWbR+OwRb7t8Kux/zpWq4qsWdR8JJu5eMeWj7bebi2/bfh8UB3Ts/X+cAsDU58
BUuCRGcnQmPL4LUJ72ywgF42bQfgI8oGuQcRyec90qnEzk7f6lmJaEHVUxpAWLtgqfi6oGg6Q4yn
m455BXacsnHkZfhQNaluTbszQcbV8ctp9M/Pas9PZtYDtDgXTGo7+hqVgPopvAGu9Usu72pNVh7Y
lwALqwq3QQBIaPXegSSNMC8gefBiYFnLURW/wRL9H4e+9CVJwscrI1p3RRibQzLQqElFhn8NWSlE
L0vwh3iv0K9dAb/ndcc7fmmV7mPn3iZ+vJ5TZEvnYI7bFEC6jVo+RdOwCVB75Y1xEEDnxsB3OoYo
NLpIFOR3PCJ1Epn9qyXr3mL7w3jvCCSTJkXyMfjudRtdZPlbN+XfIPoKa7PcXlbkfUsxOQirR1Ea
YCWOYqWr/RCwwQRuaifOtLaoioHKejYDGFhohQTdMc/unRNoUiBs+T26Ge9oNCgJO4n0ooyQfnv/
7lCkqto2Fo34OY8hjvXJM+m8/aqQPYc5VzdllYq1IIKTrgvA0fPCLvEmntCq3l/V5WHuxxwcBZU4
TctA+8uD8V7QbIMMDzpduu+jJ35nb8scRGRp19mjj8FZ/ujXpjSLKjUWx0ngiD/AfDzZnJhFCiGY
bjKd7fOI83gxPdw2jx1af9I0P7q5k7DYGOwOevY2nk8arj65pzcismi52GolgcCc2AgOFQkX5GOU
RJu71zqdlC8Tb3FM3JGEm2P8dJwCW8qhhBVcMlbJ8Xt8kvZqVeKj8SQG4PURehvJPrGodTXpwMw7
ioMyKk7d15OL0mzMUa6M15/RZ3YMgSnu3imCZcf2sJleJKvICf/zRBMGcXiKl/kqbdGxJfqJ+KRQ
4rTDU8eyCeG9240ccJ61IBofxNwIXixY1KdcbOP54IXTb/gyN+H8R8FBtyKh8zAq/IaDlQ6sW2nd
b2jLT46GvbUIgAhErStIhG4Y3uf7ve4Pn7tJu6oV/38idM7tgZjVK7E+swUp+3iXbUshvKGgES2R
HO7h+sn77QJvbeOek8L5Z/OHjXycuNRSnxg3Zqh+Nd+UzqNKRTv8yFE4b0eWm3bdoYtKTfgVkS8G
zTlHMMecJOv8zV7Od7jKKwILiHuvtyt7XXtVoTUFGEYkJObG5vVOoXdNuZ5GXooNy7JNkwZnxM18
QpsKVqGPslfItokAo1MQWX4NNQHB/UMa7Qo/IVnObZDplt+xSscZumgsjOH662dVLVPs3RGW4BEu
wuHPn0zT91FyrXBMSWE/g6Yi+HqrbqGqKDw7BBXmXRiE3wgODxyN8La8fkQTGZiOUy2A4u5rhGjS
wiIhqbrzrWLmZAVBVXIT++LNZXY49HfwsPIwVqYC/Cp5tdQs7PqqDPiAKeJ9/KyqREPnB8Bycv0e
FIsfbwhtMJpHoMAAKe+lY4tTcOQgRfYDSIDQNyia+0VjMHc7hsshTMy5cEtp12JRxpCvx1oBtrsp
H5AAgujabXGq4TrF96ItLf3yceO7rXxSTYl1GiVX2i2MKoAglpd4pfy/eQJjG7FeRx+/YEhbWgkQ
/KSvi+wZSLroP2AOzCO9GKpKcVg6wUqi7NT6/l8mplWYdhZOzH+BP/PKNvduEXHWKM3PH0ztxALU
JpoTisy94oSp42F7JrIJZKC0qAKbIFjuBpqXu91oh/PJ06kv6cAt/JBVcF3Zv3O50U/+bgyXh4/7
gT9qU2Q/0pJRLvnMoPB8Y4vTmTGILtApI90Gt+YuWq0D0+pynJmByQNHHyGtnYwYhMOCGkh0r9b1
J2KsNxSN+M0Qr3BY/mCZIeZKpeeSYI1L0ONGfvng/3I7BQ5uwDDywjQdBQvJb+0UPLvrxvsh4EVe
oVGdi5OMQxZCFkcln3p1Bcq6hjflX0D+OxyFuBS0yKjMFPW7gDHgItefRwlG4Y+RM2oMGwFt5yHf
QNafideFCG41gl5PfRDwV9ARA0VfYxoEQvqOByKoIezq2A1e4UFnQPwQbIcLhoGaqKIFUAigVOsN
Mvr8p7G9ygmWnNcvpTp7AokbVUS+sEcIEiIpMsxL4tnpspBGn9ifuBVFgJyMbbT1qOxADBt6U7kf
sxnno1qGVrsBBb+vg6E/r4XPeiCDzh7BsT7M7Q0QuC4wAJY3HUaYo3Zegglk8fEHq2E91h7j+pP1
/EOyR6bzdAVkCJz49VEYiz5WEi+f9ru1f7yQe08qth1f9NCq2aV8mdzlEzo8kXGT3ZZbEcjjpxid
9cZfZeHgfdQUuwaafhGrytparrSZTsvECjXlTsZzBLScUH9M95UyfH0kTLZiuxXF9KGG+2UYnJ6K
zTjd2wcdUXGXjCUla8OM/QPMbZTbgJ2RXrOeI7oSKprufLdO2hH6Vj5SxtyCzzLtr2m3Rx36H1tZ
IQaDuwY7UC+6vruX/d0/hm5priz4zj97j4JHgMJVQD++NOB+JgKovrW6pRTOO+zv4KkWlDP2X9Vd
luncmE19BFp5hTTHBdDfLeI4EQCa8yGB/lcsfMXmLaXvFFV1xJANfqn87EYu0Ll5T90zGnQi4rqa
urQkaMEVrUjgmAi218zXkp5GG5u+68ncD5U0NUMsT05V4mmlTQjZ5MH81CuvzCaSaelRhZzaWmla
JqZ4Y8qDK8sASZ5Xgjif+JLDM7Z1bhRHtJBlqYzSBPEflmyffcBNclZyckycXv6qroWgnfQssAZT
jCsT+R74eyOtMebzazmuLW/7OGA8qP1f5ifjQqUCYo0crDXXmHdhHGGFGmCOMGL//37w5c52KU9W
8HJU6ZgkVFB9ZQqf/fFLx6zR6yI79+ytTaMpLxqQUIbcfrMCqFGxbTL+CL/WObJJO1l5v/ZUUgUU
FvRTNXQEN0rQG2OFaL1acutSwNh9kKjAmzzoxFxsxBUtSTZkLLcv1CRo9bHdJ31/AAgvhMRtcAcT
9elE4A4WMkxyjY6fZ4YrEP7TbzvvyVGphzgN4h8Q4F6NTp133xrP+UU07/1a1MS7m0i2PqCey6/o
8j5oP4KcMQdSzlfsvQlplBeOg3MRol8xg6Bry87yiH9kNQsljawxMYDVdUZ0yqHWSDqgDSpABTFu
fFH04SWfY18uvstYyCPDTVpWhxJaobxi5FUoeX1ywAKWbrJ3NvbjQXpCRATmDtNaEI4vW5qOToCJ
S9naGadbpVpoCGNwOw7I+QXymeDuBig0k/TP7QCrunV6RypcyyKaS8o+k126+JFSKQNr35IDBytK
TpsisjAQBIUL4j1nbJIUw9Beg8xSmLKtg6AetlYNpAeF1+gYVRMcw5yNQIUuS0PX0koM7+9mxx8C
krnKMSNTt5Kgx4hh9JqkBKatu6DlAcCnO7AUx1xy++sbh2uyVG1/imIps570v5K1hQ96xFHM5LwN
XPwMDJgtz2s3Cbn3S1MOhzR7P0fXf90Kk0xy7dr9FRRYwT9Psw3WshTga5w7c/U5lUohjIXxf94n
FEFLdTL/pfe12HErdTWXnWvDdLgSop8QB2tQCJF1LAmeFz77as1793KBPQkzeMB7K8wslfgYqdyv
plDECdFjy5+NLssASowqkrajAkORWxOQWa0UpOMQWkKS/ZaMUa1lhXZjE5EpBUs33CmjpHWcLwB1
i+IMk8DuHvZOdZZ+jgSPXi0blhjEr2blJXX3DpiHZa0MtzCuJrww5hhYrnlVTpBhPLxh2Q0+esN8
dPde67iuj3vtIdVeaiKOMCZ7Hfb/ROoxsgElr+y72GFwYllLMvAwPVZi9GpRXng7RDQqyVAeoyp1
O4G0YmZWcfPOUiRa6sWeC+vZHGwX6KWy8mOYghnLnm5NcFoSI2MBmVrzktb/jFrqaOxhhd0oBFzA
H4O5nxTUg2IpaGY0qAf377isqc0abiYtcJh2xhxes4muqjDuS6GkGBVPW2On40mP5Tg61PQxHJpO
8e37U3d5PkfsKe3R41sFxUjcEOJhiciwSe4170jt/tCIYYbsoe2OOn3my1zPN5bJtTFlJxx/LZAV
nr4Wju76/n69/0ommmGUt+mdeRKUWrE7lsZYEhXZ+9EQM5iSdwtFRWG1H/4D/dvdCp/TFR3lE6UC
VMaYjHpyu5VGngl2KFkOV6XhoFDOaQEuCh2ZU2MLHEVC0nAtLGwAYOfGRk7zdeYwqmAoqhc9OcgD
VkoPgeICM2B/2AkJOTLGZVIRFcZqyDO+P0tOvWHBedqXAgxCCZUnE4YZ5NsHTARzLktuNsY6EFGN
ijzuCaIxl95brgsJZ1JWJY78YE0d8KAcExNzOheRU3GDaE/dM6eZrW3fkvH/KNDYu+N0BpIxZ+mP
HHwr3tKj2oVWqHpcjqsAgvhDxzdK/4NRq4HKtmV5PBa1voKJEovaKliOgQTschL9Qbk7DIdItuRw
juiRnZE0rAqKd8H/bCUNxQxXTa8B8Lr8RIbMJEqEFiuqGYdokVZa6vp0sxFSkey6pyoEYkrr9ulm
+wXrkLBVjnv1t+PHilVo0Rwy1DYDt8CkFw9nxVI+6/OB7ZwruSiS8dChLgcGtEKlUMJSmnLrjte7
q0FFO9cws6avwrltOh+mayX237SamZJgOGzU8DvGUnSeoSDS0TfvCxDBTij1KSnX8Af0Gyj2UZgf
UdPc7NiGtgzLVgNkjvxkxY5iD5S+jCQdTxS5l7kQgXehqQDlLXCIhhY8db4b30raSs9o2WnjJeIh
3ZtNnOj3fZbSrDGx2kKzmIPBBzHQhfRIUlPwpUBCed6ZTfFTwE4hHI3S1VE+6thvG3LgOitSPFDI
1dXXZh04syXVln+3Cmp5IO1w2x60RMZ1/4T+fjRZobPeS9yY+SR7B7si0tpGH0oRMe4on3xIwEKg
ttuEwhMNCMyA9eN0TWT9//7K/ktRZ9Q9tpUCfPWAa1ENsooWeTlc1KitEqHYBa1W1y7nndEgvmOs
8rhIVAjEMy9WxrYhCS5YNcz4BTbcaz4tW/m7FOdDE+DWu3PLHFzim2m+b1ZK0wAnfYyGumO9dNGe
Q1NDMLCKGFPw2bKu6i0b3q4wefpmRC72UN8qRt+1MJFFodTfd9OabY3DOqN4AxwLOHN6eEhyKbRW
Do2AW9jhI/wfmtySK4XhGAkzv8vaw7i+aH3wdZQU2My18sgYCJx3umIVmhn1UavxsehZNijHQdjA
Ra40AXJfjuFje3sykJ26B6Qj2ESWlX2YRTLTiQ9DwaDYNhtQ23RiFk5OlnZe81nDYoZR5/qXL4/K
LzwlZ2IMRNNfuav/adT7Fu5oRRSjEK3dlRvqUY/7qNMKA45u7SuCnmbDpG2C+5q1k1boJkNxBXhb
OLbKGoa6ahhInkV5fCTjrKSqSgfR2XmSHziXVKXArsEN9TmRsIB5AigFu1Nr3g48Kj0DkXFuJCEI
wDPIo0RiuWE9Aa20CkUfvQz0cW5pqpUl0VDTXUhVzVs9Zz2Qkds4gdYqgZUTaBnVxXaR2Kx30RlB
ywFY4zXL6k8ZiPtdBY2eckn1gfx0qz0n4gGZwWUk5iFh+JvzSDpE6Y9hY6Yl7c1g2k+pc5JEEBCA
1SOwpjOiPDoyJs1ivWniQzPbY0TmyrTjxLMEdY4NObV9ewcF2TL1nNPzKuNfNDEmSivfiv7AxX1e
ZkEIFc4lUdhmy1I8wi7Snwk8biyhQpCR6o9VY/aM7hs03iegqhYapaFembE02GBzlP2rdIKs9ak+
seifrFjS7cUiydwoOI5g/Cwkwc7o6ZbRzcds/AWaWV6ZKUayngXhVd3gJw5NTCD6bRq/fdcgdcLz
S/X/Ug2aA6x0J6K+D07Sq2ajys7+Wrxej2y87cJZCos3os9qnC73CQanKcVp9eXW7x7iWgx6mWnb
Y/Ec/mutLyPl0mUMION+D14luW1j3V56UypNrUHRc/ZbuPbOHfupjnnn1CFxrEv/r5luWCnxBUlZ
eQPHeDk0Hd6Xoj5h7BahY4MHPbXXESZBnDyutcoc6Jivixp8QyMh3gauGaV5biguHtxjHLQigx2s
Goi1Og88AC5gg5zqWRvl2LE94VN33VXAFL8L3550vgipn4WbnBCSPc1QyiyEd8ydOfO1jq5pRoPl
k6EtHgSKHvk7cCc3LyfnpNvDHAhT9YTdsSZE67FII18xVKTEvEE+ZO7GHRJ6i3x/iuQTH/T4LJcL
HGg45iuwoIhJ9HIT/FajMgoR8hJnbMVEsBhI3SoN2LWaZ0FMDjMYj+NZAu14FFQXG6UDavegzzoa
nEffZleUju7s1M5hwu3xdrUdkVrfLvQmDVjyghYBO5oi3EYphvOS6K/UtaVTswN0f5Y7Ke45Yk4H
yRzcSpc1KzS+zAdAIdj8xE9n7SF8e518zvVBB6mIbVHJWxYMz000hvLjM7YUCbxyssAuQNp9DXkT
kd/DV4HVgzPI5nSOE8EXLsUsxrfLHdHBJr71xWiOggcPhR6kHKg67saMbn6hZzzxOMpy8fZYe7Yk
XwE+oO824iczFUvCSr64ccd+1KkxfUY+Wr07I32HE1jiVViHQXIO3wjKvcrcPYJyDoEXXIUaFgdc
YrKBDw96SKsa2CrHia827sfMDmV3dllRyeUBNQpdkSd4xaxwZsS+BheXQSX+orBLSp9PaXLGV3oU
VA/B1YkN9TwjjC8MaMJoUtRVA2N0T2F5ZTrsgwZqiKAhJJsr2ATG6ZVHAkUPHXNHlT1OcSLHah6u
a/XA5Iuc5GcqnX3tCI10k7Ilhoa4IaIPpsz6ba9lbTapc+Zk7/Yj6igwWiE9NgQzWNs3tBQUMvAi
bu9TdmFI5bYvQeTOyVt/58RXK5tIeIaepU38ES7E51mNUeeWuZDBXZOjJvWWCc0cLdcASC+mi3Qv
30r7Rn9H/FBKYmNrf2mm40Sm5C8dxaSeO5OJ6fury2/Bvq4YydJ552AAVSYwTPvXZD9RQ8Sj94z/
2oEQe55GHUMwYV0dGVxD66WUHTq+Yal6znDqz9KehQvVuggYhuDwqfoLcszhOtoNaiUqMXiv8yYt
w3OCogZNrBksVQot0091Rrsf6BwOswkGi8PsNJACHS1sOinUamXmdzIYHiD0rTKxXvq+IVtvngDs
gnF5ZHCCvMnp1RlPzoLOtsE6J+iS/br3vAOnIOgmmJsqK7OnVHtoORg9cOH8fBYPq9PcBJiEFxRO
apJFkOcGltKqZQrqcMfFSsJirBMdMYHy7yp2vj518Q5e9elifFqp3IlSRoHW2uNuD/7qga7sRlib
722B3D/lf+AB9QNZJQgClWhhYdQ2EgosvrReK69X0YtxSm9dN71zoMpg2bIBqZZYf6v06HXhA8Y9
m0DA4Cp0rLSkIwKAALGhgeNuGu14pu5wpLUksIEpWXgyi+3YHGwBz2GnxlZVPUue9tO+Axd4vqfv
8TEeK+v1AM/5KZVtkp9LmoAnwhxOVaH+dEm0VRFeta+HbmFMu9Xp6pbwxXWzTmwLV/7YxRzCFr/a
o3x2BecIeRpEjdOx9kHzf05cNvIc9NltJxpkuAFQzbbxffQYSNIrA6uSdKYii/VCGzS4xwb01R/R
Gg3E2nhunZ9zKYPbSgD5nMa2iAILFeBs4+iCY0q1V9jCGZc5GNicQ8f8mYJny9oDGfo+6zR6juOf
KYk9IbEY9OwlHgTXShC1jwoZInSv0yWgFRQNypr68MTntiNbAb08xDC1y711DDusAFQIh3FNQBpz
AXOl8Lka9Lhko67DR9p0tvtpFzY0JXO2vncuYtTktHm4HnG7iGtGP77xAs8SiRKWr+dieBBM7ei5
ZKsZyxCgSSDQcSSkADm0S6jXM1RAWEcQFlIZanDUt4SvY2lkSGM+WVUP+gauOos3Cik5ytNtal5v
mbeW3jADeRe7+USYoo7DU1Wz4uWW4v7vJxQvRxFYluGdDUA836SOX8szL/15pjg3nH+AT1YOT0t6
UrCLbPHfZHyUUBvodstfNWpX3sWTkJZUWk6Cu+g6TAd9aW61FXNfppPVxbVQGsMGgSEfNQlc8IoR
Nk5uZUtJcJpCpePWPF+PPTsFLwzJqtOqGh2aHRWAXJJ7JzrxxqH+gPEqI7qogYRRldHcGwCZcRVf
LTkXUOsObgG+l/QK8o+lfeAr7Sp3ekVXRMXdiXkf39qCxzI7bSlPAEEpFdBMngZs4agEypw/HW7P
g5AZ9fqvCbQOMhCubrBWse4KrvSAoRpZlX0mDwDSPgfESGnekJ+vswACsAfxJdjVbH+Jis/eJ9Tu
XKkdHajhOjktQcfrx4AJLup4Zu3dohBM+EvuVY4sqcttWiExiT22hXMtd9UvzO6mcWoOFnmADqYF
rv4+s/pvgXoRN4kWoq/uXuqcKAV7HnOHxfDuPhFux39u7AokdKQPYYOhiUWsF9ULK65aVihQwEq6
K7wx3DAoX/hpYV3iYjBwvib2oYrnxSqV25eQqPf6sPx0DlSjLU7sxzNTKe5n7DM6gh6HTVmvN3XA
EVyYrhSwgG4MyGTlL/kcFLpapCEgoBI0NBqOq+5hYApuyifKO3Ck5dxKFNtwv7bqR/euqvOrgCJn
vYUYKLLh4edSyUxBy+5ew8RIXNk7JbiG2Ysp/JDtR//1j7QBCNXqk0PpKs1h0+8y/FOIu/tgGT98
60NeLMEMm01CHzfUIBH8Pp1O8vTWsiLdzL8VpNgcjamCCTt9Xn+IYWb+rHsNT64sL2uYMOVsjPQy
o2dYIuXzQ5jeCMG2XO/NA6NpRxcA1MhoeosVMHjKIG1OeFwRgKFq/lGnDTNPN0BwuAJ2OHCo8rU9
oER3usL/cyC4cQ7y/KpzpKD88In7/917GCswD/XHnMWQuyEg8LILQhNx30+gFNRNwVu7xmMWmrHF
owVKFOb+GttsGYnWp5axAPl//v3N6gDBuQOznlCIw1d70R3ziFDECJCmjn7AzvugcwqwpE7FdCwE
9QTRjcljMFWwf4+8BDv1zHJALGrFzGIoySeSrwW3W44aEHkM7eLuFrNHpn3tGPG5sW1w/RodCSrC
sBlM7Mg4gkKxShvymIVgZNQiEkCXFTNPwfo9/LyJ0JMxXfQy8NL+tR9j2ms6rmI2vo1zM6kzMt83
l4WXxA8/F/5nEqZ/RWIt4yKhSNH2/vG5/jZOPTqHgR66XExcLsXDbY4GZ9LLEhteU/45k3SShgei
ML8Ve9MxrAmze34mnqaMRN96aCiBklSrs7ojr2DH/weZIUW5J4hsLCXFYqRJyzy57Bqtsev8FCTH
Jj6auL5cUWL9gcs48U+//BPBaalF1oj919atvc34UN1anoETf4ofmBFfqV3orE9OuJs5V3LL5tb5
3RUWxVp1wsFlEFSWJABVp1YD4eUKkw6/6VEuxsuadt0FLYPTyuN+IS8PTcTcCOZ7uXtokI8rvqj5
NDWEu4vYeNycrbArRVR0Ru696x7zrazNJ18weURlS3BsAIJO7DQAnb0s3V2jPB2Yga4wUQv6tGXl
VqMaDIhXlTaxicnkdYb4eA/GuatwkO06+iqjXH8Xv1B6uxyKX3Ur6IURVJFogERzrrF3al10b1f2
27kMEtiOho5xnJx3dI6m7MCZqAS27hKqHwjGBOa9HNaFK8IV6Wd8diIcFT0Wz0wHcz3mrJ7nuQWD
q5Tl4hPv1ON7uVD5sqr2VdF9e/aYZEA5YtRqhcekUJmiSkB6sj7SkNwii/CPZClVyxG7ANioKSws
6oxxUbnGrX/qh9nGFqhiFWWRVmJ0S4YFFG9ryPNQQQSfMmu6t88NFcZqvh33Q1hc+iMbwHaYp/s8
3F7cb1n0oz00BJJal143WKq3stQIUJx/ZKWGZOGmBlJXWK2QHsifE45fAtYBMwoeRuJauC+XWeUZ
d5Hh6oAd4sb47Ajtm5VHi2vW+FGFLPO+zEpms76mkm6UdX3umfkvl9LKaIPyOOZXK9+URyoKplgA
64+fRLabnCvPA5tdc1YXo+mPVtOQ9m2KZmR3JcMIUuQu067m3Zjmesf/3LLolQRHS18msZ+X4U4G
IdoYjJhfJC3I4A1CMpCNMPPSjGHLcKXXDvNK+pRcZRO1IVKm6XaeSehpukecOU+oWEgnUAPPPN8Y
SKPie2KFf5k9MUZte+PJ16jXZObMqwPZNBdBzYhMBPghMVgM74btja6FRlEP/iUPQiJ0i3SUDN9a
BihT6mg3Q25tpcXWTyAbZVtdIE0ESVPgNHBmHO4pPjBvXHbZ3L5+3Np7gTEhdHnMx7lDTPXMhZL3
VhBtePJfsZsGScBFxxXkqaMWuLTTgSUvrdewRL1PbPJySCrwMedZtVfZnhgkxbo9tB0l1t27hwNz
oLnp4Fj2LC9fOTwKNJ6iJJERHOAMwgM/Y3GaJR/QPhn/5kcdNwVgwPRUdwN3GRg4ISxkDLtLeRnZ
wL5gujdgkrvLaFUcWOOlVPMuqGWMk16zKGWpDzSHa7UJY9dafvcRcXU6SprHnSAZgyGKfK189DJQ
Q1VvVkW9Vl4lZ8a0PfQsocihA1no/LqXm3cxwOOOhq5O+e39dNqttLQWtFlw2MgT8naXQw0jfmr+
Tdi7pZYdKrYag0uOkY6r8Bo+7qy3rgafmoso1Ib6DUUobzj6p8NkPOyj+judyYRTmNufpe0+bk0Q
khXWR2k3a8UNvtdpvM1MZaq3ujYDABwSiOlctZhxJTE2slPnKSohc2UzrKpiSRvLE/aylbbnTEch
NncGfL7vnuCsUU5Pw2rhGqW8BIcTZTce1v2R2ans7RbUm+pS6s5fo0RiXkUD8cXRTZEfx7Pj0K7f
sRd1h8AyD+o/D2wx9hgeBAlX7qIX5CgATCSejNwj/2Jl1kGR81Nz/cihJvacQkiPbHfKOexJo+L5
MneUqZ43r09/g+fpbvBNUKnJkNfir83v/F/TA7tmbEvWoNagHDn3ZWq1OP+Pa+58CPWckiZqWStE
gun1u4twNLAQcDOPmRzt/bMQr6izJ9xeSU1j4gCPDZ5FyyBZTezFoHsdLRnEMWV0Wpk29Qxs2rmk
zcGJZNdjjAyT6P8w3G4pRFqJRr4za/kFKp/7YfrXEJyCGotbwl+N2GRUW3cGxM+E0UirJ0sX5AkR
CITCUaueAJ1hjbVU+TZEAHWIJ6u2Yu+eWIbZ5vmfkfSZFIr6Aec97ngaylnoWMXj/oG0dzupvRTQ
3PwubYFRzL+SygvGF4wzv8N+kNufnLpK/1azcE30dFwbc10WzDPYkHZgOXwC6os1x2loN3gw6ePZ
02cpfVyLwxcp5y9vpYj16r5fqVhMsDj42MVcdZoDOxUb3Vj/Zpo6uEbxA3cqorF6cYaHlNqbSTwi
Wd5kPZ9HR7/2yddEp8pOvJlTP1tKABrCmXtijrzg8sBjNjFAEC1IJfH4SCY1NkE5HbGpiqG85C/6
ExW6aRj2Kuhtsk5iAyoclPRTjhl1HJC7f0RvIV3VH91RR7gOaKyXD2RHiin6nEhQH0fdVB02efKM
wUFhiUWGOa51u0yk4/p9cCmDw1hE//PTa1QcRIbkTF6oYVuduc5M+J68f1x3zebe6kziy3+C/GUT
Qzvo74WJz00G1HMRC4raQgY0UK+gVlDRYQsnTfCih3BDLks5PWDWj1BWFO6t9vGK6I54ytQUVD28
MyjJgPt2hnKq0YKGX1DVoq+fLmsmDKTGnaaWrwJDEim9bq8JRCqR9SaYR3CvQT13KPCVAEbX3XEg
D098aEgYQiVRXRnV4AnE9du3vgKedATx9Xt9DYXOeh2ajgqtU+7DvSliIEaY4NHB78ERWhYxEMPy
9oBgf+t4OpHdrIU73eEs9WHmO76puBMMK9fHfPw4DZwTk4vK0CoRKB+R87/irvRKS6Szg2ViKyer
rkZSv6x7h6P3Gt88IWwylaXGwMqJljVQQmlqi2vNXVPbU+8AMshmpmbQpyFzjSAuD0NnlsepR3rY
ddzj0nfR9nSHSxz6Y0xpE/LQId7UO13vKkiw3ID5wkkRN3oQ1usamL/CZKDAZg0QKFi42U5Su6ac
E+EEevQY8QD9tau6lrLJuj+5FqeSsbJlpwVYklm+w9C73sTSZvN7RVawTtIgWKwyc6tzIpkGFMYs
EbaabiSGVmIxlRpKd1ZaE/suFPfbWyqU7uOHvv3TGY1uZ97gknPz8P6CGAdsSS/WH2wJCyzy2GaU
LDCPgmUYm9EnFtDcOOF3Sw2cpo4dwNVSOs/qfwcuWIRb5gSLZ1DIovEOwJAI0nl7P20NFbZ2H40b
ojk/swX7LUHPrPsucV7+LELqIvaUoc+l3Epk/x7e/LVWgD4K6b/dQnJGe/gICIQBtVBjWta2IkQp
sUjYvtqVfHJjeOw6iwdnuTrSC+HR/oI9iHuFgpQNJdbXJyBuwUDV+xuB6wpau6GYXY9MwqjeromD
17sWw1aRiCQL9/uBOwi9yYjza5o23c2pmlbtQYWD4dpVoNWvKlNRD9VBSMAUiTqa7RKq0+MwncS5
PBtPyTCA3nh3QVnY9zqYx7M2LyZM5HepacGAWCP4rZ+fnBITmwxxh3gy3ciEBMNmIpu48Mcys7jf
9g8DBKzg7B0d9Ih5aQu5m57PPPrF544DaydbLju+3GrWp5NMkNs0+rwJ3PtbMWrwtJ4hNoRyQokI
VHX2bnLHJhMJMDkjXjVGeF7bo0/i0zMvJwXUzOvCEvQTskgElso3bWI3vi3aLyUtjGcJIb21KY/P
Darzda50Vpk+39TbweEul6SrFpRHsyzTbZKSQhPMwaAdUe2T572z691rQHJCEppjGTMAcIrzJ/nG
M8Re+wLhlmVUQZTrJwKNdN6jqRyQ2iBE1/piDDJ7T88MlRy4FnP/Bg4m3c66tIIahqwDROg2DCik
F5mDs6wVtDJP/olJF6K7p1vVBKG5Ykb+tp42CXtoSp6P6taxrsUOm32EaKw8gAcIllKOhKBm6eHC
wW5+zBrONjrSkpaF0cnUV8hM0uIIrrxIscBhYj5FIl7y4l+tSVYPAnE6P4/vVzt86PDY3dEOxS0y
O83ImNJVNHiFjeQVsc3R/Kwz2T/ofpwCCtgQX3Y9f5e+8cRXPH1X8zJOJYGZ7SiT17+2KuQAgqTm
uIIs361wa4tEpvHrE4oSq8hBkkMWXLBqo4wAqnBRh6PwKlMVlmR5i8Jq01vV4fuN0O6W1biRrlLd
Wvva58/U0/RbZ3wZu/p9YzAmsYKHc0yNpw9zpux97NOPdAUJIN8U1yE5XcA4G2JhnY83hUIafVZ1
TGKBUsEc61AejfvSa3EAe9VBT8ZAnMECdvE/UYwTF38WfMb7oksKBSiqQWXVlDHWR4kW0uUBYsh2
c1LGcjJeWE7v+To4xOTsXOJQdpBwRGDA17SZpZJRxA0k9y4OQBUYmUlDJP4GMRTyi827OqNvlrjz
vni6HvZfCYRJJpXKUj/Y9k0jwLKbpVbpK4NRmN5+9bYi82Q98C0kwSXRjNoqlKkJ/dWSuk9qmIPW
fiUaqiseLRn/RjUTSicDpbN3geC45cfKF1sweKnxxBgthRLjLOxL8ZQLxjupQSA2r2v7h+gj6nzj
XzsS7Yppo3rzuy6Tjjnkq+OPy4756JxdTyvF/mCuj3OZbfnMzSYa4uyfiXgl3elgkG80iQ3bZXQ9
WQlI0L7+nu2hfEwhr5ayO61JS6MUujHBP64B8wuEgrjNasGU0SllC/gdgOG5LvUifSDEL+DgOXbu
2oFhTxQEkYzC5xkSL0Z9UlSshDsZ0cz8pTHSyAN83Whty8BWoBhE81ZI0r4SOM5A0JoE8gFKHuKV
AbiVGkEC8y2MGBbdJk+KBez5kgvgfM/6rMXsw3qw4BGBZqo/nn2eOA4KKG1pK08tmBW+KF0GS3eZ
Rn983nDsi6FHirXyj/zh03GV78jCpFJsZ2jYIEBX7b7O0s2noeZ79jjZmnO7YGCtMOzEYTv2V3ks
xYVPEJJ9IdJA168CBISgMGsWH1B+R52DP/yPG0p8uduFYEmUP61jDMiKQbP3oRjn/uNDEordfl7B
oNfBMz+FQj8anFifwM6bTAkE4WHjObO2r1nlZ8p7cKoWCzdEGSOLQF+3WhP/BlbFslKe78QQmrCW
ET9qvZh+k/pXi3zb4JmDO3kIl7gCpKxWmBpnirVpOoKIixRSXyL4sbXCg/TJ6fzwjHHI0N5/71th
LKhIdSIsAQFHo392JCrGj/y9Yv9hzfSFMbNlBbtR+z2ii/SeDLybQKTps+U2cwNFQBMrOjE5u0ft
JFj5wF2Tpz/Y3l2XMsfhTDtXhc08p4ifbNQpBmB/utpd6t01s4NgTWK3a6bwaVtb7hIJeO7rO7Qq
lqymsC2ANmhQ//9/Vmn2Q2iLBL66MaBNyw/OYUwJ1twsBzgEuTqG7VNr2ZDgfJCsvwloSkmAnfiC
2lBXRAilIdR5X6TXZx3fO2YQSlBDBqe08evp2rJqPysOnpZFIHjCvV/vubr5cfTvHMdXUUG7p9DO
BCVLOSaDYgSb/PF8pfTVqKcw0OUbCkLoFd3Ur+ZeQ42xAA/x7RnqNrc1CKT+sGBeaUoto5xiZh6D
pQsovFWQDz8n7L+xWtCMBeMBvOa6dFnORF9WkRJFwvxBzwi0psI6+z3LRBS56zQTYzUEPLZ/jjsw
NwStxV8Jcgfi/slIuF/OhDFgAqVTLF7hfjGfalJ+q3zKLLBgoZNSw2kuvRw2gFsgQZBEq6lxlQ9L
7EbZ4mrENMkH35jpBWxAR7xKXR+WEzL1d6kSdfuOCLvJevZTG/UGokJPRVbMO7qu7xrgdZYmTD9z
uRVbktSmay4XDjN5IYmVf7M8HJrJU2rbIBaWqtokhzNwNwApqV4Gby5VBAko4ofAxcR+bq7WTsU1
EjM+ZIn33CcA/s0OW6QyORnwf6hgwYAV/SMldqEaBehBPK9dOq7COSIpirmxjLOvdcyymt1n6wfL
+ltq8Ak4j8aUpSIyjkUETYXy6U/sQXF054xo/A4EkvyXy275LbtAHdOHKFzdglgZ5k3kHKpfnQiu
H6mH1YVxA9Aml4z9Wxl7xu7pTnsGydbY/xqPWtfUEOl3l8y+vV1PN5T/7OnfGCO6HLDHJ+ISARkc
dUqpZjPtPxOSxsko5TI0wIWIT4JXY5xvOFlRoSs4zIPmuO8RmsenyEafszWB/nE5CFRBEjF5NrdK
zdwadZ32TPs2FBUtznMMWLV8eYeGOZprA+v72FTx2WvRnv4ay0HTAMnm6QRBgX+V0uZDeNKjM+tu
sJaiF9LNpHO7M9NlnWee24VadTz60UVOtPE2UnQhhwOMaoujidWzNQDNjHJri7dSC1Ln2jZiz9So
nNfHWj6OuU5zQukDRRVbUUdg+SfiVPfx+HhT8VJjN+RdkTvBUlB36fr/4mbmRTa1QUJYiyVg9uDa
hIL+DQ0HMvQusZWS0LTz6VkP0znJUbw/BUGOBObqTCwdyt8K6+OqpDUGR3oLALQKmcip/LnrHojW
PXE+gCNxBxI3qXAWOiUKYKufre0wHF3vldJHaSBOPADf4Cb1q5/c+VLTmu4/RW1HFvy4lEmKbLj4
uPFMkJ4cHYEza/XAVsL91yd9r4mCjZamoM0vdIOb93qWdKBPyN0XY3Tv0zQSCQslQ8cMvBBG4l2s
GFbaAzWAxC4ysqGYO8xHonM5vl7W/zXlS1GmJl3reZYovOqxgYXaRwsAnFEgBzeb3Xr9v0LNRHJF
rswr4hKKJ2WBWA5XD8MQi3DmT2ovdprae5lR8RTqaTF2UwP9hWFOlDTq1PqbzqX61MKCkTsx8Bcs
GPMAgakY+KOH4+KegShGueraWIgyxdBHI60jc6O0kFdPNR+vBdtznBDmjhnNHjIFDM1wSuob6Z3V
BTB9Cb6grTrru+K50fPiaaFpt9zNeVla5771TEF5fSvkUtsrjC8KlhpGqZd0+5bsXdbXUgSGw7RL
bL14MJ4iHyY/Ki94HsPF6e9xtqsuFAEPgqUdNSyCgx/lCrfemV2M9I9WazdPf4cxHP/0otnPlUKS
x7O152gIgXxuouZpMwu+FUOKXhZ243k8BrWu2QhPI5ggTIUQ1RWmKEdqOYm5kArvaQsKBBIOAh5i
E1MrHjOEHkxVWm74k6+0VN4+iOImVCoBpSQjK8t2Yb0nlfPW/MAAzOvG8u+uJ7Q22nTeeV3Fk+7U
EI5kij67NUIc1ergLaj4MCMmBlBAX336yvA9gbm/hXe03kI0iBLSTNhv/Tmp13RoFbIKQFBPmmTu
9lZ/vJh9myiUyT8EQJo+uFITRq7RcgFXUJ48eUpdLyDiWh5uYIDGn2NHyDpOtQbm8y4vcs9CeXrc
ZPv2BUeW4H0NDHZNyz8ZV4Yu5DSPGn71yzinvqsrNDd5J8NlNv54HD32gaksJEMca+xqkEgnQAfT
cj7aWkBVmg+O8MKKFQyDFCrTAxMDDrRSHaZGvtaRhRhrqBxXIwdabvFM06wuzyy1FsxyD+t4imL7
aPWect+ucOtoMj7V+dgE0SZzTlmQeWOtTU+LI+hUrMl4V+5yTshnUAI0JfwokX06fdZoc1CJ9ADn
BIwhN4c0wDzUYmLQ2GYpisNUqhSA9p96rf3bdtP1uZBgZFwjwzCXdcQq3oE0kXkFwMCeX4wwHAii
6+g5sFd0nfI5P1+SmeNlA4TZ2Rvdk/GJGn45+EJYS+lVORhqoyn3I2PyJ8n2ZhU+hyYZT1wNMFiX
lbRuyzzyo5roiAPkuMKEK1Cbxs6TERr6qyP2k15lIFMy68ndYWzjIfVLA39E0kU5oYhXbhg147RX
QRQUa8JzmCS04eQKAoBHVXOnrTgwdRZtlqgl1FNZgVRgkiKifAE1/3VlYY3okuEvwVLoyBXDFzZN
KbVww2Mx/hkssVMKkvVrUYSOnS9xIjIgXqO5wf884T/q0zaHSEf5hXfQwQdFTUaOOWF6oFVuvw50
sc1XuNvtNDUDCtv7SB7qHriMFEJPmr7gx9EWJ7OGQsLN++rpIfs6eHYEQ05ip2aiRykxXm5N54vY
W/OdQbK8MBNX1U4CEN9VWpwmASrailZgd6F9i4NNTx7mebMsrC4/UnkzneD12l/93mq4Nb0BvvDh
3ot+xLmkSDMOOuiCIF2MuCAMqXeYyvVE5zEY5vu8NBaPnWbid5cC9unQPiWdfYEW6Su0JieG9Kof
an1qOvtD4O1YfqUJKj4Ev26P0sP4CFdm0BZwiiO8WJTT6X4g5dkgzyiamDy4FrXcYH1ZOFS5yXFq
vOMLopjUg7YaM15lAyxvPsyiCkMr4QcNJ70EgkS3Hp3AJQAzvmLIrcZdapPgmmT+P/k3fGATj/mw
ze/IPtH3KQWf0/oj+sMB9aoiZxN9FhWgAxbozBoXVIAFie2n72wdhbbSeJKBzD+dDCEJzlFRgs6I
6dfpRIXO4FcngH4nyWRVRFry5cdF4aHa2mexYGWXTxMmTJuNXDpN970+p3+Nj+JuLDqHiGTXl5vW
6764o1u2dTYVC38nZRVFrtCje239DKNW0uycBqtl5ORIEk2BqHXse/HvuW/AlV7kA5D5KVcFOwJX
VQ7ySsdDSF+u85hibWJVgHmUw/N0PiYocZx6J/CIRi4SyLJERpeyl80leeKRMd4WR0TkcNpO2zyg
eRe8917ysPP6TyuzfEQraHQOS7GeqIwyYzX5ACjqT14BIreIYIN1r6enVuamXG8mi9lTrr1c3VKq
kivvysRiNtQIWHFwv8q7mOS8vaSO8JejDjUwMwmR01jViGGH6hM44d33lcITgwZzQst7gFc+UNVb
WLBXa8NFJf/2qWgAREwkcMRI7anNK05TmOuHWhAEq5wFQVgwhYKiykVLm7hQ4rCNs/ILqjczTfMS
Fhh2Q+yR7RdEJ/FZgHpSwYUgJcIl4uzWdbCxjfJAdoOEl7X6h4i2eDx+w4zLOcJoIqmBXLDDjuQ3
dnjN34ELkBKiBb48D/loZIfAZ9hhnFUB5+6uI8Sa5mXBlfM7zQWw9ysAYs2XcPLAX7s7uTqg8ry+
NIT8LDH0sJXWfLBrqslr5xEKKr6fWdNXCLIXCfoW7wjh8DOsEsISJkSuuuhotouTmCUoGBE8uyQt
mrojPSX+QIl1YEJCheX7m4hzI3lvSjBElbn0UUbAJy1ZqbQspi9icpHZitNJKVs+DCiPpn4H7fwW
56c8gOSlFII1l5gkTO0nsWCAWKTPu8ReIwTQbPdLxKrY0azgzkG70kcta1Pg5zv40hYJGu1+2uY4
49OKhUsVnDRU1IvtfuxJr3EKo87ri7pUqcRG1EL2Dz9rr9d14gUVSPDrK5xxCKq2O9OjHzoLa4bc
7up9+TVx+YAzTgJL3pTDcS2xs/jHeC8teQSwGkhvhgv2mgv+Lo0XlwFTVXYtbSVn8aLeW02iCs/z
8aRmb/RAaAK6CUd7S643E3OZQVHE5F5Mmu9C3bOcHFbszv2GJHXCcg5tPk3f3ud52mXsBxoCi4vL
/3rrNWLqUtSofH5Fe6tfoOJZtG+nw0VpIUyA7ag1BOGsq/Q558Xw6gZb7cCUGVPjJxxJkk646jbH
Hi+9qbC0wuVHgO5PGOL1SViqX7+mbBYXJJjx09AXBO4tCu84cQ70jkneAeTw0H7KqNYB4ImwL0yC
OSkbBHWwqL1/7EVJC6tU6QpVQZBNFCeMvkD+iErljoMpH5BBkGHZzcw7bgU+PkUt0KDVUcJQCL5f
QN0xAFfRKMiwSYIiUneXzlsjswhVueGrJ1y8URzEYz1BlYzKGQwjm/RRsVYWm1gCkO/frI1JooTy
bXdpBQU8VARS+JMa9WOgN/8iLeJNBAXjyo75NaEeLqWITK219HjE7FVllf4cu4U/W80ssG+eRXY+
dbJ0AruKiFsDAkYHi+omNxRFFYk5wp7dFLfZlrbVIRVe8Hv/9YUuJpJce/Zm8HMNf/3alb5FcdH+
o11kusMz9Sn53H4BAAOCCUiY6BeYDH7jO6sKUpG9ubPo135Ze1unt8Ac8b6nGfoUBStGzCPlRx6a
EJYG0mONlG4kymsLeVCx5oIBdkj13HNSF0+c4L8XhPmtKLSXgsZcaN/fovu4RyV4ftJpG6nl1PjD
QOG3yXu/CTkF7Llf5DsmOTpog2r+FX+OcZqRzK24H0PE3W/G3KqanjNHAARCaQkzifn3ZPM8gHV2
7xbpJuj/oewUh4yWVFueYsDW1rMLj/nyx+DeuIVAEoJjdi032Wiqx1ScYDUC8LuDGJNUn9TU1Y/B
VM1/ICN/drWSTLfYLWmV7/VNQhZDqghZWyyyxWSUPLeiMED80QAnJod08rELHoK23H5FdwgO+iis
VgI/k7Wv07tX3DmMA+ctzXtpYbhGh5kbGELor+6lZxiI27d++ETND7ICH3+mQ19mfGFIA8dNSYsX
uXFTmrWmTWINqOaAhvZnVDahgGDW35EssUUm8u8TqCWL2XDVCPGitRDycJRRI8VpxzqFKEqe0nar
gfCl6kLcwmhr+UjYCqERFdeGRJ46KTjiAqgnH0Aup3KCUgk6empG/Nwa4zVlLyWHKXXeMl43IsPH
PiTa2spzqLNrF+wFNllmJSwSjC1cFHWn45dxf39sF1Ce06IP+4xi4Kh4UDxnTuzBE0toMs9WYoPZ
VwNw3umzUPVDfRh+ZkBaFrN7UtI+F+3BpPY4pUWRQzXbhLYnezg+seymSiP0ReMgacJCLfg9gKjI
16ouyGLz2pthSMfKgufC9tDN2NhW2UvN2IhODvwvhJ+nQX7llYtJQPHvmAq82ql/nkA1ccSZrXKG
/tOF+Nub3vzkKhEXXuctZPH9q1rM4Y+ayYl+Kb/sSu/kwncTyVHXMKKV1PggaYw7Yc+FxF4N+vDA
K84666PNd0F3dhp/do/L9Tse6fvWhewKa+ZWqInIshY5ywHqtDGuVCiLJ+1+rDvjTVY6JU8f1l+/
ElhwhQG9A1VvlYhdBNdAU5MK+8oBOFCa/48QSVveYiPLiTcgAetrp630fBx/P8RfQWu5TFEp2eP/
ClLgwgmOWsmsSB+M3EjALBbdI7goslvnfsn2LcokuRichHv3uGWp1PlsK7mvnYMX2/7XHa1eA9Y2
08MXdppU8pqmRCZVB/7lXgUx0cKtO096RqrvdghSju5wslxYjqS93OPxQoq3rLf+VmK+j9QL/Buw
AeBhIF1P/YNi77FLuG0mFp1fKUE0Imow33rwXliEWHdR/V0k45ys49q7QKdjcxoWp4SKxdHeyUpA
b8bk/xwy/LVANRJgTfdM3NIXCnqSuRQRP3hiL8ZHL4hb25IhO4akSkxUNeHML/9g2DsrxCRatN2G
VfIIdnvPjcqUD0aHnuFnAj6915q5YSj8gbM15pIxqFNYSe35+FLBDMdOTpEWYvzF9rjEGOFDm+20
le7EXrALqfuQcFJ7uf4vlFpdBqJYBdonQXXLyojYs3Yn/YwGK97j/VLRAZ0kO89SzbPJRoXzjmZT
jJYXWkd4XypMwG9U9CRmefadDz8JQKJXNrb3M4cTZ0LJL7+2AS8ouZMRoBKyV/u7A2rutJ+J5P6D
rYO1XOmuvq9kahKa2C8KdoeM7/Bqqxq0O3JTxl9rJ6fTmo5z5ywhC3iIVuw68OBjWImZ54xL5wbS
QF6hK3q1IkWBcXApaDks2gyanvAH7rn+THEnq9/h0MXAth+0uEoXV+2lKWtYtWt9BalP8PqnIz0p
qm/QqAbrO4B1vcMMtMIs1QLrAugcF4YtH6MVXN9StyPF9GNDhoOd4yotjiSTQaVZHsUVVLCtFCqd
vKEYXFLj+e5zdSc3LfuBixEYb0YeUQYcwPVy7HQmZ0Ba8Ozf8+yjd1ag92kRfYdOFTwbKhc/O3X7
cYKox6gROXBGMioz76j0+a0w+J3JUb0W9Be9XuTDwY2acxcd0Sfni+dQBJTT9Y+RuEBahCDkbPce
qhrp7xKBmZ0DBNHmxc5XJ7tPI8WtHUYNnUBdZDEXbk4S7BCRxA/ZIr9lo94EBHzanQ049N2CZ7hT
dhyuxMAWNaaYzmyUy6lvYA0eHgNu4350CHIJQoBR4zj1pTDN8FcuLa+ikytt3bb5V1+Aoz0WRapg
tc1hJvHVT1VpTCibhijowVugLA10meoc3lXs+s5HW8VKBINcQz+n73H92StDl1JKNYAwKXBg+OMV
fpXbFcwHScVCfg5Cg0Pf8ci3v+LLyEWRV2HIxYjcjKPNuJMJxKo/wl/TALjfZOVV4YjCx0PMJExl
CbId5cRFXS5EBnbaBG72Udyl/j9ZIHJT/nchb8DBkZkxh9cgMuAuRJV20zM97qvxMU8Hv0VENot5
Cl/m2XuLewBdWBsfoxrm+T6onRxnqJoryj7CRop+7Yxb3dEwHCHlfDBHVJx0vB799p9DuIO2fzwA
v1e/Bh5qFyoMoSzvglc1PohUOrdiXp+0PFimHxSN9b/OitS+1w15AXevHMFTKzSoBgVB+EuIYAHl
d6JMNdphTk06Ejl0HEJVu6HhDif4GA8H7p91wx8F2lenvohdU3O+ChxIu8XgGQsDPVZF89E+Cfj7
wH1K94STCRJxeuCud2BHVmrkj1hRdzXLqwGh/OlhdxtuUpifjTfo0iS0/nBdKy/s3bYRq1sNtjc3
jyooC3og9ogiEJ8D533vreirmDU8x/vSp8259YRN+LM7gHVhvDpvCZhrGvTLf/j1yld6B9Gh2qxq
71UiWjr85psgEUGCKjGdXA2ymqXSac8axHj3HymycgZpxJF/DaudFGpXhFMKNvtGi+quPTugY39Q
QkMDuKwg++nH7rxhTXSLnNzp7i4tNbkPu8KIodna21ACUDp1B2Tlm6xHi1oXZ3K2kOGXYrW2rhjC
FYsGVC6C/FuNPmEFL+n/WDDZx6RFQS0VtucCx0tb2f5iGbD3oZdGIqcAIbDHd4Aj6OWM9uZ7v+cg
4bG9+LibFguItOD0/lXZyKi8UhKE//ZXmJsXsH0RbiTNsbe27pQ20337FCF+B+6KEqud7kuvSUg5
g7a3KppTc0eayhEb6KDV6b/aWvI1rW7FnWMzaP2Tr97xaWAvM8yXnWufHhdHoNiMBt3MnvxR/f9c
z/iqVNRxjPikoWwMXjS3Jh1nO61N3n6nTE6zVNjn6f0q5RjWLHhvLpVyaiAoKCpDgZGU/Wy2IW8N
NnSxMTejPNr7BHTrTz/4mu/F2N4YIOZTG74cUj86JpKh+xR3kHx+cH7yTSU9ti9v5ZDbB8uTZsHN
JsliekNO5UWFd4fjsq54h3e5iNH6oojpn2WPeBXRzOzhDDx2hhvaIzTWAy83dubYhuVZlAijGzsI
c9WNqBIEZoqLDqdDCDW6eNhWsc7gYAj0SSLhXjgLMTx9YD1/uljjO9v3zyHWTUd8h9umDhrcxJe/
ggGoikCV/zkv+1I3ck3emIDcPcX/f0SVK1CgdR/IpIUvhxYHUP22ycsFbQ9s4UeSPtvzkCzrdgDU
JXEi+Q+vH/Wm1t5FaMJMDhwiQyd+1zBPrCYgeqgI8peZ8x361sK2WDp3jCGTDP52EtRB/YD0BL6k
xMU516cOGusQCI1vT5Xwvf90RCRwO/OlefevztjDNKBAzkMDBcNw/zI4jJV6eF1eIp0kTyanVPH1
coUjlZlhpIUO2Stwv3NV0H75/LWMRePLT9mBGY5TFYA2X9tQVt5tkprrzG99ysGDOFkjK1yVkLxN
0wIQOqujwHVwSgWXZc5ROrXb+iAlK12e2htWaO97yK67B3D2yY4zTFlp0PPyQMQaCi25rtihXM8d
j7+LGO7HBrsYosFRzMWMk+haznsdHRXWso8MfuzW2RILXnvisLbbXd2UMAzZteoKZLIcCB13hIlc
PkDlxZrPz/6iCoNOBqkqUtLB3wfmZ6+8gbcq71MQZJcGlB1eAMmexGiI7vrrfKSO/UBApam/Zv3Z
85CKz2eWt/rnwNrrMfGPWZ6QlQu5eno9yXuVeBbJLutSnfqCHoELaG73pUPBeCn+eaV9qL5NObxC
dlpnFq2HzGKnwVudYEqyB5ac3QUnjeMxjqVZNutm7aZRy8845elFJpWSRY+aU54/K+Wh5jxGrQ5+
eSPYc6ku88LEL8fju9NTJA7kI5cSAGDN/M9PKTJHTWebHbDuLbtygdHenkzCPJOQEnd76am8QCy5
cQpLfYc08YeJ5JTSbSEELPrYZMGkiLMULPrwocGl9T/cRjRE9NJbyC+VhnJyRlDjLgVJcicAHu7G
SeV0NYnRucSGNDGruHUWkUhuFbjetDwgzhHo0RLheFbU3tDwDQm9/sXpiAndOOo+MGQdIdCjZ2Jl
OWVb7LCIfbZSr4KMgdYE30bRwkVdUUz9+Eq2ze/MN9+xLqivUwqKsZgudtRkYb2hXAY8sZGvHOHf
ZqIaRBWlAwC6gn0rmhg9RMIvb1issJrMFNuj1urwxzg2Vq6hsCm4F9m/Egn+jxs+Mwc8ETdxRUnU
l1HYVgRBW0ATYOUOONjIIUeSAIEYb2mj/uoeUOo+apAe0vBJQcdJqq6S55urkIAJ0a9Ah+8vXzZ4
Js3jUU6+dFG40i3bWcTZOd57thXjAcn0MTEUWFu62+MXmqo2aY/gXn6uVGjqk1D2C6qNeAMeGtLS
4X8KqF/RbvGVzVGa/gmw+LxaJZR6oIkpO9nHz7m7xioUgk3lhWVojrnPjtuJOmXbafAbubzfSX4X
oA3Ug6a6uhDO4X3x6AbLR06W1rnNlcWEAnbcrWIN1iqIn5C9u/ABFrajUIjxk1vATYPkekLzvyId
cwI+MZiWJrrGt/JTCK4aYYyeah+xz42/aKnOfpWeQ9F1fsdWl3w/JGmM7X3suNn2MQ42iWI72/Mv
c+wcUZbXttOyO2u1Rk8PnpgRh3ts11ZiepHG6V1g7pv15818KFpicbYzQaOrRM8F/oYSm+SlsKrc
j1Ky3V3KdQhSxRzmJVyRdRAg825LOmIVsbPWhECHPoYz1joFL92ahQg1NJG+q4qXACdHevZ7oPsI
1tHuMPBTvwonmp6gIAEjp+okmM2n2FNxTDD8Jfw8j2DcuDlGEQxmyFjy8crEjdD23iuchDx8rSLP
qnzLlA0BpAVo53i6WhxShGRg/fIzig0rztDhhNaHYpKnUHVqyV7zdQxvKtz/0pyYJITmWTJ800eO
//pqVZpJPVt7f8YjxoFgGc2iJl7VjhV5FRwZfPPSnW1QVGWGGcio9Ar1UftAvqZohB8HcZYICYkK
7g1BPT6KLKDuivLLbSdh7JoCEsKKCpWC9cajUCHr2VHz3Kq94dr9u52AyAxEi8OyD128HUGlYfMz
58wwTFnoscUdm0J4wrU+w4p2grYlDfses7N1seYcay9C6Xu/BIzTrfBVMdiaV5P2N7ucS2mlI/mo
0fadtpdmjOE8iCAiad4wjTNqLPyGB2pZ9IziZBi8TZ8EXztmvjqJnz2VPSPOSqe6J6tvNuL+uvtk
NVz5oOM4iJxfSg/HoAUnnlO2WBKzJyJTTA97z3ENz8toaLA9B1t6+JWjnx7XRJl5yBuZAHXH40x7
Of1Uj5RRKkyrGhB32JBre/lxvRR4NBAhM8hwAHRucYEh5BBSpF535QlBsoYSmpEKaPLkdmDd2bZ1
aABwetu3Q/enYnwUV17VyZ3yPQh3hUYelho6dgyoU3xX2CAYpO56TDpE84gTlwwuYeV0GqfkQZzq
LqGbaAKLNDdhs/vlr3WtIRx+1nl0ukyU43UmI+75DfxPXB/mY3SEKvChdtNhl2e9kv/29hXK2v8+
DTrXRwsWj2BmWk5nYvie98hHYj3LwUfxkadzS/M9ASoS/83Lcl0WYcctDgL0IVWvspqcuiA6WicA
HAIIacmDhkFPEnFgWrDWzbsnmqs8ettoUa8nQDuL1kk/JesXX7b3bhzef6dQAIo+ubALYJLddSAh
ad3xYW501b5UQAf9Ux7Fx9s0LjHVcMjdaCBFCkJ3fS2NSSGXZPU2u4dc+KeekHUEiZorzFCETv25
OczKwVpVtDOOVk7n1FFIIgTY/aF1bGUQPN7ppy+QIKYPyMqfdJ3nQGV82RhkWiicZgWRIBJyy3Ym
CfoKis7Xcz6oM293akVsvAnSMRyuXxeaTpPXgg+Ge2/C20J0xtvAJuljSNnzR6T7JqDkJPl9HVZp
6xNTSfA5DUFKsFtxYHovjJ+FmMLYhF6T1UZ8h7XV/8tz2Nq7Q7YgB3tIOqGq6SsQlZpnRfzxOesS
yg4tu0FuhhLcCWZZ570kh6u/v7kbGpUYjAzoDg+Io2sIylQOcZVdD9q6Eq+fqehpk4FHeaF8hxBD
cCzy2lhE7W/5pufXrGLovlpqg2Frww59KMopEMLbFmWANV8EkGHuOtBc+GXjYo4F29fUCmYo/7bD
by8w4OaKv2F4xz+InzG20fSJeIFeaAh6mKZ21BXvDt405Zkd4NjQT8GIv279HZOmBZqaPeaJDuKJ
Nc7lU+oa9K+c+ZBZj+5LyMtk5ZxVnBIyo70e1geSquQL4qcNVMci/vm2H0OFlaIZ046kQ2pVjJF8
z9YBU6d5Zzd2OQ3LwOL/hPOLCX2oV9kO0OfD4IdjdcrhwKsrPnFn34HlNuWN82idfd0oDvG0PvXV
MqI9KuiI/QUqaxNfQsQR5VxASwYr0YCwnM3IuyA+wUHVz7m7lZDCVjOH2RnMpbTRCnZepr41gIeq
kiDdz+qHPEeaKZUqLeqI4+YXc1uNGjprhBK8kuDTCOLMJkY6h9ZIe7ShzR0DsUwoKww1nrhVTJWF
FzAXp4Voeyz6FrQdGBggCPwD14ktoMCCimy6DoTtpApIyQgI34uNDsjtgGgKAlzrpxkTO3WoBwjJ
8jrzcKovi/26EDNbE45o02khGTYGA781tMLSKa6Pus34CtV8jcC6BJdJmfC2np515j/rF2iOe4zX
6XcB9Nmg5lnI0KpbqZpwjIkdT78gBVn2IraZ2KBxkQ7zA7TrV8ZAd+dIxfanQ0bBaC6UK/dqDsZy
5TFvoxG8cV1Rgvi0uulO3TWvlYmc/YBYouFOcdNFBVjC+EMEJegOTPThMyn6Ee/fRtuxNTBTRl49
TwCMCkgsf6SHwx6DEpKLy78IVpmu0wVaKuyFoDxYgkCAbQrQBujgwhanlt/4UBeb4tCDqcHaLmjW
DSSEyEp8wmrV2aOTDoQfuCR+287YmDDlFwU5qIL2jE1MQHTZ8pk0Rz3+wnRLJXrLWWZS5J7uCyaV
YbQXxliIQ4PRtylscrov1O/YaXQwHIM4cQVOyKQBdLcQ1Mwho1h62lSnCSkJtIbotAioENw6C+NL
7hbcV2hJgqb2UHHytE7gCAux/EpqCsjoditVjx1PmQA+B9n0JUgY8KhsCZGhViYdC3/aNInniUV5
rlYC6e13BMxmIlnFGVQPcDo9g5bimdcqE1dtHKU5Hl0GLvyhVbSHGUskrZDzdSitZPO8mICH+8+A
H9jf/XztbfXl/C50M6eJXRqivkOH80zzthSrBWwSHW5jhTExNunGAsxFmLolLnpzcs8GHCBZOhn+
bgsDdFKCtvvzkl4SWTkFspq7kZADavSodRanajKm/3FyKxhEwyKUn3tFJ3twgkgomHiQb6UsNGQf
A/7acmj7O9ZPXRiAukv/GgICCJJfKgxY9dadqedqlbI2t9LwVpxNZy0CU39CVHAr/5LADMsVM9y+
AdA9Al99GkM/aZeb+4RK5uENn5FvRTEsyhUqMTYPs4KjxQpY1XSGCWa90cMnD6yvproWnzXOzMbg
BgtfzOjqYT21o0A2Hy+QzTx4/7U65KOtm6DnQ/Eal1qgiZCDGxmEzMvRTPORcKEnqmM9yCWRPQNB
Tsuf52q1397eeafBH5q1JPaXA4y/ULz9u4vtkzkxCJQYVWXoi68nJs0AZQXQRLE5NZMoNzL9e8Xn
b+uuZ8JdLe4ve45rdhXXtowYKQfUu5E5ez6ie1QE0O8ArYGfXw5idci+y4Wj2QQ9UURTWDyiE6LA
vY5t4PyAB+b8EzQrhggIGnm9oDmbr/bHzyBYLg/VccfOPaiax1gm61Zq9/aXZHUa+8+hA41MLn6O
v9Z8E9H4K48UGP4WoZS9CP57xmLT876VXesyph3B6PMkiYHVQxw0aBjK90MtJYrG0o2WUP9vpBrX
ztRt8khqqghSjEfj0QbiRKqYHBZNQPg6zyJeTLEBy7t6wBM+XKQl9rWGxhPHqP6BXV8zbUx/XSrd
/rM8+Q2/rvNec03MVoHqlyrYwzeJExUSlCfF8GhSdNcKeCB9KvOxSEQVaHn1Cpjwef+R+87n72dO
4FgDx09tQzBjcTY5X0jZDvWGDUnQRqraltq279pbU1fd2NM7IeoCN+f35k/lk4PxU7wzO0Lzo3L0
CngfRwST/1GOWjCRtJpzHmW9KWun55FSsorQCQZwqGI5SS6IfEeGX89YhJv9/J+i/huqKvoNmuZe
pHUhuNHGZ6U/Lw1TsNAE8pGeSYd60gYwaz0uB1Is+8zno4TWNmyJrPyxRbTe1R2SjXrsELfDgNsr
7749CoA9KAbwiO217sGA5AYSUbQ44bKEN7SvZ9ZfXRyF+j/VwKzr+a/GXdU0dZoTz1QCXSdEW3zM
lYNMueuxGCLwTrmA4gKwOyklQ4pmyhD0H2AZpC8N2Y8qJX/AOLqxc5e7cPiz3q6WCKN7yxJGeqBy
A2/zBmdofUduhEJKG+b7O035B6t2KqqV5Feb0Fs87nQdCw59njHsnnuNDa+AaVG2KnJ2vDHQ470h
eGE1Y8pkIu03aRxzmsLomNCC1RjBG/Gr0HofOfxviFv/uOphnVai17giy81DeQHZrBydKBzwEbeH
irDhlynOyC+J+HjD5yEW3u87qSKpakiTMUyS2izz3n8XJeqVormY4jePW9c4ToVAYMEP7DaROFPC
cZyCTmDlg+r/u86aM8LCkGHJay39V+Z6AhZtITkkpaPntsxRK8gAmLNaf+9JWTKWuKj788Nevf6P
aNtgCx9aFTfpeixBiJcPjUjh+OMciMoo5rFf6kKE8xS+1scf3TeEcTPdWwVceHhOJFPbflXNJyfL
Qh9riyPCePst1FCcEtq7IzURSx6sOpLV3nbWpeSVYyTqph8sxjWSgDqI7cukI7sMQ3qTzQ33ViSB
iXX3fh4dceuxJUGcGKK1A21gJzEN7pmMbJDe9aqita0son4cTK3rbzi+SZkNVumQ9AWwGGVL67Nl
zJZq9YVRfdpsi/trnthrwzJRcnnkh4SEM4/li2TZHlHstjcuI2ICeGyldmrwD4wby9/6WB+vx/5P
HODPb38LF6ul6861othy8e4/DKNawiaidno1bmVst4mQ2ot3NNdq9wu89rs9fKJrtIb3hOdUjI/H
WAz8QL7GckCfkeh3ATXtw7Ne3bCk+ftPntAALycdSpYfKd2dfGrSRcPuIajFQ1XXgBYH7jzhl3rP
cWtL68P2ttd6VjDsMIfbFstJBGBXEQjH1f+tHKS0nUDLN8KbnnLTWVMnAZCONEPwUID2Xv8OwR9I
RFSVDKitIDTrbDYd6/hnGEX7xmh1LrFRIdWTeDwhtjPG6XIakXz73PJhMoguo4bndhPWTt7u9soO
WtTiSgQFSKE9LaeylWsz1Sed342CkTVvLv6tsrWKEanhiYvO9uyRewbKnpSfilAyPBmQeoH7Dyw5
x3QBGLWOYTvMUzP08KhiMzsSmfbQsXMBGDdRVzdv7ba+cRgo1eg1rnuAj6hmpF3miKbUZpBq/eIG
pjeUGFn81w2x77DE+795czEXNYiRuhwJKuM+7qTbzZVV9p3qD4y+bXw8IteZCFpUQVHSJfJyz0qh
5U/LxZ3gS4oMK44Mk9sf19L4LxKAGDMlDQ3hJ9b0NH+xsbQaro6nzYXo4rma26M8mfWuyJCXy4u0
HFxC/Ib4kq22hdcMgH6DyRIbFdl38iKV5Yg6hAmSrgTXnr2xnpGr6SjzzWUwB0/IU6AoKqpnuITE
isDdBkPbNt9y9/5Y8jn9R0d1kD0UvHkXmWkanKYYsqeslxxWTHhIhk9hd8EbMLEhu0uqhK2p/Szp
T6SCt0DJ1QS8v3KevY7w89OKPO6jEW6RBl6EGwsNpsREq9m0Leu9HdI74bcMT/JAgiHQ1tTcHExp
+CfTd36kaIufZ4PFbqQ3SoT6EX8wQfbHW2f0Q57t3L3LB8ntkvTbTdb8E+f829tkiP4rEcd0ysg2
qNfhvfLTuo3wUfG8VktC17ucLWweFdvYJ3xaXNpMcs7ZBuXunfc7Ake2EWRJVOh+OotPTS+bzt2P
aqCeIIO8EcTBAVcRnICynDddLbf3RNSkxJC3wGmE8V+5tCkcZ/kZZUmszmRAL34UF9VPEKjK2pMC
ZHHybiI1lz6T4VjPVlxoteGEenkOAGZNbxM3IfPMig8sqVsQ1gEtTtA0uw3xBgVJRJim4zx3VfEB
L5P6aIUL1fr2/prTfRy7BhG43LW3OYvF8LXai040Mg0S0iWr3Z2Zek7n8wYaCVFWBZjJqnTMWNiD
xFGb/L0FIfukeyOgwpCX+w0cwsO+FuXccOpZfo4CUos/az+2BQQOBqM7atUGxFXWD4Zv8Ov+OG9S
N7OSb+FrIYa94Ghds3g4IlkTNI1ChY2CjVxvs+gDrKRkPQwtu6MiQ3Kt9Twu0ltQsDjHpepZKMOE
jRg1DF0bbKuK4pJ+GcMyFbSthBfSevV3OiVwvyAPRJxs4h8Y4dKgh/E3g1BLtCRSweC2QmUSyQNN
eDURNNYPmfYkSf3YRsfjDlv8wvDoxgHA9CmysY60vigHhta86i7MHE0Bg4+eUWDWJWN6Q+VGUh18
HP5XsiCJNLxTgjVvUUIjH860OsP0Rv0yr0swpPBpEQsQxrS+iUyZImqF6CUIyN4txxVjkxOJPN2l
oG6FOhncMvbG/6ER52x0KFOD+n3UtZNXN+3f4daHJ4h0Kf3IGPQ/9XHj/jT9CxFahpMXWN9eqMyK
AHLyq8kbLEFCilszvHS5i9GOeLPrchOhCiXgvRCTRFwQJzyed+MXgdlzFbLoYGsHy2Gtk2bQhKCQ
XY45Lq92El6KbCcsV0IlF8vmUsSBtDTP+TQJvUEU2WV8z6T6mXN6SJ9h8gb5rlLlVpXHA91oXNMp
JMgKJlaPYmbnWdxwLrP4cKe1WkCYvoJ39l0xCpWrU9S0w5VUT0Tk8HpheOhuaaWbvUyaWZx+qOYK
ESbZBVv2/Ug8kARkz+w6Ehb4CsKzdJMBaAaNH95oST4+88icB4SHDUcUQXnNTWoJZLi/l1R/vfl5
MeBJamRkT/t4yveuJMMY+LZ9oLIQVnkGsIzVii/jjqhWwCODXHwW9K3k5S9PjMtJqNogRI5YDAUC
KByrK0pE2UDJDF2A5alumvT92J4BzwAW+XKGaU57xqzCNLIj5xzQqQAVruJaNQ3pNRw2dcpMlQKq
UjZ3CafFnK4fKr5y1Bxw6T2QkeBtmBTOgmamK4MOr6fFUDG4NrQIQEu6glX8q9iW3Bds0lx3z6QR
IrRGQz0DRDSnH3MDapqq/9k1h+ZINxuseTnZmqtSJTGK0+3khAZ0vt9glKFHAfLtsFRFqafANsVV
ZX9H5jgPNcJp07qEG+PLFmknKBk6hru+gvfPiJ9Vna1UGde2OXAu9ucQzndvJHaE6CJoisVx/BuB
m9jG/jeNeam7Ael94yCkesuCfro1++KSzXpHo3AoiTo72t4ZwPj3d3IzpnCHg5uGYVqazymYBFHN
rjcxVJ6L5aEj4MuMvyC4EcWEdQdt8ReGjvFJB5iYzRBsnD8oYmP9JP/rLkQErExYG6GRYNgJt+cf
VoxCZCBtrz/20Wo7Y7y6cxg7ffd1uywZezgxhaU1SL4LAyJM7due6Q6dosB1+89xNFR55ZLih7wn
BWTeAfvR9QhsM95L7aLdK25UVvLaPwr2TrYKjWwm732EN/gW93UOhuU2Wavc55nf5U/94oz10Ca0
BS52cbM84b+SSA6ZTs9E1QwsEklOKcZE0epODnGok23nzNgASd47JX8Vxk/CKbRYCOdKbfjC32vv
Stg9+E9Lvxq3bDSndqqUoDLd8IqiqU7To7fmUIneBOp4z0/VbrysDRtBBXyTZ5O/jjG0Z0couNXa
fiOfRDZTb/cylkYraOxCrgK76xxv7PrNTvf+3PVazphzvQr826QSYcztwgVJf2wmgBUfPiGA+3DF
hp2WGjJZ4OmODur6SH3Hp39vrZZqxeojtKxTtw0p3tgqQTS3Ah8qLgCeor49fD4fa9zn3zbV9cw8
RDD9WtbiQRYhxf0HTVfXJCxVU8Mr6op7vZsI9g3Ara2scFmzgyg9LouWxzZ+Ox8+JAGhTqgW8JB/
qPwpqy3FM8VDUilltbNa6/PgQuWFVyTmLJhfIKzyHEB4ZFyyLwhk57901B9QWzofLKPiQFt9shmM
MYgdzkD65vOKBdEWyfolhrgRWyQhxXkNxyVSkZAkjSE+RO6bWloAAASjGVInlBF3yvBBuePClXzw
7pTvqeTx6Av/nvENJaFdpWj3lcani7gSI1FcYZUaYq12cNrCMSF6M5dhlHZeBmMzwrxvLASYpq73
SjKhf64J9DFFesqtD44ryRh2Bb9X6B8Bz3C8VdQL3MkvssBtyZdmU4a+ZKK9inNAhZEDRx7s8pWg
Um6Z3gDhQ15g1viXu79X69ak9e7iv8cyhNNYrOAIrzUA5A9rzwNzmtW12745fvPmcOqUHpUV915U
6ekDVhtIQX8IZN0OTA+UQraGIeNiTCRqa/+QE1ORN5B1VPtFAHFlpCZQgR4e3S2a8IgNCZ50xiKD
yFIjmeT4jVLnC7yNbf90hceoHqdn1kO9z99iGkL/lDEcWBKqQ6Fy2+lEMsgdDYxtiQBLjXg3NowQ
0xVXvZ35wxuWo1i2j3xEGMY1x2lcpKzZFMRbKcrCZfhEjHdEkbJUZzDG8F1Tt+55uCyqxLVrt3bN
rMokJVexI8tOIIBmZBLPrKtsTGrRJts/fEPBWEKZNvs69uq7KEbxDmm2wYckj77YyL2/DjfceOhW
2zkMGrrAZIsBXb+Qk8OEBd9p8LsrK7eDfZNGdf9qi5dOkY17LPnGc5Ih6R3/AI8Q7C1GkGe5aztx
LddSERWnNsNosJCxURoAOxXyD9At6W+FotcN75vpB0IiZc35YF5gwhq/YREGSXkvyBZJ7l8m7IA9
IFT4MWA1GGg63gnZpqLr6DeaM7Tbq2VZeoHbIxKHTTr39HwDw2RKxkhWHI5pkedeHmYiHe/elhhR
/W3o8tGrgQd0SnimkVvIM7QHx8JAGNvU+h7oB8iOEkh38cZxvzBWoHR6PPVN4N/1bglHHNV3ScF7
QSyr7kLnlhzQplUuyOrnHFANL7wFkix82N8ews2dhIC2nPWOvB6li/ywXmAFweLfysZv/s9WedBc
QBWkXdSZSHVD9g7gQmQJyauSsY3sP51o9XBKPSnswxkLyzOFJur8bc0s1h6niGnJxMNUYgnLH584
6wwCC16FoflLFgT55UbgTdyVOlIEZKZs8SaivysYEJC1j01Wfgg5y7+eI0LLG3Y8JvrAL4dtB224
yRxqiFkzDYbAmVgI2U0rHiAYdcTAOUX/N63GzNE0Yc54ozxr2Sy17O2+1tPWtzOgVfknmoy1IOqi
P7mbsyd7x7XooKFYyFyDc780puFuZ3MHMj8O/20K+dB0u3GEr3wmXn4cAngT8hIuGv7Fh2JekP6N
3M/DOoWsGip624WxUOs11Oud7pQupmvpqfBK+zRVKMmzxKGTmHidAZqAFevfbTjIwlPUyE3vJeci
1B4bGMA6f3iNR7ibYGmpgoTbgDh9nGKQIMrSCSiamDqA5BsdytdFnsjukzPQnBRtMUWZxXnDGuKa
jTW/yS8Bv1PkQLvwNxY+IcrCacTLP3mBpsgScfj+/tzHyLesr+/VPdPC9QySEmEPohTr9lzdbmMC
JcTt60bmFg57f/gOSryIHRbuMz4bj5sEAQfT17Zo0r4TZHX0qPJsFpb3ZvTwn+bNMdFvLO7da+B6
ziAayPK/9abw9jX1gtKhe7YoogXIOdkkH8ZIMHroU5qQQCUEQ3QdltgpLx7MRU7uUw6O58MiaLXe
zY871wPNLxyY3Ey9upe5L1fn1xoTTieFjPIQqzhIwxKFnxJYAFvYynw7Bnjsa6b9uRctKcbb+Guo
bqcuXGYLH/YzOXUhrtzCx3Jur3mGyDDtVb9QmWPX6XFBzCdHJ9lvven7umP3cmzo3dUdP2xYGHXN
xhI72d8dxK4DrZwjTmEVFym2DSHBg5VfHLfy/qQ5ldD8jk0ofFb8OuEEEkDx1nuXZyS4zkalNvlw
KYmmGX9px124euE1IujNEDzJOmfi/15wi4XnNU27grob+y2uwX9MSn6jGnmZlbwMRxPJvDykP6pE
Fi6rLd6SccokqA0n8fEbZcubSynzSeESC1iDn9DrRMFLSiLMIs4eAyB+UlmLKv9/MnSErQ8tJ+oP
OnUm5G+AC2N40XRV1Bhi9JBmf2d5n/3+Vh5h9sIaN16/qKhJ1u7iUyXOaQSI4qwpJeec11D23hBd
26kdg2uM4AGQaNefb46mTVHg9adlhJr8CePsiGa1AOuZoBFmImNaiY4jCiNHW3EzIMnIZWqh18V4
D5BzGYfNc2EWUobdINcF8dqRNvPl/tAVc0MyDP9zTF6NAfMytgAzxxthDPE0CYtXlFZPHpT8DNhr
FEedPjxHAG1gQFg6awWQZq7FJEEP4bMZj0eMp4yUQXXKAkOyuV3auaBKmoq1MflOU48JrKcY8Ngs
5vq59MCU8JCvaS2+evlrm/6N4Zuf0BTK02NiwnyfRTSvh4GcEjvt2/VNQbFj6W0mMWUYTucCsKNI
fuKUBkCdD3z0M5IexQI4TD3Uahs63H+TtXY+fkKC0A/RN9fYeazAuRCUKSMl5Yvql9uYzKNuL8bC
dBGnSDAq9wyjcOE2a9UOVVZ3CbctJWrlveLoZpPHOfQYYB6ZJXYoazMM6e0pIc/EBZnxeQSIQeT8
AckB9ZsnuJ3VLieZy7B1HQ0JzSEknRBsXZdX5siAUQqTwlnfWZBYkS1g1VtK3vbpQjNqMsMDLzoA
l5AaC98UYLDz6pYEpskLNbMrL/u0qEkd8jGu2p0YtDObXWSsoZV7opZpD2KJakfzN3DxzRkohJQa
c1e40TgT1lArCvLppy5mR/nD6LTpR1if1a+eLGgcnbDK5aMNV+dlxoZyNJgcp0EPB/KvF8T0ze6C
H/cp14dlo6c40LpU0DeTAn4AIEBm+DK2gtT57PdlkMxnG6pK1fnB9jYY6xAahmHtUfUpOoSrNpDe
rQ5GRKegFMzgyoIRTRdCK1YZtWU+CrSjFCjb0kcov9urPTTVR8DIp3C7BXc5R2Eqm7xRUQTJOxdF
QX9MC15KGv+6TzHwCezwCcwaNrKEc3yEUW3aoVnbcfRivdRm3QzeLph/25hzLxQjfaH5jnyvkf4G
QyGIKZIkSZwrr/9vmQrV1KntbQtaU9oqhx8UjhGNypFywo5TGTfktwLzXk6qmPiRdLlMNqylXNgy
cBM3B7QPBEHDZrZmlrV16vzFCyK6048am5GZaONowPVcqQ0EEdteiNFUfa63LfYgtdHrUdZ33vLF
sWhnoJb8cXI3uOmLP1OCe7+4u1q75uKkJ6n/wfdigOIb1oPZRQz2SCjxpPhObwjoMqs7Lfi2TP3N
nlDseJkzQ9jic3KXEIX9SvoOfaskBN1MkSL53L2DY2/VD3v9TUDaLofteVEOgQoKYFw0QLd5VhdU
rzbHWLR6QMUn6LvaOlUHUKFnp8todqx+5EGTSbiIw1Q2xmPymPRVVMP+ldUDVjsMpx3px/2oaZx7
Rbui+xwBSY9bpTzUBgqF/U1Fbk49CUyOOZElYLMufYs1+sILjm2RisqMMs3tPOyMAmXPUW2V3Pu5
/cywCALuwNYIgkDmzk0um+sFj7HLzyzyhFDjvJ3l7SDtBLB02gQDeXh8F4TH6uwkKEQKQWaeDRhP
P+95EyAXx6vO6L2nss5e3LBKPZB4Or0MGBgQ+LVcsdjAGcDmcXtVMFjM7+MSPPsNxHFrZOHdtI9A
k1m/gMdvd0aW4pe0cPEdcYEjHa39X3/5/y1gLdq1HRdoSOmv/WAubxPb9Jh3ylsad6QOXhEbl7pK
j2dquRQZvhdaSLgUGkrLj9MUl8V4SMUHrAukn2X9vUcQLh2D2CKFquVZ5V2t8c23apdvASZYOQ5m
f6Bo2SWVKhnXNWhVelGRL0uIhLcYaoQL3uFV5Dji1ojtQ7C2TXLSlzPmIgiz9IchpeiHTNwfqM58
K+zfQLBpmdKPewOrQP3MF3a05XhA7S/gwZ9oCtQVNtOgvTyJzZW+ec3IqHmBS4K99YcOv6irfSO2
3iKSIK0/JG7Jq4RWQWr/GsD3Q9PMRvxmGDdeXwALYIghx/UqK34uUW9gubYYug944kHdOfEroJNi
pFxO5P5+rdQpx4hsuVu/aqrMdPVu5I5dajx2YR8Ixq0mCcqv4dPW7cONc39UK7vXyhec1Gvt5CM+
Aimdzt2QICv+lBMKRxn8IcuoGQn2Dy5bMdgaQ0YAHKTWet/VXEZDRfZx4fuzDOus4JumCKNUcASc
VWaGImiGImEXiTZTDh1NZ9lA+laPXsntgS8AQ5rDeNt0XVdiK4bXa7hWsOEZ2GXMhXAPjMobHST3
flpk1Q4Ni48C6BetXfqAT6YTzSJpcxjFG1hLqcVHy5NmTcXVpkwcupz86RAeaV543FyXXXwBrVya
ZIjHsHsicYj+TOlRlbIY7+GooAc8v9yq+1sTyWiDSD7LLaEvTMI64Fel01IXYO0nrKLeQrK20fT4
T9qAgq5e7+E9xG9JDAIwzq8cId8YdUatzBZPqlFr8dVb0bLnMvkHm2BGIYWlc7DBkUFPrVKiTLOb
e1l26yoQbggRZHyG8IbBtfXWG/gg2KvNol4L416KTqWFVzzO6XqO4VIFHgA8oYwed8SVg5BGjCcK
taNBchUPIkj+/xtbVG9HyzdCtAhuv01kKpoLteHkDGgl6kGOcXjJC3pHFBQTFsEWq9k6KUbWCgnZ
0Qy3n+PCTdZSkNV0s/g6pJGWaeh8aUSuUu2A+8ldV/K6qvT5lMy8Xd2+qNs3JbJve8YDk0/mGfVH
endHTwwMH6clZqt2EelBuPhdKBJ6WYG92106CllvBjId4Q6yG+mFJFVvoQdd9o1CYqyTrLCatHjo
bP1cBClkbFwXJw1VIHg2pLXLxcRP/RvbGDmsgo8VoZ9jZS6mAFqWtAoZP6/vxb4gjMk9ZQ1yeIKu
LQjDkovrP2Cogo38vJ6QHWjsV6HFTWtQehFfYXKnwO7I1LjeHKW4hx8xzKnn+v06aKQBCJcPXse+
ZgIiSYf1Ra135ZHZgJy+X8YMEKKTuqqAKysRsR5vtegrCiNxH/Gmk/DqMOJkHv3AwhGk/YfXGEFT
V5+BUwO6yEE0h8VtgjPhz5iEzdd17N1CI5obJHCeh30W4sxChSv26IhW8lxzf5omv3IrGT5hsMc4
H/cgdp/G7xldfBBfzFsJLOFN59IR38kwewSZfv5f2xRFDizRftNND/KlddZoHpHrujosoWH5MDEA
1OfIy+6Pl52k/7ubYEx4mUNBMeR1OQRjQrk0mI7UF4YbGpJw4BRexC2z3p9UI2cFH5nUqYvNjzXP
JloJ7KTunIeShGJK7uAAhYVeNlVzAy3BliKx1x90JCxWXOYGaZRluSfd2S1hSrkwOheWznxUWodY
cbH3ebWOnFdLhYulqbMr4TpTqKwSLa7SqOIiXBGx1ZUlJ5AaClFCxk2+BW6B34PDF5MMBXeLQwvj
Y6aMDwJqWBdSdlbX717zJWaJ82mxAg02x75UCG6BnIq0FUac/Mi/AfP4MOE/LCXuLhCt4ipcKWGv
HM78qrVGpVbdoMRUvpSZrNTY9OvaU2iWQUam5fXKzzlpd+9z3bBBBplqUEdeQUfyRE/u4ZtZSEzo
NHa2M2wAiQu4J9oSLU2/03yin0apwuExwuDZhd5SJylGrXyg61hobqkoMeoTnNwLrty43Kf5BBq0
ifWktAW8mS42+SpMo0WvrAVCy2R+WZCRa6Z+nBbJdgtGVH2oaIEwNj+E7Twef22K5Ey4j20X5Hge
MSRZKVtGX/DeFqAeUmV5hiiR3Wfocx7w59WKKPNRwMAQGmn7z+8ySzNrn3mX0SDH/Pc9vzbV5bOR
FIiBTVYbgKsGGldLz7BkR/eiY8cmFOfWw7x8ycEdn4M5KbU/e3741NzSXApfmoqmHKetUsDargql
u1xZfPeSXT6iPn+ZMhRR6oJbJdZT8aV2/YBj7u2nd/BBgNZO9BwAII804uNjnv5Fetgl4QZ5blLx
4wUfmg2Eiep3HF00dc4JxKVceEBF0f31ojrX/zm8biapYunds+Xk9MxqE7BCe9SE14TX3qLU3dZV
ufe8pxsCrhJ83Vh8GJKHx/7CPHTL3AzAs9gr5Z7LC8sAlY35O5i144E0nvf6plKSjZYFQar6ERVB
t4gdGpNIYvhD+BfJT2Hi9q8eAWLEUSuj7ryPtVqrDRR61gXDLfPIyN7qnG70ucJ+1uR4vorM+0p5
TV40GJQliLkvUiR4QJOCulXuwN2lcoIrIv8pv2oD7B4ctvtFraeIPBSmjGXeH5Z46HI7Qs1yQvne
znTXEODOWiUYeQIj3hEmSTCg3MTzgSX7H2PwZ1Y3lemzoXjfWPrdpYOsrY3avIAq5RRqsp3x4+nA
OA/zT5S1IQgOAmTtmqdseIBpa61l3F6B8mQcNDp2CqSV7XtpfuwGJ6zyG9ILLFtPHs5Q3Krj7ttM
3MbcdpC3Hyhj45BHt8DthR/u7kv96wvEj986idNh1zkxqjSE4/ZyE/mnQkI6WVpDCimqx4Dg6z4X
Ft36UuX2AzkFFCVL9kakiEXG16uywurnM6B5TL6yqFeIdXKVveSCH63b4YMNOovs2DG4eSUmmAGk
zrJ5UuSRyRimueRVBi/++itME1Wpyt2PVYQl9yk70s0Q9NVuNLMGOmiNQ/v2Z1w9MvUoEOZ+pxpe
FdM3yceDc5ZwPaYLKdmnl53XEZLAbRg0tWBkfqgEz4u65BKr04I3+zkc3Gw2RAfNd4NQwRw5CuHy
rWP8s4TcKO+y5o9LXIAUS1EnfQSWpc9OjT4VWFUADSfLJ6VyBGoWjDBFgyW/TzCnNR6Eor3/msk9
Cd4VwFxuav4zPzwbNVztHV8etLXDyGc7u6c5pOlPvkxaSyLLlAQlQX0O/bzTseSYi5El5goAaI2F
msefjZGi5/tkbZHj3TDK1DZXVhe1i+B/bABd8GhmUJ1HvCWKxnTaZR6e6Yt8Oaoo+nPVqgXhznIE
+VKUQ3nblE+XFdBeDft08sR0GGKC6zcX+bsnZRlY+nbfc9XB3WhXnrc7lLuibm/re68bKJj56PPn
wrbmryyAFX76c9Y5/Ih1PtvXBtYPVSRBr+88c6DL17cnbpujSZQQ5fAQ7AmrIoy18jiI2MLF32OY
EsRqdUZHODss2S8gAPgWgCnuKekkkgCI0ybX1FFAAaI6prgpXeTVtmUL1RNsrYA8lflrk8+hIIfs
bJaEGbIs7NvMtsDfoiIaQ9xcdH6k1hEoVglVrkOtMGGdjXJRl7D7SM1zOM7g/hPPNMSMQNEaBcBl
AJYaftPuWSjVaA+aBW8eljV5AP0vQAQTbbR7eQIEno6NIhd7cTU55/qiuoYkgM7C5WoqriHOXYsv
7Mf7bGrs6/6DijeQXY5xSNVN5dhXHTdlIiDA+SqY7QT145ym7jkeUNeND/bc5naKPrYs0yNfDsiG
CJjPGfRHKbGxx5PvipJjdU+Hqnt7n6IwtpSKQHM6Y6kpJ0jtQPMvcBRzjkHsKRpCmBS08wbEwAGa
l7quSxqvP3x64iHypHedMTqjKXBP5aFEcCP6JWfyNlK3xTAmtwcAscKuETwKL3cXYSW4sG8KKTk6
xZO9434bPKpCgMEhUi7ElHogoDexhsLA3UJt1keL/c7oONa4IY0pZ5DwgyeQRgnyUjiVLbfnRJeA
Co3H+kzAkVZgGi5ZEZpvJOr6B8fWi8f8AZ4OKzevVDnTiEPtAmVDzVd8OzLAcBa1a1DGId1R8MKm
CjGorJUKVUFI2N/bfJa/pCNY1NCZ3xDz4UAQ1CMX5sZHg9BhZZTp8MB28+LAwRzX60CcgHGCopap
n9sL3BF8T3Wn2OrupC9sKtwLEJuk/jT3QFlqtg88lkrJCcsw3x9p3Jte7qNXD2bnR8WBIkVqB9/r
UZJJDpuBXCnKS2QUzxX6f0NuqcikK7qzTp++3Wad/enXaFrdKa3kHBy8Dgmi7L6KG58eSi+WfaL0
k4gA4UsN0H4EI4KGiqLs19K8wePfVCV44qerVq/+5cK1KoPMDcGjzSx5yMQC5eFKKxg9scbMLfKh
PlFxuAUa26zm3lsWHnGRZXvYblRDyL+B3852tyBiFJAUk8DFgbhkzYObPegP4q2Srv3yNFhHDOp9
L9CZAZCKslpfvBmiyIhmdD0+xrmEv3Sht1d2t+LQQkFY7qoxrPoYz+prqvMQi8KJy9cAbH65bota
MC2cW2/nUIniWyLcRcxNxpV5EVR0f6/ywZkkcynNkGsqp4ePwVV5INu1MShlTBgl5mjx6eynejx9
mHIKFneIgSzds4eS69XrBqg+k68BdA4sEh1/jbQsCXYZCglK1nlQ2ekuPReRK5PdcogyyhuJy6X5
n5XcOJ6JAtzLVV4zg3qjMOOP5HVLola5B55qdfb25rdESmAgZUGh0hjC9tuLOFRh2x0zg6rR9lkT
ygeigzEsJSCXSB6vEUO2ZbY4WgBmS6VdhFyp+4J5jR3+WOdmUkOOzxWtzE1fI7XS+YjNaN7tuh2a
bwktneKgcNipkgpTq2D2O8UBtLKqZ8PuY8Nh8xC2mb6OLaaDdA5L/LwUpYlMzNe98m+JmHHxswBl
4mdN4CZYGIzgmGnzNKAPPLTvx1+tmy0+BW+U4/NtMFtEQELDF0hRobkEUHDd4AfQ4dwC7C/EOxMb
6oCOtXnas1EA5zvlChtnFkiyy1oL5iU6bctJAfSvfATuebnR5L94EMLSzGUZ+G+fu3tSuckFq0yD
q6YEW4DyZ3sHr2Oxw/Bx1yt5G1YGPmes2vEc5wsimUkxpi+3AWs2Bebg825gBRv12xmy1GDNQUWa
E+xnhHVuW29z+zwcCj91+XPu5g2Q2yFCTibpvzDsElVNKeJHdtj4W2p0IBt9sQsJ6RTLfbwPNP9K
a+JQ8o/fBqiSYpfW1GWA62CDIy/hFxu9PMbeeE3F/ogpgYRWVgEpE8EmZyxn1MWvX9an+fOc2z6w
+tsH3YEsKyAiXdtJsdImSTw/sEn2Ea0B5tY0EAB4p9Hp2HRbQ59DT3ngpR49ig+od43PMVZSlZNO
c+2849CRsG/BAPapjQ6pK06NJKkDfk8piyH+6IExVu8cqC2QjWzLTELjLiT7lmjkJAkKKMRMFYTa
FnuweDT+UZhNb/jsFTarRvEbjOqnU799nJiRQi7XKke1YNGlu9onGHCzSZIP/GwCPDy0o8kwupv+
l+/ZJhgAcFQt7BA2KqcIjjTxQ+TZunWtM3qHTEuK61+Wx6E32YpU4oqrXz+lVETr94cSK7qB/ibg
65iYbXrqHL1ImHyYkRvwCFVMnC9GTGIN3rPnVY+WLwMXQXMXVU5msxrROQLYsX1jUkGKX3bM+sab
F3BrIWaDa/z8p7crlx9ienQj8aq6VHXGwUy5Ckh1O55b0O4M81xnxyCk+PYDb81gxmDsy6xWhaxp
z3O/2uKS2e1UFBPtcSfynZFPfcnbCbf0x0MUc8LKROhcw3zMrwVgy4JsNyeZX587Os5lUFmE1RzM
/aRpFmdXzABwAAzSadPJtvBoB7G+OviPMNdiKb+SmKEUFwWq3NnocOwRL3U2i5tyYqXS6urs4iO8
AHiKZnsIYCleP2xNVfbCdoT4+XRzkO+KM8MYhfmbgIdI/S/AvpehwRf2es4PMIy9tgsFNtbN1Cn/
E/5UfL2ljqWNYEU+Na7oMzeFOYynpnD1VAB9aG69phf7411WacUdVoimEK+aQfMfjjzKZetm21lo
E1lKuFPkYitj8lu9No2WzZuU8RlQZlboWVO8B5gFWL3YW7cart6dID/r4/0Lp39jiRpVl/JmxbeF
7iNkPaiqeTSNLT8IpgSYfjqp+UPeksqDcppS27cAavq4mk9uhnFzhMo7CKImdehMtt8XG8TDP/5+
H7HCuX0Ogr9kS8Yb0OV6r2H1Q7T0LnXNHhfI/ltVPSSnLrmeL8MhJaRKJphf/Gjrpch/bk5ROQfC
DMTYEnytj6Eol2LPkFw8bUWQitD+XCC35jYjQzYfThz/omKPV4RKjX54IaxrXbFD27qCo1cHhQbj
Jx03wmcFk7rceqvBI/AH1CES08nCTzcaKEJkTw0WjQb2Bvp2T+rZnbzcMPN7aVnvRSsMpKmYk2Oe
YN60JWBcnC4+cXVBjJI/SznqyTep2LOxfDOAIepjUK0nVP4SpR5p+NmDNVJOLHoDb55LorWxcBN+
IDSvh9EwyIiAi0Bb/gAV+iHJyGykdN0EfhTueU+DRPELsG6ppApZ8u0L3AZ72QQ/8wOVrJ2kjaJB
Wef2pKpm9qsCeAAnhI1MPacFkrgNNtTzuct+LXi5PEWI3Sgr6gd5iF8aG+xhSr3xDBW9nIJmwcGe
K6oebrAzZaYICC+z2T8rICiLxAJksg+Bn44ihB4swyNi9Mxwmlwdew9SgP9YqpltEDLOGEhVrnJ1
WXytc2LlovXnY7TCQyw3cHSB252oNhwQYcsBFPSBinOOFncYql+EQZqv2IBx2be9OHD2OMYyvl+7
9fXTQ4s5CQhevLBwf/FYCD/w2QfjQbATHxkzr/tpRT5bBq+t0ggraxO0zzkQCR8FwMB6xKhk19Ye
VtMZ2H/R80kGIFBtD/YbkVTK9HDVQ5MW8W7cDb+o9hiTzQeYnEb+AvDOyq2YVgpZIsBT1YYGQmdA
1Pj+t5UELkN9R7a3AUoqlNDfO++xsTjvta1epIekwi/Sz4HeZHuBbFDl939uQNQ9hOIi+1YmJSDm
O4zYTeI3mhIiuqeBnbejN6YGE+yrN1btydBXEVufvWUIfUlolSUFYKYiudky4i2vveQHQ+RPdNO8
9zkXHbCdPC10JJzI6amhQt8xhw82+UUAdZK4QfSri4x0nVK0VABo60DXUMOMjv4IQ7oASD1UU1Mm
AIPGnuRkX35ucbxqFxCZ9EIvDHAR1E1eUEHPvGVn4qbRsat4Vc3EqDsmwVd+JbNN6kJUUDpxPcnI
QTT4oQ/ys2Gsd78fYuBuPUePaQkNdWXc2eTonZcpUKyIAWhbWN46WhohHf9PR1hZv9I2oyZ7REmb
qSXQqqSn9HgEd3gFiK4jhcyfAkNc2IkKlPPnEI8a+OLm0MZFatToNpVGz7QSevL3Sy71HxX/70UC
mby3iFNVhSErXj22oLfZIPIN+M6+dq04UgWDYMdlHfPPnbb29Jh69efWS3dBslgUgdKJLI7G7Zrh
h4HWGLXgakLvOnLbYr6e69HPVMSHNgf4RfXchA3dn5YfmUc06fQGlMkMH1Qc3oZSkbNLbdudF5JJ
rizefm3ojkMN1uy5Q3N1VfQGMGYC59SfP15bC4TA4+uajSi2aYtVrbEjxDl65DmP6UqXlSTla8n+
gAjiSQT5WCw/UfqSarSBfqNiPPDJMrsA2rlF9eJ/PTU3NVBncbUKhbYFjQFsORJfxR5Dm9qGk4AA
mMnkKfIUIamPdh0eFKgd7QyNRQaapmrz59dlR+qsOZlN8JX34Oeq4+7sT4QKnA9S9DSEkXpNCZVz
pUnhNVfiTOIaUrSSNcOtosg2jBtlXMVU33dOdaU7EDy34hp30B9TKnAalpreRh4BrrPTUNCgKpQW
Rq4Dm70vOn2K1En3tqPGXgox5kNezDkMnKhl1qzcEiA+925j3Jf54VNgQgpTEapRAJPFlS1btnbg
EGz71Swj54QGkhvusC0T8uKdaBvqeAPeACqdE2lrXHWnxrQ1kHk6kwCBG5TPf+TkHTX+DDwpB8b+
JpobDlc/TvbDjVbN5C+oKUeS9y0rkrI6zyKR0XvDPN19faSzDxvttE6i+jZrhQdA6oPJ/x4FAVYD
QssptGgnYT3os2dSL14KW2sksMcY3spA8v1vUDKtNV3SBpn7UN2d6B0qFeJGIzqj4UCUJ7RAsF+N
0ekwUgWOVUmCpA7aU9S2SUqZCQsMMpI0V413DzG+pssE55YTM0VejR/bMk7wgUOPMiSReVb4uXPy
3TvWERPQCYXjjju5GVgm64JvTzaaImTbqYaST9FAIEYC5DKI6EGlOENNwoorSeFYnnZCHFqD/8Dh
rTMRbHTf9lj2kWmfcMAQgAUVEiPz2eE57vla9eLjSQNCLIsXrZajoH6+ZyhKMSGgMiFOawEIGBzS
MO8io/U8KNAXDXDo6x77fkXiBxmmn7fIwlMdCRhIXOFKhV1aoh2zvkXN51qhwa2OD22Sn1B4/Zjo
5WVfO4UDdbzSmaIDlADpul37a0Usp8tV68WorGo3Q9qxdmEF9Cfvv44q9q8YJkT64mk0S0aS8pc9
g5AU7a6VARtDmvpNjXICvdFftXMZyJJnHZVkyULAL/tl5CA/PcogXXka6q0nPvnaTd0OFmnnpzeZ
IU1O2ADfFEdezosbMuSvAyeTR+DGfG1pAkGG4xh+Dg6uLbVcVXIjxQP4NhujFXqpXZhe3xd4eUTq
zUoOzJ1Mi+5ny3TqUSc5Y8utzcnSJi5x18FMPz3NsFE/tVwgYy07gfZclaTMTVRatk02m+DZ57t+
8Z9iY2MG6bN/ViKIGRJLHiM7caf8bXIqumyqz/ZFpOSuRyVdfNO7iPJrGWrZfAn/fX58mettFvKj
0fTCI7bK9qQnAM+eMzIxXYNS2ILyOu8OPVvqdsFnIGTHqyM8iVK3TwSHJH9tw33zWIMVK7jK7rLI
kH+OayN9S31t17Sbs6lxIolKiXNNVfup+Cvxdn9nuHWDmeH7dQVpRZWdTHH2GfNW7sflt5l+C1Un
4j560ib/xAU2Gv/PbidUVidQqGZpF3BZrQxq7PrXhABClTDIAyD/sNBRmrZQ3+TG5ddWeWDwUwPZ
RPC8cU+DoPDlFCWUSfsSjiPHDdxWiaFGHMjDLfP0jiwyt5v07wzWOXPBWI89uTCzQqRB6YOa1CCI
siG8ez5sVDpZ7pE6s5FSlrJIJlVAXZu722aLH27x+lybO/BkqnemUbNioWcH3ob8FDS5aYa2NiPo
UydNRoA78QEFdKKMQRDn0N8lzaEBffLyOWsiF/1feQrt1D4DzP3eCd48/4pRgaoRssyyKOEJD602
QwXb5mGcPgp2MrkTmp8jZYnWo4XTf4Q/RhajPfPZeb5dtN2l5+SCV5+hstiIRXTsZL1ueoW4L5bZ
p0AbUyg93sCVH4A8wbN/LkOWxDtExAqlRAf/YO2M6Ogn4kxrMx8+y1uolwVtHRJ6KHU7Q86fQ03e
HNxedZkCTkIMXy2j/uucIFgZlI4nQZSK+4YssmBDKNroUbip1/ANOk5CkONsoWcuPDv+bHT5Id0c
sZ0J95R/WziHLTjnjIqMF9qcvfiYJaRACp7/y0/4iCIGfJa0P4FO0cBgrI6LKHByPicBBCWeDQHO
Yds+XxH8eNFpPsTmgLxK7fIAi6BxLjtuLLiwaiqL9SUBPqQdDfnZci41A+mWKl/PEToAG+S+ktDk
82YhG4IPTTBrc13Hr6siKGYh8Y6BP9/xaKNF3XXoFlYAFi+FVhV/x6pd/hgqRnc/P/kehMTFHLKf
rzGTbnqN93jcDhFsCJhXut52IcM9XCfOMe/xIeWmJ6KSMESTICbiNyLboO6u0g8F2KzuamDXAXR2
SAIigpXAlb23FD6/ES8lNjgfHoJTOU7SiLKrob5o+knsUFelbBQ3cBaCc8JKXsVo/tsbL2ixR1Pf
ejtOK9EgrPHkN5mB7CNRKE/fPdT4V/KUASaZVYXt5zy8tCk1LX292lw7zzVeizIu7hbi/Ivdw1T5
c2qUnT2wQdjwn2K7Hy+tE0HSg/4P0ByglAFRJSaLcQRpZGb97Y0sBKuCKINbidk+E2/80zJvypuC
12xKi25MQHZTUUyux7L0vyjt3alposoMt/+pv2f711fbxs0bSil9xWCIu6Qn+KInjXKw9GXwLguT
jfeAoQdYmBPdWWv5TG0LinD6DTZmlbVyFEAXonK/fPL5OO+tiJFMLl0IFLOAIQAcqoBBnK7OPOce
yko4jn5GMawnIwm6J9Rzq5nVzfMD8CaMpHzhjsA5ncHrdlKO4xesq78anqECUJMeh6NwtsOUocI4
Qbhuvdvjd80CRDUKlNNKx4kbnGKm/9Jgo24Tl4zskMYViSbv+BhBv9WNF6z11gbsemgFERmkULXk
FRUJX1VDknFYLpJlkTsUYMbKPAlI+iDv55sVZQiHvXOwM3kU1rLwlJb451GHNN4pZgtpdaACIBAG
05eSfnNGbnND1SQhq6aZld0CaWgoQyPKgnslw7RNg7yVIx2chNdiyrBsJMIlKueNxhrxM9DSce4a
6/oWScP9bQxCWbrrHXIS5IiersmjQBLgjbH+kNYvsPtcev8oXR9dytpUonEUHu6n+kknwTYQdw3E
GRLgPDpwkwXj3uGGyuEWNobwNFir0F3+ffrWiBjaXOA94eSAubE8ZWfWBScbRHqnun7VnDRwbJ/y
r4qkA0+sf6gCIg/BaHAwzFCdRRwetuNA3OCdUOarjp/ZLoxpX0wkIpASz10+SzpJTH7r6bXTVGxU
s10agKwE2TEVXhlIIrCqcBCuPsISYmPfUtgFnDAU7wEBNgTKfE+0XLRJ1vf1UQSAoeKc1KdvfFzW
2vppHJn0HRw/CNbURzm5Ci/YbVpLn+DS/wB5A7f5JBhe5x7BWicrPDh1Ehm0Kle48jtb9yVU4U2I
zqeNnKwXeRe/VNdZmi+DtscKQrYTLYVBOyjFnDhwcctqx5wEyNdDyIJxLX+GgHuXvrg5jIWEv/fb
g3Ye5gJI+ZdkXhOttdCoss6fbl0AmDQX405VsdTw+AHgfVmZNj547NM++Njs1MEbKvxCv5bz7Q/U
TmKIHgGeYkc/m6Ijad+O/p+muxWpknLHG5fQiSr5CvXB5F/DaS6sftc8tholQuDwPm2Ir8MVTpop
65SE7e61VCWEkpZuqeDjDQ5cFynePZQ4wcgrUPBu2hAisIJmmomZYrc4ENEeGxwSW5TwSW6naXMc
hFbpo007YLJ9f88pplvCJTTfPfAjOK6wle1+G//1c6HVcgyVxiZtQDHrELb/0sX1sCNwTSJZw9Cr
9h7tusjmPUOR0oxaBUNL4FkwLGSTz29M4AF1shtZNzMltFDosB3fs1rKMUBV/ZuplbK+lmx1x8EB
iJ6C+RkwUREMcLhtAgyROvsZA3nJ0+AFjPngY6gd0MZRLrf++lypd3xxVHTqPBgEW5fmHsdEHVvh
L3GNb91RdlXNvVxOcXhi5OjkCpdbTakUSej/1B/rnxagKiM0XePYw2m3HOs4MPqGH6zuy7AG2BbZ
kEbABS/wZtNcJhIDMsJCWVF9j5xOimUoYmcgj88on+hotWiFWazm595kkuXQbDbqrxWXVuaq6yiU
D8rrSi3u/0gI9nD9EAhVojdrpS0g3ZWJVudR3G2xGkFHpHqSMoC/li0P96IZmy8SdlgCFgr6O88e
GTGYLnwnzeje8r0gQ+C2DP2cBUoeSgmM8FB/y96FMXmT46UCmV6kbuAj3rBIX8iFoseqvgR0Endt
66xr5vsJa17zCle5ulQUonRmgwQNRGWRfrEJBfZFMc1NBwG4RfiguKeTKlJdHyWVHx0Xa4Uen548
dinctVA2DK2UyNRQzZFqKO2Oj/zIWSczgxlE/RyycSQSSI1dv57XQ2io39zi6q5oNaRbTBhgye0V
zbV6Ai1/8zX1T4N064bj1/XE89zmOYsxPvPNeBCGnyXZtLAkl9Ol3FkQjuGsL3K3sMDyfQ+prWdN
10iPHs5NkEsssLQ7fLFeakeF7gECEm2wScWIylqyvL8Fie708d+yuukJGAja9NHLN1IcfjYffntp
W03tqYPEA3AsXwgzQc0jJnVV/HgaXBQKgbzajc0xtDfijffuitrr09rMCX0Qko20cIJoeJWf4SCE
GfTQ49/yOnZUzuJMMLwkB0+/ZWBSpIc6UvChUWukfvb9vnkU6vwPF8CixtbEX7KqqNhgvnpKUpMF
zmcH5vSArotPivRh2cU12ExnX2q3dV64V/yRo4Yf8LPcDcVn1Zb4YnPehXiZpPSO5UGAyx+uDOfj
Lym3uNDIB3u006LSlleq7WhmewibFSVrkyPzcIEf9abijhGXZ8dMhIDYjRcoASVm8sh//UMgqHlu
bkt0v/NwBRDxqnfd6vkbo4AU9Ecv3eU9oP2zMdG0HdyxwSdUyMC4tKa0/nVAHRGurEA4C4dz03ok
nNgaAtkhmJ/qdpWiTnZocPDCW/4pYNR1JV1AFyqLd2AepTDab63zRzJ4CmXhRpI/cAX5rg5tV+me
AJUJxPxlGDRPl0ieTWtLFhSZ/zFcYeGEDaFyKnBLuFE9+4diWyk+LsXrKvL7JhTjAmngVLS8Vxzb
nzpRSM9u9cYQUXv5QKSNcF6NLM4STaMEAJpolL3Zh42VCgkFC1FGshz5Y0taDOKZPDtxjscgXK1i
QkgnYbnPllGjOnVBHerS2AOkCBBI/mEso4vnL3DyJhjC0d311KuMJ9eJCu9RVdbJ5t6zeSEmlsrm
tpva814KL2wyO60smvf04biDbmjm4fPT/DhaXrB7EudR9skiIzOAKbMEDXSqQIJmomeQKFjxaekK
/F/CDBpxqKZZbBwPViL0/eiVA3Lwxvu79BLCKR+7exC60FCMu0LoSGRbCfME0Qi2Woxdziy3FULQ
ujG1X5vwmLzo+zHKqH5BM4UpPxk6URroQiB1HZJL4FyNyPcNCnvjG/lFFFppF9H2W9gTByiOalzj
qG+qDI6gaDkfaW9TrUreob6JvHQGefse4MuaR1i1xIAsh9DTXorYJZ4Bxda7MQqcPfh1cYjP+CgD
yrtbespeS3mznZ3xQt9IDPIIJTSM7S+EjKs7ozhhi869yqDuQqR3G0oWo8v0W7On1XGWOv88tRur
c0F+6hZw+abZJiFTfasJ16mqQco8ggaqvJ+68GEjjJE1pAsUBI9+tkN2dvHvLhROguTrfosLh4/B
rQ2k66O2UqtDvKtkPs455Ccxs7lKgb07x5EuC6Dg9PNTgf9C/imyApNFzcQRklnJsKWwB/Vx1Lnx
H9iGN8iYfD1nd9eRjkcrjS7TS2iUckqoiAJYumXkyxmnjiXdbx5Ak6wS1G1Run83JNJVozrLQcj+
+tIpvl737Up7VAyG0gCb6FIGi7RVeK3/FO07jztgfHupju1XMPnlGLz0RrP3hV8FIsqUbbiTUEN7
d2YKTTgSk/+x8oEJBhlnkmKxxe4ocbruc4aC2PkeFtDw5XIcXKo36hIwzYDYn1v3XdcsPjzxfhZb
5GfRSLRX1T99qPDMBBZUPKJ9BqteIzRtlgRJS0k9KE2aPaYl1IX6xK14ZX0aduWW3RCdEd4L7brM
XwyC5N82OfQS21WoXeYgb5A/Ell2vJW4rrQjimpBLq+z8tUh6xAEozxqrNSgHUBC39CQBk0WfHUc
Q1pOdSw9EpgygBfVR0CmHG5FCXI1mtR4zCoU9vkveo4K1VR0srP5jtR7xPyoKgdW0gk2p0/cz1MY
EWt9OL+5lpw46HzeXGCv2RQ/c2YGy3eukQoLESroUgMvz8Mg7GJkVtYys5wahE3ynV7/EEBNtoKk
xe5opJKSJ5DOzRedkg58of2lHhYfVS4aEUoOvQRvqe2rS8x/QnK33idCFyd4haFPASc8pQUbbKRJ
geXqeaMYDcIHQMiJQvTwvrnfVC12K6zSMcWweJhviFntKF+7EjbavQO8eN/A3JwoJby3NW/9JNRg
DDVAaOOxW185l44X+/dA7/FFCSzk+FuvSH6WvbxsSdl6r265SbSnJ590/oUOThQZu4YT6Jh2FPAq
fIhByC4nr9YugkEHlbS92pTWqeZK0aDdHvQpZf66HxfweKrsUuFFPOyHKjq9rTWDhY75SGIjjHHi
Deno6l8mk0Kzf8dRDjInGw+PZb0Eb5puNC60nNdgSnTyCIe+sdMSk0cOyNDB6C1NXPosqiM6mKsU
fZz/2iCUO9qI36A3MuaR3EqyOIJZvqCwlk92cfKi5/2+/6nzV14Q6mrzW1O+gVzLcN3iit+PQKS5
MmYDUVdRUkmafYgwjnz4TC3ww9nXvgkbLl+9wq64zH44jQOO6J3Bjz8cUrdubq2H3pYwnhdNhNDL
rNED6/kFKqB583m85W0tLgwc75rNx23CHlI5wBQoqpF8LZbBxGQtKmlDFRtTCZrtY15IV4GxYrKD
ZMicuP77vEYmkjJ096lSKPZARGSCd18pq1Xn01jgmFy9g2BLPWzG/ZQht9IzjwYzB7pkPdX5SLMw
oNvM16yyjkwe20BO8KFXHtEPz3KEZCz57KD/TbcAMBGXiUmBVeplCHihey4uRaOrBX8dDl7run1U
kEz54gPbOBIITtPzAyiI4hO5TAy1kNEU+7MIxV5DNBuFctkyN0P+8f6tGMv+Vq02Ah22vRj2KANN
nEzx8vOmmD0CA1KkB5doHlj3zIld4eCodV4XwPtClpn/IbgAU2yjMX5QigIzKfcMrK4G69+M3Qg8
pLyzYMEAcWQGHngRibCRJTV36HRYCeYKrGEIn83mhrM5i5cKzJBnPy5vJAoyHU/IoM2DxD61RZnT
EDm4nkJQkDbImTk2SbyHYYVW6bOTS2cyHz47kes5h9b+AE1HBOTR0fN/Ba3UighGQJittB4CTzX8
s+c4Lg+erNFiHSCrcWh/WQNnbYbPgS7dHvWE/wE0x1GvkUIkKO96ZAMnSRQ57N+YoOZFzz2wHGRD
C1ngIQlG03MDV1gBXt4Pi+jnxD/9iOydx8diy/wJzMbPWcvQCkt3yntDFMHnoMpgjorQEvxk4rFM
42VDH9XZo7Gx5YPae55g1a6wo7wf64GE4lmFCpqmOvVmLp+hLqVtmjDgeDQoIbYzWZ27z4O0JvXA
hdxAd1Sf4CerotKTCI99cErFIDH7JJ0uqSlC/Z6LdPF9gNd3EIXopVjPXwJvT4GPxBKTgCX2qpw5
PNlIg/PXdAGX+gUNEDPUEO6z8oIBKmHwDto9laEFhff2V/WcDKtk9Ag/DS4/i/f+xEj0vfABJs2x
rnGe4gWCkemQQK7V+1AdS4LJvRbPP3pa/UxP4+Yrqxj2sm7UMSfmgYbjArQuME0ue/IZf8xIRFlZ
JGk5TFQ0XT8wT1kGMl+yF0dP5pj1lJz802EEvfiOHFcbmNfL7+a5KC7PC4AVdAWKy23ZYeKIsYew
nA+vEMntGLG2OkX4a9qMbAeVzoizOT5lKLHTSXUCkehhtiSURcjVvuTmHbNH3FpWImhOubvIKnXC
4wsZpPB5ANW3KFw7x12mP14F0kmx+Tkk/sgp2bFj46CcROPmu+LFY/eH6EeZUBz59F93Puo6YzuW
I3aQTD1Qrtiy2Da4IuyI7ZCAI7L2VcemPPenSZUzKiweJLgtaGO8TjzLk9hq+2bba77T3sTa2hdU
VbMoTYliVOwGBTO1t7XZRIIkDgtMFami3iJ7w6MbTt7E/E1bkK+tHJDD61hKDUf2arQ9wlaUkqzd
NFBUMzYG+pfVcAgTq7Oy0h016vHHJcnyGjFYdsViVGmalO9IX0ez3jzfpGs5JE3XmdjiqWH8kO0b
mC4AtbIJusSUCtJ3Yl3PfM3erwsdCva2Ol8Sywm8XDzvPNRPYj68lRTXjRxNbRU+eEM6NQLQVsiH
vpF8MhmEffEw82PZE5J+yqnnNpQ+yyFs2l7ytzZqExr31elGGdf3nnxyVzmqduQTDEwHpEpnTmNV
QVBJObRC1oQA+wNYpFimyaj36Ru+e25k8iqzXPw3XBUeT0YKnjYBwwDYFsHiaAS90Z0dmx1xo3uU
APkLqm+5uONhrBlHV1dkyqlSlP90WTk1EtxoACZuK+GUGToneUPjEHqeIsiU4Vj15+vtRkF+YPJ3
Qo3tEdzg+Be1BXp/Pyl6KQqRLd/K0Q8lERB15jD7qLyebrHOdDezQ1iGQ+7FUEl/paJ6zdA6pies
X27SZU2scJLDdmDGzPOo82Ryvndafu3QhJbdmyMAu14BgE8rTD8hoOcEvceeSZnrd1jwyHFBsscK
NNTOEl7Yv1Uujj6DJwMf2104Fi8bsbzcd4HTHCqRsMUG2CSuIngea95aL5NCp5ak27umlEcYqGDg
CPexEW3SipqhTvqERg85LepYklUTu/hJgeCUHj+kr0ttrDdC2UGyjH4ZT+t2ouUCLhLcFeL/BCz/
3btJIoudSFdz3pDezBAPiQfNxwa3HyXJmy6Qe82u3vziAs24/5nDxnZch6N+j4KXq46lHvxpSka2
V3YaIXXLLh7CXZ68Bdbyka+pw9eFz0SSgTPxHoAGlQ/ucAMYYewoQsy5rwx2S01GFHaWCxgcZzyD
OpHLekbe0Mfm5lK4C7lO+hSew5FqGn2xwsg+lWBj2ljhfEHD10HUJv96YCO8jpI6T2FQ6CWeu3Qb
RbEbS6QYVvfD84SxoWVAowGEp3qYW4Dl8zocCa9nLtWGvN3CUcq5NlPoGJbcWofONkPyrid0ZfFk
gH0PKRbi8dFsW8funsiNAnNxF1Deu+mmDR8IogkjpvqQ8kiDxNr69NYgzGeEmkGE9d0Nn6bk4ngo
5WHAKBX97fVfkNIwhpKZCaMHJPV0Ld+nHwTxi/BH3GE7JPTg5/8XbY2xPxRZRVLP1hPBHKPT/9NP
s76bavPtimrPm6INN0fNSfd2Qn74KhtFkNy3x/djjNVHIjpsxm3qd/4UoyT63EmITo4lUe+XCe9C
sOcxQgW9nOn+xzTGhiEsxdXwidcmL9QXY8GuNDqYhpGJgb+QDh8WZ0Mw/JPc16n5UgTXihI4Or+3
128mK1d+6YHBepJrylxY3EHWswZiOBzE1kuj0EmIZ5Unp8aSB8Vm1iLB5HbAKeqvgHOX+lF6eNKd
PdYcyLxRBle51PMrf3QPYP661QDpTOlxrHjreniUY2yVtlQNE1NGhbSwTgq+N5PLlURC+0Y04IzL
gmwf3oVgnkHZ3dg600DXuniPctXuMp9igTkgvVd1ACsZOaeioN8aQud4Us3kRpusGyRUstrGbQf9
5TXjRWQ+r9rEoSAlKvanXWoLNc9IzKWYosKCjQVfAApe7BY8EsZf2EsamPNcnH6M+DbcZrbbAQF1
4gJujGBy5n6RpqgRxP1NVc49lrVduvQcCR9h3/38/+VaKimiywaykItGNwP1g+hLBxq9vQmozgtx
YkaoLCLopHNASnTVdeLS0MNdroUbA1PBntKe/IvRt5gkuIX0gVaNaem8qD6555Xjf5M95IUXepKJ
LwFBYn6Gv41D+N7h0+4w6LUJpiaDQxMYzVD+QzBx3v45zASkwYY/c2NKcXzgXZE05suKjZsht1Pg
eeK00nB6pquu82+8/pLTxDym4L6n8oYs1tVc0uIZOorJHVz/7oWs0mQIRKR9eumEcMb6XrGC4/Lv
7f5Bol4z/ryOt4SKZYxZBRQsxObnw2ZF9gpT3v8Q+NJ+JqNZeevCjklX9xhM6u8FmhJaXgaewJVG
lpg1XEQQq127jr5iakS1N3tlT821D30AMVv3vWeJGWDzga8LrlUHrh+HVAZ8gLgipYN98nKsmNBh
rVSUeHFl+zdpyki7k1eRKIBafox6H8s77zEZ4S7lc/48kMm8VesPeDKzimBl/tQx0bTJfJE/MpU9
lkrX3I5eu+CwqhzkJPDdpcg05iGWGkl2MI8oIvAjUZ4Wrm9gVXtxV2QrVpxZpjonlCVdmznUVXMW
KeiHWRxwcBtbF+f7Z9wzjsjWax6fuR0gual6MSqA8s7wHHX6B7ulrmmkoKH2FFK//rPbEbMQRFzz
3LHMYE0ygr7Mmt3/GHo2kDPB0tZQpMPTYjz2ezMu4ubdqqZ6tESQ5XkTzro9Fm5e36kbn7lBSxv3
1F+iSueI5yKbRfiD9l0qAns1sjsVOrO6ljmYi9KoWkyfRCi0X94pD3CLLR7/AmXvUxlOs6yfqlAi
9KRuJ3EMgdWIfeLgw/u9ITDTem5sjRYr/Ej7EkHOaez4V5/GnwB95NBh1TVd0HmzmjXggyEkOqZw
+InVkfhkC/BvHJnwOA6pxiMVcuS0Og9ReLyJUhwVyiwizh/7fmCkT0M5lcICU2Zewtqjnk+uMWDZ
zd9pUlBm7oYstxb/k2yvzdlBF3swpseFwawCmDzWWTCvTXVf+LueLc1ryokAOUvkOkfLVrmkoj8v
2boMxeN5kNTbgnArhnkNXV6LPZKAmp+3ZkYGtH2hv4TSSLUHegKNLxbt1Qd8w51i/EydVLzFF+zo
q9TXF3uLF7NHDjRFIQciEQK+EEaFmTiCegc6MCBA4n7S4aEZpGqstzTwr6ohe/+LZz6EYpNbal83
7qWMBzryTMYYvB/qSr5lVMzYioOTaj9Sc5Jz7+iYayiBSGOHqaurOLLpMeMLDFvFL9AZxEe1psnG
AjpJdZ4izRArzGYcHqFLIzNpHoLJVXOdF69HUTGCDnW+tjsdkh7fRQ/+EiJcDs8/PjUQ5zUe8Izw
3LzLS/y39UG1cZqZRlWflvqzD6GNKAFKGU3l6UcO8XNwsq35BM4d/RAOsEsB2ShUgBCSOHzdv+1A
VsWmy6jaiNdQOPJUg5mSMTULBLqyPwq3F2P4qe1zCUNQK1t4mGbs/9L8ZAcmzgIaCxlEp2QsOGjX
DCWF/ldRn8LgP2EA0+LSSxygqzktf7u6+9wG2wkerK4TkfZ00jKziAPuoXNquAf2FxnBYQfnRleU
xDSfXG4MN5dcyeYXNH7mNKBEHXsMwhu3PdHaN2p5xGQrSr7cRGnTLFLFiaSnlC9+KxniUQY9Qy+M
o8thAi6uQxCeCPscNHj2bbJIEI5UJrjDV3nv/wauUgxd4pCyvRG6qghHvcMXjf3P4sdeVaAFXYVs
k6dRAHtM2wyUxCF4LuwJlv9YLVV0qZWUpNtOlipkLS1iKjWFboQSS4gzDELOvFMHTTGhbaQXxnGp
bsWtgU1ceA9BWVYjBR0ZXr+bfJ2fz0K1Aujh3D/jSsRxswJNkyvaHX1/x2O361byN/1Iq4HkoL/H
1ZqkL9hwzu38/q6OrD3vWrOZ23ZqnkncooTBESObJ4yUs7VISu+Vppq08eqGOs/PPY7UYzVUFHHz
MT9pvfhV3NlraKXh05JL4zb/a454R6iNzURrsRX5VrSN239k44wm02b12D6p40VVv3ORsd4sZm0J
X4SQKsZNhCaiCqq+cZAqXEHY3tAi9+qe61VCGBpSHM7NIvx9scd9oFoXokQebsEq0GJcrayDJhQn
4JW+ompDZ28RgRpr1UJyULtXqrI220LHRQNthVh+rFX5S6ds90Int6Q/aXFkgMiS610kUpes9n3C
EygnCTSuZRvkwGUEpMCBDq1QV+7pdSVGbmsFp49DXKioi4mSO83MYVpEZLnQxziHLyFDrWxIWezc
kGNEgBLMDlv3tWngCmdhyILFHoowhR/II1xOTsKy2Pifq3yPbdopleXicoqKDXBfe4J3mj1WTL36
uBNiKTSISkyqoE7goddVc8Zlomhxu/YKpKqLetT4PRNBrxAC011v3qWxathcmJBvlzV/b1ySY4Xc
TI9vVKEoi41ROg+4rhbMdfOPP90J1Jq0PZjkYQbD6JMi9HKhAq8QZl1AwstbL76NxFxlJ3/mb6a3
iomET3wvZ5/FjwUV11lkPQFw2sirwJa3S2HAKFoSWf3g2T4KHI8L068OSBFT1Ho5eMcqG+sVtyQq
QiAKINUB7crdI6Fr+MQupCKR2Fe60L6TJ5WwZ8Jx+uMqpuPRfdd7BRMku/iOmN7ZqNY4TbCJrD+/
uAFCXCBGoQvNpfo/y66bc3TyOtWAsDPDTP35mxF/JtVLI8pd4FevGyXh9gmIiodte2pdtagL8dh7
YqsAJQNloxvUGTbmn9R2BugTagLhPHHeXFULkGyVg9PLmxr3Lzq+ba9PV+eirGh5KdaID4LOI1Qc
gr6VDSVOe5RSkLrbRMm32gT49hVfjE6FVgBs2IiQcv+XB+XazfynJcCI4VhishzQXXfvlHE9HpWT
pQXSCTOrcc/HPO6EJ/8MybYQHjxvJjCBkPYbtoqnfY8yiIO7pYGaNzuO5WINBUWHBq/O8fbUkbbe
lWVo/F4+Np/edwCfTjvQ5tZW/3hItd8KT7CyMRACPu7BrZp2waDWA72RbL6FO0rYRFTWshwhlr41
OSrSUKakIy9u32nIZn9Yx6mqbaixaixb7QsbqDpaGGQu71qQeAwt1SBDQueNZXzugFxD1r2VAuTr
83LjitfnmE9X02IT8XE98zwk7+ranhPlSI0JHSD7LArYsSHpnBtph7o2LUoEFEryaLaPMCXC6g74
Hfdu6hY69NYlrvYo/xcWPys5Un91TJJ/1ZY725QwRSI93WAiXWRsgP16gtDDlxyQBC+HKBBeWzuT
7M7uk6xpudxdwYybMeAIRz79CiqKkaDLxQ7i+NyRaQ8F2AepZA+9pp+3iEvstyTBfg5aLk4cMByp
FE+zqIKreINUBy0qFWcivyOnpoSxxKqgdthuuk2ZuErX//Vp5axCcCpxtDW8a8c6bLJxyI4KW10D
VSMq1NmzWTKCNF5rJIFMgsbuZC4lH5RKw7tkJc4b9ovcJs8TfdYFS+FalXbx5krR2hWnWL59SG4D
mOD4mEAu1t992tOytkYuBG1pS+RlHl1d0t/ZczuH0qbCkbDYQsRWLOS3DmHVybB7jR8VdWU3fELu
3nOMcDVu6JQMkR6OHbQoWkyPek2kbPi+yhV1jzh/ECWlbE035dGh+o1tI5o3pgNCXJe36iBtrL8t
Ex6iC3pTx1vJJBkBAJ8UOCoPaSvipbLcSzkhPvqRF+yfagQj+jNbpdPVFmM7Qya1dSg+gkwvJI0i
Dwk+WcKMoFWbNtfERlfXkemOdOh6finS0p2pAsmgqzT2sYdoDlsuEqwedMgZSc+3XcUS6tdsQYTq
182KVS3Xen1Z64OYyBwd6fRad0z5AAc1O01DdFctjfxqVZZTn8sH86poTOSDlA19UNGrqOKE2VIa
xxty3Oja7OVGtCJWAeAHyTESzE1DYkhwjx4pf/MOj6705B99U0vspeSVJioTJcYSPx2LdfKUt0kT
K2u4O/TU1oGKnL3V6nXsc0g5OvoOMPHh+l00pvDndbHEtotJiInZpUM+/c2IoHNGKURiyzFAs/Lg
0QrcFI0xextX4L0HoOwl3gI79+1AGPDIdwv01UevSSrOzcxj6jF+O/pVc/fePv6uLWgPF170UbDI
sk9kcJHIFxJhMp9w1Lla/q93MbDmgP5+TrJhm/ZxdYJjFtYlyHe3p0skIxaoLzpfetB9LjEpJji8
aHNvDC8Bgp5dUkw2s9PVHyaReW8zl3KHFrfBzNllJAgHS9BLKQL6dY36s1JLIV94fNqaMIhbGAgf
6XhaAKKDnXnmEqWxu91QK111l8JNpbjfyJLCHL5vQGrFXefwQwAspqP437hfxy24xVec6vxW1zy3
bme4n7gC83IngQuZe9xKvWambLZCeSPgpflIDFGMlXzHdKk6feBNzBTo0F24qMFPhHgL119NALAB
dx5sT/CwPwdeMmOscQThm+W3wrpEBjEYoj641cYFmTSklpIjSLsD2JeNjLajuOZCTkbnGJ6iMNIM
MrVYZvIgJVOWowmRcuE0/3w6/C1VwMDHFKJLfefLZgOeepKgbiJGcqXbxHWSi8VDNnpzvZdspaSf
V0ZuNSuDKZjmpEcItZR1AmcgZTKP99dnHokzdHtJdM08jd0/KnbE5OMjIe56PkbH6XIRcAagTJRs
OHb0o3g4mvdlgPDr5kJeXiXu7+mTKrlhOqmV1tP98sMjOobQ/dNe65CI/7LcAWCNpjHXYP+P4Ubm
JiodTHabegEL6sdJtwgE4UCDYWtDcYiDFqCJIcMx38cd5sIdrr1lVtt211OCP10uZbOKOvdqiFiJ
1a/njwZwHjvxgal8u+FhX7tgOTfbILXqiYnqJ9ZpV5WSYeYYdNiR/c+bD33pSvFtldCOupLtZiSS
apjD2LB9dF71pu/UeAgZOm4IDzDSvYhcgJcJP6Mws9a9T4/BOcYFyA4RBqCgwPTlA2yDMYNFj7Dn
MKGCOjdJGaOOiYaW5B0CT/c118ZcMM1ziih2BaVcuRli/Tx6AgTPKGErZF4I4io7Q2qcrWMYhFTW
AxxRQY7+lNJ+uVOyKe2m+75KO/+A0HTmtj6WCCNV2mR1sT7w9wfnRCIz0LWbYfOIIvcwLkvhPD1g
9FK2QXxPXH5ZV5BC/X5dDvC6fEWtfn8ckAE6Z8zoeWZa4+vPRH9HJuFMCAd3OQW8qxD31JVbkWOq
GO9RC+4FrHg/CBaC1UzlGX/+SH75Lk7HXwlHTygrJjnr8TqptTYJbO90LL/Y5LFK2LQ0ZnLAf/ja
/VU8kfq0plJD9dFO0e2A06s0A+nlYmRDgVVdoh+57CpHOBxODe8emoi539gDsY3t5oQ5vuCH59xO
XIIVjEWKYed/cBa8V+GIreg5hA7KsbLYdosbvdMQq5hJ+44GGfwo05AwnY1TG0G68WP9tZpQ81q7
nzuj/+175rsMU3mdB3r6LTxWVx+/S+Xog0Hk+AiTiaXuiV3EJbQ+YnZMBSWzNIvifFoWv4t2t19p
XoHr3VHV0jvDf/8jWl9PcPRAwmsayMEtLC9fqfthMevgQLudSRBkLBOpnjjCQK0BCUsyyW8bV0ZT
GqmOPVRIt07l/5p852HdRPChd6eGUstxgX6ujnEocii3UDOSe16Q0sz7IS/wf8XJyZtU57lhzDl2
vedF1pj3wpieXXW6HNRHuS2hWSn8KHY0CAAnUhSOKamBhMYPrHtr78kcn5sUK8glEx5h2jdK7+X2
gUtZtXmmdBJ4lKb+p+etVdU1twxqmoeOElSawDuRd6qHqqjDqotgL++bV4iQvwhGdPpE3kF6Jk/A
yi7cm2SIx+3Gcg/Wk/pOslwBL+bQOWNfwAaguQj0jAcxaFMlEWt9d3lP3qV1rVv1X+jnNYCBElMz
BiBMWJe3aJ6bnBo16OotH0zH8Dni6wY2m2RZH5cWn838PSBoQuQ3OUTH9mHQ+OWJZzG9h41JXVmE
24QHnKLOY/lUcOZydm5D9lOVJH2iWmtFsQxtO48WJu1W/QEFafuDbIK/e6T2vLQaMpO9Xvw1Qk/s
QVpyXhZ1g1VGGx1gAAiO3hdpbCVd9xrwDAT39usSYkY6UBrIY80GOwFkFTVb8HMjE6TstxQl/gCZ
koTjU1obQKrY9WjIO2277UR34uL0sWAWGbQAU0Hh+eBmn7oadjoUKF7CYs6HQZsD4ug6SxqoVoz+
3FGwG/AHsjQhiEjkkQekdOmpQ+Bkyi/bVzd0r6MvsT1Z+wEq45vXnW4K9dryise5Kz8sso3R0MAk
0OaGIQoEratsW13LpPTE2g4fcgxch4mzdEXY446jv60JdOYd6VP78/5Aum1LR4p0HfX88B0x7LcA
2mc71NhsO4TgMinOFp0YjSSt/tD4/m4p2a7Ax6ar7RIGqeHxU01TXbrUlECpabWrlP1gEdLju6CU
DuKM7LmZf0RQ3/9Nz7CLbqwDbmiajLWu8hVo4pYJm5Y/3u8oYTsmTCz5jdkJ0K+f96MvS9q6RFIz
heKTGVpN+n1T0YpTA9IimVSqF2HrLKTDy9931env/Th4b04NIwTp2+EuskBw41tK+A0X9lUmZNmK
SN4M2WY958VskXxabk0dwwzQi5D5TpscqR6W1TRPhxxSqSmyKVrzfm5VKGd811iCm5mYlbRHg6e3
IJ919NsJk3KFR6mJVdLkRoxatNyAMNBQs6JHO7LtjdrLJClkR2pYe31leqRHQWsPdfaxySZxBQHy
rcHCyXVpjwPzzizdbreX3Ia2n+uwhTFVFRy/JbAr9TNP2TkUc0PioByaK3W4y29IdwYnszdu0PfW
h59v5Xoe4NgY44dNG+7rYTRYouC9iKYnQKqSAG3xW2/aN5fC4SyVK7+VYLwKBGCrjb+hC2iSSQTV
2VRNLOuzwsSKJcU1s7rkAH1xbv/QgCzZ3v2N0qVSbU+5t6clBw1uNMKu4voHyf8yud1Rdfg0jTma
2rUFlIR00i+u28WBr8cownf0PRQFYaTA3GQQI4kScDNOJg5msrnMyAwJ7mLCaOfFBLXo4rq/vq4a
uRBJlvg0SCkYnD6vBxVXWgMrjSxCudEwMF4X4IOObrD0UsryaMwBbEuqIVJYoYGQL2j/v5py9gt+
Fdff4Y1bupsqLssBbxj804Wa1VrQc31n/Ly+ujDdR5pkO9KJJeFW3pbMrRbUA0by83PnFYTlqyyD
oXv9Js1RmI3Iep74emGSkvCKVCQHDzxegp1NTKeNM99fHTG0sz+q3tbIgJ67e3WDciuwM1yFAz6v
1wJt+JPXT2J4w3M2NJ8TNdDzvBxHFtifh3WGTUwebEoWgfpDVmeMAOf5ckh22zM6ZpP/BE1UdKA5
gdFctc7guPx2n5QBNB0mDd1RYFY108eLh1SUD/+EWQgXXTE5TtM3J0wKwy1ZEGTgClZahqBxPtGy
2pErX48fg0dZ8XgRHA1vrQhZLp1ZpfsCn8XpD8v3Rmvb/HsYvsf1K+B7CVXJuOzQ7Ov7IuowvvD+
HPuuQXVoYrXziLMlgfYT0++FvMz3d79/u+zSBvhEzAwqxRS/4MHNkFt4fM+RCy9M59BZwb8rl6us
UKCB5BAlGOxErMHKmWDSYtz/J0+DBDbuRrXyVq5kMoFl/q+2HDDJrj2eAE6GZtkdvQ1IQhqr5t4X
DtYnnlK52urxvmDZs3DG55JFR6U5J2cAT36ykjvzcQ93PSHmw77tr+gVR6QZ1tGaCHi9yFOkjcxX
+5ptDUAgGCRQcL9NvhsWO3F0bJ74nkRm6J+ORX/YoQMbzOhA1Pq+QRWrBpixRMZIvlvbX7POjmfd
f8fYdRysirspkKhW7y8xuiYvMIM/3yI4VouN48OAY9+DD5+M3a/syvnoYvLfkeJAaQeKD0yb16q6
XxHGYGa0CeTPZU2ES1EphKbJLCiHlRBNY/WyO0pK5ucjP1zkJkk/UERwFT/4MZlOOB7i7rBIMC1C
jRA+45PiIRQ9qTHhh2HV940IRAfP+gXcWjPhl+3/6a/mwdikzcvQpMhqp7keJzBycQNUop4ZiX2G
EnZZmj8yT8m6lIup3SF7kzr0kwh5vEKZgbhv5ismJiGIKPmeB5zLlasP5+FLs4ydZv2hiHinuhPm
cpyFb4sl9oFWA4B+mcGA0nQOxzucctzEQ1hpp9ccUVT8eKZKtprzKKQPX5pZYWrsnBhBKmtgtmz6
vU6xujLHV3hyZE2LPJL3W4NDtfSTL+xO4597ZTLnKY9d2JbjSfDJoUIDaTInQxNlNx220L+1UrxH
vNMei/UAhvjEQK6VUsEcmj1g4ZBjN5oqCSJg8/GTdIOS88hHglrXjsVJNKPCXi2NqVyKE0ILR5UE
ZDetsKJsS/NATIYSWmwCFdpJxJ2eP5tp96j/t7ZDSjjJRBsyzG6a/DqM57qVajfHxArrdkHEFGZY
oMP348byFlaKq7MAXo0vb39JS2NL9cQWYVdE5v3CG2rzPEwM8qmglNiC7AHzP+DQ+TZ9g3ZeJa62
Hme3ZLR2eIAEU6P8z6pE9KKjSif/8w3TnMqvAgS0EarO8cNxkJpPBAsUlwxG04KHD4d1R52F9P4m
lGMLZ8kmn91pBUM/9BiX30BW7KcVfdBClEit/IdxtdjfuxEU1PR0SNIZffm0RdzmPnR6SxbNwDmJ
ytrWh1C/jcuXaNrNwqrIvoDJ1z+zOTU2/1OGtd8yOQhWtzZSTiFEP0tiM0NcT+u6eRxiFGyXPLEj
YFZS41oZkJiOKRINmw4+oWaFYepr7L8UeyeVDmw0r8ksJ8KQILtS5PFpIV8cROPmlq4gStwyU5su
ZT9J35zosc9r8tcIAlHqKs2D0llKo8oZTAi1w268o9cxacxlD/7b70YqcKmVTvdy/Wu/xsOMKKEk
lsl72moSyoicr7mmsInGSrTTHllbS09G+yD+n/9hwyy1fGmkkWwTcGeHoukryBu6089D4RedSAzV
YjE3brrGD61KZkopvJ025nKlcZcNfjW6FQGefdF9otS6bOZOt9/Yog8MY2ndw+Yo1TakoHdmcmzh
T3TJ1prY4XW1cnxkmWsd8R1g2+N8GsesIjA4bHsdtdQ/5+rdBYu+LPL0zyzY5MhdD7qwBl7HXqiH
f4Ni3eTImEOJX/ipNUxEeFxJodl4xowvN0eH0AknbBZI2japDECuz7UbqW4HPmrEaf7lu8wCcBb2
6ZyZjp68P6Lnm/ws/ifyRgXItKWbWd/7RIf2PLFSwexIEst5ZHTDyV0teHAsQPjF4tARVIraJMq2
SsJyj2OIK5Od818TyAYmiWdHiOn7in8LCXzwHr8wYtcM+wkzOri6c+6aRjuP4j5csru1Cc53eQxt
CDGU5/KACn/eav0UTL2Oj6KRFSban5IZzju7HfaaJO/WDi0YV1C/FanFD9rGHoAmHohaw73AJ8JY
2jBrkCGD74optu6gSE3CqX/wnfa9rExGpiKtKKp4l61WiJqGaQcbweBP/yoUGu0PaNsjOd/urNip
mSAr6E3AHYHo1SmAbe31HbyDj7309cuu9GgyfhUnQ0G52N/0AN/SDhoB2aFdnQ7hTSyUYeFKZ//t
UxcNL9pqaPKhndOiIDoG+xKPma9YzkYLd1duT87+G3mVHjkSjvyz6/C33aT99QJTOtzssERP/1d8
muQ6cPT0+Y9D8OWBVtxuinow73f1zXj7ozVNKL5zIM0dHtGlPm0BpPpS6ZXjUQESGIcliFUixRWJ
G5hVVq0K9mZBoTuTyvQHd3nxW51Vgc7jV+bq+JBCwwEeHncwXrs5Hj2SgDlZYGICxSLWys9sFs4m
PjbJsy+ZGrThggURwEveaNjHiZFxmRSabOCQKmKmxf5ch9EWAEGxVgazZpLLOuOFqunmf1fjIcqU
HTC7rpuoTM5N08o9UEgtjrfK+tbaWqkGGnrwDx/903DhNIIDISFnEJ51KjEucDIGt9VxPjjLzlww
nSnREICmi2dokZcoHQZ/2xMwbgSNopjnMASX7vykk8u5ZHK7eX6nA+p3bM4//W/eBWQSPGYSdERp
A19Cpyr+p9bdqvWAAvzT8ZFBNvA633bQ2VJY8SFlwgm+pebJj5RuX1KN07LpU1Yzyx1AcLiOWit6
LhgwHpEvj9YvTCCmFH1AeUO8D4hlkXGENabAPkp5YYhT9wiEM95eT0aqZFp+UK1KoyhQi+HadRfI
/Lu0/y3f4igp3eSx0UVCx09Em7KG+k7vSxszJ3TDEQBL0qFq0KG1hb/aVeN0WBOv4q3xvbo0LN6S
/ZyQuAD/iIxRA8vHMGTF61jIEtrleiI3OCxcuoKUfpjhH34tYWhqZ5j2AsKKxyBG4aS0HAHRRQZ9
LDhSTHaG+4piIHebHr7rRkQkYBrxFweAFqVqd7YRabT5Hghsbe9fegs95VvH6gnZ96JMv68qNTRI
Gl3Cpi9Al2gFiAC7lauZ562ZsVLiYXWAWq/mEoNV2k/OgCO7f1UVvWIvZUcYWed8Z7T0FX9PjBDq
4XSvmkHBbUG8B582tbF4oVVn1/yZcfn12fpjN4yLRIylzmZS43Yf7WidU+dXirmMGoP23HgBqBSL
+Rl91FtkngUAR6qJCco5MWK2hAmQjoyhtgtzP4wiRsytKM+nts1t2JoJXS5HP/LK5ZI5PKiLe1hn
zWw8jckgHZUw+W+YUczsBsk/PtrcOR3KwqYWRlmNRatgq90cfDGDi/OZXfenby+q3pHoOa5in/vv
JkkxkMfsNI4FBScBLDjhmRkpj+oVEzv4CVZxctpz6OLZjg1jVbG6x3HVxAA60/tANCq4QO2k2jhZ
nUIDF9Pmdjt2M8YrHZlYR+zYGzVgHQEr4wb7phEiieO9f9VrCxANOMaMtz4lddGPFVSdMcDMGf/6
SWEGIEqHPmE1nogjbuiUoKPVULt89Exo74QdKiL/FVbvskSXO90hFPsXs4ntqYWg45Ie9gZ/H6BD
33bD+929YEiN2+LaGwdjiVqFSpGSut8HJbsG98ZbyOVQygaAj7E/hTOMFdWsr8CcyDVeOzOUpuAu
RJN7iPQdkvFpybMCbb2W70dYIGc9pDWq9HG+Iy73UgbzQQszvlmDLxKEIh5cyyD8Dv1vqtu+jw82
ga9nw4tKSJpera2Jnf2LM+a/sdSo8jAcwdbRMcooS/pZ5/uFPOkdFPjRvMcE8mWk8GOOlWtnppvJ
LCGUY40Xkniy2OnG3akHxaaLKMbg+RUPJtCLUbi/EmQ/Z+9v0CxV2vORQHIzVThfA8r6FCGHGcFT
fxE4E0xKIkPIEsvjWwFUFQ6CK2rG9Dkp+614CD3dXB+8bciMZFjhL1ysz2xY16xEcRzm2+2yCa03
Wph+uWZM+ue0kx69xsC2nfwlEPuaLYjlEdpt9xA1ylp3y4318ubbaDBD9KDwu4LtlgOadaqfq4Eq
AprmJy/t4Z7q6nbdtmVowWEroKHj41TOtp3tKJbrBYmrKigHbVX58VJ+KEfglxHqCVlIMVAgIZ8q
68MDDa7NhiGCGWUf0DY6NmeLT/DpxjRiRIcnz0jN1YJy7/y11M42XJ7xWO01NZ6yEiOrA4hcOU7R
qDDZgPxSVyEofJeFo1+zPqolMhH4zN3iDyGn3E17JOjp0oDonuGTXr9mxN8i4Vy4G3KsQv60aQCh
zeKqXCJlwVgOkOV5mnwb12HCTVLv9B9G214qm/jUUOgEN1orxxVg5p7PAY+VxB8eBhAY0oKZAMmg
6ln+Bseyv9WrBppxgU5DKoRKDIFz5OBHL/ascR2b60y4WMqJ+h6PWlbCsA8m/AegPxTvlVkEDaZt
LaK305lkOYbtTh0X+xJlH6FIcxfnckfENFpnBCb/bSqeplU+wSh+qVRbSRcX0HHQzfgvowfS1WES
94X0sV841+QptxTspuLQpRNSyX+QZWDIBjq6xzX+goYahgzjZqmfaHm5Qa7xGyMOrIlCewzKk835
KMXC2K6QFA/kk98gipz0EXYiqAwRuKTWKPfCz0yBhYXpvhLk6IV3Upb1spnhThbhdW+TzfkO8JRy
n6UmI5QA3z0k7Qn12aDngXCdkvPZfDh7fCWY8jnAtGEB8SHBdpce3kfQh3A1FrlRKxYwHTpi0xoC
fxNHXL7sCYRn0rWOI5T7IyyCEKgKwi0EUWLziaAjyNzd8MGWxzkHav/hE+z4WOyvqeT2M3u+tIly
nTQYNtYl3WexzJFPp882ADCRVDBoquVhi0r8tJ5WtYWYsFXn6xfhywdA5dTifhfUxz/2aiYhpIw1
O/LWcANhekrIDgFIJNWJY1R83xG45izpxV9j99QFdl4RY2Srtvp0keS0caaSjVlOJXv/mEZgnv9v
GkF4G5OJHojIyVhqj12IclmB56qOADQ4vR/aED35cMWW+mYusCURY8DgEe50tfkhZyoQyJm+AWYQ
wiSSa0n3A6iEGQ13I3ynyEy0RlwWqd8bP06RcoTqxVUsfrpflyV8GKYp4ZXluzAPxurRJhJd5o/Q
JttFhWtKFt+7p6GWYQ7PhGwHHVL1qum1J8YdOxkyM81YdSMqRC1y9NtfMltz2VjsVt2M1h0CGeNn
fEr4l5r5IbADhJBFhHvxYW5KicTNqV54sHvVgEaU/jh2z5WPyJOC/U/zAFaZTLMz8xEH6Tb8XazD
nM/ohWPeTZC0fXPNGpLIFPEX+3j4qxKyzK42waO/VCshujEQ8cCpHxMcdpPhiBjJnZotdQLkYX67
ygFC19kYlEOlGKoxbY8r2lMAffFT3sn5DMHAsaLsPnkdnKm5cuElb3XErRVmTQ5F5jDgnMhTLGmM
jSfCySNoqJu+L98HE++5g2c7JVu16OKftCSx2kBi1G+7a/69zOuXVlxCSvaE/YB66Edvklw7rCPl
ll+GxwZUcR/f/9Hmtf8AO+rUQUnzckvfMYAo4AuInoxOeDCB7ZBq5m8b5YMvldudUzNSdLNb81f3
DCbekzyRukCkl6m8dsFefb4MZoSSfLVgHH7cUgyg7Zq11P9P/dOw4bb75cQi/hTceVmIuwghMGBE
D/5pvKq3C6n07ktJriFTqZEwlzlNMuMyOVAahnCZerX8XuWmhWkGTH1wT1rSrNvTjtVtDS625/Tc
PQdEg90elZqY05NErUbKnXIXzI3H1VBA/tTutu7KmeLaGfW/Tu6VCb81FZB2wjEf59UTt9ovgzjj
/5Lq+VsLGmJrdI3MWaasOzdufJiE3+6vFizgc3rvMZyZMqVrB1PCUgB2M/UF8Dk1GTOhaFOU2T54
RuJN6mENaeYGKOIScfZdynu9LUzAEbQ4W70pPHHolfbqYKgQsW0vEzPIF1QFqgpZJS+K6N2V0Jef
djS8xT4NGatOm0zOj/nKRKVutNw/hO7oJRXX2T42d/UtYvJK+Xq784bTpxvduFSoO0e3BUR5lcF7
SnJrR3qNfECHVmOf9BJZt0ws6FUa5j4dH0qUpejUAnV2drx/zkbpZ/LXQ2nBjP75HGXdpGrSGghZ
DONL3hooxfxiwesugBDLK/VgqvyNIe2duT6od+8YZBb8mGP047FbKFt/qcQXrIliFfLUV/FJY2Uy
APSTq+amTvx9m7bb4geHAeHp0oT1BstZuuqAw82vPC3JX+uXMeFCNkFsOG04FIAAML4yG5uG7XNb
uP5XRMBXXe+1tJoOl5bRQ9fbExsEN4R0VFQA6gIGLeATVQp3TUjTNExm2WSBwhWZa5UR/13GFzr6
t4ZmKje8QPRtQf+goj0YZ0/kx/IcjyXlDZhokCx7BtzZhRBntagqXF00ZFGvlZsfbzQ1IAftKNR+
I6Cg7GF8Gz1idH9N/bPy1mEzjd+ck3zXTdhNRFE5U9NSIttWJAMpaV0IKoJhUqBJZxq0SAFvrrft
sTO1kcxmCSoiaog4QquGtX3gf7Unh/5z6uCV9o2S0hKgXvDcOXYW6MvWRH8ptolxzaAmKZz3o/Yw
/fqb613yxWenk9UQ6VZhepWNCSvbP8GFMrIlm+/xRUQTMNITkGaOwOMEsuqkaU8UwQkF1dRFHWQb
B6+kwh7pPY61Vp3TWbcOY1p2XhlaGJYJ1GUOC8b5E3yMWGZX0kg8WmZCrVtkygx7GLZOmJ9tisRP
Rt+k/73PGuciA58CPbBXGaOl85b4M5yIfrHtuBQdlm0zPDAn3q9BKHjnBLBXw2l8JR2S1GOjU0WY
b4eAiLalTRaCKG5BZ6ewp//8FyP0k6Y3MHu7KSKzvc7ptEkDd7erOw+l11GwpN6PWj2iTG1uJY6y
f31vP1FaxKfB5FJ7k512qEvfPk1pPrK2PTxtrNBNpUbR4kb4Qci+ft3o0uig5iTs7wHa/nbOcxFZ
AnZIRo8CGf+8ApW7NIUEx3boX0dPYmhmp7Ncg2E+6bTYmEimz5Cdl0MYScgywXL8Opt+tpOiMbZf
8houeDb4VJBPj2ULlCmkOEKwW+p6gSX7XJbJHBXQj39LMI7NnSbYLaqm+x3XfsmFZVU052IYzG5s
jcU5hIr9lzVS9OKSi3EMlUDymrnWdJKv05VcWYbQEZgcjrJdTFNSQOBlah5aHr5Jh2ZtdDtROOxk
wdL2nVDdVeamUYAMDMVgI9EKPsTNVf/3m05RM5MoNSFOTehF3wZJzrLBlZGFBquBqXPpgt/Yms9I
8eaf8PR+zsYObHsXj7kWYDxCsOKYbB1GRD19X1Q2rumHZm3JuC7rUqE+oQvIge+NbkArzNaVEyzU
UjNJmJx9FmukRUZD2K1mKGgsVKatT7VydFCBEmSVODHCBIHFyfuyDwWRbrFHhhWAjaS4PpURZQtq
6utkgmHiKPk11M+xk2KCdbetZJk1QnQR626guPDtqKE/9zzfxHOLsfyS//WRWHF8GPxqI72a6FZJ
ZTk6pyTDgiw4TnRA6XOEc0v6Iaze0+KTQaQeGzv33PlmpmnogyeDeg0hKYf2vBVsRbFgoV08W80E
DT69a1YbGvLOq6QhPvgGUM+tsuOGPXBNt5VuRJe6ezoU47Tu230YGGrI3i5DXpj1HCclnOl/A1kO
s4NTWe16otK57xz2LeOJUf+a+L0Ejh19/yqeqYZ5lLF92R/OSlj3gkurZfpyZwTs/vNMgVmXxG+v
bCkZsxJRI3HozqqLgtmej/Y7KJZ3kuzplxmokMTr0h1TbOXZaPFOl/q/VByJ78ojyliwU6IH8L5b
wyY7mkyAmezCwiQCTicMfJFCLSoaZlHyD5ZOnLKkuTR11sD9yp9Iphu9DMBy6d1SYFblXtNkxR7U
AlG6XDKb9IcwF+q5Y8tcfBXY5q+o4JAWJP3FqzuBR6osyt8ZQNyplSUMsphXUdRkilSutcojQDNn
BQMpivMiXsCMTZonAC4aYbbKJKUXKCE0gmi0M4Bs0NeuDvVDB2Y91uc3kQPY1xXEqsihM9z9alcs
dc9+Z2niNU6y8oA5Rh6Bb/SiOo3SsFHEmaWaB3vJtWa1L2otIjatekTPzBIEr8cFgyiHr+uijB0c
Fxr8LifPukhD+lTkEP3CetSYctZ0CKnPJdRPWorusxdwJ3ESDnfJtHuoEfXFQa2OpUPPVisIOhuk
eeI85/5g0r150ZiSQ5c4+x7sWRHcN6X19V+ralEVWuLkQ0nNknkxalJFbcvN9Kef1e/OhMgCzkXr
5J44yM+jkwCTlqLyoge5c5Qhi4gaBLR/aQTjal26jGeGM2vRMJpo+LTdWy3SxTFSvQ0TrmwWh4KD
Ys6tQEd124WArUKjPCDxdI+/h2H5kAw0OiBaNWnCPyrdvcekSyF311Xjg3cNmFGESLEG+VGGMOeR
YOjxtbux5fuDjG6yg1ezIo7Tj4adiwhKkm+ElrHRYWdrjCN3qEdk/T4gbImY11/58He4g2ZxaTk5
LlMayTUNR2jzL8Z2f9zGXdNs2uckBcFkvWW9nc9/q51YW/mniGZzoSwOAR0dnzmJvY7YsCcPILR+
e9DxEwi5GQXrZniEpbVmN+UCXJzz/M2XPfIRDLRE3vOFjgKajJdH9/b9MALLRwvg5aBkHmQzjgQ3
h+wvd49CDzba7S9/hprebk8kRzRBWExsVdhK3A7Tbj2LXGOqrG/6UYvfEUAroT3n9kirVXzRqAF6
qrA9zMoAC9hPXZ2TcTJPrOyogIGjuNGJKMPJYX5rbZ8eOV5AhCM3ADxVoZ5Xay7aQdDXItCjzF1i
B3sdDfUhKRvwMKI6j6lcAzX9hL0XO2LjE1QF+sTUGheoQ6Ok4zIVJsFKcpVods/YENkw0rboCpYd
lQMk8R5P8uNhEX+dWQgINJB7BcaW+wktQgzNE1mZAQdPR/HZAKpYLaDJCfNeeCKCaxYSPjrt0QHB
Fija5WxDjHwcgdWEfpoAPN3XSQzraaKKxbF+zE4wv4nrHJ/dX/vTEFNZriCLRzoXzZBG/jTWR6Jq
/QLH05NgL/+apYBenRTjiP6jOrMnYPsBnLcOgS95sYpEKem7UoU4ArOx08Wq0O3Y5phFF/FhTmaW
1k7/FT00FTBgzei7hgns7ocn6rPysRZff1g1mLKxOD1QpbrFZ+Dqn9+B0iSmrn6f+s949MLMpfBz
jc18i+2Pn9lw9t5nctlZNc7+OkcXUUB+jKVOoeI5OeJWwfnBkgZc7QO926KZv+Go5fOAJO2kaRBX
pnDUoxMuIWhyGVmF954cT6SRbROxc5qeIY+JGGRY60nWCfuJyuwpT2UUmyjbVn0Ds5tilkBFvvU3
emAwcskT9JrWaSEGCdgOaPu4A8yAoumqEoq/nZoRLvj8BkyV980rSdIOr53H9uLKzy8d7YhNQqgN
z8eAi60YfDK71+Xh+r/Ai98BVP01UFtdpzl93X+z8gwOlBHuvC3HiPuLmLf9j0TmSPariAVEFnul
hOacOyt0BXFKsvIdrfprxlnaEcf2ldNs+fhA3HyCh5WaNJWm95pxgN6CZ4U1KGY3i8mZjlgk/IcM
AQ+1oz6Lt6Ob4xxDZBNtR81iDo1H52pZ9RaNssqEUZERUJ14Viqz1ZrEZAjluzOzE9r4SzcKX82G
rUnpRPw8fhV7tQgj+hL8Deh8IIX4ML11oT7enaBlaO6RkRySZ5v1fX+fDArRsB64ZE8gHT8sT2af
kuukIJMYuYpJc7pRNOMG4KGZiSEFFnKpxIZcYJqEKN9X7OhyW1D97rSu0tfQaZkwLf83gwrRyXH7
7RRzxHqHkzMiwY4ebNN5iiq8UwKRSY+TEm3LusuW+ju2qAaT+QZCTS0bef59/eMhf8xzIN/weCj6
RqvK/CK4TkOR3J3ltQDyx7NuWd1SUIdeSxvH46sy5uo3vZbRpI/9mH26WcIlf02h2AXOsscaPB7i
iJS4Z78XnXHbPTEwrYu7GHyFr+y8SNeVOdmGDP+3Q5/hRuQJ0d4STG1RZMoRA7ZYCwm6D+CMBcky
kXgM0wDFYrqz9IO2qFGXIeFQjNo/yz6kluz4pjk7ULyrb+9ZknOWuDv0Rf4BlM57SfEJoAHLbPpM
4N8s3FUI7ISOWsVh0rQw9LnY8eepWfsXNMfJDg1Yv3hJqZdvNsbSiYFJfiwfz8GRYuGy6PR3qVgY
HLljT1NKO3FzWIAPd0rDY3i2W1Gxdu+H+xNGFQ3wclLHGPQycHbbYzwQc2mpcaCUnvOwO1yvaVD5
beggjvEEMLkSNxaVem2i9gCPM6JXn/9PsuVhskRa9htEFv7r8lKQkyNCcSgXtg11amOjV28y64Tt
bLorZDEmFALG+mZ+lOJEl4V9FtK9qXdbWlsjbxh6ju3WlTfZAf6U2GE3TUBi8KCFcqF4P95lNBLq
nzPKQTSxjpUOmXuz8LLbz2IcCXM/qvGjSMDAED3hZShMM4hzU5hcUppY2tXlEKDXgZ99kpKUhhVP
6Foj8XY5MN7qfHkXes39CTyy09IsD+t7/qfdcWwU6CnWKvM+BVHPl+hrR2T0GHHlUVObugwcRuRP
pjtCIfPmjCUM8FuohACd3bFSX1ZF+yOuTSoOYejScX7G2QbcSjiKkElk2/rP2A+hq1Se8wLq3LGH
pFCYkFMqWS1AzAELMe9RsUZye49iNh8Vp/Q08DZnfkG8/otvOgvuDAQfUWnbX68YhDHDdDT7uV9A
dkpXA11u3cMrQV4NOdeg3fhzhFIkHeFYeYCCxckEC6oCMnYX4HIQXIrwrFnWi0AJKkdmcopd4e0g
leEMmKku3336DCPCETxb7FXPXjh/LQ22ofKyKIPOqEPa9qSamsJfQ4iItge8wKWZ/T9MfyhIYIZL
3KLwfTlWwpV3DT9xwDECy6LYqN01nGQU5buyfC24BQ/aF870bKT3OrjLvBSJfIJmQMZggqQxzmNl
WuohUEfyrOOR7MTX+mzwVoFMOpxGjA2BY0+LyMkys2Yx0l8SXDzxNRPiHUvjRmlKMB7Xu4GGJyU5
pyEfJ1XBR/tScGXjBfaLm45SJmsQ++YVPXqZqVQ29WAXxyf1ADm4Pq1NyFKgszUzyq4JcTZn7JtT
Geinp5NS/TCdP/YQpZnew6w0UcZTFwrRVL3dueX4lO9mUf5pF7DlDkEPuymLpsoKyrzYeyC6kNNX
K9xUyAQ2l2zx5bKcm12iQSS2FGkoSrvTNc83YLUlQ71YoPobZSfQph0Q4WTPwi9sVmHFI8aKorVF
E+dL8GWEcphzqIX90kUCGAROBSgnuAuWVn163Rv7PUaAntBdwA5pUeAdFpjbYqe3JK7RT4P2W945
UPWabGLNwVu2bW9NRsvWbLNH+GmycUUJEr1CoItwdUBX1N/nT/NZpp2RJEgYKnLQjIRWYZnMk+DC
CvP1i2zPJu/ZGoCNgEjLeUPcoE85B6C7FNoKJz06x3rSSq5uS6ljxpo5yTI5nrDD4ndVwOU5+7Jz
LVSt8nkHzLDnIjtYx78Yh8X+StOsNyrMg8QNZfSzMgXAJprZ8Rc9oqhFPka3lyF+U7vckVTljDzb
yskhaPzI6we1Gk4R1U7ba0aHiclSp/icQug3gUf6bfJYbZyCEtoOix8uK8H5wAe9ziRW2wv5IbGA
AtrV2H+Rn1bpynNn9hkPtPpOp/6ckOD8ra57DsW2JnoFScLxuLBD8uGKfaguXTWQa6JCAVJ7sOPF
WdKnbF/ShO4cV5JBArZprcvOsUC6lIArM9yeUMFAV20mEe1wVH3oOSifcAXZRglrx2eNfJVKi/Ro
BHHVvkmrylGOQWH+e5QlPjLNksYPSG1E67tCnNOf5ACD6q2HBe+f69s4/mrkGeZ6Cj/qFvmtqUdz
V3pPXFNEsnFLZIyXDnxHp4GI4UB0+SpB4JAJlkp4ebvwmfUTEEsSCPT+6pKyXlTmnur9SwKKj89t
Dr4ksnHAjZ7J34U1LmOmEeZ1Tvz9rhXFbgjRYMwDAlX1AmfOB4sLpw+m65Ztcp0MfPBLq604WK1y
WjNQmk6IG+867OrWs9Yf9K6tItpBtoXBlVGwLCVMCnqlR0OORte/WqEIwSTI8tXzQZCEEuxNvuBq
GJgWRCTa0/+Tnu0dzcaZ9swNqUkGlEZx3Wi7/BHbpvIWc60dflp4oogRaRuQ/JtQfiLShsg1Hyw+
gTR7tsHh2tBAp26sjblR1Is17+vcMiiPZMt/4zN74NuX+XLHXUKtCiawPKih4ztpBkGfNb2AQ+4A
bjOBP9dBId9gKiVA3C8bQ0yT1N36sKt3k/uoTyl6LD1P8zzmape1Qkl1ijEb4jEixAD0cyq4Clhu
eUp4tMMvno6h2kjbDrtU1KKdaAmtbzp2Zb6Z8I+nTPNia0drjHF3meN5IGdLrx5ATERcC4UqlfDz
62G2ugyWEbp7rvCgwR25/uFgbc21Tyx+tekQXILkKgGpN+mqS2pCWBA096aRLD9OtJxZh1QhKvJO
ZsXqTSe+sHJ6aNb2am8ceOqpoEN5HnB7TBa1q1qNokBlsa1JqrkI19Xe13QNs/ih8uGLwb9dJMhP
RF3RHekQoCCdMXgAyNxhIvqOzLepv0VjvPWkefBwhD13xvLhiDiOgj4f4Zf/CsIJKUjuU/VgpYjv
b0LR6ZhjhMJCTNpvFkxSKTkECgEKi9XY6oRbyzZvsr9RCy88IoKNwU35PWlh9cnsBN1ggs+0hMqE
2rW2IndUmMWXbKR/yr0hzcpekKnTjRxsDDKYAhXYEmvDD3XpKoqIr2l9rJ7pFro+7YpPCMDeBOqC
Hxd/zSUZyHV2YxrMZZK7KwHrrrtlRePhMyTgEyLwSVeentwawRXn4NDQXBnrJxW44K1iQBJnM7nx
iUulNvyrOkAYPkTlGx+xDX3S4VH+6qAdwOckFZgNBQA25lC0UBWqCD24zU4w0RneTQ1hYIFJexS9
xgH3ZJEkqJh8cBT4pCTKTF3CmcOHAa1l5HCekyLxk7ieawyjVJZeCoqFTbi55VN2WKfIKp96mUR5
2MwVwWll0TxM1QUTBJH8E7dTUdgOqAutXrxHSwv1f8v99u3UGnhsbJlZh30S/IXeJnurjaxKBlkT
xu4MupJQKCYINdZ1tPehCQstRdmuRLhIFo958mLHcJVMVuFvJL1+lVFImVlnk4ljj7AQvlasWrpF
F1/N+bpCP2tVdNRhS4y1vq30HSL4lKCCxpoVxF2KRQ+NvHA+nQCxkGyzgTb2MXVGKuA0WjN8DoZg
ap04SO5Ie1p6N72FAuSc2j/QSgMb9clH7PMCCmYkJAoFIBbJsPODVnVJ19ghAawO7WhNMGk9HT4x
NJ2GcVA+C1bOlp5m3od3KT8fEyJtfmdrHFbf3eddRLz79szQXbUQs+PbFKykLYJo6DzauKmlbedb
x3xFn9yN69dlALN3BHFU3mdfdenZuynz92ZW0qG0eiwxlXJWLgvF6Tv5jgbzQrF8SemID/2Y+rnu
iA5lrHBRchw6rYUEA3xR11Gc1VA+0t53LgzuTCLbSOVySjCeep5nwrCmmpYKfZ+k2hlJ4ew6cvJP
BHltAIVxnr/EDOgj2tp0fAvgogCEckv9iSWjoR1RiC0o8ff3rgBTkGxamnUL2m9RusbBxYI+Q4HU
f0PvnNNpKOrSZqf0XIInLXEfP9odnbabB5DCaPnXVRT+asxF/FtcAQMsdo0F24U2gCqnXG3vFTmu
TWUt7UfcwZTRvJG0dxaqgkVOdf1/uehXdv5UJmrNpopFFSSQV0nHGiPrVN2PH5HmfIRkA+fxkw9d
ahvtJ263fqGwHXl/9OqeUfM6+0EdDeNKgSGR+xeGnFq6uMqnmT0BEHp+OepcgcxYR649JtBSVEEu
kf0nKCFFOd5+JJPJGSIcHMLazHhrrOv6tFWDOSOpI6OvDwSGeABuJ/z43VRNrGGWu9OBbqURAF8j
rPiKSkBVPgKA4OEhi2nUgq99zObckDE1ZqMzZ0bTvTMnao/AW1eQwkblg+Y4ZMMYKvCQwa15hmKz
t5hhyS6sB/fyLoljxlfHkea+i1b6gSjAw0rxduq1wnmY6L6K2hU892jbLc3QZp3TrVFlQuw+cWqE
3FizZK0mllWlHZxuOLv0V/h8FqL4Yt40eaOWoT/1swDtP1GX1p3e80qj6zA2r1BE4eUoYlanPZId
TnWR3dZpw+WsHUCDRp+GXz4GAdDuECY0Fd3F4xL/c7HUFjZSJUWvEmTNc7prwSuzJUoF7u7ShJ/j
2hVOW4iw1Ult33akzO0nOWnUxLrAHqODH+rq08AlhOFZsSMxWTG1/WNmn5bnvx/7ZtJhJilOXZi5
Q9w3fWvQz4kFSj3mVH8pBfIdj/crkItMRlomue0Zj6tipObrsOAk2xDNONAxmaJSszSFy7TAfOsU
PG1Ayi/VVuXm7Sswyr4GEa6zOh1JMOtmzHP0SjYPLLRz7M4QwFRg/2zSYhIt+dxOnKQRwrdWrqq/
TUZ4y8ITtEZ86EydQ1ag2l9HzlE7eSJs6WkpTD6oEIraRqAmRvvgeEeiz379vYMWkz+QiRCxp1Tb
rhocgntqwp80ow29mv94GhwUvxXgPipP2gqnVxlgw4EQECRgv6SaheXR3JhUinRI5re/nBFnEeCL
hXK9R6eJuKw40Q6StDK1h31tbyyAMTYq5Sg34NDTm4mtKDMwua/JIdjFwuJFoj6O2xRcXNHlQKaF
3JhD1K+2+y3EDD52SdDU9fAYAkBMsKUno7HWHe4gzzJErDy7N65/z7mNOuySzCvX1rOSUXgV8pym
/s2OsUbrApPCi65PK2oWUZ4jTQgktCaH+Vf/3W0SWQuJQHTLaCtqNiAI+WazKbev4tj9d0B5rIt3
zUVMkvFu0a7s5tIg349+Rb7Ev6L3k0VYUpdm5WCcnciReQYTa594IY69Rz3ot1CjSjXP2brT6R0s
38SQSckc9hp+Nr7+Ts6N9nF0ir0wcYFd6ipP+wZq3q4jCYn+nX4yHRZRhqsraBRtowJL66Il53SZ
GTzEP4myxP0RI0SkgXd+DkSM39sBohqmx3+02vl0hxyBio1FGXokp3xki2Xi/WYv9fZ45SzYCGNn
IDmal0KDKoSk0UZsdX8FbElJGqfoQl4M0Ae8lhWMtIMeIufTEPV4XkTC47TFj5AlH3dnB7oyDhgj
vXdikoxaNmJbOKD9ctROpsSxdJ8KKnHMgSn3xop86Zs/aP65fI5eANtnFMHBWvnrUGD/KqVdlzqF
AuJ2UcG7QIG+jeEiHdhd3MRwNwURcWJ7na+8IwCMALZCDM8ghuCOLRzvdq2aw8e2OQ086v3BslPw
ZlCLaLBp7WXK7J5bIQsLu68r7/lVtWwBC9vpYwOpfzBObnQ3utoZgXPO8F7ZuWHyoPUfGq6lH8zc
AbefUv7fGVf+5Y1SpPlA9f5jVUEMfgxKiJI7MPfi+9tjdgaE1fIFEdh5UxISJxdZz12boyUb8k6d
mE3lFelPLU3ttTI3mnAIVG0W3pQSM0yw2jHUAPj8BSALiSdjZFxe7So2En3cvca1PCNi/MuHNvEk
XQ1nXqtJ0OtELvesRurD6No6vsDdFs7+NR4KEdYX5wE1s+xC5JIgIAnFr1z3AcjvxMDGNKdE339N
pA9gBF/ZYPp9sMas3Va20zEJzTU1SfPaH6HoxmYzi1pQ6BJ7vIN2n30WV3dHibA8G09F5C9LZJFB
+uIE2oRNlaFd6Arcoz5UUzeSzvOkFQatJ2NKkwO+hxa4x/ZTrIbYIS7Bh/dXJ2voefNLh8s3x7GU
J6FvBCETo8fwcp3jy6RUQrYnDgZbMkcD0Hw5KWE7SZR5bcNz0FTRfBpfvkWOqczmtibQfvHfmKyJ
HZTDO0yyOdO5SLyldie6uwdgUsBw+a/WJ4x9GlAySLdc4EV0cJq8nNPvPrS/CZaW5PHs6csWJpY2
Ag2GDnuNYfGzt6cWORJmc0dmwHNWddBtCtRJfGToIBZkJtTAP3EyzwZpl6ErPbkMA/tlbPoqnCWm
FpUaKz0Me98Jpp8XobxkKdCP4iltK6X/m7+J6TTAIKxwfbcXbos43Y+UX+lXFVs1styOQ0kj7OVH
mVDdUpAS1ZCPiCXwos06PHjWeXy5LmQ8J70XRLxMpPyV1a/xFxpwq6GzTSx5NdgZd2yWJ8aTuGfl
YAo5dNyc+je22H13LhBpz9VXAhelhwXtW2RwlfDeu9ClOu+78L/b4GPqcFdOAIEm/1hvYfvIL/q+
txZIN31puvzv1fNu1+3soU+9RsQZZamkA2SnXrn1mLbx7unSUf0tUM2Vf3yGM98YvRsgXSqEBLDz
YMXtYvgxQMdTB2qYKHBHUDGd+U+h+JVRWXoLWR4crQyLy85Rt2zfHWdVumL+SFoVhbtresXPmZqK
TPsp1K0HbRdg9vCcuSn5mfGNWtjs2JmDpmDeLHSYF6/GOAiqmu8TUNiPtopCm3/FLRGryi5ewg9w
VG8qO86Gj8dLfhkWhH+7ajtTs8vQJ9pc3y0zNbI3sYXnFQzOVtPNFI/nwQJznOyizLHdZEnMTZ3X
i/gsPK2GVlNu4EK0RqUZj3in3ophx/W/13MdQcBQM5F1VRhsJCsPvLgtzZGJobChsuvwylUTchxL
QDLANieQE4wseZeSBYdp8xWA9uGuyzrKwvAr6q8wsn7A8mhIxXxGZKc4TqCouZZzyzi/+fbl6E0D
kV51GFZqZ323KKDpeFJTa2M6YGFFLP7FdB16/Stsv15q9ANJAE2Vcwuj5qeLSyY3RLgxw/Ouzruw
jQTioiTaXpJh4+jlNCz/h67dRjx3u5zTaLnOTUMlpaXJ5C3U330xs2c2T1bBZv+snv4O7mqJk/yG
jSpk7HIne9RJShTgXe9nDnbGpnhHk7I4EZXx7WpJPOpgd7VvAz/hdip90ODUYyqubDvu5uCnNZ5r
nbM7QH+Pge44lXvSOWekbJkQ5/wKzfxrTroikNhmc9MtCbogkM+xLtDOWpXUlMDKq0y41eqvXXjs
tcc99j9UzrHh4ezUwIhFxyrO5cof4BmfTTDN7X6ievaTTvAamgp2kz9b1BPd2zyLj/ozxQwAipMd
pSc2hmHypzD4rsBf6Qwx7LeOY0Q88xKuXVVV0r6Ia0vcjmY6vzoQDUPi/QEE2GFT8RkXIvub4pMZ
1isIvFPbBjSqbfWXPcri3q1SyugJNr/lVRFHtrg9xbpS6obNvjK46+5VbVloDMojhoks/XP3XKJv
lV4tVPbeDCwwp5hc94bmcn/irNv3GkDCBkEQIDfRF+isTkJxgzyygR8Lto04f9iAd8m7XokcESRs
PciyEfNJbO9Zk9wvco5zup4DydpdtxE/9n1ST941VNLC5t5s1MuQ+iGXQGm/ggL0z/aVMQGn3ABM
HRL+vRu/HS/VGy9OpxFj/YKylL4ADQRh/TdqP7OOEsoQp98gTl3GYXCZ7xVtN7nuSwsaJ3CYaXuT
OMf4IJYx5o6MmErHavRguvdfyxWbejlHG/Ek6FkY3+kJOfORxwKbcap/O1YImJxkOkUG3eDsfIq4
ogylMVzhwy1yVlfqYeU/PH2pFOR+z/z0pCTUfe0iNl2gCDiwCweQgHzJlHTIjJ/G5O6mbccv0LP8
dXz7hM1pFPROOOfarlmhoyLtM9EuYHcl5ZmvqzzFSYvJPmpLckxIYaL4lNGLIAzDz6Gw65jh2C/S
VdzAbNfDe3bw0l5ye7yNpE3UMTuGwLjoauxo12tpaDZh4trd1r5TjogwbRDmZw+N2UQh6Iann3F+
etTI+eQqZIVwPZpVO+rUthJBlrBSWKhwfr/Msz5XrJB7hJYy4V7jJ0qshvWmyDg+V5s6vWvCBwlD
YfL/u6Coz6wrD63Hsf/Y1KeS6rV3YHmix4bT4x4lhpuui2gkK1l6B27uQPcVL0+iGDkTXeJTn3qo
+wYkZzRpdKOm8gCuCJTXFO64FxraCJt+2OqSUK6NPmy5S9a/hx9Y52D0KuiKPf2Gw2NQfYCAlied
2MuAGV4zExZS+nm9GBg7SkTgbv9kQ9jMa62c9QXjd8WwDjk7+EQv2y5Gme7JaHiVySO1A5BEzocu
8PBPW2C3PR439uI2523PD7p5cLjXi5bgN1K4fWDBO+NvOvc4w4T5rMsVK/poQ8e7pmwdqs+pENHb
zRG6er/Ft0PdIEuHeUgq+rL6+MrFrM6fDfYNOBzBalkPEKTgK89kx156Qb8uaTLgVKBFpgoOAIr7
eQ4eTXErcdZSUI3XnOveRZO+rDc1HDZofbD+/5lCEO+9N1AgyYkaTqJ2/zBlVHsSuUoQhOs+XJxd
JVk0gkK15MByq5blfMI1DX+AxDtHm0oDdygk1uPAmTWhJBj3jTyVsy2CpCQScTjfpW9efdjzQxlw
OX/JT/H6aAgkmfv6cv8g5mzhNhKemBhNs40MiBzoKxJXVrVTLQh2hR9klEEDc5nMptEsEAynMYZy
FGRUijm5tEIMZK/zFtxuBC5xQgtXTU/1f6x62k4RO9FT1MdN1lTnn7m6GcBipLAJ9ubp4gJrCcQr
OdKPd35o/88O3PL1v/sFZGcn734RBVIgbsZ0r58MXgi5ZEo9WhFj+JvqCZ6H4O80Vv7k1IMuqUIB
I/C29S/0/dAVEknAIprIpjrZECH0zF9xGqSf+jzs220jSlfUpcxVuCy+IgkYN4y7FpqJN7zwH8jH
9MFrcs37jltq39MWU2SCXRq0CdONKiEVdjyrDd1kjEgKSKdW0TzAwN/R0/1G0/4jAfM5on0C1Kjj
lhZrm27Ko98+jAxibF/K1CQsAEGK7b28/8MIBD7mhnUaupW3ZyrT0rlevSUbPihWZeLqKTjW/RIi
C7/5y6pMd96aDBklzqgtbW2DVU/UsXmWxN/gDd3czsbi9T/IjIpMr9FbVKTb+t5ikt6zsf0Fv3EY
dmw5KTq+lwPv1CpDHadJFed1sQofgYFIah5mlfqAHzPUC9UjaxIsY02DviGetcv9N5VMR2XVrBxu
0okBeliAO1GSwCxMUp86VX5E4WgAFrjUsgYVwjip4owTD2cudB/yD6+Ho4A5VFNSmVf7tjgh2A3/
CY8/tS4RNTtOWFRh7exc622CTW43T6+eGlB0+kEc9qyINCTrRvTvJLfqQ2ifSHUNg3ePWMunD72q
4v3UwvS8rMT1lydXvMvyodlGvQKwEuwPnZhy3xCGdXDviyf5pv2oEn7lOG3tMfv5K765KuYMXD96
jew26WoBNylwuGNjyUmIJpvKI/KWQ2tvSgALaYBta+0HyXho838W1IjtL+h6EImyL3s2OlFnyjfK
VgZc21NtGc/q1IXjQO+cmE7lv2iFLdRussNMyDLHlJ5GRQ23g1IdTBJiH57Cvh2DIVJzPVaFKdjm
KxsamJ22TeLSnsE2/gJ11zyMWGNAobMLEK/6O+ECLYoqQv5Q1dO7i3sb0ayUpEV3+p2GCAEEJ9t/
4vwfnwXfgCagUrQ4baYKNbwuXEqKkTW/HLcONCW5+90IxzGT6NQA470mqT+Utvfr8aMC6J2iXlmY
18f5XbknLbrBvNFyf2qO8TP03P1rf75AKNkhRs0gox8OGoixHRFMKaIaTcCmNb20HSfd1Rlpk721
vhLBFNnYudjKG8czOGLMEGi5NPLWrKQA7aQ7vnuR+e2Nl9SlhewjmW5ZlOaxE496IXhEY0S3hbxs
z3eGKREGjOr+s13WTbUNU+TCnCkYPWp8psr4n1Xj4TGk8Nmu7wqp1tEFN27H723tK7Ctv7y4OuGn
SUD5Pk9p9FjuNff3Y4Col7mAR2Cfi5c74BVB2ptPH5HggSsAe+YzEyFWsvwTRHEdlaR6hohxlKDb
drItGzcEy668bRiNuNjhtkoFMBbJFeSRMdVf3+Bj78AsPz8V16mRxGh9RKco0pC+hrrG16rD9YZ4
tvjtWjKKdE40zB+6Pt5NdLo80Se/g1z6cxfJ8FlNQW4K6wm/z2DKZ4onwoXNeFFDvHaCuavk8Txc
nkM/DLC4nV28MljlPtm8689fYhBQ8n3XaJA45LiHj7wKSNGbJIqD09J5d2zI+FalbyiDcJY1AFjl
ZoU1XOGvJ2xVSXwjSArxnsJUKOXkgl16ZBSD4ft4t0B/Jy50A81QTy77ZkmXDc+0OuLUSIod47os
5Yy3O//HdqRj5H2CrKrbW0dM2Qu3ytOJqNK6SpD7rhUENtritfaaXZ8jx5KhQkZpUYz+h9fvRcrh
mHk8gOpCLCX168BLCQkTUhBvAvW2cUBP4OuzGJ9QJSpoQBD8UqrWzu9UxKrueR8D2Kmarni7y4/P
i/t8L51HnVX2CCcUPFfdJawEM+83eo6DcC5C7I9DH35DJLAi/KlmXX7C+FOgbuRnj8FwT8MZyDjq
WnOiIq2ryc9AH60eaHMxC85kD9VvLNN6lFeQw9BXz07TnjK2gdh5Mkt9CjkH9gngD15+ZjKWAjeB
UwygwD9b/xZx01eJsAHcnQCIILbZWMbecZlrYDiWYrRrl3Uj7HLLvmqORRtWU5FXQohu+croUPms
yuWS8tCgYgluFokWgXkUdvRg3Yqf3NrsbNVR4oxojKpi3pDUEyLcj9U5tRx4TG08xQqLoV84FC/X
rUGj47zz9duQbaz0dS+dRynbtZFd8eL/8tF7nhmQ1jC98U6RlpGM1WSoycNEm6CpllPlD2nxYHfE
iKwwIPVJ4X+IcLzvl7idnEouRLyxIrSfDOaNSt5HQcdv3PJQdaNI3DF0JOjI4XuyvMwba2ZIKEEB
w5txJp7FZmofMlTwsRLgnxYliOw1QTNNxSJUbXOEmenU9aqQGuKeuC+iXOu4yYk2e3TtDcxNkdXy
WyMStmj/Fjc9NJNhntWAL2T9xtSkV2ivCgeD+LYI+pMfgb9+06E8vaMu3ULKzqjafUz3ZFeeoVJA
NiYfb4+MQ7aD+Dpup5eJUnWvuUXFNLQ2emGBqjwFytaqJiu8yvUJyzxFNeFYVei0OaXcJsBvhAL4
c+6p8nEXvx61aY66owr+RBuVr2455cdYu/2rXBDX16TxLpkKRfkZF11k91HuHn8KO9CU8/hdRhWU
mshJJTbblFhCPUVfHnzU2SP2OQodPM7+qDmjFZo59Dn6Ngqj58jR6zNP1Aobl2zrwN7CPQ3XWeBV
l1GhJnL4U3DHCb49NGLU+T61JG1sEY7tNG74JSr9MJ1nsLA1OofGQMJx49A2M3n2D7zGpj+DcLKf
qgTIyUpEA0PEDCF6qYPmVTxEmeCVNkQoCPqQeUEl2mBP5VxPJOszG2F2hCPJn5qe9FnlBic92O3u
JCkutpE8Gdf34kkHgxcn2zJdUML3bfEF6/eUpaxjr3jBieFJoH1f5p+QnDYPOntH/ixEIpxQZW6g
A7RBvzjiV/y7HCF3m5Jhtl3iPjhNKwhiQ6hkpytQ3JE7/Gsp+ROUcUTyLNE5yTgEIcwCqgX3wtp4
xkdq/NVB+Rm3Pj6E9iCo7pwKxqiRbEu2KT/f7vbVe8DvbyuDxNjyhFw5skhjqe2x17jzHKUHH6AJ
LIsNW5G7yBbqlDYZsMuMsBUJxg8DXOdPBvD/2HjOZqIzbByPGnXHrhydymH/73BwW3XKUFepMVLl
GAfqkS7ETbBlHq2jqXCgQRSGN2KApL0ou3GuH5nkdCoQYgAGfHusD9UGbzxdZ4/F7mD3oDxJ5i4f
2cCUoc5cFmkH9aTFvRKrQwLTFe9VkhW8UKPI31UjSfZdvzwYdIcr7DE0xS+M6KCPA5xKND1y5UvD
FgyypBxMjnzhzyGewee9jUABujcpKOO6W5Bql/YUypScUqiyIQlYiQbLVOIHuj5DRYrrVVM1TNea
gUV+oO5U1f68sb8Y9H0C8VtpRxyHNDr1KRXqXiLM5r1E9E4P3NRw0AHgJilU5nccWpQe2r01B73T
2bcoI06CBY07X2kBOkoaQObUblpZFw6sLAEGUUpqxXJvlAKCcVvHdbxloMbqfWcUkIbO6Y1MnX4a
TI0OdfuIkEjGk61CH6cvjG8FVu8orIJzbNKA+d2sdf5OD9gNIET5Tn61i2GoJ2q28IlQBwpd46T2
iyLpEEl7sCdLgoF2MJGFxrQnvySCSL3qzaE0FKvFR8Uni9I1JP5xyj/l19KSt4sZH/HM+lV0Rj5Z
Z3wSj/g9FYNf2MelTUMN+pkAQlFVrJ0nNnXabBABA8LwKc4NRpL3132G5ME8cTWFBJzNMTuAoJOM
APx/d/WYAAeR0GayID3bcbhy02BklMzlA2ILH4Tvj5sGqcUmW8lqLeEyJa/TfBeC9DW3KFPgDVl+
R3FnxfMhhUb3nWdRHp4eWtfptRkUgyVApCVr6lZ3tjGHCAVu1ugiYIr7mLECW9W1RrYkNFeIdE91
xA8Q36MqTr8xpac0NaCZVR9ULyMTAEEpJLZPDX0ZAKMmvI11DM7NKrOl/y4JrXWlklUU16L2gPzl
MxxYAJMnlcIbVqJbpsNXRCGqNK4AkYzwBgnW2ic2n/MhwKXKgPX+1Q5KM9gqQKA9UteRlK618Sqt
47xkS0eLkADifIaE0isjV/5rKX94wAmvRCXfATcT9KT2I+E4SzUeklOH6MZh4JEuzHARK6zLFRpQ
ro9RP8uzUy4FhfJwtoI9MbalkPsx3x4oNkDlvDzJS+R7+K9nYpHUMzslu7Oqsu5V7nrhEW1QJp05
kWO1pXQJYaYbydrd8zkSTjUUoqY10oPJJkr3AmSj2Txbvbsayh8gLxedhMmzMVx/o3aNLv3wkray
wpvVUFuR5CE8puxNqTVo5pVywjoIvApy1Z9GBaq/BYxXju36z6iqwQf/YqNXKzoc63FsQ2a/8NWh
R4sqH8wYu3hbDu3Vvcdetzku+F3+muIDbhBxBfrnGK5SpS1QHXr+Pk2crm+vQja2jMJsS35ln08o
Cyc3UJT0LWM8i773xDjZpYCEawCMZFZaTV9ZZ6qn5XvDUI7Hlz72iaShaRzkNfoRdNe40+kzurgN
FRpFPDam1Jn6VhFcbVElhodLaBekGpfYP5lJxDxTZQBHQi0Ujkg22QXB3f1hiFD2DFCw+CrBUKQ7
u98OgzjZ+dZIFeCN+FowIw2+FseKNbQXD7nUNUBJxs4QUa6cgDGz9gz83zGsltlnjYRSGJmB+gH0
LKzgfa/O/dRYUbcp11JluugFRtJrcoO5o74f0iyPWfgCdtCiA+FrP+/nu70zDD/uxuIQg68YTwQA
puGqYkKDcWhHHtNalPUfyeZkGSYLxFHMBNF7PpCcZAPGVTGxdyAJ5wsPcbIWJPU78DRsh5VbehvM
PH2PlbTqREsRvzYs3wVWphI1TkZ81I0HcQtq9l5ufEAqwmw0FzrtqOWuFI/yr/q8SpearcfrHKj3
gEIPxipaq5WSXKpqZ0NqVIY3vtovvTm1jLmkkFFwwlq9yYTfeMlEUcSVBrkPQZSZFVLqsRRH9gXa
+CC1nmse2/CGM2TAVSUiyO8hdzj9ygHNSOhyWO3+a38i3ax6u7kRIZtoYa8n0qGanUcgy4b1eYS5
mHA6k7z4iUh8yK4eh+ekmgR2JnyCTkeZWvCFRl0zHgEG3vbOkzsUSitPEDOaIQYaqktKJ0F3W4FE
7klUnCiiTHihGVCtU9yI8DO8ujtpF+FDLDPfAs0a/qs+ixrsGcCCVoulC5xWvS3BKQpj/M/GAwvn
fmkQZjMJxUn9Zsa7Bp2oUV20l+NM+p7AEaN4Dy910KIL/FDrApeR6vl/eM8mhXR3Y0S8ZLCUiVNr
ULcZsddUl1YUPHWRUA4imW4V/UoWREMlmpqyUFmj9RPQaT/3yjWdbCkay5ti6fkxL/VkiLM+tm3Q
H3SjKd0jLJYALs6WC3fztDbnSDqIkk0mn8GOBNgrosrbYFjfpkn0XWdlhg15+G5SHRqpPnJh0Enc
NvvUyOptB9qZG7OQXMbGEoQ7xyMLQZAzz2tMHMXiaOFyCCqp85OGLH3mgMhlET03YEuMYn5VQlim
KF9bd0vyFGRfX6FT7JkXZv9rli14sfJ5C6RquvgQXYe5cVkYSAbu/8b1a23SGEgOxl7KqR1Um1EV
hmp7+jGWQGgWeWPu629Hr1h6zHonkhg29qiDFq8ditxSPae3RRF7vi8Yekxgw9EAYW5rT1RNgxfy
Qjz774wPh9GmK79JgF1f0E1LJayYxSQj7OvoOfR2N0xV9aw4xrh0zzHimrly+qYCmMtmFGoraMH5
3y1ofPWrblSA/7Eto74EN2p5unGKKVC8cOUqRjgXE3TlVoPA2e54lY4mfcDWB3myNgoXzamGxoXA
U49R166JqXva4lyZRi8ELpDli0caVqj55y1AgFeB7tWdqtLe32DZ2kyo98m36e0PLZuDG6c96bXA
lCCL6iPbJp3zaJcSh9ZKvxJkADTMmPddwOhzVLJXBmZTw/4mT3EdQe6m92T7Vru5/g80bFED8ZeQ
rZvRIxKijRe/6ggwWZZpkFyHnhlcUfXQWRjrDfWd6CyhBZ0FLMNDqYBGRQZVKQo7ZcMt6VMP9YLI
Qz8k0MI6mb4w+bqI18O1S3m5rGdUFVqWF5dxF3Qz/sfbC/59AXuBf/NenGfxEsXcVRnrZp6DX8Qa
5hq9s+Vb4vSVtLM8lKZSMerMYVCPb2oY7DcwVtl7hLL3P64LRz2bE3O0WQReNm03TFGYyeTnz8mc
T3xgA/4SnGU1/I0XVsUJqHhuJbEhx8Lq1yw6MHQ21AXolJVhaxuU6k4ONV7pJoKsvwrE/JR1Ummu
rvr6UOsZM2DhkC/z4VWicwjiNCuOQc8MuRAoBMpZ4iyA+8WFzA5Wkc7EGcZ6yIvKVUsjkEo2y7DR
G59xBFo9j8V3dezteAAtu7M9B6qq7Phpgoarssl4sqIqtIrb7eQFiHca6TvgkmBug1CkxmucoqzA
DYP9hOrgct/D0j7pT+jrewaZvrrnzr59R9kEiHH4j2rgLwV+xmqNQwtAgYBnDr3q+GRxLwTxMZbF
0cnK6tbh4zKkR0fGxUmTaZI6CCooceLhjwo6TV0If1XHYwiN1q1u/aMxk2D3HJXzb9XnoxcsqiYF
BZQQPH1HjW0FvUxeqVqT9aSAxsbQ7hcTwaeNXX8YWydEpWPtKQj+Ii3vRkzjbGHlafFCI9tQaeUN
6y6xRMxIj5iu6UOcMQZ6m3A9/hyzIL4eKAslX7mr5Hltb9QJP7tM9AmIw6fClqi26i8Uw7eSg4Tx
VDEAk0/2pMjL3NOVZJpxa9XJc0GahnQwB98AtOCZAu/S1j72nyu/QsP0hBcvIw/Zcl2mHj/LdaGW
2xqlaG7Q7MUBMWkm3r6W40NAwLUv70xjiga2X0JNWFCK7sYj2cM+yFoMT8bKPzDAIM8GmJC2LRXt
UhDeKUUi+S/7lxHTylGXZv/Sq+cNXiO3Nl6t9ODpQO+G7heZ4/CzqxWhndA+x3wILII5PYAvGatN
E2LwcPQHZEsjq0N3XA+O9P3/9kRv/wdycNtkt1MEIaiUEMq6jVofzTAkvL+D/p9UNj0wHZVRkFbV
xDr/k5nllM/uZiU9J5SajdOvmSTDlIVqCPLQgjL53qulpJ/N93xa92nKVikQPq8bF/QQpx+95YxN
dF0/JzKN6WFx+bs9vDgm17ZC9E4JewRP8NjD+/7dKWNl/N1xiObJcGlq/7JBB6VRZkgKA+xEkpjE
I77IiFlD/vSPFn4Viyl+i9xcDR3z1UEv1cjUJyeRKp1H4EpoAlevJprd/+r6SB/+A1foHHBQHk47
T7tDnyCf3FRNVm5N+UEOVYS4rRXq4pAkypPawLKw/2aWv1Dx2brnaWJ4mymTlIRa8gqtpaAXFn6N
qr/j1m+olC/Lp5l8vGynUD2ut3hmnCp9Q97E3rbrwws4y3QTX4tNEJ8eg23egAEyFj2NCZ3oOz61
GVS/lv18Z+IgX0pwa/t5lt11N9tuKR9MzOk1EpyAgJzrD7Ku5sdCSvrt1y6lAN8fnDn8kbzONRfS
QCY4hsRyLqq2HaSMxVgkqwbt96gjn+YzmfpvQYon0xMQYcq3ZNTE7NGq8I2nPJHCwcFPgPAp8MCB
ktVYMCORi6mPs6zvj4OnbwqpgZotAKD9q9sQKYO9l8Th8rGN032DNDy8XtMRRS5XR8JB3mlqCcCM
gYrPx2eRtdiNQvBxdr9Nom1mQNQYaByCAG4Pmu9d13ve2FqH9kqppJouTG66MEqYoenkaWEoTCTT
JdcU+iq0whTtxQ0BnO3yG/tuDgCL5Y65LvQQdIMDVAV6Awm0riNEyXCrZps5OaXJUJrz8jvRaVOc
+76D9ZPa0om89InLVzar7feZZ/1E1WiD8Km5SzQ6nmfei1UrH33wKmjRIGOzDqbboWQi9Iq6/5Yd
//h4TOiA8xDqyLg6w6B/XtT6LLBO1wsX6XtcDcLegvf55SIzlJNoiWdQBbDUEoXZMuu997DTLlHo
lG+wx2fZkyS2Wvw2I9nx9qjmM4uOIwJjTCdsFGmYXO79DUk0udIexU/hr3uBpeJg6GSd6iwUg2CD
ZoaR9PHeN6Oddqd8YEGhBrKaTeoRO57i5iX1U7vVgjpjBXkdn9GeHkxTJOMQ7my2M1hECmaTdTdG
LZ6hKRX9PI7knZk01N+aUv33bO9N7GLRuwJx9pIstGkA6YLko7TjBHavcTA8cwlUXacJIlF7nnzx
AtLiY4WdNENhbx0f+3OsOLnETipeIg2mp04zNNDx8MwG8yQ8ealCKEaR7NRYB4UBbiQinz94TxhA
4ZtAuoMduB6JtnRMGMZTYzOcfs014AjBfBuJx757ZGOmrhzBfopn2eUDkPzVAWZ7JfIKusZxylYL
aSvev576ARAkXQxlgLxFV0gkFloXZRcqrxxeeacTdTRyFkmkNxEiUGQGW6EuidRq4qJlZUiJa1tG
ySncC8v3iPq+hExhCB0u0xNgg3caBzTQHLDljJ4L0M1Tj+QWTZLsZbRkW0DuqcHL88GmOhcE22LO
dSRm++bH11looxKtaxrXS6m2Uwg/EofBMcNx83jkJUQS1LzsIZcBoOqrycMB5jltYBnN8Cm+dP/G
DXSQbLX0BHY5OsxnfNq8XHYlqh4DRy4rPlVGPP3kQT9JuNL+2udiGa+9W09J1iqPQzsdzZdQrgde
Kh+yiOTEOcOEvNluClZmSkCpJ12tj42Lno3AL2AOOo3vnL+h2/eMuH5gB8FmD6biNrOX9qAvjUW5
5rLIUWQZgu7TIbC/9lKKM2HU1JGgv2Iy7jzBhx+3XlSOqfvuaqunVENtbgCD2aCoZl/6knr7v+a3
Z5SvYrRaGWaepKDrtP9wt7WB1DM1oTEjzjy9baVyt6pJBwLPPzIAf7knAt4olCAIU/EFoWYdKpcN
jc3vamOPHUvS/O+IwhlVcWfQywvMOkaVhX2ix1JPc7XnFkhXcmVgtyVvIB9Wsgr6L0QLORAi4+Cu
mmqL/zM2/gj0XcJaPQm9JZYZdxuhrHmvoyPNd043sE/4JdVmQgmCYUWzBDfWZSGMka0CwehHNqdR
Mjlo1eThPqc0i0cSzv5Y2mwby3BxKMwpEj7v3qjpzUdt1ZmditJRM4v63bOVOsOOZuxFtso07KJ3
CSGT0Y2euDE2FRlmIxQGM/6j3S4OxlO5OpJKwvFrls0tDTplX54+SYuoZgi2t/th0tkGWjIsdhUy
CWr8cmd9gUfoOtzYdIB9XRLjBFin8/R6Lv5k7Nxpln94D+j1IXaaIGyc1zY8E+Ic8fp2d69uKUBU
RN0py1M+WPd8DSqKXdI9+1n5YptzkcFSF/c9tyzT6CMVoFM7/OT/xXdfgZTaH39/7H0y+S1EGeD3
iJPgZo7GqasYTsljJmpq9we9VDaSFcFQbtIpkc5t3G0S1vgMWi6ZspSURiD2xOPhkO2R/w0bK9Hg
KE1Jzsxkrg85VyjO8QNOkgHHXElkGYeX7ZFLZn0anpZ+bsAvvdaDVWGiNjEjhJWAQsBnUpk/3F6P
E2z1RJG+piqYvdcXY9dOLsmmwgL67TpMOTXtDZaHXNs4pJE1iinVOw7IKHQE6kafYyA7W1XKS5KG
LkmT10BkepMagqSOAzo6+3MYVIdO4PEZ9X36HKI4HtoOVxbbQwosewUCmJX+g5Iwl96Ij4A6Ndtw
KajRrbh49jaZOkQa9xbjQ2KHCZqdMMZoPXFOkrsKs1jEhQNc01B4Q6CA1DukjTm5PKk0zOtxF8f4
zk/mRjtivfpiOPiveWVXJUFssoEGP+QKJ1oTz2f1amMrvJxTfiPhuQYkHiJu2q2JZH3nhMgK09Vb
56O1NtFxs4I/p4YTpOMy4oXTOu1381ce0CSaMtqxnBD8/IHRayqsjdqR2OKDGqPQU72Z/Picth3a
WZXMneWBPIGeR4Dwm+Ts/nnypfi7UYUju/vkYoRq9FY7+8EI8+2Qlq3L94uqUaOiwQ3lueJ5l1sP
KS4sMqCEWJ9V4KXPpC/ZAV1Wpd+NfOsEUuA09XCHUZd6BJz2O3pFrgR96wHiHb481zxB9RDOOwU1
XLeF7LZO/VqkvscA4VEnMTQ7CwcKzS75+KRdnSBSIPynske7dVa5NYD0crWB8qdcuFwj5YzzKrFn
v2Kxw2vFG1Yf7dFY1DFZGIxPqzWdk1SCPmiJv9Er6FZvOtQEj30+Wzajz/z0qO0EKwt5WmVq8Lsn
+PF2MwdDs1tNrsBSqcgtFYGns5gELUUvyCOk+Mn/8r4LNWxVH3D1j3foj4kjpE56gq4Gssi3KnKj
JSdHEVJtq7gZtNfA5q7CcIjzafMmuRlr3/h3nVMs+rsDlV2kckUxsWGeHFQc8LW6GIiRwhhwV0r2
0EDfnRcLcgaRDnSIX5ryrVo7ItCQvrwJBqyKhzw9c9nkm2xuu2cGanUQbgsux/ROVoQ57w0qcOOb
lZuiriacE6QSMkflQypnP9k3GEEaQFJNAx7l/ExDESDv3R+CCI6OWzPq8AHwfZZaLVFHVF/nhfe7
+Kf25tHpgm7Ttlz8ISU1mVYYN0nRBFz6F43pfKaYcvfmBexTVp+A+t/Mv00g2gSrQ+jXijjqYekK
Pgohl5NLDzXSOp7/StkNd+czNEIMeGj2zgbh9/xWYUaw2x7eez2HV9m8BIKvPsr+R1TcT4+yFhSR
lRNUa9uBGY0AXSIJffXfepUR/uzS/u87p/wApCmy0v8Qw+oPhikRGwYaFuoOGZibvQHYpXIvQ8jn
vW1G7NRQeUgHX27aF2F+rx4IRBXhRYrD5BJAhA6zI20C6Kw06UnQ9Y0ozZfTtb4XLcyc2HrG5djx
3AxSrIn/jNPqXX0/fuyYzNv1NmHej/xQ+b5sC6Kp9UrQFmpU0MdApSWjzPcO+lWXhavUZ7mQ+bVo
p6ZpI8YZeWBr4YvP+aieULwNWyBhbLW0Xx6YwfX8GAtVl5YHnzqzwmSvB6EG7hTDRMq++p+n3f0c
oPq+jTw2zE5Z4TcP+/9UdjoyNj1Yl9cxGwYzza7Qlec6xhhOP5DVOkw4GPSwjtyM7N6T5r5SaVW4
cidU0dQAA1uyjwG143zpOH2HtekPwbg+xDfVtPSoi0ZcdmWPyQJpoz2EzfAywWR7bs5QuzKtnLZs
AI6al6+SUY9QqaI1mauvzaLEpf8VG4sLVDfOl5SE2LMymOSPimZcZo+53boPnvYAbvf3nHGA9wv/
a8BBCHRelQeu60ObQEpTkH2TTXpC50/cbV/gvwC0pZX1d4ZVpC+KFEuqEnTfk86Nl4AQNTNHyh2M
OkZxhNMreQY1eqY6uhycdyx5AwhUAI+RLTJH8MjtTpJb0FJ9BoUJgcQxqrSDl5KR/KvdX+oOarpI
TtgW+1h5A2tGMSGNr/Sx/fddE/8oyEIQ44edxmLatVtlprc03xElIuP+MpYrIAGLGuwFzOTKxyzF
mdV7yZ1YBwKe7VgIOuA7TIKFFvMHnPhpQRNNsMxAoLLbWYq7OH1dNKRMIg7UfI9q/DMSTvsoXcHt
ybmAp7fB8pWw6ziqHwN26O1eOQ/jAlrWtormzVZdn+DZy9LLbKgVzs9eRB1kVCQycQjg9k/cohA5
hdmb2/FmoGslOJOreea+cEg3yTQdzzAg0XumBOKr6NhhvviRF69FO9ZoZgAw1XZdQajNUmSBkPnk
aQL7czyAFSvd0BFQYjxRBdynnPBBFY8xcHpC/l7oqHXoZFRkRFi6SEmW93sCVyK3BJwHqqvwwORI
CWfOW2SGReHTvlW40AhwkoBT6PdlBvwu+zwPUZPrKDnuNeR35QwEIaCGJo0BxjP2F2U9zU+Zps3P
OysLxoOyq2K8NwJGT2FEx25NUOricdKSeh6/NUUGsM/1VJoCodWA9Tdu4dguxNYYYqr6c+3Oko+h
HSXzQefXtGlNHHz2iH2A+vEWqzMNoytgj5PA484e0/ep8lRL7jU1ldM1+o1QfsNuUAwD+YRoPEjg
tHaHC51gH6kQxKqkMtL22G5yzub8BznwzWfjair76LVCqx3EMUmFUBoS98nwkQmUOmQEcC18XZPe
gKBAAX8h+IO0UfCyaK6VIbW7xDaN0Ez9GFDLjA1vAphcd7Mxy39hkL6Sip4xNFH1761OjWOh16ZJ
J+l4708/W4UaQnAtdT1EowrfNci8R/WnsesP7TdtLl6A0D1N+ie1VGgC51Y8b0gd5QboD8NSMu3A
Mm9Ci0VEzErldcQhJaX9yhOYssccLW4nKagg96NdDbyWSTZAzGp/C9qo1pSrPXxnXgfqfknIaIAw
xrPIekxgysyUXCuw/SdbyGbBiKUJmdnGsRIXOWo6PSO026hz9Kl7LjJPn/z4fipAYjWbyavZaAj/
gVNPrIdn1iMqhc/3MYE67JlBpOMrUgXPI5GbeLmYQ3eko5HOv60N17ejXYzi1hZB+OYpRhY3JgS2
lGfnf2MBxw+c2zCXBoRypbpNuoxsbO/p5qnBIZbxqguAScUEC/WLt8xwMSS32ygzBTidDcckXOY9
nZXxLmcWEsTbv0F9z//42n+NyxEae6LuRKlGX6jUoGOVIGMOZaPsL3t7weEl4BbwaFyIFFoP8uVQ
PK4w2BU/vEk7EiWORqzOo2/zFl9lxC8DWsEb0L3ZYNOrtoOdmoQf+BXDyF/2Azbqjj6Z+uoboODl
FNBXuvrHXPOrhfo/HHXPDJlhIEfXAw6pSuoCHwirwhokDN3aq/My/6yQVUom1ogsgF1qPg5diA81
kN7qs19V3srWIuQ0ub8n3r+dHwju55bO7/0kCUJRy+3jV8Q9+CbdTiFPALx/KEXsXV3wUxqc99wM
Q/PSXK6uDmNt5PtItA1FyNkLRp1MxqZMESt/wShyEDoOq/pn5QeGj9NTKgo6gqF//mDcDf7HGL9V
7Qr7deCEdSLxQiqO0oAH/XiYxhq62TDyfbJeBIX8I8I4reO7TUJzUd3KoPupaF+eAJXpXFU5/pM7
hX21dvDc3ecPLUF5rbRX04ZoI98cwjf38lS01Kfz+AGCyjTtCTs/9Fdgwe6umnYwn0S51VG3UkFg
4r+7pyV9U2fAJxiubnFIEtB1PKsRMJtJ2Tn/TSW8grcfh30PznOYtn7iOZuyCbD8M1Bc6LIUQZPN
NqO6eIba8ECA4s1lwAk77KAWdzNdEzmVX3+WkGzteeUmo3k/9WlBeXBWaV0ifrAnki/0FD840Yy3
xU6kpWO1/CV/SVT6NSekqTuxGWPDQ7XVPfZucmVjFQglBUtnuC9SWPdad+Tr4pUZ4N3N0weiPEVT
21JpngrITIJYJtn0Bz9vPaXiNOHQ9XTYC8xQfgWGF/DHIhQcXFIClgUSyZzBaZjhcWDKFgK6ZF8d
vulAULFRToFEIa8jr25XrYAbht932iuNbJX47nVg21q8hdDRNNh6IZ16xVSfRBARepOts8z4W8Fx
P41F504ZI23K8akZ4lD97WnnOCnLOK1P7DZTAuUOaiWp2ljfomjgRNvQuF8Sj0p6He66QyI6F/cJ
G0xFKjFCYrFKMLko1E0504CYhTBIG5Aun/fyvOfkesrzkgYg8qiBiD2m85iWbVEV0gqHlE1y7L/9
blg8EKyef10Rz+6ksUV9bv7YPWohCvZagV8olD39V55nWpQRDYhfqRtJKq30RDIn3KoxG/UnaLpR
aYpS/FsEe+IE+emxcP4ZJ3SJq65qE8zRAEwMTCJ6JMTl694nBRUBfcT7SYWx2rmOdm331Aae8//d
KiTWSd0S0NF51Kk98xvDyGIu0svPPPwu1KFoJOnZIu1c2peYcHZtjxQPT1nfSHNekGuZJJSfD0kz
2eV7iot7BG/qAn+yzw9/3HS608hH9hjLnvnt+G1q3o4j9g3plMMm3niKnBqVm4VdEdlLpJBpP/9X
K1BG8sr4F65sD8npnD90s7CKb3CKiSi5qnr3cBhCBSNk3AXNd1+9GoK8rv4F8YCaoGdksemaFZX5
HL5yFjGO9dtM6glOMKbBX+vWLFsID62NLpe22BaSYD3a8mxOpNL5Y5u+0p9ljbWQjM7k1siIvJDu
o5+45ZiGIU0z7Fe0t5ll8tvk1USTNItDVNP5NAC82jiFEJx5rlOCA+lA3l/BoUzhbfL/A8cEEQCX
k/NMd8nfR6PyVauE2dTolbMS8Ju/SF3HrRptAdtlaFnKgKTx7a8MmAUEJEiJBucVQqCJdA9chHPZ
M33mubN9ghUYSLTH1XIN15UTq0VMVeTi6U56OqIp1PwznwTiZbSi92yXtup3qzXNG+S92MwCyhhl
pk3OfKL5oSXfxTQ1mFmemRjKrl+Ua9wvAV1+yTcq6z6b9L4/9Q1j4gTBrf83/MTrjOUtZkejzqD1
ufgNbDdJjpUVm760//2IhTsBIwKMxd/2h/R8r6hMDZFXjOeMnXhEUWokjfKe3OCdMorTa0wXp+6+
vE96D9Zqgf4YO8U2Z8aKRggKZjsTwoTU6V7Euh9KgYvqIyFCCMSsqvHZksOqDwgLZds+eHCVac+Q
JCihUGrUCHAB48DbWIJbAZ8CImGsoEi9beWbhO7Mr++gSDqTVn4X2PwieegJnb90umUQDLxUx53d
PYiGIF/4RBi70fiD9nyGjtWZmPJTnb3YEKAUC/eSnODig30pqQ7YdJCdVGfM0ch6FKYDCL8p7ABP
WSN55tF5/YtCucpT3VeZ7lYfz3i9LCpiULXUHSAAdE8E5V+1/Qbq3xjMKt+l7hRLadWcdUDRosN8
yNXjJN+XSGDXfM4iWRpFNzZQqBljIknI1Xd5fyO/A7VMPeJwTtMvbERo901J7XMie048dHfMvUld
3fuLIRnz7ypkSt5m8lXph+FV7A31n9FXc3vz4iStQfm8g3K1WU5UHBzX9QiNPJ2eZ5fA1VRvHuWj
mOFzoXVGVumkEsyxcq1wIzr2eOlW4pV8YS3GZDGQDgZMCCR2jddsj5dHQ49TttomI7dTE3UTtrAd
I4F49U3Bte4TqaZQtF3cs3ZMsUahGVN33dezAhBT7r9HzLXHUSjYJOqD7OiT0Ixg0ZNsMlbBYHdW
BaQZOiWcRfJzE3YBCpiVv8ddpWzj4cTGmjcX+X9bvdfg/3ZwN8HIuYXlXUVgSbR2f2bGV+9RN7Hu
LJdodklWJktcRgvjtyEP9aAx+KjG3+MTt7YC/Mcc+8vrUZSFIPhBIGsM1jWpaHlYwu9q4Gar+Ic8
ofl3LLZUGXIVhHTmybzPBJlf1UDQV+oezGL8HUPyFoXcaTW+1XnJO4uo/yCPuv2JVIooEJbeVIF0
I/nsILKLcT2nVmpcSaMbcJo/X7ZqMLUbVHNDx0nNzvWLWcFC7c2QY0cqvqbwTlX13Vj4ERJCRmDG
gtZAZEPuRtLT1tqnaBCJvkvfVBhJrodc36Ggw9isqCWtexq5PqCljKSNI2pFcvOpe2qmkG1Xoh6P
8X8BSnLiilDMGTpu3uYPxvo7BHrPUxe4sJcpj2cVyGPVgiARAZMFhdoZyrYGtJ/xM+zSnRZH1Vnw
H8MQDiwSrvL0dRmL8S7vZaiPH1NTx6VA3BMoasvfwJRgVgNU+GvTzDJzGwWr9MDdy4yGt0Wvi5ky
0v9lxBKCtkuC3jGuYsyJLHIVkyp54aOoOsNXuz1V9Yfg9QWd+YvuQBPyYOMfHcOHIJqTZYf5oMby
i5enmh1D/ZVe4rV/BwsaW0ggRAaz16JEJ1N+afgyAkh9ETmWfWg9z1nA2fDv0IkGUTQmVpxXk2+r
3+JesRS3V5l0MEcbuEaosLOZzr8YZI1Vnyru2wWSFkp4j7GDb9aBN8Ly0tLwvC0v2hTYqdbZb/m2
nvt9Dt4teKxvHaEZDCwghP/HzIfXrVszRXwkQeMWoGt19zry82XdUVCX7oY+H5V62xAZO0vho1pE
x+9c13wDjKlaWZbvz7Bpa+bd2HftP1pWf8km5fp+jdcxWi/7sJBtVm+A/JJn10hVuk8S9tQ2Bhxx
itj2cpZ0lW7TuLHA1D8necQUgsJ90cFbvEOARvOijAhFsoCTEpp6bvnyxReAmc8py4CQbGWLc4dS
OM5N5844prhH/VMG4SU8clo1igskx2/+HrJdsHZIl8qopnMGU2/SpFsKVbPrE9KnPvNgu3nwTPO8
nzhgksPiMlTcrTChs/Z6jB+SXajXxXPxUp6lOgULEUy2HD4WqK1/CzNWonrxJor42EQBlxiM5Qk/
b4CYEUDtpwfHfpxlGa9AknmbKSmCZssANd1eccplvSUkxtmI3tHI0ENQ/knA2NFbqYaDZ8p3gKzQ
jTUHKAcFYLg8GYIvZbZgxnGgnJ3yXmamQlDx9fWBRkk3IDl+QMhFAxpoLDK0tstzGm2W1P8yOnRO
BwUHQU7jePsf2KznSZ375fTVoAkp8cb3ovIbUWpJeCPnt1qM8//L1CYXgaOaaSNG2MrIEhkPgyjd
TOytnnRelqSTAZ+H6T7f/iorlx+YSTUNEyurePIAjbKSx6JZ1RUy7B+zupYRAXrvGVKKeAE9QBWU
d19YsocibjQCGJuATfVWzt17TeCojMRVcZv5Kqo4YFHqMRNMVXbKDL8QCTHebB9PePpdvXCDNHBF
V4PxZ2FiLYulKNGpy/vyphcZHpsQHq6CPDL//gGI8Bpj8+Fg/xy5tEo2ib3KAvR/5l9RfuP1r5DH
w+t8gtWtIDkiaeLmYbfZ3oIqU0UMol45KD2OAuC+ksXAKloVpdXxTdJkbTQgMH2sxLtG21R6w/rm
GLW6etBja6xkmoThO/bi/H+uaqA3u+d910l0K2on+t0LEYGni7z+sJUPpQub03FaEMnEk2q7shFV
pWMbFXH2SlKvFujcwE5Woz/euIC+ZHRzKBrUl5GkD0V4Msai5rIc+AQx4CfaIybtBNk9p0Nh6xxG
SbfaQCQFzJ1ZzTmnD22spdmqCYfXVm9Cty13OPPkW3hTdHk89onvW/3WhMUTHxl7N+t3gvIlcR7s
/OSnPcvad7SJI2b7n25Btohki4Uaz1gw5t0ZIigBpMlIbz9lmXQLLsRMWhbWHb4OlOdbbLUCBIzX
14dM36rSRaGUQyrGl+7XYiMDfKQn9LbT14rPzj5N429cdcma/F/0VeIWFGFmyDrtiK9/MdJMJtW4
0cH0RjbESuwRHEXiXi4zuIAhrr7vxvVicZ1Z2e3gkjxuv+R9ysSgN0RTxuT6BKrWi8VlVhFgV8qx
KhraPC1tMrqwH/RlPWlOx5POzSu8ACstSAORjbz7nYnknpjronIeA1A1tl/fzgsWY2HLuBmMnOzy
TBojtCtbe/aZafDa51qDZcrwlaMK4+cDRsAwRdMj/F4uxOuzGNv0eRwI1xBxJRTpaJfjhjmv/Ke6
TXg8Yg4RW8BoHe/HIwZj0r7ba2go1BrxFtm65vwXreNuMDjF8UQxteSyqZqsTnULZNGHwblfPmpF
H8sIxO54nQLNEQVfoSakb28olmOCLaU3sZ8zQIePu9rcs63qsPBjMMxNU0OjS8Jmx53emRYeYyy3
zvBdBU+HmtHRmyD6P6IwYa/SMpFp6NUKzJK/B8CNGv4Rwk5AoQmuaOGVl55fqCVwbTk4Ie/zXH4D
n39OqR3LxCFMa9L3wvipsagvz4R98vnw6JNjS4EPZZnmjVufgW6tQgjnc7w1ihJdm5THowN9Pymq
Bqe/Ekt5AgU9ENb2Nbdr0bTGWQIo8nDFZG1CteqqrmQRuqZ1eUUNyxIbcPLNw+V2rkBVhIsNOMEb
SOgjWkDthhaU/Ob90BuV3cV1HetV8IUTSuQw1iGcV5hsQtVogEu1Beetvm8qWMf6tE0qfOh4l2n8
YDrmBF0RPST4tY91VcXmTSOoapJ1b4VQU4X1xHPDUUfestkbu83jUO6G9wPDJJPEiz+/nWHk37wi
c5lNsZLnXvP4mhu/xEicnO6EUzhaJcZjzpxqzHWgOA4sRKaCfb2gYOecq0UGq0gRE1/Iy5JENDc0
ZZfQl8BHob9tALJg52+k4em4ipB9xq9dDwb4+J9tnA3O7TNqXpXiaZ4763fD+ym6eJcwndmCA9a7
FKJ2BeAEw6YdOew2ON4yhRWTVbI4dvIk2oyYIR7o4woNyKxpJehEnavk/hPTsIeUQNZ4qav+Mq5Y
1uAVbH0L6CEH9emIvTZOOc4Nu9V/myAA/QG3M5Zda/GbHblWHN4P6o3TWELn+3sau6XEn+Mm3t2/
fFAad+pqEn7gkt7RrgpOR4mMrG4tSQ/Fjd+uhxQACQdSCBwlS1Ohpvuw/62noEP8iI0gX5yTFzJP
/+ZJsMgGttpS1V3pb8Uo9L3+hIGNqALUczK40RziBYWpDiJSAUhKqaIyhfmWeZQSOujryN+8Z7aL
jg4xNibaBgF6vKyqxvgiQ61TEPmQnDfMVioVrvlUClCIdnSQDHOA2l/0orNAqHIsOKOCJpRirNCW
Fh0NFcM6y35VQx+qfUqXDCGhhqrz5E30xWsKldW4t7sLmUDYHpeC/MImCbr0i8kSWt2dMTOg4l8W
K/2cr0adr7StG1AmCjajP1MLSPDzK66PBiq/cjfP04PkbKB1CJO17RGnxu8akPIMHCyXWBb5qybg
J/sfbDRJziMzdIETBf0kfa9t83/aKYkZOzadUt8PCVdoPWfZYyfzNAg0EAhk4Lzs8z1UElGfkYdC
2O8dfnJJp3DXKqjRYo3yVRJSu5jm9JT7dX/F/4SYQl0wIWppRVp5T21ELdXy77B7UVSQsjHVuwp/
9w9mKlogbN0Wq30ZrgDXKTHoODqg4A7deQhS46uAAlloioCUPj/4tr22oP2N8roph6QCjVqvJe5U
PdyfT0tI3hng//9j6hocFZ707oz8u0Bawnkw4X6OKbGrG7AgpI9RWOD+2XxlxfKia6KlelAOr7L0
y3aBTtYVh6ExbmhbYfDJ8oMF05reORC8QRoZ5/tzpo2UajEXbx6kKNrxThZ6katnRtdOLaCLBnTW
HgTdbDjh2wLycoaJeoqUCoHYTMjLvSmzbXfRo/UYJUeQ1v3us/npBLoTrWMfElYfwL4q7Sr1f0a8
mXQkh4NpVXpQgVzqOcTuUiLmDONKke2a+F/mjU3zAIQnvyfrgpLAD1AkqMhk6nzbOYdVbE6FIyhp
kbgxM0QP9C7xWWFpkqyDXC43M1wJmevMp1O766mKvzE1aOQT3QZSUg5wdn2Gny+I/GlQ0gkx2zod
JPV9gaBoHpmULRttyOLyPS/TObn3LaQ0KEpGxc3hCRfjQvjXEokJtb+/2MppTmDvUXC3FN06QAs6
QE/xYQOCkb5KoJxMPHATzDilkv2UAsTX9Fr9qViM8XBlRFYx9uczvTGGPy22c5+44Z8v8ES+OChe
Go8rnIXgW1y2C12rFyf6AcS8/gXCw9yLt2eWuB2zRrMp39AAe7K0ckZX0eYe+W/+X9Mx8FDDbQjq
Quz0daifdojQd/3XnDb7VJpCZ5RVKI0jie1g2iyUW0cwqxT021X5Y29ic4DpXAbfXP1PvJpkpPG+
VSiU5szvWABxD3EeeqsyZPithFaf9qiqmYkzlKzYW2hRc65bP2fOKMhAczuFSNxSogXvd+Mlcxjk
5O729gJGBVO9fNlVW2r4VhaTawD4FIksPvb+D31kDHH86Oq6Ehbx94viVl3sfplDeILeWjZq51V9
5ud+Ynwgya11IP+TkeVbIHYibaLbjgWigq2+0xIwu/13Mc+yHCLv4VXqjaUlYfU6cFdyNxIrY/i0
2t5fEwMPt68mIKEyjLfz+jppOOM3UtT6nTaJ6mNiQtB7uP4o271wgLw/CMSO9DyHHFf5ow6wLwp4
NmE0eI1uMYr3Ixd/ioj5+G3GBddC71yYHJVTUhQgr6qGmD1uz2RMdB/3h/QlCZVk4CWidyJwIsO2
QlOQVLEV3SiEb8Tng7lB54U9Q0+Y14tcg1dXsakgMIRvUKExzERbBeWu1Z61cFUdSfD8rFk2b/Mn
dwYhJk7K43NyM/BcTaCPPH2aqMaA8yXbcL8f3l/Gc67pwTLebh+4mzOZ/dkcigG6zYGXTYe8Cg0C
g+9flZCKxu2YkQRryhEdItuyz6R7zOh6PgCGPQn8nnttEbFqMmHcWRzFLiITICcZhdn/doAEfg+M
frSJEejggcjeB/K3uS9ThzdTre9pq831e/to6k/sy/Oi/RUiTfDTyGbStuj/KapZQzmoFeYBdN/k
YukEV0+ilvDLPtG7BI0WULbquY/0rj801k25lbDd9qrdJwewNvc1Q/Ve2NIYQ5466/ND0aBYRev0
gd7VVFeBKDTap0PKbXoXFwMv2+BdJZEkVEc1c67/jZxVprWcgeWFIaDSDA9ecfnlVq78lGssmx6a
IoGtcvNMDf4zYseUwLKeChR3Kkr1G69P0ZV9c4jMlpPltEHNwHg7y3CYf+g0G44khxkElAKa0ns1
u4K3v0GSX0olNq7f/iwB9EvQR2IW9OvEZh9cMKYvDcNu8Mxj9SgCY2EtXUWtQELe4ZJiU8kXWEHW
6D//be5TS6nCQBXXDSiB4R4Rpu/694nBCdmJijb5vPYbbQszsoF3ZmBIQOFlF6a5j04K79U/H6o6
PNtcN2CzBgH0W9i7UyYAi6vmTbZKI0yxkf0xBqztuLTp1Xe8jbBkF+wxRSEPMfgAm0qZR0YK9kZM
Wd0ziwzNvDEnJBJOBVEzsq8vc6IyZRVk5REIuJIo8TYekCYJu0gn8DtoVGIZmnlveR/LqHukPybY
FaCq3Is73KgDGMLckYYCi7JzXmuMDTUS6whUMV6qd6wDV4k1KlWg6A5anurDLyo/0H5gVLchTuVk
YAH0Rn87BG1aC/tGsLwIXADQIfvw9cXYTAyyv0XnZyWbSIYb2vIdW/BkgzsyFsh+as6XcVM8LiLJ
siyXmdq8R3nRN8F3/m8gjO+vO084356BQ6/7ctEuZ3iRodOmkxa7aUYE8LHOBVjU3mRoITPbNmLK
SbhKwUwelJ9KOqe55c6gcjURf8xp4ntQ6BXpcKtjrCUhZ3fmFeEKJGSU0LTMnzGDsYrUpmiRrg9L
RPdQMNePRSP1pR+Lrk90oQsmXrTwW9oEtcb3c+WGJSSUPW97RFZ4LJsEB9+ORsKKfzTXhYZlKNLe
3Q1tUN1LPZ706kq35SrhWhomwKpKFu+jR2kN0au+ldlohDn/m8+7Z8vILjMkzR9DCmbj3YnflAPj
FL7wcukkyIrVu+mXA6sXwVQrkPonMQI5fIlE8PB144aXyKcMT7VSaNipAPaA4OqSE7UwTYKqs+n/
P88B94mx3moGEfQ/JWsmUGzhp63bUFzPr+fN3b2XV1cC02oytauG8CI44FrA/iVkFPaIncBC+Qme
SYdyU3gMZJhgVXHnVfhjhsYnWElWnOoBqCcxQiFZaB82hN3x4C1drYL4bFRog0LJGHTL3mkChAm4
jpG6Oel53ZbT5uheVy7Mi2p/WZPv9tSpAW12eAY1uWWp/8Ygp7lRYbJMipWCPqgXFuY+JJIh6vE9
dM+Ii7RsH2f10OifVxfOpM1C6efYpjXYjCphVrdBPW1VoTY9w+y3CSz1kw81+XAWY1v4SlGZei0J
AjuznnqyetEdk2SzepRiJn0cG1H1yZGIAUanfhE7jtkhVrHUYHry3jzPDDqtZOZCabCSOu13AJ6E
NsDfEng6Cj/0ne6v93Q+rLbP6TBpuDSleRdsjs2sOsQXqkG47BPpzCD2We0BDa7Ksek9EYgOQ3Fd
+Ual7v73/8ans7w2D3YvtL9i7Z/JS6wP8f0LCesIj3oIiWM9GPsEJrJQ7A0KkoMFyxxaY0CZHH2n
PjKtBTDxV8Iga/cXhiCAjow6hcN5STaILbXAckvor3dd096T67xInfuZUhkUTq3VbHXJtbaJHNks
3Ve/5oUn0ppYNUdYCo6ueO1G7V8h6NhtLU8bhI0Fc6hTVwRGZIB41PTLqqjIqUT8SnHnNHHmk6x9
q9VvZt/dUfVajre3bNgNaJIH4jFTXzryQtERyTPMAv4G36JpLEYbJBPV0VbEvDF8dBy7UsJxBrpP
ZswWSEPYoTh6Thuq22ReaWF2VrlaokwTwcsZZfNTlLxy/BpDiW7qVbuC7yFarE0iGBerX23XNs+r
DtnsqaQzLzlpsCWAfaICnKNQ+jY0riQVuaOp/Iwl3NZUArEWAj7N27t4RWi/UMF0FMJcdacfCv7Z
BPpY2Lvh8zXKJn+sha9iuObZDhUMP+9l4uBY1noSQYQQTsyveh7psQbRpQGVIcDv/d8Rr0x2xktp
yIwjz0dbHDcoIT2CijFi19zAiacxmKx9G1M89AJ5S/eICerc8xr1YA2xf8grI4PTWZeIicUBmQCz
oVdNh+HdWpw/ELl7Gz66N/43uud5xp8++sRKoqqddgD69nxGr3Fc7Egtu784FPmM4EXcWNi/ELzH
kqbhqluVQU9j6PlSmY+D0rZ4lTuFtta0MTy1uE+mHuftzXUh9Vrh4/xZsMyBQy1jwlxkwn53kXYv
jJnxiojC3Cq3rz/CacueggBCGoWJVBUehHw9jTzfqa4cbzz3ah5EpGk8di9yUpdeALZ6xY/kBBvS
GUBRzQ2njUt0yyJK0mtryAJCc9tYuZDGc0r+SGxCVfClIfgRQoY1nGHYqOpNjkbLGO2r5eRjFpye
YUH0p3QZXszs5pENNk6tg6hK0NJsfWe4bnAL443epWiCt0iNfhE+l7fMvMXshYsV/SnLe8Iuj67b
tpOIp3D4gOa4TPI76PFXEUu3Qi4kZu5pVCIEwN5QQlv6KO+vPSoiEiMW/HpuUhb7c928LXwOgG/z
RO8h65wDS/VicLENo4MVzvLPjgRNeRlYXgGQxEtSoONeiz49O/19Oi1Lzi1MoPI5HKRDGtJEGGS6
w26ZaKPODYS62frkOhInr2vkKjLFUxmv7E9KgaxVoiSMs4dC62lzpXEO1cj7Ehxr4nB7aFprjo9Z
WotYdviLiIH46zzxa22Wqg1mfKfzNHcNG1YHC1Gim4PaEN+tAX7LyC53oQhE2neGjpAIlO9BV9/T
JaHzY/yleNwQGSN5VHEIiGB6L6ZdktA3ppdA58NJCsLt80WrqWrgxlJeg8dTivenC/iJD/Ss2IrY
iWlAzZm6ca94op8a7efFeb6B5soeTp+mkETZ/D0o36PvGwNvbKUMfmWHarW7vj0C5J/rKMXnB8X8
eKVPxoPOMStqj4fhgAvOH5khNw0vDCyLkodQw5jIeNEa8d+4P1XG7bAcZyATup4Dk9DnKVl2yXXc
9HRKhAqc8qKRoOFqtc3ydV3Xu0DzXltjyRvWTPT7xhD8DtMgGcr68X+l4IY940GZHc6stfgWGTzC
7x1bYDR2dGqQKYTI/fccThS4+Bz9lSdeXOyFb6bQSLmErLCg7ctoAdEaYCGqEHtUc8bciePXLxwz
Dy32r7a03DGuRjVMtKLOXd5sPX3RdmTPMeXUxcu9biSuz/kI9qh1KG3hScvi2ynYvJSejsz40oK6
XeUxr9+7wQzICcAMMGyIU6BNR4c9stRMR/nt+vhW98kfd0uCLomx+GcugDPWCtnChEODeHH0O1ys
xGgOkdw6wdGuFmSjTO7p2GRHlFdZYmjNQXcQNghBRvhWacxk2Ho1AosOAZxQAJPX57stAXpGKfd1
tYFNEnIgt66vOFVl5HWlwfh0C7s0vvRNgR1N7VfDxxVPmtPo1M6vN2mg2eohnn1gC7cKMleKehg/
eeNHe6N/UTs6q7Ok+X4dYudQmSLh+pzVfmdoMxeAzH7Mwdjop6pPZ2/U6A6qTdjwRz1nT5DooSq7
T+X4GDVJJDCtrYcRvtSamY2o1DtnkFM8qkPn/KGJnAUTOMQiX0rQMa4TmvgdTobAuM8h3fVfMjf+
JGeXatQTbPDRR+Bw/ChfGwEnOhA6NZWFVOBc5NMD1rF9TlQza4MRjuhfANy7kGjMX4qiZ7TcmXTi
4pjSuX/3ShL81EoKxtUoSAvFgQVuZ0hEwSRMb5G0lDf0Q4jIdMXQ0IfcPk2NbLoZDDKGa+g5MWCW
C4Ru2e3QSuP0aXneiuU0Kb6DCVNXBrK0a9E+vr5+Uh9+X92V99Gkr8mDCfWMpoc4nKBIRcI5ghnO
hbq2z/SMbcP32tAg1V120TEs2kBffPrbn95t0pAbOn46kz9kcJPzTMikPIIwoQPqCXuDel4yLMOx
DjBkdNqRhSf99Pel+buTwSguc0qVksPRF7ip1lbvVCaLFG+0ZYnYcvwzy/0aJYcsGNSL/lBIij20
QFC8SxReTPPpIMwaR6HBJy+DuOnhZBlMaKty4d8euCKAQE594j5NCLGsnDX73GvWWkMjznyGeBXm
7qDRZj9U4M85rP24vbjXwFlmaCjlf8g+XyTF0BSkurq5aMqvSCP3jCUmNUXdpvgfJSBnt2vGIT5B
QgCKC42Xxi8tWu4Gersl3w7vBe8gpyteJPBwgpjkmcZzyBN6OeOyuCJS0AaiEa19laXH5YYr/65Q
3hnO/u//qyz4hFOjwo6ZHr6U5fP0PyTxdxfl83KNm5VjMPUmbT5Ai6GOivuiGWhAX/nB8g0/MB++
kUL6jwr0GOPflsPw7+4Pwk/jA8VC48S/tpjZKcz2cgi3n8rWrXSGQJ1bO+HLgCV0vJ80h4MDVMnf
oU0cruC44Dxxj6mugjh5z3/KJkDWsGX7ZaeaoFb7KTB/yJ0XuEcIuWrHrYL7vT0pa9yrX2Opb/z0
EB4qJ+o+86lYmObSotjthpoBBZzdU9LaB0rd32W7lxY9WnI9Pmw8G5Gkr5cdoyuVwdyVDNsfNJEk
n1piz3tvKpwec0e9zwyTJ3cxlzeI9NgPR0BOBkmwZJFjGsz3xCI0RYKsuUYTiHKk5O4kUO+VFmAz
W0BH4886E/m6NSeGLnuG5L4ibTtv2nX+dxExWhh7gnrDXlMHsc2j9xtZt6vy3FB0u29e8tJ6NdCx
YWRI5Ddan3ImpP2ewmf71murVNQOv5gMapqSfaLrQ1qBw+abX27tJ7Rv7rVkrKB8Fz5kGjGu698c
sK6J1P24UOOx5L4Ng7PmxoN9ESaFB8X8yGK3X5I4Vh04k3/sh+SxMjeQVGfgsc62HGfOYEvJrZ5E
Q9MWJv7Rv1l8vLPLbG44sdcIDjhUuEYx1qdg+ULD06lKIOichdKZYdbOFayVIPGv0R1OqK2t0dG2
izYG/CKaOlfKFQQfN8g2sS5n05RY0oGOPMBFtW0vUNIcqas4rBFBRyL8c01Z+zdedPGwuWlnl5Hv
hfwMR8g+uTTFCb2DTKWhsAb3cFZHb9iUAsNlULgUJ3ID5TG6qQb1I0BAVon2yHPiAD8oAeuYRpNW
QOLKlG2vLcgeLQB11Yx/BcayqwEuLhFbCItkd02XuTavnypwoZN72n4LvN2mpliSBsywgTcJXBsm
toAPX4PZVBjqVuMQ+NK/UovYtG3s1rKiPNW2p4Znt3JpYvBEhxwvtpiQLK3de8JWfXpqogOJ7E7o
JEIG0BDj//8gmco/yt+RNVaXiEljHPvjYtBFtiWwSf2rkg4+lj8ZSr+w+mbe6tlJWtwsUSrWJ7WU
CvK/HksRkMhqcKpVyp2sdiJKwyKS7vHdPH7R5VPJZeFs4f08NGf+E4XsKtyxvM7AMIWuHNRokzXg
re9RieJ2rtG2xXBhwxnk5nkVyi9KiL+K627fYAatJAqooIsCrzsGeecoHnIZCXyjABcnsBHbB/hm
gB8XzTdRzOFI4HNjmI3Af6oIYlxO92DbgrUpUrFYwSVXHZZkBsWuyo9kGz73PSxXyHOMXFsRzQf9
iwcgTM+z77Q1/uKGvObuOcanIbqV3w0G+DSFEVZhGbf3ixnA7hQdmlP2BiWUdf3RBe92xcmKvYUj
P8zBQYku4jIjNyjwv5Wy3JX2sYdyjSjaJik9rNL4DOkt2o3EQb4EhmBuC3PZCxrtrp5bnGXDBMiS
tZlHE/52b0mA55Ow4KTYZ4fi87EIAwGDuFd+rFo0oEIFKgIBUjLivupOwNHRMLRb5rgY0yk1cpAJ
oyiQEuYCyT52Ygi3O7KVfEUT7edDePWkGBl5uK6FPH9pnjXdwZGt4pLXXFjljOzeG3mYXl2ggvrW
DhG5OaKwXahOC82WibQvI5p/0Wh7B9RG2ogE502Tl7FGeqH3U4hTb8YdIQY9IAZwAxmwTvFFBvOm
PVgAbnAiZjbrScjrPYW7eOwJOFfJZ7feCeCQYVUAnR/Sde2/JxTLO/NNHBytmgwiK7611deSUMy+
wiyI5ifygq2texShHxA0HXedW7fwubmv1tgq299FJzkZ29KUA7s0P6VtGBXKfyzHeDWD6xcAn+xd
LrqrAYujY/ajrAtnYFImCdwhVN7sZSn+7qPuA2LX9UrCrGwIkKxBmVSp6H3TnOu5tG3kbVCXpX/3
+3MfmPHWkCHb9KolH2WLnybp7LIXfZ/lziAQVR/dlO8D0xEuIzi4FspG8XDO+6JVt62EPTfP9hXe
Zaeiu8Bje3K9vByXE+JqFLV9cbKcDahEkZqDb8p8lA4KRA6/sDGXQUgWFcdmtbs6/CtS+jspSPRK
lzV7yzejrNlPzLLbLzDVE3nH+aCGe7X/IkuW36SxkAGXvFrce7lrQPeYEl0KBGgecxaZu83Ak2IU
/wxUxLWQy81XEazhzV3sZU63fk95IRHhdm+2+7CwY4ZcJ1B4m+xGThruGJBr1lsueGOpIpVvUH9h
s60LU0zN3yu9+DjTszbQ8j3lOUrrGTfOem7LMCvvXwN2bGudmEDLu4eHX3YzmloVW0OriRjqZiLN
aEGeDTopcu/krURP1L8GvNKLMM3WDM94MMc8bVE1VUBDFFaCADwze6AYl8EetR/h+D3X0Qsdv/By
wD0YNUmo2OcSlyUVPbBB/CzqI5AmIN2ecfUzc6fMY7FoQbyQz9BThjYrhG1pZnmkVfgWcFnnQnhm
ATKUWPmWGCsJdY/QS+A3YvE+n/S7WaXxFnz4iZwSHp4NwMLTMxySvxSb/dBv3Hf7t+qd+qNoQCkO
3+vmdrFS551ljH4Ak28ehcd/kW2Jmea9gzSdV69IaN6VOn2IqLw7/eZDWdafApxeb/LNejifXd2R
CsD3+lPOcc5n614nnr+jxUX8Aosa7COOGTl2YyE2Jx96ZcFmCzrRt7CvuWommXjXe+R7QAruCTHP
nn4b+ptieZJGq/6YFYJGF2OWV3mlRzSUeJMGDmV2pzXEDR2IHxz2e7x7L7JOqLuPTrP5vtrgpUnM
2dj5zZpT7GfAKrxJ7/jogV0c6TX95cVhW13CNufCbycekJwRO9hPCPGs2r8Pwg8+C4ZlLKTbbF0L
T1r14/UQKSV5G+RcQLQRaszz8KoCFzpdZs4htXjpoiL/vqwGRDuC+Bb1poO5pnMqU8TU0cwS7AOs
PmejIfrEU4hdjb6UAR0owKAyFvRKHQ1HEcAzye9cmmR95amA2Y2/EAhKbBz8/vOSiZ3G8nQdEl1X
69hUd7QxCbvk+g7q6fLSwCzWXFjwZTDhiE6SYiWHnab4MhhhwDQcoGt6zLvTudEICbPsxSYm4B3C
IrHiK4dcTZTmCAitr/ZkwLneo+2ZTEsAY2a3f//rtkO1VKETQtZgTUH5QhEOGoM50iYEkkGrjWNo
tixUckf8zG6O+yZz4zNiiOJImXZcEnksCSPCc363bp7biQUPo2otzbA/d+qtcTXH2WjDEiUtyp1+
OC4Hao1NuqGdKmyCi/vkI809GNeP5xneWuZ0vZrS1lA2g5xFrc6q/wZxXumodeTkf9rLfUMd0I2d
P9qBHE+mGq0Qjq5jKjU9KTLauds4PAp9Zvcd/GNQfPnt/snmOSKR/c2wGNkyIZe/AQQnM/IyAvgC
q9TVaKrqgsBimBffG08+MHtQghFZKnb+NnoxcXJCHauLGp7Ptup8YOfN8Ww2K80I2K9MIQKaJi4T
qNjbgYJm5Cjwro2QcZ6swz6NpN3Dc9QpxpH7vgmWkJM8oFcdCZBoQtF+cVwAAoOaJyXh4xSmaXDS
oG6zuPzKEaNIMspRkYle6n1cdxDAfJLGuiO7sWfd6uS7FN1unyMe3wHpTGlfsr/JoR10mL2Ar8ne
XNUiVlc/D8J7DIQd033+FWkughD5VXFP3AJ7H8cF1XgwMHeXf0OLpmxBT0aljyN6SYOI1hfySKl4
sH2DeHj9i1VBisxAXUmO0wGZnHABa7gilFv2i8EAuJcqb0vB1WtCOwwxD0Sb1YmB48KQ/toC5/7y
/aUCOhiL270cP3Hc/Gso8pl12lmLeXPNT8MWyliUg4pgj3oUQ7LOG+020qdzpO3J6BqmJvJ03Ich
Hfk0uahWlu6kos0ApuOJfkyVQAxfxuAs7dXOztZ8XG2qkl2OUDZ/1bIde4owD0YIPizxUI9ZSYH8
DvzY5mdqTlq/4TfVlIm7EnBubziPBbZ5Z/nLYN+3KOgd2Kax/19TekslZ2s52ArHEQECGFBUVk9w
UC0BvOTgBCHkEIblM2s2Sw+zlNofm3rGsABawAQfT9dcUhE0HlQF5Ii3BSENvaNJLok6Giq5YbEK
4xljM8xD+/PtP1eB2YXwkp9fQCJBI3kjsKyAlm4fyoEDNUXy6D4a2i07Xi/Gj5YsLZei1VRJ7JS0
zn4EvrRdwvpVlF4Y7vbOcHxfJ5rYpk0WB4e63VlfoFuCXiB7lskyWjTs/QgjNvTmqKAVwDzY4wc3
/HaAwU30zsCZlPM14wm26OkMvRsi0IEkAhwi3CfaR+REzRlVcKHtewnWXmbYMiehkr4NTq4jF8uk
9cP//SsGbatuUZRoTN7ZNCC7+X3bRtgP6FfhopVPIcMdClWmBEaAEJBPS7iBwhZgaL8EgVbODU2l
qGB43lEIBH37tUBs0dR1JjOGEzy7d1Y8FIhC23JhNCyaRpL1BFH6OB1sSZtXEtRn+TZcclD1hwMb
ia5cjOsR0FPNxp5aAHyFeQFZWmi7dEBqjVUubOMXNezbe4JkUV0jShXdH7nYCXPqrrCsxbkPJsf3
EegsyiR45vaWTOFZobQ/7h9obtX3HMTJxHDqMUneFoYet/2N6kMJphg4RKycnGyf0a05c5C3Jeas
k4rmM/uTGDCXI9aQ8fDyNkeCxYswFLH20UPP+kE73cl+ZHgMRWe+xMFefs67OZIfTt/K7h/jlwbI
7XOzDH47RCBshRNgacncQ1J/uoH6DoG8sH0ev0fPVbRaZ5EWr2/xklRVfb+nF4U/mObP3ZddFx9y
TiAUVTUEx0RSShZLfDFo2zG4ZtlX03z0TNGvvib7e6Owl1qk4bbnlOKY8wDPo98lsXfMZfFK92lC
7zsnTPOe4PtH6CAo0FK1+WFeTN2p9aMqFJuitGMZVEg+wSPos9cCf91uDTliMTYje+iqBY5EE+rs
74ZJb2WK9Utur3d55furP3PNdgnLeiRKDfqZQXLqbMRYYuK0GHeEkZnwTdoHh5fAJyKVD8g5WptM
B7uPxpwLh1FjP0p4EAsi5/Q0vw373GvuO06k+mWhlnJ4gWit5h5Yp4EjEnCaD/viTtmSz5R5ftJI
gAgqgOQUcyXfuURcyKPP9JvYTXgSc6AR0uj3TFnaVKgotbPIGHwqQaZyWjNATlq+AlXF2/hB4wpR
v3DFmdDzFuZiFh45Du8vgxxrkq2LqJ76DZPwsjXvZfXc06oet1RBy/JAQdh53l7ORjIZ/hZcwd3/
aIMqa+LJd9XepLs6/dAOJBc681cbGoOdFMZy7OFQYdpWKUlOk1fxaCjnobENQc2mj9OJ51Wrh2MU
LQhhWSlnkRpSBzIs6K+QAf6SUz420Aj+b+4MZH6vO1rCKN6R6UoTzB4GXivqMdZ/9L+XD1IgXND7
nEdlScguQzwDrxVLdewoM3edn+OkJ17s2yg2s+23f5QUoN3FKDNDSbyan5FfYz8NIzAjQtNcIBuA
TTNf43JIXHC+WSpVLks0qturrGZ3S5uY7WtPwy61sw1nf6CeG0whhaC8IElX6o5Vydyor8O9t2cl
F8A0FEboEtnS8cSKl13/mWinl7s/8yAx+hLocw+Vlkw0wMOnReHHKwuJALbR5IH6+CVfGB9OEsEP
UdtPtKREAwP/uYieBDlxOK7c7rC2bom26gQKq/bhaSYvMWyhwPnK6s0jJAiqFLHl42rZpVFW+5++
CgHdTVc+HUL3/tNe6ZWjUKDXjJxv3yCjbTSoxWkVTs/a+VNFXg63WshD/JvFsO7vjey5FQ+Q3VaB
oPyYLGzHO0zmxAX3lg82g3/xNaDc7DeWzIctKOFA8dR78WY8ii/CaPLwS7LLwxHEIvo9l4kaZd0x
arotpNAYGcBYUMQbYWWuRWASQrJZe/BIUploeQwdM+1QfDJ3HNWhgJnjaJgehVKVfUtn5rEtWJc+
McEbGuqQjL1lFqQmdcNpZVVyxKcGEnMDHKTldjHibeCHYPsH2gjRVTGY/ZGmcHe88g7hSvBgaHDN
dNHe9nAOuAiDXO7yMIK0DbbdcP6wYi9Xf/erdAgObU5FyjyEkLVIrw31IMZC9XLdTiqjVWM95RtM
5Lo6hKas+U6TNL9cpSkKe3wG4Hd+VXW2I8zMGTBHHY+ee+1d397xzTpvZMbO6yodU+oVbRcgyrzm
+QJXZWAtGDdn3qixQros9WIOsDBH36byAAxfGzbKbajMkHuSvtrZ2m8dE5Ji10dHDW7WfXVFEcr7
H0GHwbOARhJ2eFz5dItrloHFi8Au+X2VXBunKm0gCFVkSIdjPy6GtazN/lk57PQf6wHl88IpvUMZ
wCK6vVXWPmeg4XuwZsPmaRLcmsHvIrIAvf34+YlPjpaB5cCt4Gg+G7PA2VyBDxWl8CC1V2j1YV5S
gnUlVokeQESpPWP1wvFS1m0EDcD/xt0HQfXUp0t9IKntMdTPdt2ybqOUq8XA4VlynXG3ir/Wo9mD
jYceebhTmG6dkVTlpl16GapXMVzv33BxgWmR8nANJCrTURG4P54G31Id0uQPsEweWTbACuLjrBy7
5ZKT/a2FDeZB3AoUR3vpAwNua/Gx7VR09EbRbiL1d6N+Py7WKbt8vY9rOqdZIrIuWuQRJBz4rDPD
xwpdsGsLYoChV+w2hd1xlrgszDjLC1Q7OXnYhQjpZm44Vr9eQlwrVFLq1GtQ4Vc+ozn6JI2w1Nj4
22Tl2ucMnhNiqZ23Ev21DUD0mTsBBJ3djehdCKclN8xD+IUP+NPThL2Em/Z3AKmzISsIc6lj4I2m
fN7b9dyyHdhRl/reFa1Yc8dzrdmh+L9SAVGD0qzgpLSx3mTe+OMvoNwT1kLUcNugCktIC0rvNWDg
XUABeSJiVSjQy2Qh2UBzR/u2xoj+2ydz4w6C+X7GMgufKf+MkMy3K4OgbaHJZ/kdVx8G2lQsMZpZ
o6nBK/IeJnLrGU7rHfM3qehQxEL3F72am7p5EBEGKi4xOO3wez1IboE2XCAwBi2zEkbgm3D+/f1u
qygeLR1xtH4ZJlfhIiXCIJS3M+ufUNbeqtlc9FTQGeiX4aeoFoAHhFFZPVW2qd9XF42Pc/EAxkVL
/UsQ5WKJiwwoS3n+u1SQyGuiUBvfVD1V3lDUZAztyGGrGG0AJ3xlwYLY4AsaGZwrrYe7CJDOS3TA
wsWjojLpyIIAojJWJ5n5jdt5U37AAia4DUTgalOU6Vii6Kn7O+RBuV/uLyRRCbRqudQh/LsX4hhf
vp87vptsTM8PUYrIj2SnrIQN/aI/4wX61txExZF3BbNNSsEsCGMNf2hDspAxBWiyD171FuaLemwS
gN617tBRMMqfEEnbToz4zty1ruWuF3/8AD5DNLndkHWSfWlJGm66VlgOAqwnTdTGUSczYROrudva
ESfqNecYMLIWUcGLuLilXK8++FtoFTJqmlIlvCkmwY61TtGfnbDqUqJxzE8g7k98uyJ30GLhq+K+
PI3TTSrGl7+YSoWHj7AcFgYOnfPnnS0HhofFp5XcT0slciXuf8lMfH7AdSTejC24YEaup0jMECNn
H9jYpjr+4UfdJ+CU/xFaVbG8ongXsW3occeYORDvkoHzTIsNjbzpu+5CrFnFlgOAIhIj1LvPCqGZ
Es7zfvN3hZ8TDQwv9ndD7xUgfCLoGKaORVtMmcHUwgxqpaB1AZvNQM17zxsTMiw5cYim280R9Gxq
fp+uJe10cEE9w25iKtn/JBNludsfLhYPkbCstycicn2jJKAX0nKwLyKal04btP4QQCSLXvGW0vkV
gwB90dDZelAMnYQboMoCxdjzoPIT3eexYzA0TwqA3JN8o2h+rBmSwpMA2WB5aL/I3m+2fiCWCOGW
Qgbg3sf4gjWd8dnYZKCsv+TWFk8+TytocazAsi2x+hU4TGGOWknjiAAwjQUU914QBmAG/RX9zO/5
SRNgMucrwETGFPhHu8aej3i1GIK+UUqIwLyWTbWEjt4rjTDNZJLiUwC4L1ojcXziIiOyhlM6ypIi
WIVjQ4xHp1yVMcJQQ3GHNuO2/8vA/gbnu4NqumPJWjbhUGNqYe1XEr+1QNkHpeBUsWRt+y3y048f
vytNQZA0lNkDYKVKPZcTgq6YRtj61vWwxzt7jp60jtaXemMuqvJKHihekSHDyjdyv6Rzfcj0GWGu
YdIaCBYgdpcgCTcl8t+fRZl+N5rlez64kzPlWSEkAPjBzeJTipuqgTwgfklZrVhfU4zhC2Bitkqr
DC2iQbuL55HDIKnjvvOVorENbQ3rARKVTRTyX+tH8DPobPRGqCBzvRGcfCNBh52MODW5BWiOacHF
B1it4DcgHKIjYBzTVAoVulJxUnzxZjvT8mCI3JiqIGQEcc6n9gUyyTx2dUCtknFkBcfhTLHtLqRx
P/GrLsicSXnHTN613U2qSU6UVCSL2zeKSTt7OV9PGUSM3fdNgkII0wjARSfgSUFt2m3rx1wJfiU3
FZi6hqfU0oMe62JrQNOHHY2NiGEM4KZKtPFm8+HX5W/rasBYcwzwtoacGJPdMGa5joiqJ1XOsTTG
8O5q3n1V1plAdvs6c7uy9xu/zXPa8lb/XwJZn70hW3yCIF4zCJ2E06KFnYAOPs7zJ0oWgpTF6mt/
awhLueTPjmM+64g26wSPx+u2Ygqh51fHv8ynK88EgrWhb6VzslOorVyivoL7EhnveSAZg38ITksl
5w6bADb+k1x83JK2daveO/DvE+MKr8VQ2v2oXFIlYP2jt8cXs0vQp4JO6PJOp3xNEs1/yfiOmiGX
yxy0CdviMSny72FkNETMUm+5q+Fgi+flPgxqhi16xo4WpBQdyFK2h4PYC/1ecBsGZoHo+/9cKfQy
ch6EZIAK+lL6lGRcrHtrVPyqCjm+/GzOLG4VLSZanP07Jkh1dzzV9SlpIwueWHGXJneY6wxuVsks
3SFg5RWIryKnTZz2n0kjGTKoUvXyliw6HikH9msnpvM3n8nhb0ZL1dqS9O0tZ1724CA1tjEbhCnn
A3NwbtAWGxgU9EWxXnf/astgLJxfOK9txxCP8AEVGY256J5IvJSdlXWFtgfyMizUc6hrFcFkQQYu
No4tK0p8fCSAj0nbtW78euyLqn6vtuP3VQbz6SIUa30+w1shCMd5Xp/xGbfAGKXiiAD8AYbXCBOI
4Chop3yEvnT+ynvuZtHFWZLmOEPXa/KGPAGBIWm3UfrKhlMVOJZXGPvfAxo3gXVJ/fFHr4EIVt4h
JV7XTUoaXDWvt03GVDTzDJgAQrVTPEjVkZHpxIp2cMjFP/MwoJsnUEt2XDkbsjQejQk9z/VGrLe6
VE2VY2m9PNdXcvaNFKd3CoN8XNhFOIaxcVllyXte0qr56+mvATntJMhZ3TqrDB2al27zMBLR29Zo
oXt494DZqp9bacXVljz53sbUqb++fZa0hc4ubW4dER3/Z5cqg/IhW3DH4bHr9witklGYYByRgm3E
g9GJDO9kgrPr7vMi6AeduBPY5oeFCa9K24MxqwmWq9Q+pQPU9oJE+g7LIBB9HirRiE1SE7Hom4+a
Fvdg0OiPTrVAuQjGehVZpD76mQ7e9pYJPJWRSpPbVowRfKne9Sk2v3GL5pTptfxzdZBwGgHRqUNt
o0azhrtuEF2NCq5LnjdOW7SpLtZcWvRCWtQZh4epYG/XIq1UK5u515DA3p54soeLh5Js5xyUr8YH
xhbBX2SderGk3ij7jKjdogE1htezgHL3wHRNMWp9vK/VZfmvnuK7s1IhWTerET+1+rog5gjmJ/kc
Y75+3I1HmIR5i/POv04/QbvLVsU4ufCk7wrAo59XSk50OofsSBaKWszuWbya2F7Z7o13Oqgg+elJ
NXJUYMX8rKLO6dTUd3iG5EcwNhtJtnMypo5Bby0Cbw6kxX++BY1L2vJC7dHb0n0dUMB+mi/pRka3
L0sb0CaBWy3Z08lm+gtdvjVL3+mWc/Ap+ibp0icSdAWrGyF3/bFROD8m9Alg5af8dfgVwLQ9CeiM
4wsaYISwoc8NZ1o0VkMGz++GnPo8vFc3ThsosHhccwLu+l88M/OOtWIBZCATNmGBABZU4ykt2rKa
egorHCuMWxuC15cWbVEN1U1tkHgMeCF+zVegiRGE3QhnynTygCeUrpmh54tbeXaeFCg03/H7tALY
VA+j4+dMuVwRzeOtIXAggeC4gUDh1ZslE29keOJCa+7RUu8J2FkbiMFPfVlB9ACjg2LG18DEXFqd
t9yDFARqFBUlOtxtjOsTqtK3jqMtd5y8AkZjSAEZECiHDO43B2iHvQpV+NhuQcHz7fKjaapxM0qu
1xlIWBeLrlWf23/8czarTRqwuVYEsN9adqhE/5R3d1gngdUMkRq+XshLCnO7wlTLyya8QJpNYkYF
zyGJpR4gs+5Ha80AzeWQ0tPdUjD28E1hFTVtErvlR6+az1PMTks62qWZLVEAcmbxG6nJI+dLIHXM
brDeuGAFHhQEMoinrthf7aQuRxIt+aCmRJCAsccFTNPKZW7OjG/YtQRoaXcQcRfHsd8zFOhFQsLQ
BCr9543k4OmHKN6eRc6qz2T+mvxpdB54a9y5Wn4Sgvqp+TrMJl6BUI2kxtQfGsIpiNuvQ1ubGlpj
kqN7SAUXar7JvdoW2C07uSyEal4FUOKKAUBZ85qLxUa/+rad+whGJKKWE9RVgs3jLREZBuRSohtg
nuWsjkRz7wQpMQZbY/wcHhZNPeKP7W9sM/hjHV1KCtfvKPdKfyMHZUR1lhyQ2X/mXKd/xoJn5Kzb
rPJtpnyOadHgefXWvxS58+Wzkrim4YjwImC81kSLNRrf2dq8VdwwY4tRh2lYpTTuTVB7A373acIw
OLggNnt1OBLV2AxpcGo5J+k2i2MIe2Uzux4076V557Sso4o9mNeFyW0zJyMHUOCcWCyD/ymroV9f
Q4itcwy1iax+hBbiNigu5yymyqWOhbOfQhFQWYyacUHvUqX6/gCmBFZsKM+F770ZY5nYtJNHsBoM
wUuao/oMHwGPqdIXdPJ0QCLPQkM886j7OraQXnj4R/UTnzuOdtS4rmRt/aH6aEhl4TYnC07wOzhx
NgoHkKk+7UsqmX756oq1O8/kw6DrztmfkxT2LsUldEAQEgmj1o5PU3fh5W+VvplPU5hQyVQVycFk
OxD96UYXeWUfzXfvEcmsg+UujF7h7s8HEkTLafxyvGskgHDlX47WS3N5qjc0e8VqFMuHHEXyvpwQ
1HgPaOPjpxjQK+fpS0e4g8/Afar+AWsPQP236nQufSmj6c2DbWCyu7SMNpIWApwdjfpRDybDyj6T
/rsluZuk7gtS+PJ0UMaZm7bNekVCQ6d1YR1Vc4Xl9AGbryU3I/iiRf//EcRkChgN0kPM4Jq7hKOn
dDHKnUuZCgf1TSjhc8WEClUOcV9gbewR6sa62eODkPJQug0FJa5yXbDuUqCPDo+vzip+gBu8GKDf
RzxtV4W1oKFUmlqdlFKsuTBkm2Xw5dXtwHNF8n8TM4+Kmo/FqHhjGtcg/EV/tTIGJnBEokLWQDlN
/IJ4usRIgPmRbWUbuxfNhDHfkVwfPvqI8zHJTDpfh7gszkuKjlOKosrKiFcFh5vmXbB0jNVHddF3
ahQqIrYfUizTxsHrsOewxajirc66k5KtqvGXjX4zR9AIUmzDMu+bgUjkpFIALjLu0CsoXG/uP2bx
uWTYTqy1XAs38WlJbQ2Td4NSNBcUaY9Iyp9tFuodtgd4IhDTPJILCLQUvi0YG5kFvLd20gGZhHYw
meu51YMO35XzGFiD9Sil6WYoKcV280QP0n5Zcv7PPmuJQhazgdXGmyVg0rU4bNhvvIG4yTQc7Ca6
g9q8x+ZaGBsqCTghpB1fChK/VZwljxWLrIeXmVH0s0YekLcANA3kuMiykybBQHp2fyIhp0EiW0KR
Do2SRi09D2DDK4YgvAajRaJN50iSLgms6jGpl1HFTz9FZWx6bqpNoBy7EMy501kX0MUWMOLMbceZ
HBTpUXc1lgc8Z7vb8pu0AxxvLCxbCOUjfLwxwl/vraWx+0MZTlO8QE+CbRfcmYxfvSJiw7QocTCL
fRYohhwzn/r326iMDpFm/GGCRay8wXm939k8cOkiUCtn/MJ7meuUtukNDmmsA4xKJzPvoC8fkyzW
AY92yLUurMKGbXuMaWSNiCrHOEEQuGzom55pYm/nPdoemgMrD62oUfCeCVd5LV9ishCONAk/MFYB
mJr10x+QlyyeXs+a2OsFkq5+g+C/dknLl1xz8MnL5uoYyMQjil/msPx/vgC1uTnRf7Xl6Zd5jY91
SyOI6VXQrVo3yMR0QmIE/+TDKQeXNnBSi5/1q8dRra9T/L66v70mym7bXLE4RM2ZRxCSV3TYLSjh
mhDiqtS7vKujWQXsGltipwGBp71Ig0x/B/9WmDQTlLQHhKsGmoYvdOmSViDr85KvS5x613BKRxlY
jhx73RymCWOEmvFkB/jiw07Vw85GObWip61Xw6fecqc4yujU4axRvpKvqDTRspsdO/cAhnPDgKVU
k0dvSrBt/Y5q+rytaqFyAbDPqZSQvrgkR8cNfxOOeMIQh5POB2o3L+W+yhSK27CUrQhwNuDFqGqa
hc/oaMpVH+Zss1140k2LUCLxsYWjvgqadVhArGQXsdKbPFL9l2uwSk83HCmWmAMUvTYFr/hPeoar
Y/2vk47MiBYTl3pqTdFaIvo2QWog9H/v75Ba8V56Rh9wrFkx3dFHVMOwPjGI3n1JnPpfsD6LUkwT
hbBeipFMud0ifNU2Te83nVygnydfKqn2ReqEqlSoa2g/MzbWkMcxqUnJvf9/nTuzVlomfJNDjPX1
W9I8SgUfYHkyOQyxhZLyaPGBIgPgTlG9BzLk2SAHwL4XD0Zd42U9jfrjmQE800JqSWaHfvNcGCpy
IED9ZEUsY95jpY8Iq6ohWHpEkWubaOgm/Qgq3lZ7kM2SV9R5Xq+3ubq+8ylbtF3Jkrm6Sl02+vFM
Cxux7IzlSXhs1oddPBMQ6q/9TWF7kYsDsl7Sn32LR5Y1stNv7jTMsdACRbir7PzS4dMuEuh8CT7D
lPp7OnSIK5fio3LUdGjtBxXJT5fmnQgVIFEn1x2w67TpbhDzeTWhfPM2XiPPVSVmSH5YGUNlCx3p
LAmzGjlNms28BHMHTnFyQrAoDugvgYjK+L1CsuFryh5cVF8pDd7xdSDfMaPnZCQ6yK+2N9liZame
CVjkWHfBAwtrTTqxSfushQuj0f/uvDyxnu3zcgQB9LK6tv/ThnH4ap7O5ZUidwUcME3lzm5AZBgv
L9m8EtyJ9a/Xzq++wSi++HoBU9xZmjfG6d/SsjAdU/kLkktedVBJ1XqYX5+TAH5FVd3q42wF+fxV
aP74GRzfB30sWvuG4Z7rKN4EI4giCsTmpGe/ZRkdgIyuHzMrocNIpAN+rGe1gax0Pl/cFUAsTTa8
D71pu9N92HTqm94x6suShM9Cbfm5IG8EmwsmHu+aEoMYDPdWHROD/CdWmsyG7HuGxRlfh4r2P+Dm
FIU+TIAeBZne4FmnDa1GMoGcBv28y/ebiWdyonP0ie3xBdg/ZMdojFtf8SRndAV43sOAsmj3fWji
MxzYXFNqgxksUVGoLQlhhdIVoFqAkZZAyI/kS6uRWZmCs3teYEkguCuFk6cnd1PMHwGmkqtZl6AE
Pt3e7N/wJ6RkcVdRjdumjM/9L+QlB5XFHOzI8narMe2EL9ljZ7/yUi+EABKRjOti54+k2QXgD24S
MS/H1gxgTQXt1DltY+Y4wFsMwbCNF4nxGQB/hUw9bm17DjO9TLdPBmJyn/jh79qukY77S+Aht2zW
8Yi+BxDZFlUMA+KfqNpyLFb6Odx8Xe6T1tyOuaZn+yVDmFhDJv+3UH/Yur5W574ae/55RGEH4reW
KtsKeM0XlUhcRZnbOxvR5cUqvxS0odubaW+lDKzUrEdOHFqI35UlKl+Oog5Dx9a+oitbdz6dXIJK
YxD/PmMtVse6sdk6+CoPx0ztRIeM3dwSVAmouhmkMVLT9fO/UU5U1EUynuXrlAjVe0e0QCkn+Y0y
vnOyf2rZ+JiMa5ObG4GfYXD6o9ZFadI1fRGMXwriHQ4cHA0xPD4HZq8BBKhJS65gc9n+l7ggj+I7
MM6Tak21r1dX6W2W2gluIxQXOmgZy1a/hsBgi8sMR2yrD1cs62gP21yxg4ayCoe2W8rMegDhUEQr
wujjNaxusAK+RL5I4zx7nY02DauWFEEQ2dx38R8EjvD8bHtwgOoCyUqL3NFCHOlvHoFMinRxyoDU
/5pbGAAFdmnGLNEyWLX7XO9PgdlTDvNDIViqaKT0xTtqszUtG7scAA1WAapyNFfunR5dqfVufe5m
EJrtM320nWeOs3D0JZShABPd2Bqbc7oJl6wMmYS7sziLfHkFD6ALK21LId/5PCbl/VKjI5dEmNq9
uLQRYcCkQP1afTkfhCa11cwQ6vRaAX1LKdBGEQyar+gHov5L0D+PmUJjraJotTgG8VyDDQzGKCNU
wc0N2e+xV+j6fx3cC7u7HGcDIYHfLsvVqbsMdWoTkhQCPwGTN6ZbIpU9cVaWwwJaJWfvzkzKW9J2
6sVmkVlRdzlqTFfPjZr3zpoUgR66YZRu6px6beEWdHQOVt8S+z0iWSGna2w7QH27tpeSDZ8auaNU
phL4y19KlTQT1MKeBs/2RYhKQ16BSUAFz+HyF4hFB9wDhMR5eoxcUkcVnwpSqh/DCGffK4bGyvpZ
214BqkCCqMINJpgWeqyr8nf+BfDDqC7Mp042N7Ex5J/48PxBT4kPDlMHjErum9Mh17scD9E0JusT
ys9rx2IGGZJ7qvwgGcGom8xJsCVjWByNFE/IhGVTkMur/a4z8kOVvoxJUII0HgR7ThF1OVXoQFc2
Qacz2a5dlzXpJXI31AgdfEazgLGBJXAPxEumhCdC0wtBwfAUrlIZqoLnNDARYT6VasDy40AfHPe0
TsUXpyRT67bVJZltHaKSSkX4P9zSsR8t0cDjpF3zWOosocvy7XqF1QYVpgfHQSsCtZM3ku850qiW
ppQ3QUW7mY69uTSemnWoO0P34ULqe9C5HNlMPdqA+IEpReI3UZpgF7N0G1F+wCQ426d0iuQx1HlF
Tb6IpXGKf5A+lk1ftDd8EwtklRxnPClWIsIZt3cxmbdDl3fYvvv4hzwTroPZKxE05MD3nS62+HKe
hz6TlKPxpoiyW0po7fUxv3GFSXiXgC/PyLlSRdisWIirBD962VR5bUhP/6Mo+bO4+G6esrxU8WNw
VDFHZA1nU6NHYXGJu9heSdUSdenqJH063CHQSjLHTQJJpAolNZPX3VGchCH1dA3rKi38t4gavbC4
AO1WLjP4klisQPHrbDBqcv+IKgY6x64ea9VV5sA9yAjPblUWbWFtxqAC729kNOGWaj6x99l2C9PG
CjRMwh2JNIIIZ0exfCLtR5M99tdkaBDdED/Vj5MEM3HKFm1fZaWz+06t/4CP8HuaSTsCdFVqlmgB
9N7apvOOcCEmSQyOjHtfcAncNbVVBShB7mbpCQJ2g1nl7BlywJNRuvz+y+0I11DAwzWtdoLi02MQ
VQtJ1q37sExluLlC+cTuVnJQ5l9HdVQURbXgbZQSrDDqFbB6bcVFagnenmxmpwlZ7yeZ7KK8zkOZ
dCQKVpVFrRQw3ll+g1lD1RZFhcCtryxc9V0vwYCte275QDeCoqrBmHNorVPw3J3yD/yFtvrn7kfL
kxPgLYRqAqM9iW1qbnigP5os2zhMFQirAQUuSAvxvskyGRfrT/EZFZL25tlH9V1fZxkbrozXV+bK
nbRvHxOYu7UZS/ccHzUDG41Ex/A22prdEOUp4DKKBwHelhGbuBi0JO0JBWNBN3oCM6TlgUtP6OOF
yXCpQQJ65J0cKg4FHK4ltxByXPaVkhyhLx9yVF3ZZb1Oe1nlGUsoq5zRIHyTyQa31MDXHTkhWjAx
LEtNPfozFObzlJSfMVVTUfXe5Oti7ZlPg89eKThfX736Jya92SOaebmc1WlfK0G2c8nt+zi/wF6T
mwOe3AdQLhd41BEROu0my1+ikZ5D7UNO8QzhalvlCe9Trg9kQ65GH21YnRUM+xNd3sjt+0hAoeKb
eHZ465TyJ0I/uataPZ59JvmfWZ374sIybSSh7zSj7BN0kKa6ayqM/7BzClpsps4SU2PsqiDeKNso
IxgX3yKOgsGfQ9qAlqlvnJgVP4byzNVkUSKmf73fjde/Yh0/6z84YWaclvGwBPJlo9Kz95zAqlZ7
tWqcReHCjiZl7uDS5zcuuwMmrP9lBv5QVEaX1FHCm8rChAWwkpMy3uZygq96Z2eVq90/Ey3QoKvn
wdkDs6thN4NjhOy2pcBEk7SPLXwli8Mvv7nhxZ5BbzdTMWkrZFuQwuDQxqISaLZjpavm/y1yZ3PT
NiTWAT6Vj9R9SmZkSs55ZnM/KfrtvofZ2C2K90HoIFkkxBac11oGAlvlJjxN4gAY+7Q6dkKu1H7A
0o3xfGtdXH0zi4YARHxmWPGvKYOBh+RB88NBf3jHxkpsPTnN2/gOHfdEfDlqOXikz3UC916bfuAy
uanB5g7K/RmCBWiRFtOLcIBAPfdW7TqsMrynzIEdQDlicyJde4TlxBlWohbZvuMD+1iIlYiRKGyz
d5GtU0JwmBxKuz2gXPGDgQHPOLMZBHXdJb2BfoWxawiY72R0V4uG3PYvYGD3YHB7LXicudenlJnP
LFz4V10hmfk+ZRngDRz6PzTojOt5f1Svc1HqrmO+99JfcXe+a/xwac95DhHaCyQw1DyHxwsIezFE
rPkFz/2dgxGOEBw8E8A9k6T9KqCCq90HCCmXKckLfAGxMuB03pKbDShmRrStIjMqv3QTp5ZgqgIy
0JGXnxdAk8BYi0/IWEalFHaTmJUS9FPCW3b7SNvpgm+u/9pYSgA+61Jh7JZnS6W/WdY38A9Vbb5q
hKGgvmUp4fISWxAicAuKw2br7ZGlJGo8aXxMiZ5Qf33xPDo/z7oLageDXPlJQL3we8etpvCBR4UR
GEcfRdUMjJBNMHEXrD9Po8fGFXZHFTjTbM49ifkcFJnO4886cvx3JRLrlApKLUivCpiZK54lNhi6
3FhOqVES693nd4ltIflvfl8hDKOkoexJVi9dq9K26oxKmaa3F9hRfBchvFUeiQ/1YrBvz2P+Ozl4
Mh5Wh9kCQ6XxLhDugaMYYmcwHmrmrDngPozYW+GbWja2tHBu45Kyl5akIV62/YCHrmpFZgJskKy/
35zAO78/Wvy+BDejYp55z1MkS+67WS4B1eX545FHtxANyd15FApg4t779kAn8PRH71OqkOf7NPHe
X8xpLfREHN9NHNpJ/h3K3JOwgmDeM8xXCJ6vR6LCetIkHbfmWwYcBP5TMQJmqZ3EyDB3TP7iwfni
kYo7XzoyN7zgUFV3Ifxz3jqMYV8BhBnyzZRwHxvwdsiWJnR8N0PufXb1luU77dPIa3EpywP6uNiI
13gDQhVXsK0+Uh0PYLMzv+oMnCexOfKKsGCdUyAfIR3uqyf6wJ3Ktc+eFos1FHJWbrJWN5S5ztzK
Wbie/NgsQSBxtcgrhAl7TSO09KidrRoxgOTJ4mMXzhd9rXcP329dIyXFw9CVJwxFos/i8Dixt7pP
neJdaXDiUyRGhGS1APAu4oVXzEqRl6P4Q8CYx62fk+hsZz/H1sG1q7pBWOkC7QzlfUmli22MhUx9
rPZNqehpU88a+WTiy3HRHZ+zERA6uRMcQ/73/lMP8asHSbx5sJYtaOZEcTW6NJj2k/Q6KpufoRHh
tPEPi46pxq2mHs0iKxhNlhUXXv4L3701jHUXDGAjqJmbhty5YTZBUX1hCT1vK1Y9ukcfYoWEUgUv
exbWkb6u5mh0gNu4hsBDrn6BxDsoACZWLJl4cPGJck6cnE1SfeVlS8v1doC5xPmsUeinHwlouuYu
OR3Z0HwAZbk62Z18ldQydETJGNmHRVkEpRXxWWw8kZ+l6uBhXgLviNek8pyOjv15qlclXOYSgf1U
iDlWLXL2q19Hxnm9pfWKyFo4kQLZOsCQZJS1QA8vPQ5w50K7AN9xBoo/WsQVaz4vJ3+Px3n1xEVA
TWA0qo0ML4zAgIrWG8IawGhDN3Y9EAbBBiKHaSj/ug8GznDWRsXQAAU/m1ZA/PxjowIwNK/8soap
Dr1ZjHmJRFLPM6aXOv+efcZFq6gFQx/r3WQyCaV2d1v3BfM2O7Pz2rV0nuMTIyAUXY+NwDDNKgtU
n3ldUEU2YpcVIXMrQkIVr/J7MWdREpqBvxqPyDfwcxJ0Rpc7y3q+mEc+dkm7+/+QeQ+ramKbvOMY
xDJVTmwFGsLA4t2sSSLg4vO8M2kzn2mMREyrjFNg0SqCuwJvbNeDS+LPBA+vJPqdLP2GfJmZASmw
wM6dtLTtU1J3V5A5j4wDTu+YRWjwmsP8kko+6wf6qViKA/lo5RqUyCxOzqSEFvbAvCmxbI8BwnxW
t8OqR+jDk5PBOEAa3ArX9Ng8dV4Z2vT9svloQjLqY/lPFd/QIW24m5NciTtq2dwH/BlUFCdVigdS
bj1zpJ6CtbLOFb4rHx+jSsStDjQ489IoDdd+mX4I2s++Y5vvQ76zUo0CT3h+fh9cPfZnLhjq0EY4
XQlievKEv29c0WFi1LFpA4q3uMt7VKGIfaHbQfoDYyc9RUDLcOTbcPdVAOEfBDB49wivlzaEVxJC
rompDLBRZT5beA+mQqYgv/OZ7dS/BLp8KL0sFvI5LE0G76AoUZIupbNliQfSjd9QAw2hE6/vvxTZ
oJsAv9VxJOEKdrUW4vLJ9E05bk+uUOVc+3TleQclrhtwfvY6In7BEv07209/ntvsqIzi2mdFk4xA
/hNWYtSkWWgOnti6JN+Qgp3jYtjubpFa95djM7k6fzdFsQC2+P4kX7ffnuHjEk83ju9QEwZY6HvV
cZUVlvirossFKGDN4ZA1EoTqmURfYB8fiquuhYHxlZu69JXuWaRCMoqumU49Vltz61mGS4XzBNqe
A/JbxjFPuRyCk1oOe1T8juKO+eKOHha3iQw5FNT1ZHbcLeRH2gW21y7eOjAPZJI/gfmdS+9ikqUa
2Jl8n8ix4f+kdpRw6368UfUBeS9PNBzKVockeir6ZWlTW45MoAtC/4sjGIRG+nBxsy4LxJZgAh25
Y6IsMVpGc711pD3sZcEsQjuNydUHguNiuIYgbu8f4gfuG07/ODu624NN+U3AoRcGX5o8o/5D+opk
9uHfgMXn3dbIBNgWuJ53S+pYSLMDu9Ug9A4c3UTiSgz0Ec57yfUJopwHfsOlI8cfRp+TrzR0ZtNt
sivFmo/DmWSzZdyqc6DRf6KaJm7HDQyk9e+0j52RDxXSVoh6E/G1gY8jbp38g5kd00ubyG6M5bUG
OyYe8ftZrNbItMaLybR2AvewYVSgJBkp8PEdh41xwTbwPWNYU1tPUDxtQRpaa2glhzsrd/srdlqp
caHtGIub1y3zl9NQtfNc0jWQ5zfR2bLNwwRUTgaCQTiBBrZYlkxgKT17NKDnf+E/+b+fWWqOZ0VC
j7OoHWc5mOWSdu5q1oGYn48ZZI7dtcpEnIxxHk+fOKsJPeWjXJJNvDoZ3fKnmPDCeELFtFoOg8Nw
mNIaRz+yvJKsOMxWxNdwKzamnlRlYqYqqmjzZrj/eRJ7p+EI5PMaKGv4BIrRTXvZ3KTSkiFkhSIE
THNjyNhAyBOBvBXShZDpgB/nrZGzcv2DmykjvL+Hl4To641XZ7fy0xHzgQlDjgvI0veL/1sdwBAZ
DabiDCJzJxvIiP4Yna+jdwiGLkcIe9nLqQrWHYeG6fyTQmoQ19jMEpoqtv3uvPk5VuqfdYtHh3xI
xw0Gqhxyhyn67ts0qcODpNc+AS0tTiHe6KH5Ac84CdR5PZOVuJ9qMIKsTjBIV3J8QytPbE5ujUG4
sIF+PnHs2MDg0xp7CExd6j3aklTh5XGRje4jE9FVMscTWAkBCHCZ9VGbxe29noLQN6v1xx/+U1SK
Cx73jkeWGHK8CAZ0MnaJ4ISfswmlAy8OewzIjEeKDT1S3xpmnbOrYim07ionCu54Snf54nwlh1j1
BH0/SrdarbwkCV3ttDnU3wOuAlqQDojvOx63kYszmHRfpnMJAuGZR8449uZSHe6qL0bdhf4W3Vrd
Qkr7+zovNlb2X9ZT8DqrxTX776IrO9aQ+0JfgCPuOToa1doqt7gckQulIWtKnLA8bzIXQh+TTUv+
nllzvQ94ggtaC6ujI3apSFpiWg2oht+4A0sb/Yc7nmdFIVqHVqtprhKVxUjcnpP/wW0O29ewO/dt
6CX1bLIIuo7nWtFzxRqYusMLolocwg3VQaDJw16l0RVYjamoiV5jaWV/R/ZmFm8duEm1sb1H0/TJ
W6+rD0/+QDFW8CmhNT9bMrYxspRXq78E07+1m9Q8HA90DcxKG+KeRfhcAm0PiidIAPsztI5CpF6p
1TsPHHdNxKFstFvs6GzZJGhHcPby1legyuTeOO9Ms8ACOya+Bb+vbKYdlqimXo5XGwqNQlgd+No/
QpuIFg5zlBKGoLrgM8zyd0VBTM9/Yjaosh9T0kTUXQJ8qJl5hAXbWQOmMyQsXnDEpilLYX0qxtiw
1FBE3JlGPBuaxjAcdS/tSPMXWZMNZ2Tx9FvmZOmSlCX+sXoFMhPTWGReSFmlfLJsPWvil52bqz9q
YelSDeSGZXfJ5bsZHxSg8/NeHSdx13+/y4MaJMDNUkllsk90/49fTbc0NQK+GoHmC1LAX6pATFYG
9F/7Su/L76JFJxkh6u8qwK1yCZ5JbQASOq7qiHN/PLy6rbD0Izmxg+9/NMJH6paoRqw1aQ2cJLGM
wvWqjhyxca1AsZw0IIm3leRuztksy/omgfHsvFCug9cxq26lcYvzmb6ntgkwRfz57rVNlapFXKuw
gBjhbmh8uL7Yrl/wx6r1IVs4qGMXL6426OSwmJj9+4AOpojMQG7iQbcLrlkkXSFZnsRtFMEn6JT0
vz71pvF0X8tzbGX5TXobrWlvEKl62U2N3PXrq6hWINFHmGGZFVg7+DWCj/+tfXT7ZI/5e9j+HSXV
WIG9iLtjgs7Z6IcLV+KPQdj/0tuLCJ1yvZJt3LT1esbAvSzrGkUH3F0fB6coJYlZ/dFmLGBvN/K/
3VEe9+Lf5jzt75IDRfYo4To5E1EeJiZu8A36L1RdcxQj6OOEpCa+1aEaTlks4FcvUtGswOWQY9uK
Uu41Pd85xnaoLno+UI+pscyNiQHTGX2fRfaZiJt9mHzYwvYsCuc0SSjqE+avjqV04LdZBjZYV65a
B1CMKAou/OldK/r5LJSXs97gvn0+eHPUbUi/N9TOIQfPr1qqEI9+oftA7J57ZBlbZQ1cPQGsc3dF
aDPxt/E1z2Is++2UBQcRbrPJQaLty0kFQURiqCiPQOIRLPQFxDc2UYMDJh+MyyRNgSG7Yc7Df0G1
eKQVRBGpeWhIvRvcPny7TXrllLxeum+rOtO+QEaaVocgaFFIsl4Tfxt3V/9puT4YKY26vGTneETz
pIOkXHAoqXXmTHgdtLOqyPHo00Rb3bb9a8s51mcUpzlh7A8iBD03jfkAtvUWmn70iG7Hdw4SvRp7
KD/lDv3EhRqMdMD7ULr2ZMo5OzpmgDrBpkLHGeDSiHgj8d5EnLXaUUUqye/YeXltz7607gC47K51
jBQNcpiUZmf8D7CG4q+te+X8mcItuPhKKA2gmcE/SYS6biRJdYU4Cd4/wYkP5UEK2H0A0FFLaRvh
KWYP0Yu91QLkqBmMKqPJ/3wxGnIQjUt6s7KYEHEk3+ANSHq3C+d9ytNEEDjeowCK2gRt+F3q31z/
dm2y8hfTRFXMn2P+CaGpwH/X1PnW6xB+N9qELj+hqv5bHAlErOuq5XJ1Dkn9Yx57X6lAO8A9kbcw
lc+4bjvVNFWYrnfD3yOwa3AGLG2vftZYmddU76xoR/OXRbIGcL98unbjqoPbZStPVxye9aTN4dIc
0CZttJsLdOkcLmLf/NRTOVXWkMwKLHZgcyrKeIgc2Jwaf6JhKXMHD+fwhtN1AL8E4tpNqI0SJxnv
fpqRj3X5RM0DOpfqMInpshcoGnrsS3iMG9rrsMS/Jbf2Z7nXa3x8/+zrSvpk80PyAXMmJiFiRuPN
1k0iBjX+bJtI/rfidlaArMzhwErcXFGq5Ugs7/p/hHg4iefl1O85DVr6jcANOLEaq9Z49Ad9oF0R
sHiFDa9ERJcmRqYmuEfJU4hKRpWWOBTlDGzrnLmrKXwGSHhxfNPP3MvpSH78xT+9Pw/yOn1m8qqp
OH1DlqqElwOpTNapb0sZ5OztT9FQ7apuNJYr1ljUX2XoiqgkOFd9y2pMsceGPjgZ2lEtsFl5ay8Y
2qWj7EBph9jJbOcZud7ra49ploPBrfvwzbx3/Ikwbht2q1RpkmYURXc+L6GLTjEUpGIL0C60rYkJ
9pgVxDHY0VaA5VPlNLQRaSQNTFj8BOQjKX0B3T/d0nCM0d1W3Y40woPb33zXjI+mDhRmFHRqhXR8
gPSh8yhhzqeYPIFnXk0fugQXF4XoSZpN8qVCL+ElNNPReIE6fTmTSHpr4mx3AsXmpIMMLyAwn6JE
oo19mcRkJLnehPN/TKzMEC6aNgUl4/3D271Xan/p8bqvpaGFFNqzHlurqQNLxoRKXK31R/KdMULE
WbsgjNzYnXkbhaVVBUIiZSLqznGTjJtchwFOqmsWlq0AadFY8bVKroGBYehvWidmY35lEoQDHssD
piJa9ls/G0dBN2QMCkTSfdd/dh9OeCbhLNaui2IZMtf8x25AiCWDGBvfeSDc4zSp4VEomX4Z5DF/
jzSNTSZ6dU94CgDbkPB3odgqdNk6/OqNqriJndQBMpskQBSoWJPFlw0d+XgbUVxztzjqhGMMV/M7
6wDb5t9FuNv1paF7RQMXRzd+3RcdOEooB5ISXeSQDIzFwR9yWmLmLUlTh94Dk9eGEqLRw0kpRPKy
ImIIBAMLAlMoo5flsShRf4oYFjm+pgkVQty1S8D1G8nLse534kjxQDM1+v7ERJ3lYOIibO0CQT7I
VtsNzrxfay3PshfHSauSAn8uboVNvRe1kpNdIFtV373RfuoOW9EYVQmcETq2z8JqDV6whowKm8CT
OLPGD7Ip1RRoWd24DPQHKiC883PFg80Ps6Qq5u4maUa13P1ZDs6cIQtEJj0/Nr9fCU2gr2Ps52dx
Ahcts+9DIHCpv/wPHz2OGtveljb0u3uVU8Wk93KjVnd0taxp3rwu1dXU7FEM0xiIgVsJnoc7q4PB
q0DDTDKQiflDPHLe8P1noHZiuW3nieg6S4uIB0LxeQsbi058NbOlPb+PEi23cqX+2HUyfq8QoHSh
KEirfvsHa5WCV/l+gghoAkqktjwR7UgelMe+CSKlWE/DDJmkGKCfVyYtP7FME+CGXItYoKmY7rs6
g0h68dn4FOFsO96qch1bKo6nnlEtuWpbKvOS4Sau4rzxmwVJDg4UB479pDYVVcQ0Re09brO0Fu6g
Na5oCtDef8rwmqo7cG2HLGVFBgc2tWmqLemcAHZrMY46rhIVXEqPmvw+dTtC0DGfZCUcPxXFReOf
CW3Qvbr1vebZMlJckvRHQCYU4nag61T5R46TD4WZ/AR05+eW80UMiGrbsVb3smQ7UJw6xY8yZwAa
6W28sCiRpfk0a8ULq4nV2esjg8BVb3kQiXFYXHHO42pZ4NvJzwuyq5Fuc5408lht4yPYyqqP8L19
OU8TGtINIy+T09vKg+hWdtd7gngt8X3rvM+iAUsT1E4/czpxNenYMPcLOEbpRMBuoS+4LB2C3rWy
TgpPHYDvkaPCJ6YtxNHY4zwiqox6j/NjXzPOc/PxWE1rDi3uFIKGmcfgDnx7pe539OfP3RxYUEa3
8z0gHXOQsnEy5TdsMuq5rSIqAed4c//ufXYEQgBEAwtilCZ08DMfX6GN6Uir2RI7pjDBqOWgz4lo
ADm8lPTq/g+QmN7StGDyoc/KTmKGSJl7uKCs1lKyxyUOs/OP2kl8JjDbV04yaFVkCgVeLtwpvUTG
wEkLaYZJs3j6BuHu7PfX2E84OWMkiEVEA3PX7v9BZfm1ixqhibc0x1qIuAby/c/uAhMbvu2ewsfk
whcaUZAUxokDgvq5DPPJL0ED9dzD+lbLvEaaD3ZcNAETS88bji0IUHnTX2q8dnyebKBGTgpRtO/X
4gzbNPh8DHhPzWzjDaOXMBwWK87st5m57I1e4rPuyrrYD68cHguuWNhRWiyQEu1IS05cZYxmMWs1
ttsX9/BZ/NcXAjZZqfTPMCc5Sla4cI2KihP6XoK6MQnT/5T0eY+3e2xW7+khNUAlV8i5WOlIbDH8
OGpu0NKETn72o36oGC8HAJ2vwljko8nG4Ww1wb+VisRDDpWHkInMhvfLNhbZgPq5Zozp8xQkmovZ
MAEcMV13Dql5st5DqGQzsrMoJLi4dik0Ps7aC1KS2vzZpgKZm5sOBtLLGbcC83FUQ9QUiYHW7TI2
C12aibWzTo8I0sbg4PYQo4KLodfG5V8N6D8l9wWB2HTt1i8V1keh8qwB1imC9OwaYFWbnpqf9Kmz
bbsePmKDsjfHGo2PxSDybRwYVuN0BBUikohRy3U2VaKJv4c3pefaK49p9kzilNEeQKTsAHcePiqW
hWVvDfCn2KI9ZexjzsWVGhKziNY/88XtHrGPcgNO0fVN0txV7n6u7gqwieHUjp2ppuYHF0tPtfc4
erXsuPKgf/EldXVZtAY0gr0rE2iBUH2eo8sXGl3qW1vt2wVSm5TrwAFftSPguu96/jf3jokunt5H
BFRd+yjOxcCKlLZ+a8uxg321GFHWiNenTzNYTwA6JoWZWavfI+s61I/yoHYoOSa+YiWjGIJc5wLZ
29c+ogAb8Mm2h29GaN90imNGMkevVgJNpkLIh9OOqcC8CfK8QbyXkaeg1UHSrpuO6Oq8iJLDZbop
XE21e4NnqV8/2mL0JBuQ/D6qvm5T4VSbG/VFawJbHndMTDoo4OlXDL9YT7AFOo8gkF+kXOHv06yb
9mXGOxGxG3V+R5/oFdxPg/15A4qF+OPIB7SQrZvB/KdQ3HO/9HbsQzPABghYNCU2HI+ahqBbFjXz
xCQgx5hF8vuEMrPx7Om2jx4gVYH5z1KPPe8lgrdIuLZHvY0zUABAMs4zMksoOTbhOzj8fiwWtVhX
AuWRBxqDnVSxipKQjEDqHpEMXHztNaYRpBX5C8g5uDHqhT0xmK90RbDzLPUMpWcjRTSpEy7tlgxm
th7fctfI6G+XC1m5f4Y5rCdF7/dsIzSMqHMQbTKjcVtCtrez1jhMJ3OnkeAVWK1eJCW08R4GibAR
WJlc3lVcQc4ak/AZTiqhXpDOlbdNHmNofLXWWWIIVQjikseXg1OvlcwkJVS9mcjFVHyjrBO5sMla
LLqpqnvxrlGQfRNhpMOV9wnPFUH2/Z1QSBht0Yq7dPadT0N5lXBsCAMxIGXDU9wPKYBIvAOT0bOw
+7JAfaKphJsYcxTvF5qkX4s1ufaH6KuHRtB4LBd2hOdh24IoV/e936NpnI4Y6PTt5oZeRZGLoLWo
Tu+FRk32ljlSChclWgJ6ubH8rnYggQALiUYfYAA3DSB+oTuNZTdKLw9BLY4So50bOaBurI+OTgrm
XMwLmk7DHAaxhKNAJ+MMR9ObR5JCI6uNplyyzn4rDqwWNFycz34ex45N5LxK/ETIjSoAZdjgFRLi
3K/Lxni9ob7d8+0DndgCdtf/+mT+ol8OO1ap/fu2a/QnMj1tXZS3VEJqMwc9HepwBg5Sw/ekGzFK
2JE2Wky/X71wznol+d0MpRfHQ1kfwplxUc0TP2SPRv/KgkPVcvgPkmSPOslYU4YLQR4rxe2580L6
IndhWyG/M2SzQ4CoXSo08QSOxMhiMoZ95yv4YeWfs0GlgjdNfsjJ9PFPiS7Hay03k01W9mu2u8s4
qQZm1l88wjaYV8xK4ES+7TM4VIyNEhorvjaNDSeVl2DwOIoBai2Q5xIOYC6OzsvHPrg94ZvzB5SK
83uQxsS0sDZ6BINx0//w9AT6eYyJGTQT5Zll8ELndr9MEDjB1RR68ucKtKzNcdcLV9nDdqFdIfS8
XtnDhANNlkX+fv87cyLY+ug5ji1Wni1dzmGsApzq0P+CKWKYGFyQxdCeiWIouu5rj3Yy4sOM18VY
5oKi/1J7wjxXWoDG6dE2HHWlP5Sj9IdjrxN2DHeOzh8tkZMcViJqqziJh0rHGnrRwSNiq/ZePnaz
in80sqhdvnoRTcwBiMVXQFU008Hk1tJShfYRLA1ZgvTrEor67PzkarFCeEqyJPacjW3ujvzB8uuu
18K32nu2WVO5gyNRFLzoe4xljSgvACElKfw+UuoVbZbd4OPG0C2ey2S8Q7f0Eld7DIYN6Qy00fbs
76f5uuuQSqWiLslgdGSp71KUmxR5vIDGOc/HjP39M+EdbXpqQznxzN8xoZzsvtukaKWyDF2MNCnI
K5TuMNRD9AINudr2RZmz33uFD8dDwMrfT1z6LYvfNiFMAnx5LwD+EZgppgULwCREPMNve2Coset+
FXalnDqAzHcM7CBnvc80qOpBNI0l6LqriFihDGvqaTC9Lht8iKG7/Y9mL5qPyRnDTmTToGW3GbV9
bQjgGHNOMzRj/3htFSHQFvFJFzRthTeGAX2R8ODNBholgxMxjFutRw2JQChx4Aui1z30K9rYyQi/
Si/eQUVIcbW1W5uXrRIK7s8fPFFWn/KZAQTL6COLwc7idnyrRifu+VIjydKQtigBC7A93L839XYG
S3mmVnKgjABEhFpteq98N4uIN64biaU3mneI6rmL7m/zmceQlJI0t10IWHelnGBNgmc3w7/4GwSr
idaoUrt5lHSSWejHHAr1aql1QphHPZ/SriVLs69vxzTlhvSaok+bd897AY49R4lcOQcF96XaVEOk
xH76bvqrmpGT5v5TUFmBVQl60runm2wk4yZV0jT27gu0rwaOUrP4IglavqL0U3Ys/gcs7cvqO93z
vKjXwVoPctO8SQuQW08WeFBkjJn5vqquZGYT81qrJuFBdNubLcHvTnpc6iRpqX3Wsc8JM0lU4VCh
PF9Y6sLMlFZUsibflNICfRgWzpOxyaPjTNQTplN694gyXkO4Pri49LwGpEUMFzow4yAh8Jpxs8ah
3l/GKLjLH0Wxkm+Dg/F6TYOsN8yC3BYedZB4jzZj0ET/jjkgppQ8VAUTFIVjBQ7hlFPcw2Lxw8R6
wkpPBtNek6qjK2WDFRD6y8Y2GYcnhsha3kEkE6ZkG6TSLl36TWexqGwW6BxAhWPzGj19jdwgtTOM
LoYnnkOGJN8ishc9gRzPKczVRtIzJ1j0/rG/I+tnOtuoN5oR6IHUVpbE6HFpqF4zFzQk0ljzMV3l
7Kax8oy74e+PzTrhw1SWSt3dHxvxFrEbRYKLSLJoifFpF6c83xRD8I5q+k2eM7mQD0+/j1kYE++o
+rbjxIEI9HcDeWNfmfnhn3Cnuu40ZNx2IE0i3hZqeBWs6t7WcoFiDR7wZQ+F9ojNzANhw/0Mh1J+
EOZcZqAJslvDIfxd9I7+Vs071jeSptrg4a/cTeXlppAPfygpjz0kxqLBaAZS45RdJ1m3+UstiSQf
WdIiHAxB9Omca3A+4AVC6l7qnt6XMb5wFcpPbFuYPg8Qb3L6XrOUkYR2sDYFYraI5Ue0A6XSBg6b
9ct4AcA0KMeG7BDx3E3j2q/6FeQNdYi87EKO8zfKXKMy/rR/EjHLEDSUaw2lXWkaTr0Nk22Tm5T9
uOCi8sKgDQLG5xklsD4ffH/yBZRQ+Cr5Kggw88jMSdCQJZudoDNpctVNw1yOM6d44l1U6d/3mu3Q
INvfAnu+pt1vOvyCPfbaJoTZCNf9KRPTFKrhDMS7RCOa2KUk47e/sGWnvAAQTX4YRWoxybP7Ak5y
kgLlsRzId0lIaD6y5SMxWvyFwhau/e3Rg1xkCoEjv9tXI2N2NrPcOck9Jq1/l0tIbdO0RJ4nWJnG
V/GB46QO3HwGAMQUYqU5ZQKNbZaTiuCsbB+KnOdgesPqVo6URmlu4cct9ccmfUdptJ9JVthPpv7Z
jr7FKIQ+HmqMnmBvrXXLReT6EHjhwPM8KoOrbMfgNaSjkAeU2MCvf9SW2gPYxc18HdSJX0hAX/n3
0YTU8WOyqitU7hsUF04FBwfCFtC1qBt2fD+NCKLBtqRK2ghJ5qg7Hvrmd4Fz3Ygh32jo76T5ZEa8
u8dTcWUHQ5HVFYTBJMQe1Bj3W7Bc33R4BtbFIMgiQBtHCCVYAyQ20EOccG8ZGuhlfKbG9pzh79C1
+/bQ+ZEhOR0BCC2OFnqP1sxeKeghNEgOeZmZM2Tz0kAqHcXCcqUYqK+U4CkTymenM5q2uq3xVnrY
hIVGkaUG2azYrK39QaqCqQkxYFrJFTuI9f39RRGe3ec0YudPKYdtZLEIwFSLOospCmIB7mHW7Pf2
Fz20qilvOYRHvlitPTd0qpJ3ASbSzs1b1CG78Z/SWl6tIKDcBQ/FpaueKrZfcoxqJj0yZ4t+ktpl
cizycWEKDU+D+/1ZHK+atDB5Tsatff47Of6u2sFRyngE5ZcQ9eYFr2bh0lurQBzDmBV6WgV/1DDC
7WUxRnrN/nNeck1ZJ4Np0J4Z7wx3avdslx2I7fAOkdbi7wXTo+A4glX8NaQB47YZ98xxVSGxossZ
Si5wlmCs59HIscVKuyG7YRHGPw/kbpFMI1fl5zWGTKAujraOuoqPynvNviikqLOJqVKLWEYAUd/U
7tmV0sIE2APWUgDXhLcbhqqnU2/ICimGy7WZnEGHeXMP0h6XmPc9MDYrGv2X/7Ntq1P9AXJJdbAa
Hj1Rc6fuHhCQ2REVoYStuLADmWyJH1RGlRvUPPb9Rfuvi8H4DMI8yN0FHUjy3IscsHf9rYx6amCS
p9kwSHWpDDTkEAN5m1+pekVGx3NsUE5w7f52pDsFwWdqdJjc9uFruJ9f6/96kR7vucYq8PTD21XW
1CdFfT+mLs6DNPIHN4zTaO77WF/+hJlcEZcNZhbVlqibrk2ZeRIiXRHuCAru1mlCAjldWy3eyKww
fhuCSgLKvftNb2T/fVpwRuHd8vwEHly2vrEqeUfFtNr81AJd7RQC1sfUuTh0deKjQn0ofif9xzHg
bg5i4BEBurpFR2FnLlavgT+weTT7iMRLqoF9gAAPN4Sm4QZIVXwJjo8KuDO1w/rhqZO2asBNtXNb
xKr0x0DyASXEFLahkVWpGKrH2HiWsD/B+9S1wHokUIbkL6AArQXJHpcpTe8+ygifehGT8r84J+no
eAblLbjxoT6fp/d93rv1D8JBVrEB1CGL36b9NFMrGHj0PINNFJlEy9+ymXkjol9IT8+EFjpg7jVo
w3x++XL7O149VcisgCi8IDQg79spSJwzAeh4JRS7APZ6erfipGjm+tH1NuYi82q61Q5rDg/gXKhn
wynZPkk0nzf5xAlZqQ4hGgU+BYL85Lpn91TDpKfrk8lNtDX3P5tBN3tFxaTcwYZlRyU31wtMK/ew
ewZRL5hUTfzqABQ7/qgN7YDIVBaEEtnGCzx8854d2oeQmWGm1GSJJSychFtYscH1J5t3uOvjOoJ7
1G3AqaMJduitqxpGpIk54whE7GGnZqxFjRMVyq0Jhet23c71CT5qMDJJx0jzeW3N1fLED7KkTQ07
WbkTRLrsg9k9foDx2/fkIlNpYKS+lSZ+wz7BG7FDhlMb/dGO8aUsr0Oy7SMht+enoMK8mIxktlxc
yUaUu8veDUMwsodh4ltY6aBkoSGEvVGYKB2EomFofWkRlWzpPYZuO3+UprqtIzZ6dqYvj7XviVzx
uyFNTXUbZICLA/1ZPQyY9FWf/lyYWQNnXz2EWtFP7lyHFGBurrwF0JHB+tcGBfA+Uy+KD6dlXW6Z
OqAVw0nSPSxNRFH512hHs++8itnYerh2kmFgmJWhyO0l8eVxZXuDsvEMVVIyCS/khTFv5MvP4kT6
aUKEJ1Uh9XuJGEYQmiFUsxyvAMwDFr63xRooN3Sxt5ujubIu5P9tdS9FvJnCVXWwGTkBA0oeDsab
q3Zek/6PhbGoqcUfhQksXe6so7DobCrFaVY3v09ximBKNl/iXH2YyLXIATCMMsPJ/Fn4JbZD/jiH
LLTyWheL12OzmGo12TA0q+YaUhNblqOEB3Gc/GfMbFt5tJI5vnhIuW5XOSCze+GO04+T079Fm/Mo
JwnItVjQ6qOvdmPHDiiSruDWh+xNf1+zpfv6WWO/IUizlAGgAaStx4GIHr1ibHj2+oG2ENyO2zUr
Nt96iWMZJtx1IYxynUZ/7XGE25g6A/f4N6AKn8zJbGPgyk6m1NTRV+WXB/NDMZoiNpF7bFklzanA
zhqGI4MTmNme9nPagYOIV9yUopssb2al9i6Be53cZg94WTa9/RNc3Hb6XBkygBRhcr4N5Z+N8+PW
s0c8ZcRomGnzCKQbM83xRAySyj8uRUAJxP7iydHxVtPcInzQgU7hvQcSQ0Hk4Wit4k6hZbhZql+7
2gVKW3t1kX1YQniaE3zy6R2+p/G+YRkbBZIhdpJ9py+eye+Vx/sUA0JUSRYuehu0bwZOFqJASrWh
SFwceiLJ/5NpW49gqAHiPwP5T+sEaFuGng2jXWm6t72OAzqmDbb2GPdoY4BXMrzTuYHTER1+N0cQ
qZTfwWZBcgXn9mlyDOpGZYQE3WZCxW3uXj8Cx0z0a+4ZBWLKhSko3QGTfU8hKMaRf3alioMzbaPz
aZ9t5zLGZXCXWGaM5tu3FEUXzgRqoSXAL4+BbrkPPVTMGLDpjnyFtnanaBMaZWD2lCuDKCWSlWai
Tg5rbc4Dn83AONJT4yJYTEiO5r+72lE//0fBkoSeqazE+0GH3w6aWQDzRYY1tNm5Gzzk8q/nWlxK
Fgh/8D/jbQfh8Py4wFZsFG+3qk1+3b9frwNkZJ6yozYMZhq+Lds5CANm218Apw+9l271dtvfKpmo
/XaomvnKOFvKoEqZHKxG4wrq1W7pisR/KC90kpQ0sFsa5VvkhDuwc00idEd0bBkHXJaHuut0FgFm
7NFX/rzlVbZiuR5Ep+r7Gd4tke66ZqaKOk6Abdw3znocRRPiFqIjphdrhrYtowRUyycdvuZjNjZB
8o+2fBtDW/QXIxvTy6RhZozGbdrpXzSzHvAqksfh+8X36af76kTwY12vyqLnU33s9wTaCYpZ04WZ
BhVDnieJFNwwW4GaSXoSUG5KPUfP/kBjrPnC9Ignp7GVSrbQJkf7vVXxb6O7dHVpL5fQtXn1B5+r
4ved5ZG2ZJ8K2tYayiKe70+/yc9ir5GavuXrWAo1agg2G98bgpBpu/jCYGLNObf8ewUKCmbPF+we
gg5+X7OOev2fCf6q2AJ4M0Gqfvv2OB5ifjWAp6VImai0693A294Bl67lYQt76VI5cNsfbXn1cvGp
DrfMXku9u0C1Sk+q2APCfF5qNVPuklCtTUCvMSDvQTDLCFcqip73qOMdzGUZt+RrLsxvcgGtrtei
LGut5DfK+cvP/jYm5QEbLN3NQ/BL8xJyVQyEq8bpoktcoQ9hTkaSuqZazLf2pFv8fxpsDt9DUi6C
WHeZkpTr/9q7jn6SSCxjaaLraF04WT+B9pdJ9nS5WNwiP+deMamXJacMbJWyQIqUys6ZQcS6E1M1
3wYSq6/noZYKJe5YslJVqTokrU2xWpDHw+arYmNAZF28YYZ0PuqbWl0CNTRhnyHcdLu/BR1Ldsln
rORX0XL9xrgfd5ZhG+MOTB4IoL7aQs/LLfehQIXsbdRGLoS6+sg4KO4bdD1UWEfOZfYaVz4PToXr
dbPgPsniZvcoUfhZ8iKHNI2yoFBUKhEI2kKU5IeNj0316WzBieWYSP5fD4zDcgA73LicK6d72oM4
dFRx0+ZsWoSNrFrQzvwe/lzNf4pRCm5WWr3/cnpr3B4WSKOqVgkS1iVLjTlFelYnK/3nvHQ0X7No
qcJXvSrd+p/oqoPlKzjVTJsHw/siLAuXD+2zsoyban8WzLIj9GK3ZOvzcs0yrh20YAzAEbEi9DOI
Aq3gZpUJ6cDuFDT0eHeWCXut1KwbshKsd/k18EtRJ9UyLpb1snsInvLV6PnfSnSxKSI9BIsmUJ5z
xnKGFyoI5KVZFouYJHOM7tnyDtXqERy5R8sO6G5pCkKqDISjg9cdpMcs6mYqRw7nUClKhnK45bG7
rXJlpMfpwqYd00pL0ZZWwITQUsMhwsBDwhuSqfZc4ZoFwyPm/fYVFYsigzYICzz7YxRV0/ziEoZg
Sz+EtJoYWvOx7B0EkdLAGpWYHWRb8/kNP+p36SLwcipRNzzAhDskW0ZR9tgPQWJmmikeWncUwugw
s+CMPNxY6/hVPOOJqLx11CMvAaNBhoNALSTMib5hl4ntP2R4iZm9PBXcSgUxpp/Sm0xCMuTnHWMW
mRbWsxeR1CUbySTDHavAfag1EjAcDq3SU7ERVum1Y/5WdfoHfNKNU68hdD+lwON3YVG4No29wsVc
B2wvXanHbO1+iG9TfZ6HKyfqquB11xRekdV2ir1OXTAbybL6OJjo76hzY3uyUFfd+OIsZTNEto5B
sfiHomF/bG4b+2REd85MTFHI5a+L22eQm0azMV4tVrAnNqSmc2Tld/2USdyWCNHU1TxilCbWQ/9f
6nlP7C9Ke6W0BlzCDXQXKG7H7w4fCRU7phhspJZgp11Z3m8kKwkrAyLFLQybf02UcKK4jv+XBEVg
qXLbj9JvJlah6vXIwW5TB/j93HaEaLQhQw0w0q/Kpk5fGOWmikfEvYVh7Y2NX8twNY8h4+VUx1Nr
6qZum4VVFeAzRJrnXg3GmqaBpSJmMsNbp+eaQsUHJpfAxbvmOaR4djjFr5EE1GxejEBoBuTj4pqb
STD/hdfi5fZWbBmQ6OQsGmBFK9xKrHSNdpVNalOIAOHr0IwYZ3ByN+UHMvJ/ArQoQTnyFpXNdOVd
TySpfKP9W94e2yw054Tv8jTtjuaeFYviRKprIjxyUls3eXVsg6Hj0GrhqT1nDztwV/BQmw+qfOFd
PBUbBzKDmDeoAJ8qdEwy/6C8T6VYRgt2ejyvJEHIFbvpPB7YuNwvE4g8TfgM93L8CUHn3Dz1QbyF
LtlavmB2tUFfOg+wVfey02VYXETZMC76ax8gAyhJh3Ltp1Ey/OxYJHCrnnFTSl6fPsaujfzFrnZc
8tM4fhy7QTtUG2iL7izhf75RB+NiTe/y7T2fagpRJtlUfFkXpoJx1BcUHvda3nIIp2QkhoKH6JpI
8QSpk/lhEKR9iYC1vapPvuV3lidTlSikjrSrtoc3VXfs+W/bVEetqupVz15gs19wjjSeg5Cjr2cz
0/+YVfe5g/saIIX8J+IUiCscaGAudwDOqL228dpZbzR5AoJUQSSo2Y3u+1FpHK//o7qiI4EwVK6U
GSUNEhIHAX+A+4IlbrvwkR8A0U7bX6pCaEUdYzEaAnBJRKpMiBGqiEZu1Nvuuuqo4PhsjPuD6lu0
byAeplhJoBao6syLRGtky3OudtjPp/FvNYz/4d5uRRx5m8llPZy9h5OlbLB+EHjudP+/3vkA+gxE
GoxBQGXtjGqFCoUToK6DpgxGNQcd+CGztOLaSMxiB6cdLR1A6XWeVJ3+TkCT/30Irlg7vkR70Fxe
8jtQsMkLYPhi193NZvHm9QN/7KZKblDyf59s+vV+L99CJzmVlgvGfvm3Ib21dsmbnpPLZRgJdwYp
K7Ce7EzPcucBVK+k7TAT5m3WnhqcCw40ss1NKNiYxKqs7v7p3tPRkjsMFIujWJ4tMB2ZnEyKRfE9
tojPWMZ+6u9NtZ0Xx3+1bE2Ud/Sy5S6hHKarTLjfzdH3fH3F0wn00EkxlLocz3O9VlwqYmZ8cZN0
lj8+1C4r9P8pKJXhx0GwNMUDDW4MmDyO1+wywd2zho/SRefcm6Yd618EGs1tNZ5OC4jyVy9svXl8
Acw5zK6BqSAXkYYWiGLlXvja3sx+UvHdxN8yAoIFw4e6sfbrw+F9k4iKlONKt6O1ha0quhV6/s8S
Lb6Uf0lboV+UpM3F2V5RzA7ApjzurFLN2XTvxcvCKsNcE1EjpNFrU63Y8y+jwSohOLrSOtEwy9bS
XieoSf2/D4R+28JBV736QDxgXs+OPiiny4x1k5nmleckYkR4/0wLIlbKXun3K5am5o8stCmWxAeq
mtzTWOBdA1oZvo4XZmtoC2RbGEzfxuFVQ6KCWfnNrjH4FATx8Gbz41r6YPy7a7GatGSmGbPA0uhl
M3G0O5DHtjTEXoidx4Mrgh5pTsOOQKdaIdn/DEnULZu4fHf0pcsl5T6K4owhHm3rQQ2CDxhr1+ut
GQ8b1WMic1ZY3PCUo2S6zWJVI/QNs3mBgB8QnWKrBF/THD+vD7iiwT1QfAuqCfVh3uEMQV5GTD3g
m3TZ3bFIxwEgWQ168IyUtXcISmzNB/Aw/uLU6wg73n8skv80QjS9ca4nA1inWxXqKldC3l4NylyH
i5+yK331l9NaZyNY/aq0qGZNiVi8B8hw/VdivmYA7aB/yjkRAtBGlFOXW5s/tlX8bntSHdKHrWhG
8U/sTJwpfKnHLAQxVWpT0BG5Pt5KolkKgKCbOKRbD/aA1oQsPSsu1Y6o7WtPJW5AFu22FNhqgF01
/ayjTpWelPaqH1IB2jcrkBZeU0TqRdntGDzZZ7kVqxa30B/00CVwXjvPJ2Od37ngvi1AFfNfVCGH
HrMgco9xEmJ9t4OeErdI7geKpKviSHHKRIGKaytg9bgINEjW0tzgrhd++vQdtqkGEerOWTbFSIx4
aVCbfJLG2U+NWUha6R/ID0VLSnz8Ka38m2u4wNWAz1oUynyOQfzJ3rGkLFCVRRHrgEwCxyffYWRK
U0H+Qr1Y04SQUOD+GikhHIGfjtj9/L5LJW7856mn11p/AS2GgPIYy4WF725Ogu9GH6Q82rh8Bj+W
fxmoPTOd1TTMllR+8UF+VVOJAMX+rtwqZpMoS+4TlXLjRmK611sOJMWMvMKMWGh6sz8JF0B0LTlS
NNwagIwgeNrL6IpcupnrolcWYBdPUaXvClh5qyOaPxCdZ9IL8BbDSga5rmhXnIO4NA6Yi0svIiVT
6L6TxbibYehYDpRaMVO56xQNB1grjNNqgXRdY3RGNtDl4sJq8jWAcK7wZvYUgupuputLXefzXXEM
vHU925XTy/xVN09DNj6qCAyWA6TqgQdvb+NNIeRnb793TRRzBS8LTsl3uydw4FJDMjT6v/pIN0NW
84z0DR3AmfiM/8m95Dza1ijWVZmC5xNaSfIAPx/u8ojq5Gnouj8nJc8/gnGCkbqPHjAbERJm6XKG
aWx9vGyjnZ72IBsgctbp38Lg46mn9CfsVB6szfcoCas5iXT+PinUm8/8SPbzVrxw+zt9i3KW1yZk
iZJ0l9u+a+ejRmdr6fCwEZSX8HWO4TadVDpKlFA3OQZRPkn/DKa+Eo6oZGdnbT1JgqEgNDYIfVyK
8WOKUELztjjGYZ8+2wPqmoTgPst3AtH0CTEhArId/u8q/0qPjJZkLcB1OXCqqIEmgbd8BUFJnbLJ
bgtswWVWPPxBEqmlKvhN1LCf0PabopbMoh6jYZb/VBHamIsVCvCb/TGQvDHbcgBc2dfaa/3l7oBM
FfNsGD5vOoF7qykTrLefL8wdHARENhkZgU/vIvAnhcKVLpyxzYoIjqa0rozD2H8PRXkjjNGAl1Vb
OH1vp7bPhp00QfwDuADJPikET/bxy8NncX9Pewi/JbMqwzOY634ClcMPvhaXKbjfDiOWexkGKDz5
mC6jzBHQOMKjz0MV40YRUsR71VQMk3pKd/u8FgdQQCuJTHl/Saah8S8P2gLj+7eJCRG2MdbAWvNx
UJVe2J78l7rRglz48ZrAZa2UBR+JuMu/OSJ8RClyXzwIX6izQ966bHHOH8NU3DFox3DvB1KwO3Lh
4wZdXDW4CjE49Eb6rNNVi5/n6S1vBwVb28f5pm6yqh0+gVtKsMSA0Jpvv6Y0Gp7WTD2cvdoEf7LR
nqGzotGB/Rryh1PJIobb8BSWN95Fr/LkjUsVc3yEZjMqgA1bEy4WbFL68EgXG65FlHjeVlhkbDKk
6iS7R7nziZ4OxtBrgFbTTEOak5DI5id99hoREc/QFGjfHdmmjzVJt/Aq9qJwcToGkPoRxsRzuR2H
QdgAZqpzMw7uAlYT6c+sZKHmVQ4PS8EtsoI9pond68JxsB1/JliipgiaBoCfuIwYGBNwaJiLxuac
ygKoGHfrBEpOLdwFUt/VFbLIjny6jkSOXp7ezLb4j2ZQajcJTz+bKvdu+29Dt1dXnQB0/S5RxTuK
7keXW9GG76jjwZVb/1ue0Sk1KIYDQ7fn5ebr+nRwZobdhXRqQkUBN9RvIYXSt/lD2c1mgvZXHnAI
OD+oWtlGyY6s334MITC/zC3dMHUNfRwFVG5TBAtiaSF7cVEL2qEYntMsivA4/95GzX5fJEjHTc5c
ziv3rLHakSoXTkOINTzbKjEYTV8UZ3YRMYOVAEB3StzLiAko24Dw195WkstjMQt9N/7kcBCpSK3+
Hzn+Y1BiHm9ARGQOxHOtxHVyITmVRsCc0kQ1vrPcCmWAWQFfeH5XB4H4z2Agwr9KK1TdrxEFPDZU
EsCB2lmN2e5DlQJ1Kk7BC18VZ4Bpbx2DRSZD8FGOQruE5DUoRMggOm5lz6IYFtpM2OJHXiHuIgwn
xzIuvTmE/1YfCHM/YNAMF+2uBNEmzzbfCDUjm82pe7DDsvLFXhGp+gqcQSVv2oCG4vQPPb9H0il4
62D/Mj3AnPsdTNM0Q3BwoJl206Y92n84B6Xfrct2qNGAFaNStri88mdpOXrTdp578/YM+1C8rBYz
JZyJ+FdoSUdHgmS7mvVHrD3cJLTkzdO6L1JIiM7tMbbf2R8PrD9hpLmKRHGDED6pSnozQPD4SgQM
6cFcumwe1AceZENnX9to/jBZ2VipNyGfrwyIxraabgQb7Wqq1hzE9YEj8Bbws6u8QOlarnYF9hm4
313GNl3CMx3kv3YwmePwF4h/3Kq2Ud5gZ6fNdgk8ctdELQHawpiY1sb0/09tZL7iM/WxRocmb5Tx
OsvS+kaVRAYCyY6hpMMn0Dh2g8PSPrXqXBHGEY9CQJyl1l7ODurz06EfTYB1pq5uXBNLurow9QyY
Yn82R+gzgOhBblB73/+bGy+9ElNztrxCdANgr03MYFXY0RxePWSk3fiXwbI0Q1yKTEskDtkoHbGI
4NLdGricD140F1yxsEf19GKvD0T0ZptTou0np2b9y6kTKT8qtASD8ugXvdoFDN2lmzLhlpu/ctZb
YBAu7ijVVC7AIagemZiOixWF86UfFlbW6zyPBdefyNkNow7SUNZarB0tuaicz6Rfp25K7TpDVqed
FgmZq9P/1+vcQTTvyHUUT9zFkeW771q7SSXZgQfZ3LX7/ZmrWvBGU1tKc6Thn3l14msbV1sHZxzJ
oq0cvYQKjcYEXt1zDAg5fPKBpXPreWw82ceqdC24RHWN3lV+1au/9uDc4sWPHhW2ce4CIBBCsxil
uxc8HhKzuujFuYZ/FSHvJzYjvjp9qN8/fx5onxvSXuzqAowaiAI2IWlKDok24Ac+y/csLACbN3UJ
Fie4EUazUj3TpNFEiIfTHmX0bm47yIDQA6Q37n90i9b6/LKWkHtmMNYLiS1secE2EHXwjXwGOPUn
NGNkCxXqABxtOpEwWE+GEoq5VpGfz+9qLtx7O6nTVSjJ5lalUE21JfWJdKGhVjrWLNWvz6qCq9el
c2dL0x+KpHYSNDzix9ZnXbav3WtH7B9i/yJAkvCmzheF802JAMY7P2ANcMTj1c384+UheS2fzMp2
hzXwRrlvlkv9ht0VcbwgQA+faShTAF4PywyrK9UrwBl6G2/rPyfVOszBVQIv1Kd7bR743BH25Rtf
ZaXqLwHkW85SPIBkKKBwG+YUskv+n/MYCISPhq8EehvwlzTVThYidEldcnXaVRdK4xNSn6YzfDDu
ZmqBE5YU9sea6m5+/F6hPX2oO/GibuQvGHFWKAX6RgEtjKd13ADIMV8QKid0+Uz9+To6Y0pXsYnr
e8vitUJiamKOehtpgR5b5wvOhQ/kGDK+jSAmrfFGPIZrdhJAZMOCbIk7rZv/SqMKggo7wW39P5Zr
2ZYZt6St/prpKPouICeqKaBxlda8fGAKSm7oKgUubo0reVY4YRyCkktwL4ZYB3VDpf8Kx+bGX0a3
t5/0aqufw/abwupolq02Zst73mMUSxgm8tkFnvO3Wx1HcYv2Y/QZ3E2kkCAJbwCMA4MTBxxHmS+T
rFk+/ESsw+7Ic4FiZqKSY+t2XxfSa8Hxnr9sR/y3d1+BVyEo5FLndNqamdW53DOdb5UUn2YpHfB0
F8P2V2HPH2aLfaw3mIQc32/eLUlBvaGr0qLQxZIMC5sDTLaFbsG5vAHmqTO+BuJcVHwCDUhEaHbZ
sI1D7RAXNnb1WAYGi54+mXfsTDpZJHzdCSxWB3Lg6J2Bh7MlvUZFsJ/6IVMG/zZqTW9rmxwOdTtO
79Zar3xWvs2JWoM1PqR0TOHXenbgJLdaP7s7zz3LO+agGRg+d7ypI1/gWnz7AJkmpSjQ5jceCCmz
JwRGk7BNR1+TenHqOUBWgNlL7w/AskDATP2neEQvXgZjlEVA/QyMF2S7QiL+jBx2ggp67CZqSZIc
NhmK9hnOl5LmlPI06EeAHIXaQ2d7Q+GZfVdnVhUti2Dzo62PFG/alVB7FqQVgh+tg2AGzmndRmhM
qYpHHZ8c05RziMDuX50i38XlTFUCMJMVd6xdh+GCn2CxMJoyFcVnGbSV4BMvBDL+UCMhseK/SYuB
A3j0ZZcFao/LxcAliNV0MWwUpVR7dHAghKm4sYQUMoT2d9Hv9XW+2o6ZCW4HJLegl+RHgXTXW3Be
Yt7pcuFRqldrR1XbNKqIFJkwaisBwj2Qyn2DCfrWlszuJzXO9qpRX5DpFIT5VrPMh4ES64T/nFdb
tKse3lss/UrLAZqfS1rdrv9wFJevOmG+b8L0Bi6fvZcJGF2BQSMv7A8Bdp1RHMZrwfe2kN9FjbZr
Tq5z3GQ7KcSV9u0oLrkHnfWC2BtnUps2Nlp8sDqJokmHBxafbzAerv5/dRi8KN13cdhgkNhGJeWm
4Q5GRIU51FPkT+ky1gXqQrgIRgtW849b+o68AP39Sflgf37IGaV0W07eTZZKf8TLLnZ9Hl9Z64JW
6bPkrmKqZ4YEyk7wHNEyU4TGv9wk1vbGf+DUMbUodEHb7qqV/itD/gW+3Ytci1toHFzW6Hl6eTMG
LpgY1ottE5YHSvnhqotEwcNw1MtkPpVzfguSYkdcoQUu3gIVkZwPhRa5oECgDDd3FPDhJzDheOus
VxnH5GeEv9u0Y2C36QPA1VPEOEoLWmyQ78tf2NtTalbRFgw08azWgZQB+RonvSJW4Db3G8ih9889
ze3v3MnwLCG2XguqdS3hBJhWheSNo1HsiI1G7pYTIrzpCXYbG9E+DOTrF7UASMqClyzHAJI5vLcC
Pv/cwnI+Cs/lAEb6yJg+igSFUW0lp01hQqIMVEpI1tJ/SzY9qvH3KA3M3+Qk/zdXT78gOUR6sqEO
8XIP52bevGS59aivCtt5JByqATZ5Pe+LdqvTOpZOFA64vl9kpt/dLBsTe61uHl5kxvOEVdVYojcc
vo5wWWWFc2eBZx+hdC5VQrMOAtj3uNu2v/FFqzDGo0OkIvIZ9KoEXV6RhXWXki3jfbFci9Y1/P3x
1xkii/L9vnEJxxA9a6kRqq3y3R5iNcGb/Sbb77mNFvuYpKsQdsyqs0kozXFZmDBhttelmeGZY9YT
PdHJ5cKLK0w7IET/IQKj+fMny/TH+qkAGqCb3VfcM/4PN0KwPgjVZYYXw3OYUfBsq2n6/InxZilB
aL0tsccHa7FlU41ApIJsOGEN77wGNbogZFPUWnWl1tIEhSfOnoO/VMXLvctW89AXWSBHwhMzT/0T
K7kNGZz1X0lb37mdF/xR88CzE69C5mQPaFADPzwSElLinKs+T4MJXdiuKNGSOykCtlJTQuGqZvv6
QY55pzCXPGsJfA9CPJPGe8RIR1y2gX9a6ckNmH9eyLvLn1nM2tDU5+Kftoo2OBnMwIR9+fnM5dG5
IJFRECSE5IfprTLDtMuxywtign0aqR2Ju8SfK++3G50FnIblNh0CM/tluTxBnaFslOcPPVQZv+X5
kl5JZSr1JrjLKgrys9ghojNBP8zhuN+dRRuf6PwwQMryo/necgH3kck/Yd9Xh9lP5mxDt6SJ321V
yJ7/8eKBdJaG8rmx1ILcFWUIAhAC6j0lB6mtBAh3BoIfDyzJp4KGRxF/eSRNyN/mhu3JYhsDcnpB
fOxw5WsIVKTCBP5QcDqJqApbXvucHF5H+tohk4GGDklLkTMSjUq5gHn4Vz8DrLmtooxPs7e06Aao
v7mEiHkGkYNQxiPmZSP6Dow1hmBtv7hBbtfSxnjKuNH+05/Vm8T/cucGJxN9L431oAzQn8pWTPeb
ueD+Qf8J/7/LWvn9dOhdDGz33xk5v1gkbvXpcmmNDSa+5emo49s95qy3Ojpd1fmUdJF9QaH/pgUt
GN6YZXpYzg89LFnssh22K5iRSwDTU8yNWjUhP0usIoN2Yr0+o4/zvhfTNnDVPDmEZ6zmQAajPwp3
a78luweBGdLfzTjAhw4grnKMzVDMidfo4vGIVYwfSm9xKdoB8jPyy7zbfRg48dTY+p9FLKRbwkgd
2VQOH6fPZwZUwnpJzNHWyzYkHdR2rKQ9pnsPA1HD+9/5wbJXd4JxUgYX1DljusPWDRuWBFqFR24V
DynPDksvxkbq89fOLozq5//CnIBzW0uE+KtUUTn6YmvGKiZXByhh4/BdhZe7cWo2sso9oS2CPghJ
bQKh6qL5FEolr0L6W1txmB9hk+ocSEYXx27oL4cervfdxqv7i2cdHV7Qqb0NlmRksyZ5pwoAKspt
tLliqciR0rcnimPgTh4dXs9GarKt4mp8kbhaiswolVCzhhLR1UuIAn8bqIOxtSA5IB3pJ0j0tELL
+Sx34r8QQoRIgykHj5gDrosRd0POXgqIcg9FNmo/ljlpiKUPCHrAbxrTh3DFJshKmzkwsFhEkwIt
NejxBIXp2BOh1Hd4Y740+Gm2gn8D/DJB1QdELo71Et9WMQgGyktvz/OTAZrJa6fyqDdJuXp9prbw
aUsbViOYVY1djiiQJvZyM50YdjDQnSFpM3sLxWDJimbPV2dOeA0SnVmZZdgWaxvmBJjf3KR3BW+C
n3p7KPSfz5WiLns/7H9cEUnp5RSb5yNTjtexIlKmgtDz77icqVdhQp3hwgQV+h7HD08R+Iccwd5u
w8LYIiaWrvwSQTJLxHdd18lPzoyYtWokD25T52mmyL26Cvrg2fuBtKqz2NALhdAdRMT3n7XAD2ze
52EJaLjtu0U3JCebrgEHAX//svwuqOGCkIGhSXLi99YKOGCK6xuwLw/br4lXxDX2Sq6szXA8wUPA
0EJ8rtZdlpBUO/KqzfhP718/vHTxaLQ7JS6xHnLt/FshRoTFku/gEx+v1yQ72ttDPgQ9lAcmccpg
dzMW8EpAOcBwSnEGkTYAPLb1cSTVLF3dWKqxGSqv0YTE3RR4Dtp8QI8T6iSZtgNNVgMEqCuTFQOY
Ow2z1t7Q7bPAGlGzg7FRCswL6l3DPSs9Df4SVt43jdlvHFAzSvAQ4+ikY19PU0in7+jQ5mI4MPrD
RIb8PETlgA9tLXJ6ybtFXJgM9k7/HPiGeuYXc6S9nSrbYPj3HURhLvH3ASVYMb9nya2/GjCIngNB
gEji+3S+gUSICDETG9HJqJ8PQ7o/jcFKsEWMYvWxsIMMmyNtlFZ3fnZ3vI4roDQh3dGcNFZSSSrC
mzQTmpJTS7apeU75je/i5xvERtE8I6u9ZTDxwThBFScJAwsv1lUFiCjpp1tJkKjkdqqhEtVuPDih
kpq2zNMeJY0qYua+MqDdP9iQiSFdoy3Q9EWAXfKTsGASc4NdTaGHgYv7Z9LuLoCS5FTQvcviIK9U
djBPRrG7gXNa4S7AiYi1ZYxtaJ0KSEA2mP2Vj0P9UA3ciguKa4IWjAtisLBVBbv7qSaWSeIOLSYA
OU4Dp3bqGkP47QC5fKxPiX2+SrOc1YxWbmpfpHHGELeMM5gMddUWpc5GeKhgizXSgONWjrE54j4H
il/MRnZT/YONvzR2wvaKSBnAK6ZbMvuqVmDEQeY17dK3YzFT8W7/h+dgyWumLKNewBdecCp/WV2H
626CSdSIH9OE3Xtp8CiKpmoDtYc7l6ZNvsVdAa094bHuYrrnJpS20rB5k28+18g4qM/payLl2qVQ
bOLlITN1cYpjb5Os0fp4h70oR/ZD0F4fteLmBOXIDRDqG6NP2XzW355h51IHg27Zajm0GrMxqpj5
nNfa8/bxkLu3LS+MOToBPCb4/qSrq7AB78X4RBSKX2lWUwmHS2xjZiWYcgzlG3m7b4Z7jPVA9GxV
55XlEFdvcG9tBCnaL+Q+ywnyYoNZJXRmotZvxPt1eQWmEtbtnhgD24LdZwj68eUP+MzMs8sTYd6t
KG9uTP5ZLTffYK0z/MH+1GgqpB5cQAULCN7z7Sku2KUbohUUY+RZ6KRUo27vqEwD/Hccu+ISXsdb
ItlUztmmiUwv1ObcGTvlvSvJa7JMrdE5nDZRqJefXCXtjCoP3qxX3zqmmvau523FcVw+2Z7DP0SM
5XDmA4wQMb3pGTQbqN8twoE7w1uDJyFQp6q2Pa1uyqBCpwaiPnE0GWnSQGmBpSRgzOWCAKQ+e6nR
8REPX0Sh8QJt5et8WkS2y4LEl1F4PgaMPn32hhgY+4DnjGxjtbFYY80GJ1+dcTEh4wtxcxRpPy/O
3pqAnKyVxAtfH3Uiy7vrWVKOlLyfOSpKecRH+YEwd7JZ8Trpf8JlZmTEIe/Ic15gBoU3vfZai1C5
yvEVi30P46Rxl/+8GwG+nsmYTRboo9yyr1Evm0dgApIhvhCF13tjgjySGsPvawDr0Ke5vR2OunBZ
HEfXBQswOJGHVZGYz24ETF/MIzgaDEXqQqfgcYA/9Ki7nBflV4hE+NLci6UhZDGeu7mm7+i84whR
BiBnGd3rdlHZcd9sC/Me1V9ifYq9HbBDuFyoOkb/DtTwgRDX4p6GM2Xgdtj3dlE6g094CmqRIrz+
Q65MtoJAScJhz+J3Tni6LedkuUkpRI3EqAVP6ANe+CEdDo3rwdqggJpb2mGkOqMCIvWhyYp+iVkb
aPFCXetG1CEWg0zlzF10oAd6VAlkRo3dKFe/t+IxGR1kFr8PVbB1Eh1KEN7VRsn481/T2yjWMaz4
3JCkz5hZlw1+pddVSwn6SWZgpWnvBKw7TXhSwhz+nKicz/nhi49A4nbVJHl29rH5H1TrZN/hlxSN
v1Z1twjqtAF9VzlCfxaoqrFFHUkZdFwuNqfu2k8WFmBeA/3g0gXmwZw4JPvBqHXANEZWV3IZBLqt
jOr2BlYwVbtlxANjaw4l0z4AXPX5vz7e1XhRpIToY/Aui0ndJzxYdsBnDdTAYnCGp7tjog3YYnTK
4x3KOT1fKC2GwxvLrKl7D69qg+1wNPQaggzLTv4NOZqgIkoYBnINP6xZ6EaWE/XRrN5CmHKi6dRu
pPZdHRJbaHVRcgnaLbnEs+9McLEgqr2vT2iCJ6nnbRur2ebb3RjqV0qSlEjiu50yR1ZdIOKKTET+
CoHRKneF/JG8m5isc9IkVCRsbUzL9Vyl+qTSC8KaKyK7dtRIr2JA7Dv2eSZxsZewQkXDb99aNWsY
eplovGASVswpz5BbObZFk0K+MQCAJR435UHomfcM0J3W1ew1NNDug4vxYIV5vB7KkQRzFHhmoOmr
h2fqkZGiFRYBpj1R36lONoogMDF4TbNd+6/L+89uRSHHEHrE+g+7h39Y8I0vG5QAqs2aaDvy9DUX
LcrT/Nitzs8adFepb+gCWnkISegRnapmKHcdhi1BWfulfBN/dQvFucs2hVKHg9BtyQ9J+NlOaggD
H2ezhm4Sc+nexYqYpOqplm9CJ7MKeDe6+K28k/8Sjz/vZ/ajKl0wuOf5irop40umq26SbHG/LE4/
rY4E7+4Kp/i+AAbFLOzgIQQ2daWXvs8qqZkVuCANEXUwM3tb0/jLKEG+9DjSCRJDYfsMyw4sW7Ud
HcvRQ8e9sTloeIxbSfokEJKngYvYBz/DcUrQaDbA7oN31a+hHXeT76u3zFuwIGma8BLLCrfdk/2K
ib0o4gLY5PmiH0da8AUGS34GhLw0VzyJedhHNf166TmKRiM6ifyK7JMpnWCBj3XXFRmFQTlXpxtR
Jg18avFLhewpq9pY1oORQl1S0gQHxhT5mTD8xROqi1PDhQc/Bh0/aTt0FdZz+q1DOr2ukm+5SFfu
Z305JyuBB7UUlY/V8AQ2+B0HULhG1Ama9iNanpU8fz8Mw5moc7ic4VaB6j4W/fsrCVR4QBDPY9o4
HZrYm75yMGFhm+aQwH4V7oyYa7CUMsi0ACM8WmSY7tpdpwbkWqm4Gtgb4JG/OaRNJshWhRQKAtLh
9dZHB9puyeBa1UNJyoGlWTFg4RfjMwRaRSE40Z/PMdnbvinOBvCSdH8lE7KJHUgvTzF5Z2xoFEz6
0JKqJWW7STuolRMyaifIXbZlNFWLvIYJgZLMplZZx/rtqEIy0mOgtwdElCi0AEjFCb7erHFbUcNn
jS3cFPY7jHO2o6ZXcyUKkYl+5lJ8LogwxWCLX//9Oa4k4wYgeBqSWRNDN+fxM56HjXCFQ4RHPq2K
qBHVeRtYtQ8Wr5QZy6kbImyM+re6Lqm+ImiP8ahNNYujZi5j4wk0pPRXs7K9kt7X4XggXS9sKAoM
6eHMTUDGx+U3+AzNZKDdcRp1GFPXCVihH+IRNzZuMtyWOqnmyBg6NdW30t2swVRATEOwLIfcvvQr
TOXJ3O17sSL//gZQKQrkOK3xI39vRo+8Fqp1/Ub+W01nb0se9FuirNLuiphDXHYmLXw8k6vj3ymF
dZCD2CtCJTfXQE6LGZb2kA8qB6KLkkdPyepAQPF7niv5jy1O4LvQ2Ze2WprUGSI5b0vKqzxBqjBg
oeWvRxHSXj3tMTP9OrCIt5OWeo2y8a9mlut2E7+TZHMgNQnVdxkTG5AQA/rS/dLmFiyTkug1Qkaw
ME2hs9IEwZo2XuYSRK03fq1O26hz8V/4DqxJwLaSALZdJ38OD4EQ20S1EFxIxwY9G6HzQ2WNtwSn
/mHCCorixVHUb1p4FYEhYxMfIX+CHiaBA4/n0C0TMShqx0tP0O8uh76lweSP3iVsbmjk9vgA11uJ
oa5w1D7Rt8u1bFXmQ9Dm62pNI0xjhNF93C0qjpsyqPlQAzmfiwG2rj1/uYwvJmYa+0XthrnDFg6u
8GTu0HlDSfJYxGZCQHEkYdR25xgt1kQaycbHLQb8CLsYlsdlauCS/zId06v4WzZOAr/Uib66ZPzG
SKKm/J3SF04hUKCrKoZPIcwslTeeVPcJPGfizfaDOAeg4gJS4+rms87NXz60cfejABomwyubis+M
sRDuAkMzOodZwOouoFYYC9NMpkF5SDNk+th3TjkS7SOxiFPfHeEG0Hfr+SlMUhqFzznqYZHOVP6R
MyDaBAAB9wV6LSmI1BXJtB347GPJAVqAdk6AbZBoPow+TlXpglYUnylJybMdxVCKdc6APGYxTup/
TNWAjJ/MaR6Ore0BxUnvz7vYn0G33urI9zmZi6Ch5BLe9DDpsF/y1jBTHu2rz4z5Ht8DXzJdos9l
A6PBlO1drwalFg3DftIFIc2ATdenNdUI7/U4VL/xaUUD14SySOjf5LhIn6mMaj/u/dRPH+sZZ0Bp
ke/F87BvfEG4VNBmLLwkAy6/EmbTqHB3O+eEDNqWLgnkxq6sWh1QmX7RB8Ioxz8QS0FK3S2QjehY
m1UNfZQUw0vprXB5lo2cAhZDZtP1WwnBX0cEEZ9XQ/37VbkantLIYhrb7QMEbp56KBrnocGoMr+B
GwsSXOFXqcotSKO03ll1l58tC8rp90W522ZNpJs9wFps9agZhgBSnSJpTGd3bSYO/n8tefSSOX+7
xWG29INDorWtvOAq9PVIH16VoVyX1rPnetR5UFzy3lzVG+yqkeB7EjCbaBpEWyaKoAsAlgQ5ERHF
J7wd2YdHIGbs0sLqf9GANHCNnN5jmzdWYLFcuXifQHfuLenLNCdX2cfzKTzi5ZeigVw1k19z8XDE
fEmT+XzfQekxX+d65kF79k5OiOBkdB3IPDJDHBGWk/Pm1iCmsB8yr59i9lzXr2hj4kaok/eCVUmC
noKja0Vik7IeMwLMubbVqUdA/ei6p8e0UVD6hZL481uabdDogKHTI1HwwyjhB46d7C7RdDTcRZPT
UE6N8NhUOwNkXs/XJCEM0yBA+L6yzeoINHj6NiEY8qKKOiIkETLyIxjdeTMZFXcoPkx+pEs6fnkZ
merbejz+2tYIq/6AwXij8+IDP/kwRkKQAXkRc6qYChk49ueDMcKE/0a4hnYrprroWFP6sEc//Iq/
C6ORkkGpyZotL29QwYMfgqQ/gFdEAmF/CeumnBFy52tIJ9LsNEV5pLU5VSyBHr/eWUVahyXv64jY
xtwOz2UdWyCUNdZ7c1gr7XLz+MZ42q40dfi85meCPxeMHnWoKvPZKSbsLFTUPRWc8RmsVE4p5Zpd
GBbztUycrF0NqG28d+9ixnZWhf9HxYEEHCfY2bGQGb4wmlJRKAxL9Rp9QIftPhDWckaziTcEu9fm
zrwqf97TkfiZmruin8UWMva56LnmpZLHN3mPo6sfv+Tz8d49pWs8YJ+sqpehOlTSzvm5DIzIDVmp
ZM2T3LV3za/B5MoN6L6RGWbA7FzgwtQEvNVrR0QZOK1Gtgefwzt/wIy6oh+k/otqfZXkwLPnzoKn
2Gwoc32m1sY9JThvbt9hWVxc/vLI4okLMwi5xz9/tsUcDLMhXpuskfvC8WmJtqojaIMCLjUvmh0o
mg5OELHvoaQqTnR9zTJb6eQMsmOphyv66z4r3ypqkZMrGxVOCZzIMBz8FdvIjmuH61d3UiRYHFzN
9QuLp8svxqLzdEhs/R3l1mITsfYlDpuyvyv2Gfq/vvOw3pdRynKyNAdVGvfGFStDqXS8l5Xv1bW0
AjI5yTKz2a4FWni/tzvmsX77WjX96bI8OU4uJITy6FZ0JFBE6Icl5W2SbIhWMPrgaa+xrsmep8v1
HDzYp2JY4dUrPykkTxHKF57UZ7czjsBHg/lhRk09HbJYRIqpHsS3PmRl34BPovqM+uFwMYOQPueb
+Az/Czvoo7YOlHj8Cn16GglUopMMxl9oi6j+jK2xgQA54EZYBgyUG+VbnJ9AdMqd/ifmnYLXWv9J
7jl/xwaMcX7Z/UFmp5Kx77qWeSAkSC/ecmTyeIbOgHd2RYW+r5YLE0rTaDgo8UXCrqMsvBd38TRB
4MOobBTCqCKYBbTwDeFY8xk0rqxhWODd2tJ25LpyNum9NJ/DGr/CaogvZC1tsYLTx1fQASGXTnKj
8NHrqdpTvRzcMHN93e+ECFb10Ya6qgBVQwUh4ZXbRSG/vQu8/OSIMkythIvR4ygx9NnfyyI4RPkl
haTeCt+SRLb+4lJGNLaDUXKeTL1QbBEMIMZjsx6WHslGaa5Akln96w65MwCzVIXVoEHXHVVbfmxA
GCPZSONjmOXuQQUFveR5F4yiimVtgXqHTet2WY7a91Ctjs0TX5u+7JKta9Dd7k3a7F8G1FCDifzk
ugJaRGESa8l2kCOz+vWFbjex0MaTcdSXS0PhNmAxzvpY8DNwmpImKaHGuoD4xv1FuZ0VMDdbcwbH
RgRZBbArdCIdHPKtp/8CWZEI4KZzbcKi0QA/jONlwDevaQg2UG+Z8siz1ZUYCE7MEIqo1psl24PS
7qMCICT00YylAWk2MEsiC4aS2iBIovUY1kXU1qhMl0hu0SFpXR0JqgDPk83OY2dom2r4JI365vaj
IXu/RFyX+1Tzz4CL+9J/1t0PzWKgFsYVnBQT23w21NEb4fd5uuYnSdt/K9egIbQXDLthCPXURTq4
Ls4ikuySDgIjwMs6k+m1iLd+XxZNXuk5wzgPqDq3LB3U0zVfYgO4dIFxZYaMnH776stegmBrdkzn
ognmX/Kyf/GAGcFLnTYnKqmKq4U4T+1IWadE0jo6UGJylqcU0rYi0d5Q4RABORm1ZPY86NQxfSEN
8ZLb5NKcD8QsOkEHbZMlx2uJ/VqDEgenJkFS6PDohA4D8o/39ZhnZQ4C2nTyJkvupOVygR+u6gkr
tbpawmrkIKZ2BcGM6YsLvFkb93+Z5o/aIgieVc64Pov8zg2gUgyCmjtGQuhlg7+jFZUzeVCz90Kv
a3doGgcLcrm5gTjXGM8cRg7ayvXt3yN5LIh1CSr5AFgOIDtvFYCbDtihc+9L5X0A/1dsXB5GPZXj
slPa9ylB0R5jLMRj4Y2KSlBEWR7il5E17pGid2NqglWmtVvVYc40KUu7SR14fA4Jwhm0PIM7VgsE
scumYrlcDb/ee1CCpa7WqclG4G94Rld1O8WQrnAy6HxSMGKj+BZ0vTL2PZjz+hHmTrmY7R7qKf5W
SDrh+iG/gufEbI5RcEuw/Yw5HQtotJ3Mp6lnq3T2OtV7rGBaH+bsNyx07bFBAsPx0JA3P2XvLIJk
ddTwhUJP+dRE2Dd46j8M8tdY59cC3DQ0lHU47KwJNb+IpfZRXZVPaaQS435V9j3dlariz9FLiMDK
HjwUZ4I5pEkMBaXvjbvLtij4MtGyF+hAYTzJ4jsukdEqLKAGL+Ofmo+vmSx+9u3Rd95rmRN3MlK6
VKTWuQj5e9L50o6qFDhKGLMK4v7EOjXnmtUpv8OnrJSrJSNMx/dKNMY8bnZR9BD1PrtKFyhyWFlJ
rU6bM8OadjyGfdGqhEjo1vnw0q9YGq3OBsZhZ9g3bDCJ6Zg9R/symq6dfs64lj+ETJI2RRTiy0qU
LAal9UWe0zeze8gssNCLIqzqDSvvYtSr3/i+ju+zMBimGjPi322Bv5xzYL5cLTbWp03x4iT3B9eP
Rw29YLAaYMXiSNmEduK02rsjMwt0/7sX8HG9CcWB026oQSv+Cq0Z+xwu2WCY8dFCD5vwfnzMsowf
HSLmwusul6R6cx7M6XoXQGHMJ+CuyD/IVSar95ziLjw0Bo/b2GP1URwOwgQFuCQYEMlkwX855xiz
g2AZGezWNKwgx/mgnZUr1PLEtVjRDAqFMF1he0S01XvburYoTZvIP20BLKM2hliQ9sK0JTjWlZi1
BfTMoZ1VrKwak28Mks0EMWThm6rUj1X0LFmLU48md7jELt6s4iPJxbyC1s4b13NIXZCeew2azLPA
A3ydQ/F98/9ie79fBH6CcSR1mw3Ldc8H9TCpPE/2SuOZaefuSME73kwfOhQqHft4Snq/b77dCRXS
iUiaUzwV8IHEd5QqW4o7j+Lnd5PUJqvTCkqZrEpeugTho9eXCTqUjK5YJIA5PZilxdofedx8XzDA
TiEmrsm2+pXtbjcj7cWJSTk51MPXnNNLgi3hqetzxvgK1UvzWIS/IdPZbY19JHr7z/D6Waa6cn7x
ILmizZpOzXAyBiFFM6oU6TlSG6ut3oeCy0i1acRzzMumiUaJ7jFNna8/O6uyPYN7hNAvHXnmJXyh
Kqr/yFZ5FTQcm0zUJFiuNX5Itx6dctNY+wM0mVPmMv0wWq6q2U4dsS1mvlZoOLjatnafGawQrNiV
oZ3NnYrHwLWBBo3aVws4eiT74yYhmQB4cXqUCFxI/6NxDV3eD89uTmnLBnTq4TfZoJ/yvvxHsUbV
lZlc+WRdXagZ6aVIZf8aLKjxfllECB5w4yf6vWEng2Y9RSDtW2eaRjRbtmmho1GmUjHTlsDXpD9v
nzjCNHztBGfOXC+TuZLiK2Of21+pUticvyq09KmsnWGuPQNJss2jMdLRoa8222Q8nWT7rjE8OAjj
l2my9O4MVN7V762MDYcXQZWTR2VtvCridpnqsh7R6IQPzrZy5qZNuxkccsrAQ8yZH/XnXWPV15hq
6nK9OE1xKJZRI0ctGT72hBJF/LvaW6FnXPYSlqxr9iFgQ4CsI5zGA0AtLcZgn4LdiVA82kxDLzZ3
wqPA7bpBX+kRRosSgIepnjNd0iZUFjoqUfEFwcroQ+uCwNQWwt4L804+KLP9ECsT8Z02Dp7Y7n5j
uq/m+WE3Oz0h3OcFY2EYK9AOx7yX9z8Q6cvfczCtxq/3fxbDu1bL2WisM2MYBitHKvq7gkIb/5wr
jKu0d+z1BeNIGq/+0ePmxzALekqDRw4nvrXo/rfosHZw6guil8PI6TvjNUHAxqIGcNCloW15qT3v
J2EnkDKH8VeN8Gs+nWrx7fPILcpYZXlI9RRyUjbV0EFIe64Q9kqFUb+y7Ic+Er3sa/eecoE6YP0a
+6jAoUGSdin9q5URL3Yq+SDuv1IwwFEB9CGZ650yTClKrmE7XjemsNe49tprTtqBfUugktnntpPD
XfE9n1xF2GdtfADmcAXZ9jPXsv+tLe1pZ12vC6HYslBhzyVaegV5DvvlrZj5rmvP2wMO1/hiLRfb
S+D/DNl/THZICxlHJoDMy7pMfUx3RszId5YttMNT9RNBclebwTbnhwVYXt9NlH2pQ7hzt7XcZofQ
Nyr4C1Vvibmim4E2Qq1TfVrcTL/PEl8NOIDwavN5SQTwOnmodn1blsK5lsSu5V8cNBNP2rKFkQE5
PK7J9gQd5j1QE5xOAjXHJ9xF2nL06yrYPAKTVYoKEvpreR6XghYpnfM3dO8oujTcEM/0qEbRhE7f
0ifZ4slgmmVyiBHXa87kwq9ig/eESXn+EFdoFAEuCpvjtQp/9hoFIRqsnn8oK/SYU6gwXB2HIhTi
MUPAb4mV+uZ6v1mkpqQm6cPEQEwPqLCd13KVL0FXU3Ep95NlBFJ/v9S1sCrVo/fGfM7WjYRmNR4w
s5Hi15PP6vgddV4LHlRpsP5CF7G3if/BM1b8XAGD/16fng+7DVwwa5UlOsfrhgGAsqpSx5ehw+qr
SP+8/nr1GvLgeUXUdpFuG8vB3l7Qxyn7N6xIGyA3wgMTXEY4700sCB6mERYq7tEInUyggMal8OyX
noE+kcOUEVi6PKIaL1ZbcovwXRKX/5VBw+3D+OPPk63dwO4euSlLxBm/cpEGEqXqXPBuN8k70AcG
H9IqQXlHLYHXnnfYFEiCMY5yrlI6OP372NDhOLhWNY6T9rcd7ciyKQ4LKCtFsRxnU3Uh+rtj0Fn9
Ig/ryZA+8+Ui2LjTptkyT5D+eEDdNDfgdDv3BfH09gNJsrZ2EiTuHk6/MKVFl5GD+7QZKx34RpFS
+XAr9zNYQ4Dse5+K10Tj729RLPdGLmiWVgj0jzuqH1nP8MLrVkA7gxjugnyK7yt7Ubq7Rl7HCH4k
/JOaDSGX9QRC1UAg/tYX23fcdlIENlk4RvWvI3O3tBGqEV9KrtEMXk1WrwvNUCp4v9rrWe1DxAcK
ogEb3lallIvkrF5PXUb8va5JomiQRFLmvRBfGYk0rB8S2EzwFWUKFsQuFKYI/bZG0XYnnGmQxHdS
CfYG4K1scXiHmvWelYZFjP0EvD/RXbgU/3Ykx7kouGOs786KQEntv4XTPXRrIgjk8z217ZI9/eb0
1HVWzraTJfeo+9a/ARdgIbOlXpDpoPruEGHTiftKArB8eF/NluWfvGVtZczK219i6I2dSsMIFxej
o955DkBwRAERNQoc/ttvFkOgMZ7PR084ndRrSsA6Q67Q921uDFx1ATF/1SvMUdhT1+yL0au9EUYV
MLj9jHBN+AMnoVuipJ6rTMdZYWnfxeyZHPnT6bYfzzq4yEuLWLOaj2oRawq5CwZnHUd0WKc/MAzE
zUlB+tpWfHLjP9JaQNEO5AeD/A3nwUkHm3qrAYTH7abUkYNc3Uzu++5Gt3/2vd7VbIOXCZIp1ghM
aLejif2J/ldgA1/WfLb1w8jyc7ZDKyXDr3I+3O5QBiayLlpH1aMLnVfeOt/dFUoDZo44R9TF1PTx
5VBCj3boD0vWg9TxB9ixU7tKYN3aogpSNHpzFSriCnvnGQdtdfDlZoZRPp+Wbzbj2oYWXvTokUxu
3LlOzFmiCpArecEPcTjSnqyRPIpAUZKfvrR5rHcL5g7CWgZme/gZBT24Sm4OCflBV01bT8uxrxvQ
skNDdt+37/sRvPwNvYh+ca80CuT7mQN6OKzyoTB5uN33oWdr0bjOHyr2lSUv4NINNeOzJ8G4NuB4
iFLhne+UO2ptNXJSddcS5EBE1F1sKJRQTp6jN7mLMdYj2eb3PIhbxXvRNgWA9pAH8a0Oi+/tezCb
d4rrzG4gIe4Mv5HAtYwFn1j1zZPCu38VFoUyISIEHpFgufadfGulwSRi6EDuetoaPe3ibx014uij
7eX9GN8fHVh3n6ZdQv8i5O25ONp6eAYwFC4Gs5kxL+qY/ejJ5IKgfqNwGPrAPj3s1cOssOsfZqiS
VGTmTlTkVFXVEKrxu2zF+M9Klny6JQb9Bywkkf9qYgApBjd9c1AF4waOKKkG/XF/NMuyd6LQh3+j
9o7iXNqdpRqMcIRlZUcILGbS9wcsZdjdDPRYzOpsQCkNv+pgxFfxIQQi4w3gR4eP+jR7nxwQxBNQ
wQ4UawmFjLlT8eBp0unXUDgUzyevZpLQHCPJT+tKIp5PlaEFo0sceDTHoye7O/09fVhpMKxIXMdD
5ngnv/ppUwOPgpB+ClyYA/+W6dxNjegp4hThF8WBB5knr5Zy0QWhejJw7NuMBfxgePDnXwMgzxTR
ZV7lYDRcjeAf48XvMu1Kt3DXi0OKldxVDfrBvUcktSvs7UYDg0VxyoG+jdu9c6G5SRnoUF9Crys6
SdBKOnmGg0uqBhqPCiLP/54MymhkgXFB/bpqLra3aGV6J5WZC7/m0INW1S8i8tVWeAgvaiFdX1Lm
abXdyGE/ugdYtvJO31drpIUUwtFPRnRPbkfiEfa6MZHNUE3Ij2GyMIZ08jxUwfJDw1PMG2WHDuqp
lYav5STjKHSUcaObtF4dVdiU9tv9D932MizCEPoCBPe+qPRAsKpUCiqj6bLE8ocrVp8sjhuXNWLn
4qSerePwUGHHhhbTi2piDdPAfcTIjJonltqFLsXSNrBGEgZCBzAdGv8ACJcjpnWegUO1V2Nz3upy
iR9kNH44YLzmmMfRIRmqR6oBBObVbTcF45RbaYVIQomJZMkRye4Mz/pGblUkN5xf8NYAdZhPpGCD
grePUvMzujVosg1eomsGOD8oslnRr39FQgeMMYgVliX4M+eV4MvkN5w0q5YSweB3SS38MEaSMPWZ
/jrx2K+11/dt7hxv5S8XtCVWOYy2kLvDqfmh0Z56iVxdSfZEpNcALiVhZU2Wgdd/giXmUz/cx4HC
ad5y0KTfZq8ugc1Wrxl4XIDHQA+qJez2pgPa7N45aS/XHhWBhBqXRz9RayeRDpmqizaxuOLW6xLY
EL5g2EMI04gLbogF4EVUIxzVw38m0IVXaa12KmoKvnutEJbiVuhM6kjmbEiNLTC1uHtXk73+PyPZ
ihVjgaJOpOqWLYBN9lPYHCgXZeDywtvPlYJpY67xe8mS88ZLdCBzMDtlT1QODM0A7+F1z6/1eGfq
QLPDD2l+Ij/t1r/jv7hrTllUAC4ycLxm6EKi1k9mFVgyMVhN4n7R7yRfudxNJkWQY9nSTbDaR0y4
VgJaeH48PtLeLAzOi74nPnjPQnOXluJlqt4rIEdqgHmBYFB4wpAqrXGxwfGYXSEO/Y6uPa1j2QaX
FS7Rpb/xXKZLBx5Csmxlt6ci7KMQD2IPSNfPsxJvLblFvahJxID/HY2A7QZnrczUjpUzvRxixLkn
TWBvjSzG8U0YyIkUbi6bizJ7iUU86+vTeLgbBiV4BGusdsAE0ZJBaD/dJ1AehJ+xHC/F4FSvS6TL
SEv2pYnlHr0XVja3aQvT7yrwdLF1FQ0kKJ3azB7bohYWFkLQyw5i687uuYF1VqVtzHiVgVWB9lZ3
Tmhh3ymupGqIch7eE/CZgg/WTDQ5uwhnTys7dsCZUYLAc0tiDTNVhFbKHnJHKxxtRrz1azZcJl+3
7kRrVzTu9ClyJ8uC+UKbUjhQ4n4KZmNaFun5u3cjftbfU1g74q4EHB9yllhqy23/KG+Q/0OUVuMD
AvnPt0tagetndTSLQ2iSzJST79JB7kSPdUaTjAAge8il2EQ4UjrbX79aTXe5EbnMt4LHDYnTud68
g+oDCKLzEv6+U/8ixV23QUCtBM/dVC9ZohfPioFKOzZEcK6ovwSCm2PNFMDWBMeDmIvQH3pvoIjb
vN9euE0I9ZuMxcw0Ad2DvFGi66OqTHwbnakztE2r0+I6SO4O4CX3VYW4G7qaJxY3Q56x6CzF6XUz
9nHe0YEocOZ3qCVv5WDiLtxN/yrdjaaWeGsfUYZpDt1uYgsuzvAaIQ12e6JaliNK28CQwJmUqvhN
pPs+pQov3qDIvv2PBTJcoG2ONch2dFtp4HkgSBCMnnUKgR1ngzSkRkZj34H+kj5WRwm/nsufP6BO
xE3TnWfZyBIPAUiJElNJkD4OdTgdHRG3ze2xMZHJrDkqjCZo4NYWW1V65URCD/mrLuzEuuaFTfu4
3z/m8t/hs0ivac1z3LJ78rPQjAlqzyijlVTPSeh1GoxaSsOEyQZPQ+9OVw7EFNdJbpEtAdkBBwcQ
+0kO0zO6/ypzPHuelK6eDDuj6pzqNEUveYKGutfEYzm8tHsL+t7Nkqwr5TpShf0VS7ML6leL1xnW
gSH1LeZQ8DIH5R64XypnP/eS0xAjW38TBQKReWIvmd20zsprbZOaNe8xTxRrvZBMhlFc6fkEKIfC
4xtFukjQYLLYaOYDJ0syq1QmxegpNXTJxCtnFrRaCr1SFkzoerZwTl6f1Fj72pkNjWyRvZuisjSm
x85vnbrudi/OLQzlcHH0Tf1Jg7juoCuxHjYOQ3ctynzLrOB4clALZ/a64N7uU6mt0XhkLx1CpNYA
c+PuTV7XBH1+gkDE6/MiXR7gND9Ld/jJgILWq25wWoTBfQGdyFKuBZaO8Mc5reFd100nQF6ODvT7
SBnIhAtYUCLj+7klEuiTptLJT4LIvva0YGpMafOH6UAcF/rit3raqszhdlUZG1z9QJziJ6QnFeD5
V5qnanRsoqJTA4snCLXYDFKCOO3RrQY4PLJWMKDZWrNtpEFYPz/zg2PleOINgmM+qz0MXD3JPdlF
QjLWsUyLBzbbjzrh//LWKeOBvv2l/yxzwBhu4UzZFuaZG17N9dXxVlLs3gw1fT/z2JP9Cjh0JjBi
XBEZLnNXmJ+vCbJUpH/NwuInlGmc4mMOn7oolls74TVfolJ93abefKkz5kN+ZO12G8jlh+cXeubU
cRTtuHlVYX+eirbe0K8Za5oSyxnE8w9zQ9One75DxcIE2kwo0lsuTqsc/hB9dh1j3l3fGtP2kyvo
F3sgCv6uc88og2pwLBh4Uz0IPg1c3j4ZbRdDoGEpdIrz+dOtdE9nNUwiu0s7yeZicgckoT5zrJrP
Egkfupzwqn+WUVlmxpc+rUGomtvoBEMIZCCwMgGdnJW+E5yTI5ySM/mbs2xVDccYrSmPB9r48xLM
HGJjXClUqC+EkjYVd7xE/AHOqGUzF2yv3Hs6Gdk7rw/O69O1bQ6EWphP2cTQMVor8I/Xipk+YOGE
GjqQUAwly17dZI73SozbPwl6X/aOXifpgEcxi5ivouOE7r06Ty1a3Py5fBYTe5K/Tt8pmvZjSH1L
jDrdvEvtdZDO0o4hR2kq5oFxx9L2PsBZngn2AuItH4iQ50SrXq1PLhLCiYFT5lHPGfIEZQmHb9cz
m1+d6uIQj6Hk7BxUfGAgnRD+bcdq0JSPmBs4k23hDH1QZxJEh1SBgVkUx0pEPW1KyMOzAtb8aolG
8ij3OI8AdKdovJFdI+iMa881I8jnyk/XhY26HetW7E3Bw0tHh8S6EFa/mbZwps1zmBAIqXiQ8fUI
vZ1P5dYOb2i7TMDGEsS8JNWKu6XIqojt1cG5rnhPtsmQaC88R/7Mjh1OllgqJ9LfEiwgTdV8+JI6
+8LB6zdNtTbFpRNg98NXZxAc/mHVkgeS5IO77ekCCd3fPMd/pxtSufOu35QX9835hyb7Mmm0QWl8
0BRNJQQcnF6sWWAfoL7yBQKHTzviQojnxi0aMB42J+kiINOEw2X1BS6XGvBIaZkkn1MZDnJtyM/q
BV+Z7+qoS347xieVBzV4iTWwB8pzDxxBRMuiEDwQ/l7cdKrSp2GvBGSyLoqJW6OqG1WUb/ZHRdG6
QZFLz7gUjW7ceseieFYINgTzytGPkhREzplHA5XqLCLHDJbN3ymJhJvvVNuageMAX9znBbfBc7Ui
U6p0VtEEsaNkimZwtUqY0Goli1CFrOtu3/5AL+ODnaGfum8CmKLZffGJ8FKt5CZpQ6j0ha2SLgjt
eQkdyWUhT0JsUYJe5FThmt9zmWcCIYwKw365k72saUyt8OmKIH7REyXqiaX1wfEuD2rnjpfHjl6b
ZfnZXRUw/wvmQNJy9Q/9XVlbm7cOmU9uo6PrHgkYI17KM1A1OmE3m5dn5IrtSQEfhk4/DxkK+dYM
LlYPi7ao23rgYrsm1jcvSUU3MbIj3SMLQ8eTPrt8AExLnO/DM95wE9lYmxlKKVSDSPgwkKOXm+P1
3i4TLPIPdY41shD4hcfyAGz5QmOyeaWH1puqWUXtdbMOVFfYHzQedO4ZYAgVHt038zZqYQ8Q68RI
Q7Tuqy1a1S8YJKLVte0apm6EyxPfpyA3IOnTB+n8B7vGtc8i4NCHiJm3SVz6mkZzfhCg76ls6OyB
kzbDlXJuDoRrGP+zJxXYyovMIFBlps2CVgKQSr9rpsQpYd6tofRNkymns6ejijE4dh3ZDpIpDEBK
BGLnQF2LpeooY4kIoaF6VCcroZd1LZVcnM9MK5yAxQlHhPimLIxuuQMiSbmLk3bnWb4KjTXYn44W
iK0vKaPCliEMFCGZIwmm4olajWbPS3rrLsrU/tlw6/gmJlWZughvb5XGX508pNKbP55TTR05lemy
AEOpJ6Sup7Jq659YQIApwTyMkF4z4FeSMjKMq332vUUZglsBrjArFTWqQacpJxGcseL8uxeK6bQ1
2MjUjfU3fkQ7sTC2z9AI15IChL/KvxzAwCTINSaL5zXt/ePZusZpHH53jiSeH+lwY0lhv+sAdXoy
N7xoMXGLuuFhv9m6M0uX9YEDQWppTxjoA55BCgevOnF+1Uz11ZjlWRB/7DejMZlhBzET2TDOjKlh
BWYIDaxZz73XxNSlj+Yo0OrLJvQ4MIcUizRQMBMc8Q34/l+AMAEey2y3W8kRM5NfqGs1QVmeCWU3
/6YSw5Cf6ZRO6wJGVyeOxICVXclhYWhI6Ihe3Ch2owTSeb7UFwKaeAVSreu/mE9TT7EKoMBA75cb
E+3aF2F1Gjk1166HVdQlNP//SzCQltKhkn5Oa1Mh5kiabCVaHIaz6HAXYrHNmRXLWHQQbPF6N/S2
6opsmDtxkxHPByofNmpc+w+1z7vUHKIY2A2UmeKVO89gXb443sBlqGCC1JUVJEHgMSdGeV2U1/tT
d8szbhul2wW2SpyFJA+d6si1lMZ7ige5AOCjUTl5MV1PWwNm3EZqgDkM53rRKCt8p7mWiR7mE53e
cLjo9wsfhcVas2mL4T7ESgUnKX8nU8lS3Yp2dzUqo7pcV6I6apP3oyTn1OduWCtOHzfS+2aS2vo2
nvlUPa6reVUzXyzlRoDQy+l7m5006GpxFU+90ldkc/lQ28gp35W55T65Pq+DelVP1Kt1+qqyL9LU
fdHqAiPfhpfrMZrQ4Yv830vUi+cQPlCQs06HcgelLu5n2pHm4Im6ly0jYz78l77dJuwe50hNLueO
nW6PVjvphmaLU0tgIJ+oozt4lU1PqtPElfs90GM2dBrn91hCYnt7Vo6BLJHl9j2aq96H3umM6t65
X/4NNNMzwuhEtYVb1XJyuPzDsy5CICVEdg27HJWrPy9UnJec7mMNSjGrYttrzzYRiEy+GwI8Cbeh
nQVVwVHtojjLr9lIenTkGgL2ULVTzUk22aQjZLG0ZgFKZmVrwcX+AMCA6GGx+HuqBVOMvHWHXObz
CS3o/lEHU3Rj6URr8VnWnBy3NWD5KCxTsST7RE++gcCewFb/7j0Nn5hOJt54A32kACLDwECNTdll
5Dnl400gth/6AX/bbdcZllfiRAUeKs0dHOUMvK+vjALvEBRyo2HRVmWLl5mW/2/aa2vTRTgbAGHI
3zDqe2WNctRhiDpI8zStxfAfODWStf+Uxfsr18PSGKAu07SQDRxcccju0Bw1T0peJEP9aZv/E4oK
3v3thcexVvtIX9TE9u606E26N4uHZmPfwrXjYFGm8gWcJjGXlWHJmrUQeB+tL4RkWuX9sPbyTz1u
Ty7qAEoF/d6eT4s/ypJzuCF0yMq0aYrVvFIbA6ifmSbfKBjuNitT10m1Vhxx6BIC3Gkv9NOHiDiI
t9W7MfNTSw9IxTzpa+UO4fRrVDQZK+3gXLrBtwa80sDNnr5LMiyqZ3vNCwtISW74vMq/ynLze+vc
X6X2SSS6+CqaD8bTrptkHeGC0Rtsq15EP+Qmch/hPJUc+FAkRBguf1qtWHDpClKG4zdryTCyVzG1
7rQFdKppOy+AGw1anSDyb5onm298KIAzQCXUcI9oBtJO4bOp1cLuyg36FDpchRoMjHaHsH32eT0t
Bd8QnUZTDraE/jobfakEjdDZ2dHkkHADVD8fXdOaBRh+dGd4KtaVTrcvHP/NeCux8PTuj+E2V2Oz
GXkonwgjua5MUBRMs3pKn7lIv2EFY4Y32l7O1bF79Zwh5mmJv8cwPBpt9e4xWaXdIpADAdzNu5g7
Ui5zazbwQvy3SPaWAu8xPJlM5PvYzZ33n1Hjn3m2tfmoqH0PXHk3tT08QSJ7Rc8YAb2DbDz2i/Pf
cYqzG0fOwEpH4ujjyiiF3RavmovDp7FzxJ/cm9l+714DoE2clU5gZg8LGr5neoGdXGP/fG0Mxc7x
51kx1f6cVu3k8U1RC6oZo3W61JWMruKrBoQRulz42G6U9IsQ20gi3kO4YAlt2sKQ7kVgpW8Exs1q
AEkYWm+C+9Vp5W7A+KdHMPQa+1vefo1126LZxMJuICf9uz7NSpMlHaiu2TBmZWDBAYI8AjXLUvSp
w73PFLXQMFT0T+/bpH6m64Cdxd2tEMvgWFGqYEd+KlUJIGCObQoipkUYwzyN/9xd8kaJkN4WA7aa
nAMjRealeu3XHvJ7AMgWUsV7g8mlWUxbtsSoD7fQr48rzqNZVGgdC4nInnDtElknnKVf+/edgK/0
7X4Ydx4Z8iTuMZmI10jIvMoBlMxCQ4iFUS6URVV+++o81VptjEigRW1swnrP3GFmyxaO7ps57lK9
JXDSpCimGXBQQlIJaPMhD4TcSFFFNIXveigS4dyjiimKHCObFtKqnV1bT2GjYLVC1S853f9m1OL5
NqzuR8OLFbgIZeihXG9rcSHL6qJXSgt8e6Ftn+wdIO3Od5lEdAHn60f+Rpu5TTmDrfCabgrdisve
BlEbMUPv83rFALrTUazYBn295gRC+XybUsKCOfomt0d0Ztcw8c+DRK8k+7x+yN6mBspeqe+hJn7h
OHs5zAO6kd0VLAhhkmjWRbzgOZrjN7thS8Vvk/R0XlgHmNHHg9W9wGOtXmfZ8xexK0fsaQHonmeN
cDrmZ0X2hx/plrlonHMKUWExFJsT/iEhhu6A9nelCnHDCBa7WcPZTrl+s4QbFlUsOIeQJLE5O1sS
cuuVTPbicOgbj0frd2zpKqSg4Sm+d/XzuXZj8lSYTbxJNmNXZ4reR2BIOQw0hDVW1y4AgZxd91pt
leoqlA5rRNmz4iRxENd9SieUaEecuTcJuv3M5YnqpZXVo11lPg+y1CFxmP0CEVJMONPC5CmQW16I
H7NoU92MWo+rTEa8N1iSJ0TVtErBDcuo191wqL9o7wi92UFBvGpUgNVNPlrfYsaQGfD3WbnH3yP2
HYCXrmgeai9Vo/NZHtZZlVN88fOkb8mvbd2OKXrFCQh4eTSki97pX2piJnKQEFLZoVaDpUu9/qKV
j0QrSuth/bxaRaGWOWfExV/zk9bxtCijhAVCtWmW6L1G7PdTGD9Qk4DUIbpx7NFL9QRYHAtK3XG5
MAL5J5+rE+fd8wEHWOvkB+JkWvJ9+7YrdR8DMEJVNI4IcE9d3Z/W5S1o2lDjPoURib1ZboL24Hr9
hCrelPmz3p9UR1mr6FxSL+H7QLuUevEgtUnbXOYk2zJ0b6yng9dtxONHYpxwe3TSrtEvyXw8jIDK
0U6vJQAayjwqprrzYiOCCHXTcLMwLrHqelhmq45pIv9VgUtSNgLupDWPvolj1K5KaVu0U+9j3Qxd
Rl2qfH2ddmtn3K8IM9qQwzKatfFppoI4hZUsgn5nHAU7Qff3SXelFtMIBUTwvBB+12C0E06+DzOW
0rriUIlDAEpEH1QOvmwUlUKCcIOqg8LvjAcAXj/ILAfU24DGAN0zQTZ1WgchawkMMlFeuV6+WYtx
w5HE+rQyXu/CC409xKRcaopw6UyszhApZlDLBZ1y2YghegipX/v0M68NDCTd7/TFM4CahBrqQBBF
lVqyCKno3h2EZmTgIRwfI+z8jH3kqJBSmxrg9wudoRebrN6aw99QFJYKklFRX+XuvSWI07c63lRJ
pfl2y9wdeILHT2uL+KzxsURPO69pXIV5uG3xNbAqj8qC1gxhfDmxqUDJ9jm/eKta5+pB4BCE/GPi
/feAFSPcPmWgwsSsQG84YIcP6lg3Mk+x4OULPt4OkaGZDaxB9OXQl7UYwWA9mYqtuBhaYoX7xIZY
2cg+gHYxJodRYF9axpsoC5dWpPeVI81IO4l8mE2xJF4fh5acixhy6yVidRutUVunZ2OfY+JO9Iml
Dp4ZcLvlLhVtREy5dJHwZPKaTjYxOzgUkOYM+p9QCLdGS/GlmpiLWuZDTNujP7mhQc5PM1ftEt+p
ffZM3SRM98lNUQ8lJN86MMfENLzwSBw5y70Txa3piFhT7WDpHRt5AbKT0uEuGhQ7sZeGtvs0vfo1
hZJU+k++YZ3jqrQQ4vpi0hsHp4E6FdvlywppREJgeAVBYt0xtyR5nOYOYOqe+xIP2g7FW2x6BzQE
61whQpX1WdgqGK+cD429k1VtFE+N3WxytQ9Z6qcnmx8jfGqpbkRHkfi94OHBd0mFcNZx81fpOHUN
mY6/Bc+yhdD3PqlMDabJmU22/meKBpRT6YJKa111UU8gC5CjHpcoiz7ncjHFn5M6TYSXV1d0Umn8
vJ6ZXP8kgIn78onhB4cIdNDr3CxxcKbAG36HOuefnjLsF/gLkf7MvCa+Ezb4QN3nDnNJopinrAXQ
y3AnI9UpbexVM7cBvVKXDdZzXfZsTCCnAtMSPHsXv7/UgPbcoXEzKxCE1LnNLQJUlevOMaM7xgeG
5bxijGN5/3Nq7iZgnOVJAs2IplhEIc54hgu06s0/ZQJ54b7PM7yZm0nygyhywcwcJiXxFaOq0UOt
Xiy294z9KccjRifhbr6L4iUI95gj89ganFy9G86nlCcTdbFhtDgGkMpsvIx9C3yKlk6BwB1B7JXV
uTOhYaKqC4YBb4G2+4EiRuID6SM+KqpZOeMH5P9BoXlgj/gjpo0AOG58cJ8LXddyvMgGw5FMWRYF
GoIqeTXjMwQgLw2N1jqF8yJ4UsM1LZB6gTAGdtfK96R5HAm/Jltm/87rIC94fxJRj+xvYj8nQxk/
BBrn/Nv9heLFqz2VKJAnfeq8h7gEgcDAvM4OYaZdModhBmmC7cdtz+IfDeskEMkAIuJKQcdaNIjN
7cW+OPNoP21nIibAm2qeZ6TVdGVtxm0GClvSHugN0yAQTnVdGapbkWaz4SPjuuo5T1kBL56kF39C
tOoPd05LRceEDCZj1XB0tvWr1tInN//epG20Tj7y5BD3LRp0R2rHRxT5rDxSAzK3/ardEDuukC+t
HqDGcYWGokdPbs5yut04z6FlzQNVPP9mmRGMkka+1eFXzSUQ/dlbLTqbD0lgmx/b+NPSbksZVaRr
azwsL4xEfbPd0l3PnMaEe7ZO2L+AkEUY11ChmqE9XPLOGUX6Y5Pz7Y/aSVEPZfjoPpBvZXf6IE6g
vARjk5nhnsLG7S15Wsh9/I8XjOMmG/iRPmOW4J5vhrE3KboXKzBZNCXmt0XdZPgoNUceUkrVLIU1
ZOqjAH87t94v0p4pnfNMOXsreZDCDrtZAa1NbDsNgp+AwRpQkD/l7eSqsf1oaYd/bmb4BrQ3HARi
kNBdKoJFw4BFNmp0U5emiZpHLQAGcQU4qDdp5gzGFSbajb6A4jC60vkqiZjAP3TCLEuMkmeaadxA
tbWi8qlsEtbCCE32mL1gQ3qOsGgh6pk2P/n12xrjag4cszhdCdFMfkuElCTEOsI62OhR0MDAnM2S
LlvrP+MIkQloDpBnjNbLASbE6yHImNAEnzqH5SBlpxbCoTo7KE6thgQNnxph9RUriPPQr1N+TstP
PHZvF9vKffW8C7ctqysy6XkCSTuyVwFl3A6JjGDWjHO9Zb3UdJ9Pi+zMeAXKl03WGDMUvh8A+x/H
zVz+fKFybsuN/Hv6yqKxeds/0vvL0ICNvcAqvEtTmmsT7v4nveb+P4rPNixYCoamMhKUzppv+AET
anckUA/f2tF3UCbCcnJnjnN4MmVWCCAHSGKF43yjn+sWCJePry3+aKlxnpOz3fy3AXXxFvL2pBrj
z/4wJhSmftihTsmEpV2cjv27htsI4R2D5HsMNXrEGMXnUV0e05Xl3jR4Cfapd6b7rVLn6W+870mA
L/3wt0qvB7lbYpZjG0q9J2x+opiYeOePSsBUgR6P2nE2jFIcvFJIdbhdqDugU8rlTuLW0bcbOaUt
hIpCythQDHvFGsiix+m7IOmtetNI7IoQ6iQbRm7JtZsZWxzH0Gi8wyCSNBccOU7sBzSSl2sHvyGq
4SYKzENuXjLgU21L2pJZIQeCBdxJj311mgR3jB9/SFpOh4dr4FzJwu9E8zmTkbDLv1YWjkaBaYYy
K0jzVZDl3D94kZRyi7qgShOP3TJhjxR26lsS1AcAfd0sziQzIPnx5LRdbsP6Eb91xss0YaRFw0p7
X4YKSSLacD+DH8yifLYxQcuGyP+T1r0IcdnXMJ+OMdijMbxRXIFpJxu3Yi/fIv238OgUCyL23Ndk
CdgWJt5tj8T5qGzBrn0EKDhlqcG/G5Obe170mjsBLw9/dyezinkHJIRI2UBLIP46xMHr5czRYJyv
tPpfgQewc50CvgYIPL2q5D0cQ+7lomBukHwlE0RJaPiZj5ll/xO6LmhQWykuBh5thuwxU/AloZxL
FEKixNtPg5YBcrOmWwpm4dstT/fKTsDDy/m9Yx86i4Q9DssEm4KGrMqdmGVujfRjaPPj3Xkx28x7
t/4EaQOivfuE/qaT+ih1ilEOxqDk+u2BgUDzYRa/RA0RadXMkrHJLRSjTWcUEHlmYkIPdgtibgPv
zW8NK8K87UWAP3WJyHWqguWNYcOK75i9LzYqyTPnaxtBJH6GQp0yxqD7am04Si9UIPDN+/Qxr2l6
xHjMwNV3DrIEEvi0fxEmTF6jNwRYiQLH/gm8C/QWmg79qN7KkQxzOtD4PVJ+LKIkPdU1Bd7AyFOd
IYyK3sgOwsT/UR68WRMQCbER1jXU4/GKTHTVWj/mB1UDnKcwsE3h8jS/kAtESSEXe9weBaW0B/Xq
xGOcqicvO2F6Z6tiXF/AulXZNcvSfvH3eUBtmT0ObFrlRdzSZQJknTyWEyBd2SQnpKhIDAA10sde
Ef5+5LFLyRnb5kS1I+hQQiFsLVm68hRX6Mo+dmmZUNhrRJDCk3BwOyedV46zVe8LFfP961GvuqHn
T58NCskSyZGDCQTufUGo35ycn7MFQyYlhKeMbHUOHqdRwfGcghx5pZxAy3cg9l5j6Oy3jbHPxx5I
I8vzvLTJZKnaCRuBn5nhhr1yHnDmAVEs1S/YFuHTb0OfVusHlegkzbSSkReAHjn4PGNxxLNBsAht
srNyANg9V2ulga6XVQEsTtMJmaH7iv4YcGMVA57BUFU0Ek5KXCWg5lCe/mxzo1cRvfOKadJ4dx8Z
QacE9oZPZ3ko9vRhMvuZYGtSoYpXm1NxivKywO8A65xAEfoOmeUZT9dpDNuiR7LWEgm6RaFtp+iS
EV+O0XvWab0y5EA2i5Az3QMx5HuEAiRMK2MUpVPhrgeuyIeL/sdXawMwuS+4BtprJ1sXQfiDPCtY
u3xgx1Uve+Oz8EQssuu9PxrGmfFuHLlKF+v7oceJDLJGznbRzXLAaK3B0MvhxdUF12k6mOY61eUw
tHIKpBOucgedoNuDbcg88RPP9OYQGrs1bEhbqtk9ng6RXMNi+KtRQhJX+xDgKEo7EarJfXK87597
L56+bJO3cVXdVT/Wf7wtkYQY4KBy8awpT2x9vDda7qb2klkxak7k0KDe4QPmRVt/kyadxO0V19h9
9KbMQF8gmJZuRhKXrg51Vjn82/kBMqNm4jA6anFHTIe29nPW0zo/TdbEAHgukC6IcPn/8IoAU1Vr
zllNZOpLCTsEyUvJvXJHMDU8Jp8hWvcCzNDBfmMHMEfBBwbpw5BbF6k1KNOUZNWFkXLA08Uw3lX/
ZHrIJsvYBwZHeifFR3O0TvQdDvBNmj1vNyLsOBwtZrRScOnBI7DSNWNVVC4ft98lszzHFfQR4i47
rjROggNdD4vS48K7XfXgP4ERoYBvYGOOqvRhxgvvJwKKiB8rsBLpePS09TjPhGR+LMBk8FH/Xz/k
7SjZI18dA/e/J+aZA1IaGSKanUWhccpbPZVJ1qgJoahzJQqxsnamP0is3SG1U/35vjIC0hubW7/1
PMEHKGCyjYawPFWTSryuABt1favwZtsM0Z0fHAw7gdaJo1cQOUVCUIAMOreB9tXthut4OruIz1i9
lk3Z9NUzZQb/ilgXWlR5qSAmkNffdur//KdHCTa5/cItN5Vok+UsQCReRCx9hrth9Ep+TCg/swxM
u9pFdr3K97qJAbrS+jnSGYJVajxbGutX6KreH9ZzdM27Zk5vrd+8am7LiEFfi+FmRwVzpAUb5kco
7D9KU2uSX7BxxPhnANRQ83UwC5GTLTXQ6fW1Q68N2Aj4VPaWq+4HpzQ0lLXeb46h5ERo/PMZZq6g
uMLlGOnoy5Vw3TU6WD8exqVY5EQLu9UnWvvPApsDJbObJz/yS/fD+sqI2b7e0YI2miYOtdpq2fJ8
nIWwXy6FIeCUYNA8zI6Grde/RXeFd3EAysgjdj8nEkDhatND7R04kmAmAVCKZr3pavC0l4J0BZut
asZxjiyMh1RtImu9PH5dMNe9Cd8vjeGsU6Pz9rLsV7WI44bDLrjomSdmXAOFfUeyR9fB5NXIqGhS
AM/AlxE8YKpB0wabJ0x+OkhJEPSGHoubB7KSn0G7a7p3wu5Yp3qkOUVMyygLX72EuRcD7zsNPfWQ
pM/VDbfJXz6T4Hxcn6z++xmiO4emzLDxw7F0IZpAgu/ySxpikBI8JgLna/vUJIb1VAGptO3LnXD9
/7Z23pcKb2HCc3rC1xQ+MZY29zUak7Z1rKJlngPjvylCvqHGjylECRao6BLCOWq9EP3NeroXmTzJ
qqQnsN+JH/rAvEbraara381xsEHpobNzSXFPpMip5MsmEyXeR7rh/FQVjKkKy/RX/1hQvR05uZkZ
DuF6ukS/XpDYosfjiG0ffu44t5Sdle+ZBSDI01dYokM46jJB1uSDU7IaGTTQQosLwUQLomwXhN0Y
0L3J4MqDAHnvIGB2pDRwnRKsim9HUfkZuhRd3bDYzfA4xBR0nl+duAhnB+6nuVTcDu8K8I3JY7jO
ED2fqVNvVwQqhvVnb73EbEyLgp8Ou1DD3j4574wYLhjbSWGsBm+dXk50oAsQ5rVNqG8wu3vARcTX
R19KRd3KYpNd/SkXy4Z2zRLeTH6jgrDMRh0AFlYL9LdYR+EuVM2FZavkjxC4JvR7Lr5rRvrrGN4z
SGfqhLbM5YmisJpdvD8DjnoK83y4m9ZX8i1xeQzz0n+s7VojOM8cVEBVVf6MqPPY9mwIUY+SXkRt
aOEUZbCj0ESafvv9N1VFAAPhshYW0EOCJ6ipkUAMibPjBfseOYOg7NlzblghVSDRrx5WUlpTuJM3
A3gXUqPG9ymRfjqU3yyknU3CAPUxcnoyI+8qpnV9OqqvMkTDn7zbrfefONdIoKZgs5RIbWuJNi+G
Yiq3dBtgy6zyNYmGI+ovRq1KXAzLu7U9ebzjRtC9cxHf5W4u/Q9+HOfhLeTCVSV5tmfVZMB29xFl
FLteuuerYZX2hZRzEtpz7EfvRdTC+9oV6VX69KRK/RidxjG7oPMvd9iJz3AG68BhhefYRAgygYC0
sciRpyGIizPtHaxdB6XSbPfvf77V6l4NkoK3bGMbXAzKPO0yzaPyg4WWuNnsMBubdG/TmarNuRGM
ZaW4WWUU7gYEgaOHznQgQ0lFok+HiIpnEirm7QZQlBq22ZcAmFhIW8W24qWZ/7279CV/Mi2n5R1y
y/aT6nRjGdcbxDH7Y2fmqjBd2naCCeW1Z2NK3fMNYNuGvzKg8Pk7ySKoZcj7/RGy4llcixaF4Ujm
f5wlwVKRYWyUGs7D1RXozQqKj+wdLUzDkK3nKAKR7vvrAZk2r4gdDSikgvfJSKpFSAQ9skkHu64o
+n85l35+SmNfc+YckOPTDDOlBvNkBfMmai1gqIMvpyZRXY6vJFd+Y6jlMy5hB1ryNEcF8g9jB9M4
ko5E2ymS0Xp+GZBVy6el7oml5lIJBIduxV8rpWNIRvG56mpF4j8gSktA0RpVbyBakSfXsVSJg3lo
8e695aNAQRgLAPewOMtK28df7ASr0C4ercps2CQNRsBjVbl1MA5vMX3sReaSaVShKTtKEtM0PgTA
IN/tF57vFI6BmWwzrYx1QfJlc870jzi4YS0LbnubplRSfpX2rLxHsrJq2LoohidyxAfVJgHhIYgU
1vSjOV++Yoh53ZX6qugn/s0eblWlYt49rh2TeEl/6vXLXCOs4OMCw0WNVzLgCsadq7+Vi88RswFg
392plecbV6w7qhQZEgKevUTo9/dpebkMmh1U7S/lJRl3CisCQ70hLKCaRh4zpI7HPA5VKi4G2IcQ
gz1+FztyXkZBvNNQFLQzyMOtc8C2iPTcDndv9w5JwzHcrs90b0ADBjr/tukxyvpi0v2QbnZLfWNp
1Ro3Wemlzrt8YJ6eYEEedQMnd1bCOr7iDHNzHoqfOfjc5Es380GHuG1lb/ESVgCirNVnXgk/2VOM
GQdMA++PQ0qQDIwn2pFyky6XotKSTHxRKO6IVNKB484Q1ry5W4QwEIpPy2QAPfcsdiDzs82HsQCJ
WH8WL5eEanzDct7cYvv1RqN4pqozutfy5CRtCuyHcmP3/yuGXNteebFnD4Fja2NMR5XG7NwbV5ni
jbcG98HlIPv8Ip4Dk1wmIzwPK7aqonfcQrsB8EM3felQkDGlxKZZ1HWPQ2EPii7NZ8LntK40ARD2
p2tiuAkhJEoz4B8cBTnXnKCdyN0EddveYff89IixMUw9ww4pURTiPN+BdrEN8T6Ur1YxEenbTMeO
yeqHETkYOXupox+KP/CxF48Qz4jq5qcmxTJWeUuj5jmfg0Uph/qkkbUWN7HegP3UITiiB/DvExA/
b6YeavAB2PmKrKQynUGPa76GANPbHc0k6BUtPKJka3G15JKnPa0EPOa6z9N2moawejkiTlvIp7qe
5xOWX7HJNE+F6cHquHWypgbWB//oQN2U95MdX0G+R28tNXX41+dLvNE5PFxH72t6WJk3RmZL07eA
Y6Pnn6dWW26yzPwnKLSAaSNwnmAPToEgYJhB6jOmX0cDboO29bU8Vnz1ED0Kbko0JUt8bX25VHht
bNZF8LDgZZULRjhVXGJUMHunVQcD68yeqh2rXDwlmQ/O6b6IT1SjX7bHioZfaJWrMvL/EvaRL9xL
O1jxj3DW83W+ijUAq3KMue6qQHE8JIupXuhx5Os5PHtaiEzh4sGIJzim5BDR1OYEF+DNku83f8f7
It/H4wbxalu1yNtyX2cV1ITTPELD+398JtKGHgqI9+MCB5sHn8WK/H8ZBhmrkgn71ek627YR+COJ
7yXF+ivyVoSW55RYDmVY35Ktnh9eMee2/bXkaRhK/3WWRbFfXeyDVilEYqUWV94/mVfGO2sBRE0g
L/EG3VHWlta2EyOtdsqkmVH4W00xXkUUzS6b9/G7SsZTPMkBAo5ZjCiYG7GmywaO4CiQt1a8TDlX
UnYMypdIQLRf6QmeSWBRZbx61o92bknczDIkClZ2RXOvO6EDAKagHnO99d6ICGK8udC8A7CAZArM
JXbQ7N3cn3yG9okfPOHnf8c4Evk7Howy02YpR72H0Xv5EdscmHZ0+vYt+c22mgx/d6gH+Vxe6NX6
kI0u/x3/UQeun0vZJsYyiUTdmlXRV69xKMGMI9rHy89+bDf0qqeH69QEMM3Vd6AkI6II1doUS5UL
d/HJJE9KiaH94gHt4ZnWUPawqeW64g9/t18mC9g/BVqYsPRhH9CQZ/FlRRhsyjd/W67pAob9ngoe
uJAfy36VVh3vkL5YgxY1wSelZf2+u7TmSk7QsxXm4LiVZ6qBmZ1tBNqi9XTUeT58XI7l9OBK1tRl
x55GNY9Xdz+688cB0lNQb4AZD0JKsT9yjuiBMhIWMQwQiTteM7RwX8/jIByr2ILBueRDelgKICt1
eexPInDE4t9AJq/YiDzUJdaWfL8wTvsJAevI4f9Ya2JDtoz4ez9PUF7lsxe9dubFWBu/nEDOHbdT
TLhwtApXo8K05M/L6DLUAbFdmVCbDjYqk3bKZ+vK8MLov1WglTkPcOTEZ7WoKDSBOPlSYnxfRkrg
dupm72GcY1DKGJ3+dta59qKCVUJlnTyM0xZpht7USLpiY78ng2CkEA5thNrw31hSLsg+t3+qebll
J2JPzxmwB5zQuZNfiWCZpmJ01wiQKEBs4D7tCE85FOSfEewh8192H0HbDNb07+qZkzCf86hIqhxD
E5qhLy8M+XmkINgFH7aXqSho5c8lNcG2CgAz3YmLPF9rNSeM2VW3gwkeVXmNLnjrK5nuFeJsQRlB
TGtRiE43y8c2AgRzpr3NymzmrHEsqcBk5WY+7wYxQwb4CXXR5k35su/Ht/oZSNvDq5KFou7j+Tyt
ouWIW9owru4n17KSJ+qhISIRMO62Pg8+KTTCFPrLe0KckIr85y1Kl/PQLXMHd6r8nzno1bJ7bF0g
gOHC7IUxy+oMW2ma1sCj309H2s8y75lXXuUqa4j/ylB4O7dOg5gHm4g9e1CwV1pouTQIURVC2tF1
mDIgmm0qFVyK/+lUiBtl9IWVJSh4qJqxtJKWNhKoQd3qmyVBSaWsfNZLBgvw8YI34dTbVUJt8Xsk
/FkGibVzljchSyGsh+He32g30k9FuqSjzuqRkxcQIKwYpzfvN9G1J7esSukTlwNM46TkHUq9GyiE
anU9zG1DgJa1Mol/vIXZTQuF1d1hU+9IdPqBDbzPmoUURAQD7TlOuehu6InXZmTngGe2h32A2p7u
Qw1u4r+SUH6ccKMg3szuyEeYL1OjwrtgoCk+vksfJa2R7VbJhJl02hzhoI3qJfqYqDe5IQayXWla
E2bI4SdzTD46dCaxRLrbAbGS3sjb+L+p0nZG7njF6UVc4MW0OhpVCgjK/12uqirpwU5JDh3R3fku
W1hyj6wKqQ0uYlBM+sKJy4USLMnTqELd9czddFMhs7Sg1Ox9AiM9TuzCxH/B+DqiNSAkE61/LQ22
wfv7GpnMHZDTZFeDMItsgZnrX54zoeMvkoUiFFs9Q66ZsV//K6OLdT+reH1Yd8P3h6/Ccl+4DF5Z
oz5jOxqMhowQEbvT4jM4OzTAdva5J5t3TJMBzTK4gPPluXvWy2LBi2a3ygazoXyuEzdjm1ALpAa7
M8HPpj/FTA4goaM63sETwzHKITxG6FKo6QjHn06NlUE6sbMsyg5TkdK9diltP8in6BRL01qek8YS
VrT4m9GCrFaCPosFmC2q1a202Qn1CRStOfzR1gX2jUQCKkv87lDVdYNXx/m3fmbkHgE3wQp3mrz1
Bmp5pAcnekE17AvrF6fSXl6x1D7TtI/peci/b7xHMibUnI+/nuHmJbjpDm0yNQEls0bbkz8aizWQ
41plCNLdbfmFtJbUKNOt+Uai23r15zIBdsN887C57pK7ti7nI7e9RFgBBvk3wzqGQxeMFSVyk+4L
r9Zrcuykg0ZlSy+3x3dhjSjiLSsL0B5Ho4JIYFHSd9MS8znPIvMVr6/+dz5g2/aBEqDNtfKYwWxo
genLixxIqPYDB6i96Zw8bTitAochc1x8zvu/V4+5g3cHjqCwnuCdeyhRzpkHxWmZfhqdsye12SeL
QZiIVYvZ0zBhZLCCNh+quEqxGkS5lMYSj8r+NhqK6HbXCHh+ZH6j+3WeBZCmnRexYRLb1k8FbY4S
C6/3uwbHrzq7DmG5m8KZ8+seJ5smsLBHspE1uHQaAGfLK38MbU5tLjuSsrNeXbQe+Mu1499hvIAr
PZb7XBlIz9M+rLVHNa19PS8J/H7dbvVSHrpDMFEf3HQoqVyeHR5Mt33F0U0IOpFZYAea/FoVwX5S
+r7zP+jMmUN8YnIdvlT1OXvHcYShBp/mGZieHRfqPMkawNH09ihcIMM4sL4Pyqy2qWNUrp33vSCx
fpRtsK5/Dzzp6R9G7qPf5xySzjIRGa4ipNUmffGy9rb9xQJ3JTcN6t32sYE0HapSzZXTUzv1Tfh/
20EQ2EfLr8IX2oJbY2g9Phq63yAtX0hv08JISR/yLB3yvuBQwdHq66mE6jMBKwIEfTtVClz3tudg
+9KcSIaZZ/7+dVSD5wpt+jc9wNte3CnsOClPoP1B1ZniublCWAywpya+pZKSSjRzEAWszzFb7DD3
V+L/Jh8aXIxSgMokmb2N543eERrr9mQz+YFNqr865SzLreG38YoAyoUPPfh4Ky0vWmfHo6cqv1hp
CUjh++lrmMNqTdmRPzstt2TtA7A3E/9+g8XbTMPlBwI3+00JhVRchouEOZJmd5/ARQWNbVBHNLlY
zAA/ht/R0pg8zA59f0lbinfVGlc10xXghzDA05juBWmWbkfWZ+0pcaUl/hRgSYhH+KGCWhScpXpb
6VC9/xEV5zoqxcC5+dHOpf0D5wdTh0mIp3NUluM7L3MKnOlRZNmGxbxj0CigXgLt5aWrZxY/3Rus
Sz4esCD73J3/Hrm6ruRMK9EjGFQp9E9ZFcAgkhrKuCYZV5surkE+1N9ppbumkSEt6N8TNjL3pxE6
6hTZQGMUJ1oV+juy6HMX43yW2tvhYXTMPdvUAMS9kN2Ci1Q5UUjkORN6MuSV/4hnXWSRAPbbAsUS
wjeeuNoA2FiQQ/Xp6NNSBaQ4lPUeFt8bJPpufL1P4rd+Dcv2C99/jMc2P7c1puvCR3AB1NsXRNbI
aGWWR/CxTiWnt1P37UdsJu5pSAUu86grcTKHYjc/miWCah+qGtYjVK8b1kpPiKIN7K9PffID6xRO
Ib2z3BSoTYa6lC1n15Gryw11X25xH9297Gz2BJ+Q1z7xGo6r6UjjCb+muwwwfxOq9gGFth3cytIU
hsffy7bxglTaTt24EqJRkJ4OsQsXwx7dCW8QIYlJyqiGzu0oDin1nBwP0bHm/6Zzpu6tgQ8q3/eK
fCdQaquTMipU5rhmwSutNYnmKKVdb9+2cSN/TmDfckBlnbtPCcdk6KHwV5F5fSPnRiOtshX01t9O
t0W1NvrS1YtUxOeVRrNcQx9OqS5wMR3iASN2FFVLGHVhjUGBUCkMurE+ZaOrbC4EWQ8mkNbE9ZAx
EveweV5A48lt3RgQAB9VHU8ZKskLhAsfGFQJZR703YnAzZ4C4YODC22PweMzZElG+H8n7BLTNGTg
M/wDaG1zS3kkWf12k4kylydIaML7/EuTVlJVKkjnYvpdfK89kJ+jKu51QqavoxliqoAXIaZArKxd
E8dWKy8EWzP2LulV1FOopUVMwVPNbQZrppp9dp2678lHP/CUCepMCJLkTbjfs4m2RYGleeWbbO/v
B4W158NrUhZa4orPVKyvK8E4Aj9Gt3ZSsywDo//KUJfW/Npv3GXk4+SzTFkVQU1wr5JCADhwti/V
lZP/lhnPCutg/buZlk+iN3rwZIGU1GJ8xpopcvzidZg8QQ4Rf4bwlCJzkbNDkItc6fnarwcSjAFq
wZJK5kYQoZVrMyCx+8WHLBMdFe2dqMKZE4OrM/Ui/ufhwCUH7VpOskbRtKM+eUqGESogl6K2IorG
QGsoZ9iiuvgVYukfSpT9HPSDS8cVp3yiDV/yn9BlH1stKgemzmkeVJVen83s+DuLWK8NFIPw791e
BNyRHubfATa1x3e7WajuLVRgbSRGDjS3MpMguO0a9FG7OWolAsBz2PtxPtWXDE7S0IN3I0MHGzfV
cl3zIvqJ10QwFXSx57s+bXnevGNfEwMvQxA3JIsT9GUkF+KYot9fz6wiEp5eyD3s+B8Lc9ec8Cv2
+QwKgRj/qNzXbxjFOFbei74MHsPgccFhU2UVacC9b4Nti1iF/Tbe+JJWjm23Fwj9FlOzYolkkv2n
bmxn68C+GwI9qFqpCrfZ2XEdqpSHxDmr057fW7ErY8sEO10ObiiZvoSw7tW0TOED2OIDAYzz2+wq
e8yG1uFf9wVeG0hPOEy/jfPQDFq+3eTL+xze12Nyyb00iDGnRH1NrpdOy9D8O2GpHPmUx8HsO7y8
rrXYSson+m/M5DmPInvGOUkXIF9ffRyO+TOfB18pQoACOvEDYU32aK2KzgQweH0u1QesIg9ADViX
SP/+ZqKMtMJhU1b6Px84zGp/C9Q5yonjekB7ccHmbE0fBDArSiKsJEZWoS9LF2AoFuGbLxywcAhf
a51l5shgYc8X6nmaU4vA+33jAaa5GdU+0zTwkNeLf4CJcMP6oCBiLmvE0IPeBhrdXfyGrWq7JUF+
xhkvfQ/wq3G4gwZAzX7iHrojhBSH22qG37zTdvvnotSZCWAssxhfn68yEGVS4OVjiXO2shUqDIlf
Oafefn5LiAjENqksH61pvrTEaEWoyEffRA3gM+8vM8Fq1YTZA8nhzrOE3JdlEvUpUz+G7qSJdv4e
qHA2e4PcOMzeOBp7FrDUhI2J2sYiAV42KrTpnSyvaQaXaEpRzM9ITXLZYC+GqPM5a9FVdnPy1PWl
6TNkFRrRldQOjNrFF8KIbcy0NFVe9W4cXb7Pm+X6I8nvW5jYFV/ttnUqgFEMCpBzZTA5FkLEBTnO
VAHyMjPfzV37GDdJBW0HBxCL3YUz+tt+4pMqGJqs2Qsh85G/RyZKPpEzT/hGKtKOzmoGdTvHHyQo
RMevjvM+GjMWq2PpX/kZm582Eq44CEbZ3KwKbyIOGLF6PhMEo+LtxOehFHLVUmLRFA5W4GIiTOrS
t4/nT8uUbqy5wGKPrN+s126xi0h2Axn7bpiEOISqcRZ2VIKt75zSmTtbfl4tcgVPFZIlGosXCXoa
S7o4vtb0e4MoUhQWkpmkNCFW7bOJAUSd5XmxMq4Pai7qp35Zw7BvEux/vGh2xNcoBlfD560r/Fji
BSaEyGb1xQBmsIcWvWHgx5qW3IzVvGQAvdtI1tIO9AN1vmjuS0SOgPStVxesgwbXH18OdFM5huDx
a7LN0Oan4WLSC0Hg6oiyDKRLwntUOTnr7dwvmluElMd3tZ+v/684auhZnGJQ/saMuJRisHEGxyo1
Rf1sJMGItynw2+Dc3f+5Jc4FM1SXQj6nvN6gxbR7UkdQU3x/JsTWEq6U+ch64HCBb8KLzGT9HaaB
HFZ94NtBXY9tfawyXjVFTU3qDuD+c7CC2nGhEeW0ldzXr/QNm3JDdcHCVjVQKtQ3k9HZIuuaU8t+
tAnr2iSIum/z2TDXO0OtprVZR/62kJfQslXWRTmZFfcEonu3jjnDFAdufCx9q3TRhzbGLplIN175
DvR5daNVl9kKaQzXTBa6G0cbtkY2Z5dCNd5H4ja//vIuYJxmV4VSinQ+oi/8Jr4EF8ny9PD3V9aK
rrL8vtmt5RKejGdzq/1ICQTgKxWXMfTA2ej0s5i8Ypm9czy+BDL1yGeYlQONGMVm/VtciyyOEevq
nX9KlCS2PUJ455fV20UhhwskkD32mgmzif6Rjo1Wfgw2stBtFYYl9cnrmlS6zFzz0XXS2VFdecb7
OA1gOFdlT0LNuWfHxXwkNlw2nACVSpta1tRkLJUl9M7SZNyzMUnZ8DnSokDMz/D9CP9Bxc0cYyI3
8cmfd7Ln7vXehWX/Ub5EjsFGjay6N9BPck9jpmesXJKb2zYsWEDWFG9kHFrs0ppT4qSjJh6CSIYx
cg/Le1MQslPE3a7TzG5GWkrCvH0OYAFWtJd74vXZ2zO835PwZtGpSNY78f9ynUx/aSfHbOewMUpP
5boJfnFmJyayO+W/VWinf9DsXunYCm88ZwOQA8AIl1pj4CvQTCQVCe/EFaFD74p7/C/zVoeRuLVm
+UGQsi4mbPlepuQMdxao/6S+cMT7bbEPc4WP6eVtqy7sIEuT5FruNcYMGQrFoHBg5oZdpcuy43bg
M2q1GSVqwwL/+VJWzTSHW8a6A2zAot54RTjIaF0saO6ZkAOG1SiRTPFo5lMmx1PCZHU9H8mxbkSx
YBNBzqSwIRd7bxqYOOtBN0l0QbLJiycrN/TlRuYoJUu+qzcNAeGxCpsphhaZ73co4df9voQKn4Fe
4oQZtmDu41b4OeesZi6mJz5dOBvL0aDnU4KwzmHj1TTJ2h3+X7hSqTwWKbfIugoPSYstMPfcQ8u8
v28oEpfqGBka5fUSO86iMyAlW99hgOJQdmX2iTX10JQyXrPSWISigESmdgAfqPsiqw9KQMd8p+Ax
u+Ke65BbYQFo7ZfaO0US4Qitzn7n3MSGVjv33lZlMg87y3jx/8tlSKhU3qh6DQOcpxoWYZWnNMsF
k0Cg3HjI2BfOzFXyQQAzCCJUm/juo2n/oGoD22H+Ig04Zn5yBCW+DY218eFkvwPezXM2d/8P3j6P
7pMbvaQi+zfxpaLluu4oXinkbtSofWhyG6Nld6hrNCgzfDy6fhzOMTvaZ4lYRM+x4LIWkLs7lsbR
fp8hp1lSD9hi+UmLEAqLcie0gkk0nPqlaqjW3z3n7vRUOhoOZtQKqBdzk292QuTp7KCQKpyvYSJC
AygbEJwVUB7yFZOAOYIbJgDoS7NvzcVHziqsMziZ7zkFE66v2QgfDKuwTBovCyN6rxlXVMIYrhWs
op60wXtv1+CCt8ej0jxfM8S5Dh+kjq+9ZE9HG58olaUz1fExyOrVocHySaMf/6AblAr6sBkpYK7j
T9kMohL0GG1PdLbPwZQ985+FBY+iDb7H5OtA8izFOWW2SK1FMZQr/kWo9lVJx2lVi+3vsAl+BTuC
i25wOVzpgxidBTeEbrLR7UIg8YKDWaM1A9eYBg9Oikt/R1MQYEUO3z3l+Vw0fk0sOQu9xc7F2xRa
PEJWwIeSLtwvaH63OwHCsB1YwyJ3JA4NKTvy3AZ+cPUbucP+rO1QHWo30SrQfpEHwI9IBqWVbCfb
ZyyP/Au3XyGDo7NcfxR7noKTtB5zYuO9x2dAeLneAjCl6cZq1dj3AKOIO8+UTnlg2tVu+BK6eW9N
dw83Mdwk9D/4faXOl0ZRsb7UrnsByHq8SXVv08FjRik8RHcSokH/M8UircWH2PbUNCgcgvshD+9Z
3+SOwdPqXLoSqjC+u2KLdqCmIKz/b2E3pgcxiATIiwGVb5AsP99HVl23SgrVNlkdgMnHpj04lx4Q
+wh6v54Rrg2RYClCrIP4+R7av3cLSybNe5ilCOiXZNmoK94+m3Mq8Zb6SDHWEE4uA6WInwexc4RC
3PWNYetqRcDKSlxnvNnfo7ws8JITSs3ydffTZ5kGh17NTC4W7RCKDa+Ie+rsZvP0msUVbP0sqs5d
YA01sgXdWA7V4LhOL+G76kwnIgMPQbftCX4PxHJCR3zRf0caCenrCIebCKBtSWHig4QCavjEXWYW
HekUmCdI5E5LfCPyVYx2IOx77gGmAIdWrNNEZkAZ7bo3x9oZTgD5kDhXLGTke2XDOz+c9KAtq71L
jQMNh7jzgFnLWsXEdYee6fpY2w2pyWLS4x9OVqmX6jIOZnXflrxz4BYdcL7k+a+jwyZ8RgEsct6Z
YTQm3jdJRSWQE4ZU0itVB+tVG6N49wrH2R+bxJW7cHtwgQ70Kfh3njMv46ZHgb/PWylP+mBVfoBq
6WBU4Xb1T5y4J+YVbMvbSfv4WVGIUXusuw39/hUreZcDZKUEhxoEfX6FDAymAQ8F3ahzNUwq1wJ4
D6tjTdZw3B0f3Kc+d6wtPnaBAQygPpVHmaBKgdSmAd8VrHYXBQJUFkP/zgVlFSX+pK0qckU3JdgV
A2Mgg/RWir6AnxMKh7HsS+wo8/wY2LDjPw5v1Iep+HAPu0VVuQz+Qmo0MDqWngQrxTaWKESdbsok
obRQzhPpn+XMUMYlxUfTuCsA+mYcEG4ozFSABq6xKf+f2j9dgLCcjKShs5ay5Lr7ntqP/NRIvOii
OJbUm1fZM07hthL+GNcc9JUAJCEMjHSQh7MoOBo0MFQ71w8ZxtiRIoeIgZXgo7es/aZsb7mbryUc
mtH6jQMRTr4h0F3FlbSqpfXHs2NZlO5V4pk2aGl65V6cySI7qyov7U43A/KMlCPGGrP2J2GtrKH+
S2QUZ6bZZs0mbE2FBslUKBNkkWT2oIUt3YkB1jLajCjGM6oiUeiGayuTQJOoDLFHBtH6tDTlWRft
FKw4TSTtio6UnWr0xRrhn2QCuvSeq4KY4XyN/ccJkaUwAB0i9OzgXE+rWm/FFwhfGm1MhmUxFtEd
ePXDQvfEZQboVzcm5M7kY1RY9km+Th1nsv70mIcASLoCy+Sd8g48A0ORF3ADzbdzpAglT2XKLjgQ
WpZvhygzHfMQqrS1Y5uxbT8I3P3MzfpUKytVNb1+KAiAKNolPTF2OKjCS0EcaUeIdmvOf+pyn1vc
1+R4uTXRVY03bwFM9AlZ76Dl6K+7Oj3V6DqU3FSzY7zzQSXSN/mk9voqkXA4ZYEUxtapL9KaVmaC
LteK4dm41L/jbiKeHlsTka1o1Hg7WwaQaktzgYl0fMHKa7R+4yIKSJDBHKmsluZXiODrAMhlpWC5
Og1WMQagJLHlkMmbzHTrK9xCm3ZrsM5PtyiaRQu8a2OK8Z6FBBkSKPztowpL+bOA6fOKmbH5TzJ0
2bfiLlqK0czI68cldiUKoE16k+6IvPf+e/1lsIyxJh6oZzg/zCG7Q0PIuisccvTi2PUGk96Gf35w
5CUB46JPNRmDfHjcT4Hv0yCHgmQnP56x+IPYFSjd4axH96Dr/dAHpT20YzO6m/HnORa8u3sDOw4v
6/A+b8dblWGuWC/ukqNLaas2w8CD5+0mNDKorrehRYjn2Fp53UiILZ6L7Bgwqv7XOU1xZVf6wa1q
uBdsEG2Z8Oi25c3PAbcxT9Podc2VMtYPUAquA/kM+pdMaJOM5+ehStNhpZjvF++hKQgRHxRGQ/oD
qxDVFO4PNX18Psw4QGwwH8lnoZJS/GyZaAiGMEkOilwMvH23M6v82/u3NtQgeaA1wxr0lyElyK18
VcRchF2wjW06GEptLgNz0SMF+I4KcFeRQx1XGGVbam++ib+YHGc+ho9QapqZ23QnwW825nRf037F
jYOhKKYrIgvhZsBIHJaVORhApRydwhbHfHSKrFuTW/U9YiFw95wqcHvT5U0jMtSxMfXWfmQNreqD
XzHH55R0OLUJKbDmjOZ2nxpw4PtNI1a3olZB8EmPxiJnwJrDH7m1Gu5txAp2i3JiavmRna2r8cu7
FRwRIC8HOrZJSFx44YK94a+dSWdlr3ZzKU0k3+Y9o1q9n4Tc54AWuqlxPSLLMpCF2eLt9ZkmastA
W44XaXbr7E8Ki0UBdMb6ZEjBN7fe4rYyvcKNFyDSm3twSkkeuSsKjOkhx+uZEUmLULz4tJjUAIcx
BRl0cmBuq13tU8VKh7JR8PtkUm5UexufJwC+kSZTwXZ8wtdFyvwNi6BNb6/UiCBJWfpA9aRxGUGx
ECLn7Mqazkn30nOomPNvwkHTbi+t5NPgYca4fqxiHQfVV2htp6x1o8aHASje1mtUG9D9HJ29uwrG
OCDnB4N+DZbiPAVem/D/+9jG5zBEQTK0VTDSO8siCweF792i02/44fT5QyW2HUjLcwaRYXhdWGWY
t3Okr47gXIHBWEyI1zdDEHt4wAIIgi03iQEuQ0kBdXFSpFyOklOIl7nv6WpuFu7w+v2N7aEhfaEm
9mQHIA54nhw/t24mdAwIdCAb5xEAWg1zd3fTzjsWSDcm+TxChokefQQ4XL6Nhr5iYHTPClO5da9S
xhP9RoPjc7UCe3tJZ/rej1hiHplSsjWJ50XPF0od+CvEruNxBeZrnDqAJnOoXhhma1Fi+IYO7GKc
9Aqx0suO7xLKbaKiETuNRNDvvuVvNdD7FmJEewEyVL74oP43eZcLigWZDUag8btKh2eU/F6aVRH6
X0OqYmUOZbeaFfnxXZefTaoX7lXcI1Mwk0RWoCuNSxR2KMXTZVUYpslyO6KbAUf17BI37uVfWyRx
IMZz+nUXKPwn9b6nz0zyixfhUqAlZjfXLKDyGzMeok1TkReeUmFTw2amFc/vfp4jGckOMP3gz1Gz
Yp3nTuBmKZ82lWBDYbHi9FVpRgO0/aqXNrdjSD5QSHQ7RTBGpakpSPd2DyW2B1XBoOCRVbLraN6V
bN7U8L/UAwL3Jt9533Q0eHfFQJgrFhiLUjTyWydwM2gXRTOIEPN5YrtTZ8KcAFMCxs1CRCSZHKiB
kzalDzyGODzqbLN4uWgOBQ7pfpKF4tliiSQ2UCwYnGCE05jTZlWqtQnbSfaIdvoLZ9j/WDHwgfsR
RXV/XoaFNhI60aPjF5nMZqWupvtLzID5RVTmxt1iheb4vf7d/nkYDek0oQGXyKVkgtL0mLDO+kCX
32z4GAx4DVATjszEiFRB/c+wcUbb2FO8fD+YbZOEBpRRgz+hizJuCSN9LvTwfcaPhd/JRXD45Tb6
n+t7vFKfVklQC1xxGRV8/5VA0OkJ1kQhBbIWYpX2XChR4Bm5LgkVPhay207XT/FIgg/tm/09iqBX
J9bceNKf56XccaKKGNeK61wK+PCc83K3R8vpPQubt1jRjZXaFUKJiQUj8JleFhkdWl2D/lSC0K4G
iYb2ArCn0w7RvnngLmyz8wm7RC+GBhFPQrcn8nN+kisuEEq+emTKaO0I1Wmh4qBFh5bCPh/xfDF9
+9Ot3ihG+7BtFiwk+ZiWwNtczBnhM1TquWBDYJPpIj1anYDErEVr5s2DXXf2b50j6iIp0MUawOID
b+I+64fMyimrpDZD7Ph0mcfaJKu4uTg4KfIsrEsQAuo2ssAmYcG97ef5ZjjP59mum4mDPf9h1mu0
8Hluivpcmkmt0340s8RSKLttHUvlI/77wp1TOSy8MtEPEVjOFEXmw70zZAvrsiT3u19x/DnlUgzy
X+hW2CLyoLl0Blj26FQdt30Z23/R7BzbAF840++uid3qjsQZlvabc1cNJRRZNQ/2rnJ0AzgZYI3g
aE+m4B91GU2ML+RvZ47IPwmEHXNZgvClG58s+pr9Mp6WsbUHeqglg1DlJskCJnhGDsU8I4uS+JzH
OVKh3svpOkCel2S8ofZsv+BByvezPC1IJIyjw/17Ak/vTUWhzo4QFBxlLvZH9ZS3SixXyWlPaqPl
1QecnAdPTLbG88DVYodsmC43eaqWAf0oEa7oNovm2ZBkD7Ej1Jri/zzjU8VegA8UQ4r85TkBIG6J
k0x5uSiTdPrZ/Goz0paGAA0Zm2HrHOL4BEQCGUr3EBek3ob/pmBG9k2LbGr+FiUzAvRigzufGogu
rjQEkX3x1ko6XU5uNOtdswgl/dTWPv6WhkHjldBbhEVi6rkhiYkHrZ/NEKjc6sLlvEx8IzXeAf3S
nec2iUvDtm2o6WT9SSekClkDLV3BHRm9CpAfIruJsY8N3tgM4LGwzAQuQGfW3fa5xD8M3CrR5n5n
t+O7107oEGiu3JOqmwhYHBNzYT+Q3+CZp5pBpyV2d4omlVyvUc4PbEg7JZDzAK9GjWzpdoMfIOVK
oQAJ4mwCG5djsKVGoZsLSjmRCNZO41b6wGelSzERGYAye8KmKT2S5/NSpu8nO1UE8/wu9y883B36
Jw9F8XmIXRbA+VWy5swvPcGNEVTmtAKjSfO3Kfcey6j3WFgnPgO8qywfBCN/dj/6lBiWp3G4RMrL
/p/daDmEdMpHpeG9+cTxv4A0jkSCS2ejQqBZtNuWEKtlI1c+cAZ871rKAoYosUuf1YoMRvt7kiEE
ZdWDnKr2olAn6uan8K+aZ36tGQhPNzoyKs8sZttwlR6NaQoM2lZvx8YaS50WwR0yIo3yx+bfQ3uc
Vme8qsnxykDhzqtxX+dVi5kxcBguXUhKiN5G9gDGijnzRMh7LNz7xz4xEo7VGIqpQTjTtZVNXHUM
KDCKUCaUrpQ4dbHnlMAmatC0qAjIuh3CUjSaaxQ/VJG2wzfNQTydYzvOT6ONvXluAOUS1qtSA0oS
k3OqHyp+bGui68A578iq8O52gMkAzkXoCcvTnAZfM9A7B0k4XQ4F4LsGKgfu5KompzoDMmF+uHM9
ENocWfzhmeEkiOjvHOhuSyPgaPa/5Knf9+J/xUHvkla8OXrT4d+LCJAxq+y8CtMLZZbNYHfCVunp
d/TAIxD8DaV33JDmD77jIuN3x5S6D9v3nIIDmxl9VCfK9yx+3firVgjfYgKZIzNbW1mnvDP/KQWL
0nj469L1axE712S737Gpe9EBQb5S1X9Smc5TZJYMzZYr56j1kAXHZJCSIuORQL3kFULXMAhqj5Y/
CEjiAiqfu7g32vEH3akeuQ9AZlrJVom+McwmYQI1aDhVsTfi7jy1oNLcSDvVaiX024eG4f3bo7I+
a5Wr4Rt7cjovHxbKAfb3qmZyO4FWf0mAGSi3Xut4W/UGqPqDDuTF0VKA24n84npYXeouHAZYYHiQ
dCJOT5SesbG02foj+z0kNOYEk0wcoR/Ph1lSTKBr5vpapxv02/FhsId2YHhYk9EM0FVjtuVtlKTK
1+as1l2FfeDKl2zvy5WB1bk7iqi/mK3S7YheShSFAZVXOT0Bz1kc7d967U4zHtWNy+OG3d4ek5Ss
n55DT4vU8ulhHmY01uyVrDZdYOI59AYYS5Q2qkHVa6uneiUefHna/NDx+BBMISicM45AsaDJQ2fo
T+zWCpJEt7mMqUkwH9h5BUsHMlgP3p8Rn05vYIZ2mbwIa6C2L0rijNa1QXqphlE2kUNQyjZ8gAvs
4D/VHr/5g54A/TAvvYvOMiLhaUsjQHSWJAJgLtkJO2tjvKnkhbyZ1N4tcmTGEou4fkouqj/XFoNc
Pu3veBuCKf0amsz53bElFgXDWHgzKoRGJhSROfaXB7vXKyCpYyhyOeVu+0Pz2C19hAoL8QbZFpeq
jg+SYyRaLemno6PAFjV743bJ1hTpn9jRTqfYtt/qQ8JfLHTbnSbfiUwK9FUlzjqvV4WRcoOfu/ZF
J0EN1EX4uIFzVMyRpAixyNoqVXiKaqDwmMqJKLI+lFJueCiZsvjTv6Nq1OGQJMsrtMbP5FjGrOKX
V3YP0ya5+2TJE3AofxgUeLd31DZuGPnKNUmZOb4hZasgMG7gs57wx/sgS4LV6u2kXD9GmqfPUIzm
t+Y69jWf9ZMmX4u0WmZiK/BpcBIp/igPSx8iVBpI+kZD7wSB0W7sh8fsLpWudPrxXENbourdRywy
xIH9/hIzDhbwHXUvOLW5WEWFiA3wWZGDXJEPjKWXJeuNdMUhRYB2nk2Q+wFiX0p8NL3ki91lhUFJ
Y2kZZ7mzfsiog5isXRwqEBs0T95sGNvMBr//ot6z3gfmWIIcGvuC/So+/gs8201xwSFhItxECT6T
XFMt7KGjjkLjGfuI54DMYQZY/pAkXen8jBH3mygBaNe0IWFYYYjubSk4HW2pXa+hzfszx0Eu3KRv
WbBKdS4AKqyy8b0FoNr+SVQJ9iL/YK6RgBhEoCpbVU5MwxORT8s5yPZ57ogFsIEEAeanjX/lpeLa
rIo07aS0+CF3bijEg/zA0xKB9INeqCQMoVPw4cSAaPEh2r8zWhu0jlIjh4jaQfoghf0FI/5YraGv
C7uWWSIgik4/Bco4T89HcNYX9fKpBcmdym+Y/AanxexkV7wWPyRBEipnKrOf0+Ym9OT/ZH/5ZjRH
vm9M/GGUBD7duGzul7k61cjfkMS4S/CH1akfX5nPDCAQeOWpfmXNxwIsQ+hXL52H5r/abVLhG0Px
LMX+6iajy/tzCmJgZ1aYmGWHg3pHU8wg3ulFu7tsLHaKYBJs0mZGtyEhGWRXsY0FWlVAX1YnX17Z
zM2W2ajf6fQxShkyBRspqL4HaQrUrwLnVOmf02uSsid6SvGzCzZ/KygPWLJCvXaiWeXZ9Ci5IwdB
8dA1cK6eKEB5JPKdS5NaY8IBQQvGEMDFV/0zn5oJ/zzk/fNfuB5mNGT58/6hskm0XS0O8hAlG9Gj
BWhPFf7OWPVo9an3WWBx6LTNaJXA+62HiHUYK3suD6bYum97ylumdnPFkMg4ntV7T08BFPhCyyc0
TEKq4e89NwtyxMGXhSHmkICnh+XeLoSW7B2Vc33g4Ebp+DhLvYyK8rq1TMno7P12VunY5+x50QeQ
18uEpKTLdjPdFAaLgrGt8Y5nm7cPz2qHECRDSaXQHtohDDkQvjO9+WPsWttHkXNNNJlaBlxaJT2L
89Oq1QKjL+j1+vlnRmkAHQy5xolzZoHl9J6ZbN45a7J7duQFfIDU1pg6ArYepm0V4HtbQxt0dNoi
hpEgbhOwVpQc8pwHM4SWVAIkhEwRrKq++IR82p29ZqSxJPjRIhb8VJQ3m7BwC+paEcqauhBdS/oP
HVsO1Bp2uBsWmVW8Hp/JYNQ+XGevkDA+d340mNf++0kNF8+Zv8lLTMtqQ87ovCAJcwSfnsXd+ptZ
qygsWH8YO8AXhtOahMNnOyHmDVl5KCBBycJQ2v4YtuV/Zs0ItRvGcq2hOxJ0Y5/mbzQs49jsM/1Y
TvoyQ/jApHqbRwTplf2OQiN7zfPzIPn3/w19Nr9vFYIvqUDykGdcaxeK0ZxVW0jRKUgNgi0B4HBo
Ljqu+S5YFwDOLYRNniD4x65qY8piGisIigfRtmAEgBtgBXkWIflxJ0ERc2EroYB84IAPCsgy89oz
rENpCayyKUJ61hdxN7YmCiQRwlrVDQ+cQU3SnHthmqagkO9cO1L2lWt/UBcn89hgvZEirYSYPrOo
ddU3WVc2m/mReJpjScK5Skoo9B6nQcGp4wCeYBwv23HrwduzlU2BZ+bbWlLGl5BXigsoUOCaGugJ
EOp+6UCZAQM8trmTg5hGYA8mVUFO8ciNbegTmBSR1bzjxDNimErk4D4lG1QWBylXC5K5NgIAIr6w
cXrgnDwIs7XYESGROywCPmDgiuZdjIcGRJqS3y5LiQlR5gMJFYp7GyCFtRz8FCSX2nJsctNf3kLC
RCaWguFR/0/sqtc5UBN0pzQFSrGS5yMmd4jCpjWCtIdz+eaSBMkGwLPkbQkJciDNaDwUrXzLDFPu
PCP0gFV4z8vyz89ZWTAk4xS+aGC0tHh2tbSUmC8fvazqmPnTu/bveBrzD21CNS25j2OglOLqtOiy
cqpuMuU7uYmyl0+WpTZ0FNwON9tJWWLd5PIewkKjq+Tq13U1Ei/DzrXvs/ireYPi9zJUZ+uOXI/8
Elh6LjqX5KlxD0fjeg0fRROEI99xN5ea8z5ZpbOVm38o9ytqHw4Tbg/j7VqaPtmV+iM9PtoZQkJ1
Ywc16KuvVPf2XyT2szrsMqwf1rSFF5MhNTsVsBbgVjjGNnPWELarSG0GLCrHFQWvw00QBxpS5nHJ
UNmWKV7jLli7DgqMAHQkVMCgjFh3FkJu0yWHxDbq8TfjwInTOp5WT3kXS7o96QMDpmGiKM55xJo1
fG8/lYL/s+CfGZ0T9nj3xEzbnNLOBmd4z7fE+Vx6EoT6afe+3kC/wWv+bDHb7XEleaFtmoxo+d9O
whR3wSjsE3ajUU3Tuqtvh12Bx1xoDTBjbMW/tfvw7GczxjHnGeYh8LwKjIueQl8yHK6a1NZ2qppr
ib9QdgRdCtiDjsZA6GHP57GkB3VJAjVhi4M41kCILXCrDJrFpyAKfAmF6Ur58eFvN7Uu/NurVzVr
mMQv8yz39vEUB1jpKUzrGqButgrM2+1TLlLKz5F1BbWbZ1+wg3+vZz4Rm0ofgrnhpGQotx/JoMJB
PZnbytx2nCxKFUrj1sGNzqL0mZ2H7OD6RVeG4bO5cg4muB9O5k8svyEkRiJdy5pAMGYgsb2uXmSX
w9BRXTHqnfXKsRimZfERlczaH8NYg1oRF2s2etUEcrWGQz/b2/+J9kapk6CDMOudP2gL8Ys/yeTI
YEVZ1sf1KFWZJgfAXDKu/0huxUwFn4IZ7t6LwwTpZI9b6tR4QdwI9Y/1jWc6LUjwQVX70DxGI2Mj
uw+LjNfNVDc/2+wcnZojqJDdubAMhZuwBz7aVSEiF46HEfyUdKH6ab3zH5wC1jmc86TsjSKfoonT
qrOkDTn2zdTLRhBg8Ew30VKFcGn2UHw1fccu6+XmwuFkfKUyVxk+c6s9tsBlYsSWz8ObUgv1ZU7v
h9Sdy4EWtydpaEQBhwcPtW3IUMQhuA2SELdTVo+0dU7HtECPVHcrKqKSrzgHmeaG8XE3qc+Igrdp
2pp8lSZSnKbR497MFggqPjp+RvhGgK4S1dmtkTe43gZ1qO3dG/7FK+xNxel2W/3ikm98tKnYi/uG
TkVgCtqYSc+bn2bGqQZIwOuAh3KCpM7WBAxa+3hDiGAnMlaVhzZKcuVlrUjXAV4liHmpRffIcT//
Sysalm+GFPJWKUyaPaJlfKQAzwQUBlR1Al6VWqyaXNxkA0eklsEY36rufMjDLukm9ppjHfWF3cAL
7oB+vFpccRVn58q5GrPpYw2OeGPypjotbYPbW/wEUBZpfp51pr1W0M+e7w7XnKtRp26HPZ0qZmWx
oOUiF+yeG1KiswLk+0mB3J36JlCElwCsaWJ2TVQeskA9l9wAMj/rAHMV/CuqZS9cD2oLgx3acdnJ
6Kab6mdfaA9le2/O65xkKbLe281e+mcfWtOjHEEUWCoODx5KVnSdieffJsjAUIGB2fmhRtVg9CmV
FeVj4GKtBL+/5ECQltydFg2Dfe6Apf+ebR4s7GkqB9up/IasBW75cRHt6DysT1ZeJYPgPpqLxeIb
pEX6iUvL5tGGnweMwxoPZrpxMeyp19g98k5TMP7h9Livi77KuHJSx37BilHed+WomfFEvhhlYTXG
eF20oPHi4st0B1xNMhxI/GhCsTSuZEoalG1+WRSF75IYLyiRaVlozKfrKCS0xBIm1EeXrP2rItn0
0UkCHFDQEh661sxZRjCaW9iQHZGTrH8CfBvOvEDgyGWGe8yWPJMFlhBd5Sx4oSyTMnlt010OHgPv
OJYQ9NLIx+2Fi6M06RsT7R60KvYEr9PgtilDiTMhzdHT/Cs1XLdLxXHLf8eElWsU+IE1oVIyTlMi
1rl9j9EGPmWCbdXDrMVlHMg1vl7OCgckEOVFkJY5wo6KF/DMnsLOjk7ielCa/WXU8yw8BJ7IvRwA
nVll6xc7DSblh72Fq2oKTaoLnpTuwwqNmVQkhpXvJyTTBEed0q5ZiqjSqsWjA38WGNhdKqf2PnXp
Kmz7jefBTFzaFG5NisS2qNRh5iqB1urD9i8zb2RCoL5senryI0TXwg1oG1RC9AxSJY1kZnt1fDZl
hAbzsxUy977prt13KO2arAmxwL1xyQLXW6/+gfqZGPvfgmOuKF28WFh0YjpG1WT/lFVXPusPcNHc
ARMIbWPVS3ZC5c2WbccnLIi5Kb9TJuOb3bW3QdK0+Y0Z7iry8OKESc5elFbLp7QTj/+XxQtxmrup
9fExoAkeU5O5rZ1pC0164JR41KuxlVAPkdvNmLV/OnAW+CWoCWYcssr6nIxArw/k5DU6K63p++Lj
pRLY2f4Ss+GfavExZuX/gaOu87yTZKjei4SbdviJCS726NCMYRuy/ufkcb0SqTg8XYZ/dqukuKcf
ZTXLG09U46XdH0+Cj7g9mK0oHQmQwDpSCKhMbfFUr7zFR30thZTo0AAMRSOE/2BjFbABHJxghUt6
Bh2dwcmm+9T0/cKFGqBYUxMRfHv6MlWCuSZxEMheUM3RSBRA09+nVsKwgVKS/gcsf0afiGC9z9vM
od0D6T1OJpzi9OhWj8Kxuq87Dm15Wb1cuYQwu5URxA4SVM/vmtaOWTMJzJULHed7BdjNg3aMIhVD
+XeQq4Fa/r/Wl7Os9qe0IXDvp91ZF7UVRObtK6oAnTHtAAeR7FzwSdX9B0gLDg2x7LgTcpIBWRDB
WlfkEQy1OvdAscVq0rrwpvQz6XZ/qlMvbGWR/Eww5OVNt6/ril/jAyqp/SB0Mw+GkbIrAsUfF8c9
QYiGMpZaIrAXbzzXVBkogse4O5UQtBcio3R/5OfkxMOpOERUXNPXuvAsSFLZknbaaG2fVeAhRFFF
+nsZ8r8EW2r3+l+cxpjn/bvnt/jSDDSwo05yn0LuRG0BP0uSrVODkX1NufIBXaYNNIFjt/1YU5G+
PzITuus8R/bH18qI1JIPYWN35BLQdzGep5SJ+//p0oiq2eOWrXv9PXscossrWf4Ce7CAoL5xcR6T
+wsDkECJhCpMQci3UPktjSM4oqq/BHxCmpmCaZ05C7fYqBucqPvvKAvJjoHr8jdoVveGMoMcmpha
IPw4tU8C4wItYqkG3IdPJCdnI4LjYTKzlbmn+rvRwfbSKEvRfmdsKvCrfJcuYnBzssVHFgdxvZye
DqUkS0qAuRb+gRkF1JTiQbkoOoPBwwUx8OaKYVSX11Hv1uEhGsH+T6Au0awkt0LiqV9T/nXCh2rv
4IeonNHDT/1jep6d+4am2DWQe8K3nxXDNPmy7MXsIWd86i4OEeJdh66vC3EMPAyG5mQtMQ9OtrlS
gqOZZAmndJdT1mTaqvoTo34mnO8F4oUbZj3q+W21hBqghC3Qk9C3yNcfYkI0O6jvECc+VJJadgaY
bUGqFUicVcVtTmxuRPMnm8al0/nlcOih6cjvQV8GEi2dBEcaG4FxxlsvXvgdnvMztodn8u381Iih
TfofCtMHP5V12lcgHJPQXHfzOK/00V7OtADRwSePBQ7up8PiVWbygqOD6PmzjKNJZKQoWnRU+KSj
aYgnsRl1ez2I953kVIVnTN3byHzGO1ZPia9m7ANRwzuy13TMDg5RwXlOavW5ykWXzh2ukwEml5e4
bMPDDOA0GNKkzfTFLojOrxOSa1E7PFIeSNOiIbVD54t53ojMtRiRLXyFUfKuVocPr671YGG8G0Td
e1r1OUQ06w+AoBTezHk5Z8rdQ6G4P6bhootO2/x/T/ufCODiBKuuyg1f+v81aHKf4PQxZ5fW84ct
X19uHOIFwQiTP0Zw9gZv+Dae7aFix4n3FUdiuCMd02w/faGnwGiQslQZ4LA49qy9rLnow5ColCsX
dCUa2YHfsdbzC9gbjVn2H8y4jb36OpC64XE7jXa/oOTfMYw7fk7XEGV8PoTPBo1sv6ONwyHLmsTV
g9N5tgNP8TL9r8xQPQ3vsgvtX3Gdse97z8/laRNgGVxH73kClLVTGpYkIzDjF/jbp9k/XLEivNUi
m1iXp7mIrg3jDh35WR+h5v8pr2M2ENtiI1o/A4sJKxlxzLFrLDes/S8WUe2oxc602TYeZZrdvULv
UH93d7pUi7Ov7yPsFJ/h/rOUubqGZAe/1FAB5Jubs0SWwGBAT4Oyct706dVrmtPjqtRQJI4duVnD
6sTEXRgC5CZ5jyXtHWJw6Z+Hkqx1icd4mkaWSkPPl4ifgewsbYws904gWxV/wiPXPDZXb1OC/45/
RhkofCd5fqJfdpFgv3hwIMmlUns5TJ8jcnyv1weZEL/oOKpx/62FcN2WAfqpLg77PkgcbQD3jYnX
pgW4i2tDJESebw9YAkDiYz5MGoChm4ahpD9wRmg/iWB5nRSjpHFXiqTLpzoWvm83JkIA11eTw6gR
0/tTbf1MMeAX1wwGJ0FCJOYJWND08QEBcrm5GNOJyIi5LFoSROvUSPHn94Lo0v7YSxd817lk52RP
/OEkYS02EYIG8CicefBxWheJa4Qk2NfQEZrdZnHCSuEugn4H2fmgSH3Ivd10yoAcVCjvtN4Dj6Tu
QNDYr0/Cp7sOeWaMHa6cUCXDf/mWWuoMilstlgjFursE683WLafjShjwddyTb3OWvbDzkpq5Y56E
v9LKsxCxStHPeSQypaSjBPyHD6ldquwJwRnJYkw+yA66Ck55d/KuyUGjTDI0KcGDuyhL6ETEXqIa
tBkhcO31X9RVFYwxtLbfkm3KUEvgKZIkfyFivkOMCY7r3ruivRYJtLf6Kr9tnOcysB4+XGJ+5kNz
Jyi1g7Qx8OT5vgth2CpzEd3YYwtRRFMGxQAgIk/KcJICvr74bzfWQrPsbeABnWGy5US1uOon64kX
zLobbBNZ9+9pw5TqYDn/YILwUFQx7BUnyJp0zqT77RqnbrDPT3wse4nw0Nzi1moCZWOZlCvwpRsj
28bNiERK99GdQL0LRDXPwCuEt+17JKYcUBynVZ4wrR+t+/GEYLe9YMbrP96VtLmquEpq/2w93xEm
XI9NXCiHb9m13BAYO3gn55be4O8+oyyGTsr5D75qEMuHQcfn5WiJu36qvQsbgSj5If0sWWF3I1Rl
yIm9V7oH0wDwOfU1Jfpi2tV+BZRavTqpruN6wPvZVENbhTplgTBGcoOpNW0e2aUUXMHgfMODD9L+
usI/sKRRNbNtecb86EzuZ52tP1BZfKkn6HgRcpJuceQoRQrxKvMElKpSBRxk/qAvNsXdhm/vLA67
+1orIi/DXBPf3sr63v1wBmEQ7/H8PPWkaxldhlVAuX8Vyb3U2VyK1ZfeJ1mCIJgjcqinvKcEDR/1
8rtvS5uCUc6pPoVBTQJi/3fIUuXAK67/P9IBeArC7XuXXF/zEyUz9gr+elYAGCbE4fUCUTT7r/pN
vsAGrpOOyZMR/3xno30SK13xjFgzbILv/dPjnLxiVDc/Yt1kBjEOXUtL2xpmNZ4tOD86o6/8aP0O
/sxzFFZ4wi/eekn3YwQS55BJz4JJB76VZy4Yp/IdvDloPmiyMxAwwEB5HztyN48wNGmcfd+wy7Ic
aUFXQTXkdCbvmOYQ1s6Ydap5fAa2p5VrMxbzK5YUMVwQPOS40jNLeM0PnLq/XZ+yTpCYzn1K3Hvi
FURSdkQSnMhuyqGY6Wj/EK8HAoEy6tG3A0ls7uPrCfGRfipB0cKff1/tJ2ehGo/0YxCq07pTmihV
sKh3XnpLUbc4PghZX38fRgw0KOE5AOQ4WWsYs9BOND3i5zO+B24y0Y32xmnEwxdxn+tjnRkmZca6
hWNqElEKHA1WgnxLC0/NmHK5f+1UNSaTAuG+mDdVU4sGu1NFDo5ikQBLKT5gDVSA1o+DxcfA36gW
gaGR4QXKuUls56FoFF5ofd0YGwFr0kBhbinESX3YKq6P8dQvmeLcEN6aEAvlw5X7J0OS01+r8Sev
zQMWKNVPYhCRXAIkYMnAi3pyYmea7fFFZwDaZN3ZAFKhmNTefhpxFBl9uRg3Vusq1XJxblXpniOj
Gfgh19nAGhd7hW0SLYO4SAvGf1tD/K6FbtxVAwCNdIpfWKI8Ow4z+6vwaqylbOYMkmvFsoIOsucr
dGExT12YFL1PA8K1XOPR2Vd6mZtzcQG09bWDvzu/ZX7fY6h2/QFQBtIkWRVHaLM7xDMm1v1esemA
ptN0Fw4Qj6BmxdBOR+oyYnko/ZGGcD/X0FRS3yO2PqUgQY6yMuxzslbIrnr2zHpsS/CLhWCj0j6g
fMxSB5VTiXBL8eFGEC4sP6lRMwfzPR+b6fzh91LwVo2iaMhiEvtBhWQQfkB1G46hSgYaWtecWC15
jX3867St455suam3xF+n5xvDfJTZQM+KZ+6mj17xU9kJHKfTIRmfiwsiiYmLNBr0nmlS7rLkV5CN
+JOkhJLuC1h/Zh7sh1fkqkq9G8zreg30FATTeqvGZANk7eWNziikx+EfuzMdcKiZeQaoaF/5tWWh
a1gK5OjoCrSK7QJgv8enDdxi1QWoVhsVbALRUpS1LvVoioW2+0xrfDJV+XvKGPIQ6FFGxh/WQ9si
iiTjZVrRW/pEk0YCJ8iwYOCDZWhg3ApHtgneaoJ5HtP0NIdMBBdk5NFHkrKCmQcVZUpQzQhakDFb
UIj9L18HgVbijDg+YILb72jyAR+GCBTU/gXiz9HkAHqnE0aI1E3GaMi1oVRjPH+vxZW1An7jwzuj
rReEbNOOXo1rU7ywFs6ycclQErNdXH0UIVPJ3g1oUKFdljrDZ7nZTSolFvDn+Tj6DT6zLrrauCeC
URu6FeP4BD2qSId5kVLZgYx4AAyXHwGLxwSPMscWAMPCypyGGHwAMEA5yBTIGPkTG7ctVAGl1vJH
QIsYekyr90++SsWiNlUmc6GsCSnYJ2Pu2lvQIB1YV/QrCLDUlRuE6S5LjA2dpIn3I4vzh+L8Yta6
Zdd5caI5g6DI1mYLpxlysYo9tkvhri1zy+C247+IqxGB/0NfLLpeYvsbBiG2kADxesuRxCvSmBCS
zrBQr8KbghChi5EGFZOpVlMcJf2rCZt1fKsvF+s4FG/X7g7dcTksB64PUyM54Ryg9HLpDKFoAG/7
VFnT+OJFWdWBHPBVVexBRKJ3F8UX3t49r0d//43o7MfjkXk1LVKm+znrRr9FwJ3y6m3wPRNPB+r5
C+3V8QtELzxzC+VluysDWREgnQi1hLRJysPqIsEpFgWSPyUgRqoSpJigCt7IbWilNHJKN5QSG/rS
yfj4uUnlUisnHYkXFgjQHzv2IF+8htHLGCoGysucUH4+HRZalWF0I5qFbjKLfElOieDeKWBMxqbr
jUEp55FW2AUuow5S3516KGK3mtK8S3O/3VB6CqWBheFPCYyVckGLuzt7/rr/itdDYz3BMwsuEIp9
imMdsxN40k690ZbGkJZFOuArvcElVcr0fCJaCl5PzOzuoi0x+qrc/XhYmsOSl+dpE7S/QTvijcQ5
ZF4lVGbshZNH6L8TaZnbTzeVwLLDCIqac0I3riamhQBB2fvoXwDupiWu+wo28ZVcYvbUUJFoPmxm
xybpFR8qY+JLhOnz2bkKkOLw/YOOh48l8585lMJ/hK+RSik7eobk8dVDPTuqQyzIWfIa2zmP5HYG
iZUAEr63uf8WCoULsDX2roN//7daqRytA006bNkaQXSQOW72TnP2da9RvKYcTsf6zTDpgJjn10Vp
x6snUajME+8W+Jo0+U8Hw8hnDQSiQSG8qwQOZ4isA9Vlih6p8/dipS9+wtdV4RXy6nsG0zY09cqV
B7ZfSGjjlQXKXM5KMyIJPGxeTW7dl3a3/oUbc1deHS1/X2N4uRGSp5e2pEYFXII3CksAF2aww/bt
c9ZeIImOn5vjzf6H+wDd71AEZp968IZxpWD1gpP5qcYLJzN14APUI5gsZVMSjrMw4JviK28Zsj6c
SGtCTwU8MEKiBINqQY55HGUCgCMzIf12diTEFSF+SLCqj1JAA6/8BDeXNy7eLV81EFBFvzgLKJuy
Iz8N7HQUEVrgwRbXYPeuFMaw0alZrZRmgTbRkfVKuQ0yxqc0G6qz55m5xKNoMA25D3RwyFenVCFQ
EagB/zrc6G6lwpowbMj8IrBC2ZktrdCa6B5WkaWPQFin+u6gP+NdIXZRQtsESirBq8OAD6Wac9DI
fLNs/rccDRgASvJrVJG3YNo1fD9eKGgFuHmO2ggbao2QqgxFk2As8FenS9noSur98vb58JJTdGMR
Sq3ifpL3k9W9ZRU7hw/xp6cMyPdymkLUIcJ2gCj0YMDcl9lr5jCnSJohoqc8AmiKpatqyNux118D
QrlYa1wscLzkbUVMqsSSG1psuf5CE2SDmBYgDHdxPn0Dd59uBgze+3Oi1wRzSanD5CEHcKB0wAGE
LSP0vi6LccWFCkNwewYjVoVjKBVh4qEkUi3hX36aSWlYzPpeNiQOWyH6eCcKpr7hFe0lQoE4Lqa5
Qo2asAIc0+qGnTbpEA00J3tbDZh00YS6t2hIac8v5Gz+nb+W+HSMi3KUTSWfL5q1k1ktTwF6YPKN
UMjZqlVi46njx+GToZQmTv+ZdrOFAHZOGbKd7ocWUmNVqlrszCCBFedJI70F4rhKRjvFRUga2KKP
nJH9WBGQKLjLvFxIBgGSQOLjc7+Cz/rrAixERpttC+m2qbWFy8lgN3g/bMHTVI6SOWbK6+ecqrTo
k5yHvatpn/JfpAHMM4BV99KooYajSVh8iD1ULsxcS6WEEKGavWRbM2I/FPdUpUnQeaxnGyH84QaZ
wjCcN7lMARg0P3SpK07LFoes7NPDVGeTsr6A+MMkD1QYpq+Pj7sLTZeuwcGpHfYg2RKBEHRpT0IN
0r4jV3qNdGqn38XUpFmx1egncLJ383scFVR6sEBSzSC/cJ0gNijV/LG1OBIidOQP2cXylYSiwdQV
hHoW7yPpSo3hmftCBVUVLYdlMMLMGU+Mw9wrEjAVL5wRba+UPJtsIYFTKRn2hAf9kLChPTl3/Wfg
/pBdRZU2RnsoB/PHiJJra7UXXxp9Yzcp2LEXDQA1tIODhlgt7N3YzBKX1tzuGUYxwdmT2sEoJcxA
L9WexE29imF8fMwQyE4KLOs7kDHk9RAkfwI0778NHKoVY3gEigYfAitaJ6h7VNzyygtHkbGgov6S
l370Yp6Eus/px3IGE/7oFiOS7iTdBPmuEeAkq0NtssmtnaU3CbCNz5Vvvfn/2qzRBAyCCifnLesS
OClXHsOgMcqf8YVMPyboyls4gbQV7e5iImCO423/fulm0GZUZY8i0N14RnpA6NBTCY4HNEhzG3+0
9ZAu3L+WVmAsNzlZgQi/cCbstOSlAzN/Xhj1rLFQXxWXthr8bcacWYtdI+vLJ6ePqaxfyBjhKIgu
Y1WAr3Fl2BDgD1rALGUnJ9tfKVtqtP0urY8nhF/aKna//bKlQs3AYfQGGhmKMzkqVH1xjWK2v5ZU
YQxBc7qICTxah8orEj6M/61IEnQmHMNsnkd8k8KGdqRkQ/ErzHIrzIn8cDO/LUfNvVcZw5JSeD7y
1XHT/Ps3VY+6JnCLr73RtNHGJIoYPvemNS+HrAhwLavflYDzj64pqvy+lLMZXMrNs6oFVhLp3RT/
3GdVreVWEwgROac0O9ste1tBJtSj1pAooFnZSJQJFnCuafmyOWrMls7Kb32D7eST2wFPQ0PoVtiQ
bhUsQXTeDOJTmxTq4me3ukqjPCHUrXt7iC5tz9tDmnIAJbFJm+Me91Jn0f9CkngKWPU41m37oIFU
YMZwL6Ou1Sc3qK5GK0ib7jj5hT49y4yQjrJZZqyEd3iun9MxuvInSQMk9x5sW0YVCRsrCeKQObtD
KxkHbzVnK0JeJW1zmE0yOZ2Qrb4sG9AxGzxdNZbvJAhZbyGzcss+7IF4ru5ksF8c77IQa0RSZAjb
d1Dt9MUUwVZtbRyBCmPklyT5TDmdS7hG+IWDVcaXwmkwm8PMMg+5TskgNOSerUc4uYaLXkBqjFai
23X1+ZJmYZUqpL2oDHnuTu2u+t73qBV9WnysY6ELI27TzIPj4+/uz18GeCweNinV4Uc/vP18s06Y
5HNgpJdmTvUgoMUyOXhk3UtSIKuf9tqQvJNKzlCYTOTaycJtyCXEaAeRjexj+DWR5z4eyf5cPZdA
slMWXeNP7kvvctepRohnF8ClgvxgqsVmFr8eNrKC1uVqwhWZ4GdGyNx/G0APLwgGhvhlHJbVSP1R
5yoxt7PPvH2cZ0WJb0jz3Mkn3BNKDQ4uSRTUmxSQ3xhdbm2xsVGZAz6NFiwF2gBjpjqu3bfAlMap
rfjJC2OfXqV5m9ji0W/80zl2SBKMP4kzxC+aXRNKEJ229v5gzD48ohGm28WspvpDUOSYfy5p0AnQ
Vjxi//RsPwjXmltSpYBNzoRIb4lxEyxZiP46aCqwOPpffsxDqcciY4SQX51CabqnD6ekX057PSpq
8L706+zlynuxFJHpnwpN0INi1ZHKw873Qh5GEZxBeEHAbtwS8FbxzljJF1/YMEpQntikfpIONclY
/A9dO+TqoPSLjeTAjkjkxGwtnkfr0eRExVhg1AgznKi3s7HQKUltfKkdx+3mzH7Y0L8qSBoNRv/C
N0kvMmUZ4NQPJ5Wu1322QW84Vd4ndrtID2uU2VkyH2YE+fWq/YHPXCIyMA/uvAdMl2R2P2YW25Ge
DifopWdau/IXnaXEV8c6L/1CtoO14NbyneOSxRk91G4RtQk/51GXQET5t1rhsQ6eVXVFwgcn2Un4
ic6Ca3c8/U9Glws3HpCBfO7+rRFPJL4BJb9tV5rBOGQKlsvDc8hzATTQWy2kjlCNuDY1gOm0yIeJ
XNkzfoe16Lx2hgkL2XLfS+n9PINXwoIPAp3x1tLT8UbvAkxDudCLavncj7umZDBhe07gNBH3TXmz
4GCICaqWxM3iMorh5zGy9QZfdUjKAuufXrkCYBPnZOV4iUHU19VAaFCFNuWA9slKKhkldkRllYkd
rmWxwUZBZr5AOvwZk3opaaqptEw4+LyFaViT4ZJKP8lCL8PkRlQGeeUps6nAidMa1+U7d9BoTudP
Ok7WPZCO7Y6cPWxLlPVbRniO+f1zBxlJeC9EsufiVvR4Pj02Ps9gn3OXhaRFUP0ws5oyZAl/mkEl
BYpxka6FK6vAXcBg02IGEHXG4rSopEwu+Pv5SowOAGzxINW4qaxHyhuGaAiFFGC0MjlS7Tl/yenc
B9a94X5ebc1iZNq6yHZ8sp5Et4Z2GtUqaKHt6Vk8JpLjoncy+x7k+nFPecbpO0dTCgX/tXHOSc9M
M+TB1JRGu5I5wvnZKyQkxgoq7K4OsnmLNhlouCouNw/e5J3m3MiALQLnbQUKa7qDehwubdNnQskZ
jaVdXdSVxlHLYZ1dVOzkG0diBWhm2UYP/Dbg3nadvX2sQd2dekHrd2doPjA5+VyRMi9QF7wqz6Xj
AB4RprvFSTFmRRFBih+2wVuOz+vw/+d/edHgdKPVS8F5DMen5WF3wvTlufh6NfRy+jViUZ3iIi7r
ppCXEacQVv8NoQYYtwQlIIMVqENxFygKZrdfojV0RTHvZz8ApQXdJmFIXETWnyCu+Sl97m3mgrUr
48NMtHXGjwCqTZu2/Neidlxj16a484oyT/AKUdg+XTo+w3FclRbnO2mMUEj49fLGGYt5e6jwVDZ4
DaJ9mFBOVFDX0f1MWH7+7dVO2NvFRSgWn99qHjzoJYwI4WCyPkA+vc5Tv1l3e96YhKQAdmITQeqL
x/R+0Wr1/L2TsQ4tiXWgBRjs+j6yYa6O0CGB+qtLj7d0/JPW+jIpOxl78LLSLPZ8k3Re6nW1XoyD
namspLOAidsBkIdLYJiS4yXfjs37Z1VeX2xHHAe65noB0jL3SM4U9q7Iow/MdLGfeI9JXV2MOSMn
mQFxgToGnCdSML5dXiYVAo635sWFuNYBwV1AehvQZjrkK56d9ZV07deCI5TTPvpYKPaB+MMbLvLS
CeYY4WcJ//4/X7gH62xnxWC0LUPLR7vNthDHQiUUmNb1MoS+w7Lo3YWvRrwxEI5Ev0jCvVVzmMBO
RYNOdUXUq4ldCNa7rL6K0Z7TeQ8X2cOQgZ4dqiVT2S/Kl5XW/MIR4wJbDsAUUgOpKkeJrhArpbXz
CKJiAJIaII6spGlQIdbOovDQtr95kWDvuhBqW19b8tXwDZJwn1SLsCzUZzdpHc9+R1Uso5it5aHI
5sVVsNR0idft8RvaV4Xlq+Uf0wmbY5Dbfyo9z2CsE2S+r6cA5SijHnE9bfx2UKmGf91j/9j7TACF
ielYwD867VDtKK5/6O6/PHvJK2CbFJeQd/5N0kDZp1eKnrPa6FuIbbQ+kEtG0IBjploVl+E1M4Zy
fsHClOHYDSDaGzJylNIW+YHZcbxCUEU9w6Ff+NenOq/4swUWbogtSI6epKTLmKNiS0JjVYAI84kS
T0u/YIkGUx8p4igU4m777vM3OmzjVDwObw0dEGV83DnkV25JbWwZ10T4FU1c1osfQtgYuddnN9b1
pY+u/jHje9bo+945pxzJ7/znpjpWkVQziut+uo1iWBQL8ip5EOERXb+Sr+V0qrJdv4z2Ls6XvZhp
BSRB0lQ8WZ5mCQYH1DjSgXxXwtzvdJhKEnwmq3GFdIHcFGrJ5YfWsnAgeVwHuaJChUV4edV86n0c
9ql/CXSZ44pcDDMkCCxdvOPr5KqjUcHyLiMULmrdN3YckNwDL3X4ffEBdOAyosw4DruOUfwv6y98
uNHuf9HFUn8/zqB7kQxW1YxnCoqZLbEYVP5Zfkb03JqB/wQujv/R3pu78ghoS4px6ODPsG5wCH3n
TiXaqfvnKafiSTSeR3zkLZ2sW8F+fyUdejwq0LgOhXIBqcjHrELIVNMBs+DkfzF6e/d8IPr0cUYI
T5/pQ4BpShucT8vjpHqJFS9uTVKu3Xj8D9z+Vj8pg1UHt8/NFJac0d0juZxbqPvpXekaQG5A/shy
CA9JcSoMI3IVS4MyEHq7VavAhHk6bjhHdC1KbhC/UvTnq7/rZ5nCDWNaaPJ/UAqGew9BcM64xutq
PKOXXr5nud1VUf0hkXUqClWfc1ol7d6YLSEsGZEflt2ioR5Lc2nVHjccEEwv61EDuLs75Ufcbdxe
hPRXuWePAplr5q7ivX7utUh6XFB7rtVuaLFuCZN7+lKnsJQOkbF4uhsYtuJrNMu2PTGEcNqRaDok
lq0F5br2b+PR/rBOn5etmA4oJfASH0FxNsIBXKLsdMlLTDSMdFem4y7c/xMJp26TJ5I7JBUjI20z
uG/V9hgkLxYi+g5RF/q64n89Z6THBxEbBONiXWUTuOoYbaroxC0AsYI0Ti7V3xv14qWzzi5tfiS+
Qx90qH0WGqlFonHq6nRaULMchChyl5uHV32awof6SV+M4NpCyPfU/UIsLlnpfVg28KOc5Z+doIDw
gDAcAzyAUuW9e/4UK822hwYopbMTdj/cIALvPJuKbX94WZNtcRrfHx/6fFSAGeQABE5EmiHcADyI
4HA92eujTQqqySwZXUhAUjnya7Mj/AmkO3O6e0/QHf44sObXBnLallTvTN+Uwzp/0JpzQaXJrevm
NQ1GJ6dc7t/mge67wCQ0m5fCft0NZCQRD8lvKw0WiAzitOzR6GTnTEXYMyvmj+zedVjtjlqp87Hy
owqHts4e5D7L0KdU9wv0BJzTLpAleiVMZczRddC+rr0VbZ5VISERUIR8lfgHsQy2ONoCgsW8NjZE
uF6U7HtUQhAVejZ6OrywM068Il4QAxeTJZOmYYcZTFYx5ADFtE62wlO3NwbvA6t1Q+HtTTnGAfK4
wco7yLSmnNUr31kaR/ywfJGheckzhRMplYAiWuS2cQxLdOA1oOZP/gcpKZhslT9fCG9sUCiVG3SO
qTfybUq2wANxv11RsXfBtCwAsNR94kCRDfCIT7WLspx9If0K8oPEQj+bSd5taCwlNiWdEXMbm+0Q
P7CoRXbM/KIlBLy8BNxB0eDZX8M3ByiwPKz1b8O03yFJUX8OmUoMnLGSJ40E1BRGTKwD/hpt+zIG
+/c4SqAtbChDSdpsYWUKrjF3T23xVRzeBzkob/T2o6quVin5Paq4xFS8PYO6fcXKk7BKP8aMd7Qq
q/OHVcvfQTg3vXNFTDdkm+cQigGlO8g97nZ8c2PkN+YbpYvB75Xv3X4ehIi5Px6v8lD8gXedA4u4
QaqdH1/HRRm9FHrmphs/1ckoYldwRGT1SRN1qOX5eJlD7v+R+vjBkQ5M5qXqpCbsTIYuG7rZ/h2L
T6x+/ikV1x04k0rPDBkND/fWr/zxp+aYbBqqyOWNuZwtVTZLWv5jwbL3sECkayrUJKpvq7YS7hjQ
RWGmWTO+U2CXp/exlWk6oGBIQqXNmct7zNtNwQhp9mHO900OiyrZIDdeKIJ9+MvyZ9zfOfeK3cbv
DDPJllO3475jKOI6iw/js/eUpoUcDjtTsclPrp/3mJ2Ptmnes9AbEKvhVzu1McfBSFNQcpMYp4wE
Z9NHnj9Q111ElPnaoD7qZ+7SGsIss2WvDcPTdTcoQYiQ9sOHVS/mTCIBApN2IE2mmKxlsTAUQbEp
zadb5dOYTFQxNAhLDONg+ANPT47JlUq/ig9Qj8TBrffrfCjyvmZXATL6e8Wic/jjlhIQ1BzFk3fo
7B/sbocdalHZ3wV7ErzHnHeu9BO40TFlq2OEFiyH45RQ3cdoa0cjF7zQofirBeTiSes7cEnShsC6
E7tcD6ueFa7wky4R1HA92i2FZ5DKkFBwe/N+p/RY6YSnccVh/D5gOtaxzges2GwDSkxSMEbR6Ifu
9eGOvF8+GNBL69nHHS+zJ+NgEVRQWb24z9rncj0CWs+9pXVVt42Y6WbwtPc/I3D/qU/+3pW1GiNN
k55mXkleT+2LYBKmLeYaY+IT3O7WmF+r0dtcAyFy54goBDonKkl2wg5UdXdn5G7MFjH5k4efdrR/
P13noWuaEOyiQr4CPRr4kqlpGpOL7zdW58hnvcUGu+bYIXS1i0dXU+OPTB95yGiFpi+JtTAfkVxN
X1aw3qMZ2p6BkHp7VmH6oIGeZYLkCri6FXQgKcPM1UWarfiZSS9yWi4xqZ1PBwl9r5CXTt1HQFAd
e8VybVy2eZnhL06L10jY1gWvhsOUFW8ELukeotCVHZvUWEAJQ4eU7z0yYMUDRv7UEYp3/frv3mIF
R4GeLpH2Rc4XTFd/mZN5OwyGkbp+P3RSCotMfcR0XqoSVRUdI3CRe6sIXC0wBWukujAZX+Wzrc8z
MiT5u2CCOFiM8JC2RUr+GOifQVlX7WaVhuMEM8mlKjcxvgnDEkGNMrVBXeEY8mAXTe4+RXXLcj0x
/KrDG9RmB42SQzpvi/v1rCl+WGfGGXgTW+i9sv0JurhuD79wI3LdJkgUzGHrvz/q14RCeG1tCSsa
8U89qugrMx33OKhdC+12DxHBLE/EjqvSO4q4eG7w17DDsN+ELU+cbiO39vh7ZxJFq/WprjhA4Uc+
pWlMP4nWLwHWEtwz8yRFgTO2wGNsQEi8YPCaaGFRUuh5j19Jbm6SW2Ecjk0Y2xqUWrWciofwrlla
Ayd5kFlub1JvXsboFam2NE6N77KQWzk4thveXJKu3bDuLzU4jfD/LILF3LPLUMDjaBYyggQiyxTC
opEPAo+lW+YNT6nAl/4P66/carcX8mQ+ZIL4PNZbrWHL9t/mVxuizcXbp3mNWumLrS6SCq02DGDR
FqXCXRUlnnwQrS/UZLZo9jF7TH8GgeAqEe/2hkZRcgCcNC0cO510f5y1g9EH+b3sLb2D4cOAEur0
yVFNFE7QFl8ue7zwCquArvPM0rPsjNbanAskqvJFr/wl7O+U2h9arIHDw7luPgQnfTvUbxxkdAJ8
O1ItA5OSiZBauQq+4No0sWqn78EM+gHrfleXNmh4ChHh9jVcuNPgEdpogbtEtBubLimwyJvHw4e5
JurUvkW89tMY+99ybeMUxUcAM/XL3wYrsQc84V6WjTkGpC61sZkDjL38ALaIvuIm1ntEE7OxNCup
PFLr4J1IBHmh49DbnWtadOOioucnNhX0+qZt7oePfRK/uMmleg2vsHpharh9OytgBlEdLuVmsU8h
j9aKIqIrz3YW7H+Cx1RGfNqzDGEf82YTvZzHXQssoVQEAS0G8qoiuOuy3sBf3/lbAYs/iUrhQtmD
IgTn+PuCtPOdqL7aMem0YUQiPDTeCFnr6NusSTG+59s+n/Bd/NWi5ylcNyLPG8NWkX8jZd7YiIWm
73qZuTuDEKge48UX3thMxQVaZYMJfT9t4LB9lnfllPQbp9CTa0iwobBjZ/yzcO+1K1TRLwzD3bo9
aEECkzz8pVeVuvwMD224xdB5RoxyAmyOqu5ZtX5e+7mTSTj0wVSBIMEFuSnnlYf39Qi059jetvfe
Feq1zBQE1u7yuw2adVl4T08jE//JZMjQW56Uk2yXtuu6yw0WN0NAUNZNbixTjdrCyIRqy7aEamFB
XCW2OhpLMZg2JFELUylK3d+ETrH4xyOApFcPUxEBCgtpWyCeDCcouB+Lf/pf6uyE52nUZZqRZCiE
hEuIs8uME9mdjJiGRAs0zCyoCsE8suB22Z4qxU7H3zU8ZnQxxFJFZoxXYvIcT23NnX6ORJ93cYfZ
Di3KK8cZeE15y7Uum3qApaZmEa8EJ6l9ZhT8LYGbkA9Evr7TCMO9Y3S2oLbAcmkdtdgleNBlL2Un
pT/+aP9TAx61hFZ/7/9/adZlESGbrznBH4exolLR8oEOIoJhZ+1oU/REmR/lWKN6UB042WlKzvke
4NKFg1sdZGTrOnkKhktx41QMKaKPTcFdIpxrg6ITFm7Mvc/636mSsEJgGhRWKSaUBC9WH5qwy6aY
EyRAsZBMoSkbrnD255V2gD7fOdZXyFB02oqv1uGRJ+C1b0MAA8OXbfkKto0f0odL3EeFcPio4sKO
0EVW2xM3+t0YgZI2ok1LoABFwF+SFWY1szJoa2y4lmJ3/3xeXzy9VGN+2DaVb3erOpoq1HRsxMRG
G8CT6gA290CDM89TUNkFEn3fDpzGxWd6RYZOweYukXkRF5QFRdfPEPl0R4rFh24dZJALP3i0Gl5z
VpmY4LjmiQ4QmUcyDFfrrZFvMHMJdhvFQv+6oniYks2+Jzq0vRPOSRASt9A9TC+fEZwdtrjutldk
JT+rqCYv1XFJ4lQqcw1k3GS+yPOZd3XGLqvTJHG2LQa55qeW7YkGGVGNGLj5Hgq3pgAKv/AWgT5Q
i4+KnJDlYCDWnWChRK2c/CELMB9Bi2D59U8N93s5E6wi4PGxbCq27OpS9HOFnmt83muMfb36QNoN
0YwZo/ic1LS06Bq4F4GxVM6wCkP0KEeGun8XuwYcCspZx+RCab85OsywsXuIVCbIIaMKQsRYjsHL
sbuf9sl8OiBFryh/E4J0Rth3vVP7KoE4GFyUgEubF3CyS1S0Tubctkt22VyXDzj9whkZuCDwmtQe
1Bm/6ZWIezvda4SQIhVM3Js5uHuoOtXiEz2/HSqnk73RPmi77JbDjz91o6wVKOZKmZAdkk0SMlFc
3h6P2JJZQfSqNJFXd/11mNeKj1ddAU/E3IX9XDxk8oQq/A8K1l9dy0KsQHdNbTCcLF25iinC/sQM
CAnidu0CFkJmwzaWSiFkZPZWOd0YVD13ZY86hlb/JhxO3H455CA/OdigiOtV4f75cgKNGbqlXEWZ
KfJFNpS07bXHiDlKsB+2ZnuFBZG2TfM892UW0cVy1yru4SB2weCH7R7QZq6vuMLtUiAerdE797Zl
OxtgeqpBroF92G0/CeigpwE8MUXUtteXtTU9/x+IKYdwvvITcnCX2I/7KfEWec6sPKuvt1GJ71Ab
1SRmUs2gBbPF85InF1buf282QNoxFHu20/Ig1Fw1pCoTAQphiJqhgetFsJ7JZbeH+kxWUrPLem4A
MFW0Cpoqp/zYeFjTGrr9bpUgPd8ytzRnJHhtS1DuHj8500fpKW1V0EYt8cJWrJ19o9amRPWxxcBo
jKsBCV+gTsz0EPUFbQ5IpXrol4X6boDlYKsRCODSfsilAeE8EY8lBjp0bQtLL0lNyPUUmAaTBlk8
jUUKureidWgG6eGgVUueVUJpmAh7Cruc2Dl+Hwk/hVA+EbLaSA58B0Sq4C51IvEkGg2bXx1BuZf4
p/JJh4fIW8Sf73prIM0fN2j5/4BKJDTfDiEXsvk0KGvgXWZIYODBB1RAG5TAWIRmueamYChO4joe
R8OmkYcUF/yuQwq5lsz9hxBE3vHCV/I8imTYCfkU+lJ0BQTwyZUB9r1doFIxkLm7Qk0BxxYEiBFs
6pYjIP1wO8zNKe/wEBF295boHqz2CAMuZsR7YHBVne8xIgp8LKJorSaEpOw6nrPX0kto55JL2j56
oQZdgWtgd1sHstYxmaYWZ/tik7blx0ixa+YB4epvQZsuLtqC1PQ2pIJdOA3vd/VIWDmPeB/6rXoh
c3wXjp7365ub6RJhdjrR3K7caQbe1dNohajwPQicPQWV3whg0TTna5aRsLP459uLH6ENrUcWGB6c
CP+voon2qVBYhBtChJrs5+MUKyFYS3OLPxezDP7BUv+iTArLj4hN34AY53AdMTEl+tuBTM9vHhf7
obxGupUpQ8JVare81KACBU3m0NC1l2SQiDUiYEfGl2MQi/dPwddkzBpKODY4f4kG6F7onoxtPC70
9DUwNAFKt/iJx0a4qUGimYD7nP2ePLYLsWC2Sar+wR5qFmrazOYhKPFZ1fuxstayUH0mnojJSn5h
X8v0dnXrxjDcqfYCS7AJzA4TnBIaFLsV6IlK9L1ruqKmlHkCDDolnKsg94r/G6HD1G7lVWRD8WFo
sw93gm4e6PCvhtE4N+hxlJdPJ2gw9naP5SQiII1+DxY8UGxaG33e590xqea8zAqQamd4d250sfo5
N9IAwq+Xzj7gOdimORPCmZh+4Cp8Vu5ZufgxU6uedxo72ITcT7xwBWvzZ0V/Jkhd75kiyAPN9T/i
x0EhVe+wvBUYJjWcgSkqVBgKfp8Hhr49apvi1Nqkl/fMCcg9GmZHH2zxwE1wncOYghwKEFg9ktDv
3fPRgQuJeszgIfCgZ1tZfJ952L0005aPMR8FKscJ+DnGqQ6Bz1j4hGCDqu8FVByy973/JRjFQbh2
TTPTZ/lw0VtbddrIKGnnCVOeJkHNGl/rq+uqPuL8X8NOCUJdpVGG57ZswoFT4NJgD0nKdOzILoGG
jlbLT7g6kXqZwbTwNsC9sw9PD/OWPLJweZ68kYe9TNDyDImvYb/R3LKFfD0sWIX1e1OPT52BNbDM
l48xZBUeVUihLVZ5dEDUoPLApFp8I9VFlXHmUs4ZgrK38OiTBrlSzVhlhK47Gtoo77PdBGIvZ1gq
MzBlgA+695eRF+YHMHb7HO0cD+PI6Jw1B5iCnLKY8RDZccrl+ns0rcrTty1PqpJUnAavfYUe8UTW
61suIrEf2meCXRWud3XEfCeHUQlq3u44Yu71tbQO9rECv8C/ApzmR0qnjc1M4nVkHmvxXr6SDlzx
cf+6GBsQiBNyPYPuw/CKwvC6A9cNbYObS3nmeIBbEvaKUHRKoY2Ac5L4/Md26RPP7dbk2K5SAHcW
RbxOKEKoV2851zPBaVlK/mlTx4K+VkWnQ6ER99Q/5TYkIuIiP0IZoY27hrtHvJef9ajGN/il/yGH
7MIIQ5bR1RQgLtoJ7X2SqXaw+1bcnaEqHQxwPh4AnghJdw5iIGL1e2Ai03DMV7YAp1nBEQhW/Br9
9xJtx2ylnT0wSSedDsSTtQ+OcJ8qheB7JKjKQuSl8uzU6RCAAKyZ6cjlw2YVw1xpKO0llBppeXSj
m+3bKWO18wDlCzbKrQqtKlhzVjqpc3oe1wPBoJpcSpgIn9G0rEzfkr/zaCjVWXD90/Owxr21kipf
61gZCaVJ4axtRrdKpT7M/1SV2nYKIlaW31aoBymgNpfTKMKeaS6FIM7bCZIcrW3OBfk7Fo1NilVm
CM41wAP0Tnljrk8lY+3C5zqQ7GKTbT8vl/4y2e9Ae409yDk/UKBYIKmLgK+vT3adXVdOsLhE4uyB
SuBQQO8WMnM4XPhafP0iOGGkfpayIbwC6PImN+Oq+XLS7mSe6oOWgaypeKbvmzqOFJ+O6JDD8roK
OXcSGpgBK0WE3FL/7gTofse5dI3w4bX1iT3D+mapsXpRv25I16MIocMuEJMfOP2FSK2v7UPe6PV8
jQFbW4eXEqL237Q2ZL2i8SJtTzXbb4mkDyUO0niv1py9w2t8YmM+ojPjVnMfhjMBPBbC0V4KzWDG
BJxeXNSfaGlDE/Nq+QPJIUqw48Vod2yhPp4lO8UVkP1ZMYqNBSt7UzecSms+rb6DWyiJODpSH7wL
gDOstwFYyezoYwGbOdjvwxg6IYkZkV94+IQGRJRyIMywt5oZ/a93agFHslQh69a0wVOq+BnGkM+2
krx+idLoGxTRr9hq3LGKR+hHeXy6+8PVekhWbtNOlIfGm3snKT+TFs+f7bR1ubHQ9nnwUUwFu0ep
mtGQjejw2/b8bogIRc6KDynY6hyxwBxLFy6dpLeKqR88VXmEcrEXyD/bwuM5jLO9mSQ/TsVdQsNI
xsHC+PeYUbNdR+lVF0xgNRojK9uVq34jumoxWUgOWMvcOuyklIl4POayoUPEyQrTXye2uQdGKA1X
NmYwPBauubFweddERIMBobxLw048MpII9MqN8188lur97ZAQDhTIgTbnfuRYDKohmuosGvLR8Gsj
9RUYJXCCM9s+gEuPXwyHE5gXoKGJ09QiNtqB9EO+gCzRVcAiMaM8w8ibzBXbHMPPabjMhuWvFvCN
uT+byrTvqUIzt8OIGBQU7n1cp8W3Rj4Dka1SGZSwVJaBX6qYqAGaFfj2jSTkaz7Yext8JmLqhkj/
vQLSwRHyIyMBDEsDCpXO9785U/+eSnC6/zhMTKmbhwRh4VKkZn3k0Nm7BbUNeU1Oi/9oUdHitbZu
R2XbiKRpjxncCMgrpkyMuwGp81UjFNyjvbzwR8tBkQ4dA+lqpU75OSNx1/pFijNK9uiQz1SBkB59
kW0goppWMVNapl38lxg4eyFKsGOiNSNuK7KZi9Rcmhm6eXEyXyXPjsUvf8VB/iUWiZPmkyc18/W5
EDnmOm80pePFjUUyqvxMXmbrVaIvr4KJIVnzDpFEDblHTH88oJXFsZwXrvRw/71+EqNIYsKr283Z
wtMr4cj4g8ChaLfOpnkqUjTu3iuCIT/FIr3qwvIITUWoWknhfuAfx8QCtZrRlJ3k7Rl4dcvZqzso
F9xyAuXyekkgiqFlmDaRhsCHyd84chpJSgygn41qeqrNbydBRat1+iJXP1RRRxYF3cdY7lrWg9mY
7g2BukiiK+LV4+Ow6BpelaRHwLE/hIzv9CAuaD2LonuSKZyMa9l2PO8+CyATpwoDTgeulIhHRxSe
0pC0ZZHi/q18boxlFnW2J0AwIpKRe3GA2joWxINsiuUK/9o6gIvP6KPbkt99jfYSPTn0/z+h74a+
JmNrB7GnC2X0tFL2aapw3C8TsmC3j4HhMHCN1MCUCzpmlh6uVhpHRqhELiHI+8UZ/oYKtEg0Q8ND
0dTraqPdW7bsxB0nsVkmKPd9f+xrw9xjRjGMBxRGiSRAg/BUqSNe/ne3Q+fFYhPdj/hK2BEgAwE0
9K7LBUusnd7gS+3JU2Cy5kwEuC36rw74YwSLRDvMkAiZr9RCc3BGrqtLmgN9dy7u6J9K4Seu+ZLI
bXNvet0+Vx4glLjtXs3CIHx+sZk8x0g1h8Z1kVwvhvGcOjGmla8BcinaNi5epy1j5XG263UxWYzS
V+0cIlfS+kv7WbJ3rxG08kWRzoRf6TN6TjLnQ2pE2hZE0afBPnX4eVs6j+R1cjjvBXMSHVGRkkGG
u4DjeBVGxbY311ZnQmmrYNwJb6Yy326gkuoREFGqgQgDm7GdUp4HWfiAATaoBzeyx9kk3zRuTCp5
CyNzy0ivH9t2+TwWtSw8kN8VlC8L8uTAiAxvQjar8DyC7xjXpkxJT5yf122lfxNUbpQRAdcYWt7T
aSF8FwuuwndOtr66Nmg/qVwh8gyUbXF2Ea3jwAH1wogmDGPlq6nJOXgWlnuP3qvQaXjIFQdHRKKD
dcXoHg4v4h6feCy8yEJVhp1do6ckuK0du14fpBl13BvChQtB3z3xcs9yzQ8wv4ZOy7XsZIwzsmKJ
8ikSYzOZ8RRCj+EL1Zcf8hqF0AiMUG0xS//txakIkghIARBMigaJK7lISZ2GU2faGBwAwTWHJDF4
D2CLK9zzh7QPYTcCD7JLa4gn+nKQXHZ3cvk0tXunnXTJ0WiXPMJHCiTnf42bAQ4omWNzztqp153y
OEGfzaSpL1a0L/vjNFEGvkiFWzl8K7cFfmZOjFEBcSePDfN3pgQ8yjRd3M36Z5t+dmpI26/VqSSi
K3nG/SZtudJ7JNASUTyzMMB2xXUa833qAt8UJh60uv8lo8NlOnOTymYTUEXwzIxz3khVv5olsUEt
LInxy5NhdjRqoGQK1Lm+L6pTOUv62Ta8sMAuR1sifVdMU8wWOOBsOpOypVM8K3ChI6/kESeutm58
9xjJl5naTfoIgtIXXkryZkM5erwQPR+LOrbkV1BtBSb8xMzNjpxwMSfg5OD5Z2LgIfVNJ3Xcb5Tq
auPDMJY7LSMmAgZGMJXlZOetsIGmA0wAMso7FaSG6gvZQKRaaB1dAcmr8CBGNaRc7QMbN6Q4/MEi
PgZzPgAASRH9NJXz/t52jx5bYc0cd1lUkgeIzNA0cNT36nRgladcAAQ/Wrrf9/Cz+ji04Gcu4dB5
C6ZstnbwE8Teb9kG82IJaXCeoqiXxxzaP47XGaRmXVSbBmN3EbclEpIcAjvqPh6taL70R8+dYuoW
nymZ5gTqlnNgIcn+LHYI8QZmRicpkIbSmnQ5IoZI22o7FfqPRqYiA+/mY0j3/1MxmX81+zETnncs
jCQlq/20odVmSptOPrEW/QQLJy+wsWXCVFQxb/G3XLYF5PkEwYEo6YNLfzYkuNJCQgtXGjM5xWjr
B0VUCtwyC1be3EgbdyamtP/QWjUdayZS21plqW3Npke6VIacKSe7J9gYnyvOVnCAgh1Lf2adkoTM
n489NxPTIsb9tL4A1fC9rkOFCLrhMiHTJBJn0b5edzwVJ7yygWdSpp7+xku5q8B1spLRTgxb/qxt
qHazV8RX2M4sYtjjjORzqSpjOA/QWqTz2sPxzp7cP0PGqsAwsX1ZtmZAas+xZ7Of9t4zfhnhnjfI
dp6RuzlM90oVs1IwZ8QSjGHJu1QUBRqVgj7jHj0VHom5184z+mE79v+bIlWa2akM5gWZgQwQI+Zt
HGWVmfB4zCdr4c8RpSSYxzhtONkUzcRG88+wedXrLRYme4xXOpyMSiFMkD4b+zLVIC6T8ltswzna
6Z0hDTps0MfvXbACdFZmizSari6L7xuXCH1AKvYTf0rhbFaZKxhdPViB7AW6sa+QUt7n4SoySSqU
qmDoZ/AVXEV3AwiPM9PmaB0xp/6gpCkJCEwiwP1866R7bertF8Hholr2qOr6mp5Oyf0LlaAKJsSj
H7rdNl/I5xdE38kUv2o+xbTDgZLgF3iA3bKY0SSjHh1MuuJ+UMeRHdSJUoVsMwXbnxGClap6WNB6
H8lvWUqbFNpKBkQKR2jbxmYuelrWgVIh5ql8OFAMWK3SXAU/nKeu1XQsF0qaOhCLFmXl78pg4331
rNB2Pf5+KMHtl16+jgkiMIRGlciPuo7GWSxL/fK+kxmiErJZ/vHEVlu50xsr+BwhQ1kHSiqUSv4S
dI8ocwsEZcYvRt6kOy67PO07RnGulT775xh52VIeJI93B7JkHnqwEaCc2u5r5UlR+IHYc8ARqxK3
JDmmYYx7Kv9wtz1csDBWX8dl+4hI44iAz8aN4H9/cxyCmcOl7D+KuWkL/h7Rv/b7FRkYqQy6cwh4
M6TSxj9nsfbloLBV9zuzY0/n8dWa7P8CcWf1m/C7hrAmQF3OgYm4ilKnIRo/Xeiv0ZmNzdlPU6CY
y8OP4ODtIpyDc3ViXq5ndpaIy/79BcV/QOJ1pfl+xiLabwS8U5CokGG5tGiDp3+ZJajijK/tZpA3
5ySlgmpb5+YNRCKGtKkDUiv7nS3QuMzgFvW+z9q8+BAbqv4jwNScyas7bkymrnVRyievjLTXNbsX
tNB2bwl/zgxvzcX8AxlqjdQKXUNbDQtO+7J6xsCs+JMkTectKjW70ROQTE2SYNqvuAK9FDZ+Tk0/
RjC/TM4rR8wHViWIT6vKXu86ok9WhswgbKhFdO3onPrzpxYfvbmS2S4fijVTkxE+Vh9Ab32tpUzz
FYOIrMZ0DDAi/GB20rELZnLfVh/dU+cwCkDNB/CmvJ9ifbOl+htFMdrxxzqnXkTyoF4CW32rzPOl
5wn89r4N0PNJ5iu4YQwO592gnChdInwbHmUcY18rZreUq2VuSCAssJXaELrCybE5LDdHY+ppgeeg
Az0OPioxoc66UgxXN78vO+iR8GamyjnEpY5TFY07vHYsXbeV5OcETazlNgI8+xKrogx6v1zVj/De
j1u1+x6TjQ1QNhh8Aty1VlnKiYqwFcoTkG3QQjXQIWP54pHvmVyC+mp2HbfcHP2ZKsTi8yo1BgQ2
FBle5hU8HuT8ejomHdVRAnM2Q2IYs8ra5nLhS6qqKB06fXWCrdizS7nGg8RbkPDvQ088wWqVUEhS
BIQxGKjsAqq1AingmgiP6XpSLAZLSIQ1/uymeYejiAn0Ee3sWRUmUSSOVi9MYUphpSBiUNjMzY+m
a1J0WXgz/8Bx87n/HcvJX7mJTm8nv/heDLlqMslfD9+O6MwoubgOHyPECtedkBObpi3QsRtza0MN
nZZE+VRmW7GF87pDhxwHBmd+7bo7+uw4X0dXH5zto/NPcYX1H4St0CI6cKOVfs2AniVHoIQgjjuw
bKW5h27bXCAk+4Fd0ZAmPOJsvvIW/meiM/LXykRbRjgYqek6T8K0h/YYBzGtPK8C3Yfa5Qy/unud
VKbNs4EYMkhuzHUEEIT9QSkrU1Upfi3cGbnSo2IrQNS0WVUgTycWjO2LbMBpYfQ1x0FR9ohlToBG
gLFQQanilV0olR/Jqr2c3TXUrbY2wVRilvtfzvI8GxPD4w27pSaTPJfDty3ScdAUcBX9ejeHtph3
KvWBvFJ4bSDOzkZfyxhVG5G/E9CKbX9s1BWwbznYvIp/ftKbTVKED+F/qgnqScZklT+ZzM9+8N7C
b0wCG7OBFwI/daJuvxCX+A8SUHNszw9FACnTQbEJQtpYvfFnr2pwTzTf/SQAvG9Jsf1hmATCUNM8
0Cmx2UzhOoPOnhs25BurcAHapSsMVyRGer/21/r+Bi8O13b8X7dxuPGaaFIy6qsi92qe/az61kKG
1T41KYzaVZCXFBz15FGlw2SZdGKtQOjgJJKKuzzmCzop1dm9tpARGJ8ZBzra8mJJzxI8s083S8B6
jCsCVwfBzWruRkFMnSONn71g8DT8uLtHWUmTCRzIwOMjoPFYLA5xppne0q9Ze6K6G6Y7O0HANdnR
UDUlYNgN4ptOCwohfjM/iuDuqqJP7zaqr02W1g5NHJuXMwuHS/gXu7DJ98LCAwkIm0SAbfpRkPjj
l89JpXj7U5q+cwTwQlvpiww//9MOxOXQj2HQA1fVkdT5qlv2rTrutXiaYzIH1BjEc8qga5NJ0o9Z
ylemImumCRD8ChL2RcWgb92jJEJ3Zq73jjtCV8E4GfdG2rmq3QE8a09lutmIvB7wzau3/oeQc1EC
rKU1tQKRy+0WGFW5GkIUfMEzsE+nDKkoDgRI+PCbXsxQ7mjrLlZE2qh/7SW7PtOH7HfGPLwTvzVl
sK6K3EpbB8u4J9Sy7AnyKQN7M/V7sIL4x5hLLxYInNFpQckVA6m64DtIp9FftoMHYmX0Gak9tjWf
x/9oJZRxnKpKweQzWR3jgq+9w1EfiPsb6EPC+UG8EYQ9RkjBGGXZZspOi7DUVm365OjXtRzpNsRJ
/UnHKRJDAhsEuz7bjVPUd66NtMuDvUQMIFFC5sdEaCsBz2sa2NGDzCfrpOkHpC58kns+lfLu80pm
PX3YxWLH1Xo7gcwuI2jEmF2daYz3C90z304lh9VXEgNTwlvRC0W/Ohc1FqJAuID+LcP8iaS/DtB9
FeLJWWeGB0n3aA5/JQXCj1AtWg/ix8yZh2uTmoloTe5dmcQOrbOPAzYtk1voEU0pI/cTee0jaWie
ljYw2kamR+OUULed3PCmcnR96C0noKxBEOkBJx2HF7X4mpVMbEpa+cy5/I5CE22ofceW3E401yTw
FSrQvPZbTvsoDJJmFz32LMjdIhLBH+S2mrLfN2zx6eW0qGzBG/Xu/YiL9hGlZVLQKEQIvXIAEoxv
mIbLX1LFXzXUXmfV3FVwN6Nry4c7nshzhuczZfmmuxNHTyJwilwt4jqkjhE28if4/PfdnvbCEOiL
LSLeSjA9gXJ6IEfxnOL40f+ObsFQBVlTgj+b0DM0xQ/rhN1kAVBebqA20kJ4EswRcRvd5ArrFbrW
MRMDVxfNdjKk4U07L79q2YurN1QIulQDuXbkq9I/0prO7x1C3MFpEmw3RKnIFiM/SfwxtNCnxAi4
YslOsasVQNGihKnXB8xLlJmDxrQBrH72OeCbzliWFrz2pLlfNcuB8VKTJgAZEk8JuxXjIzreM9AE
ovT/6URIor8ypmAEcTFPCBlHHZuyyFUtwY24X9hghWet+Jmbp84ma1uJd0wsxjMfbGWBkS4/Znq2
TIr+AQtzLBymzkYe4Z6+UppgWkaqZhpR2xR0CC+F5WhetiQ8RcHr2YCd/Kqazgq3AlnPetnzL2DO
VA8wQjKiCAbodGGYEAhKPfuPFkZoIOV6FYGy3L68i063nvTPHaOB97D4XvbKqwvMKsyw0Cgl3fVD
Z+AcHg7zJSCSZlncMBKD4drLby3EkO0fW3kPPU/+25AlsV2jju63CUOK34ZwtNmgooJlGK1zkfaK
aRMEqAP6ufpKpzcwnlo4vpLNCJy384nQ7U+lLeSiydwNNMO0Xfm33083kXJFR6QbjJDiR0czonTG
IjBkKILDAn83YXHyqkxRUyxI4dxCOUZngTmEhXPQheHFNz0UsV5sLPFxE4z0R8q7Rr3VvXs+yEFf
DD6DSAmgl/11dPv9KxwiMdl8D9XuGwyML2iC65Dr2pO6dgexRhVD5sr2jTudM7nCJmDVnh9Sq25o
I8gOCM9kY3N+KLfK/pGsExMLoNwHyRRije5klZCpKXHnrmX55NJLITBAWPJeuNx6FqZtgtw7/LFL
tgpjtcbRLNKRdGRuhzVfmpAn7VvTchSnIUp74yMvZ6vXRM/JILtYCZ4Hln3869W/g3B39clBqOXy
nE52+W84bKm2NvHr90nx5X0trjjKOq/mV4CfUoDNksBgb8rqjBr+a9hxyG55PyLbvOWA+w0oN4Qh
5Pio04DKTmiHC6+ajeTX+cT8DNl0rY8YxE5j91lpZcx3CirHdqDqktm0rDPeIEsCpw6LQNPGedd5
2QC6A7KhSlVt1hZl7xUD7uuUjvGuuLdABCA9MTX2psLcUEJxnIN7ZMDJ3hau2xxbgb+rXmE4QOxO
7QI/Fs6PL10EcYKdRY52YkYByEi1m/3OSPfJjwUTM/r4VhwFNeLtvXDWKt1ELy/+zcihDy+xwoQJ
dQkjjhtQCyqnIj44AGlE63liDsk/IWLBTRJpd3CUIlnevSFXHDRe1Vzeluqx5+GbQPGUnNe1aacx
nDqmJsOP5Vl+bfH+RJTHSV94sXi/YXfA9yrRCx4z5+Sw2hT1OZo9t7RN1FoevsRb0IWu5awvFkSn
mQTmdYn4x+Ii7eGz77eSUq69jqV/PMlBCS2pUwoiZlcC7spZmD5uzXeKFldTeJqMwJZFLuRDwVd+
0ptWbPdcZmP6HcFc7ltlTuYDdVmFLkBtod5ihbQt1q88xdsY9BxpfK/WhIxBHpSMMbdnPJYrH4vA
w1C/ZjIZ0/Lt7i7JMO/rk1hgxc+OHCKULwyYHIKEfj5Nwhjl0a6gazRdEkFz84lZWuGCSAhFPVl9
6E7o8ISeAp6yVFYRQU4sDc7dNSm1e1TMQA28kX9j68dYe7NCBuUCBEhywfVoB4sH/+ipP9IEP0C7
+EQXnDgREZdiMvLttBFqOpxGyZKP7va82+IHZoueokgRQTGqaPD52nWjLMCT6+gwT8IsjMkJUF+/
UomJN8lABXKyI7wt5kzXOIXruAwrd4zLIBlOiKosaMYU5KDAW7JZGrtLVvpj1EOkLvalShKXyDRN
ObYK1fk5E4D1o5Nvchfsipn7GjONuEhOR4WnVbzaM22rnHu5WEZ3sHYDzi9QSHA19QJ6m1Pb+5lx
FFAqr+caNJe85Pxv55s943JUVWuROn2QvBVqn4ThOBHJkLib+1ouioUoL1RgH/ldaP3gtGcbs0Oh
qC2/2xepl6T0Dc6oDIyjSdf+xrLI2wNFn7zI8ZT4Ka/HfTC0Gg59PdogtXrtEKZRtCH0I6EM7p47
KWwB0DiTSXvcbHk4TPftCyE30BG5izZ5lfgdyHo03Tn074VBqJAxX9VZuNQwap862ksO6vQ9lGNQ
xCXnp7Sj8bmEHDrpVrmhs8+MkOSgCcWo0MQQ8PblRlMst+aRei0Vk3xhNng8gDg5mS9RU5v6GraZ
OJYYI31P8DBE0cYtQbB9vclGr0ArkurFz9B8dTmxcB4bh2vtIPK11NDXuDR2aX/IsZJrOKT/e6nV
/Nr2U/H4hZz27P4Pcq4yivNnlDBkiQzKemVPUWDEbxfhpdVl7UhKCEwjocPaod3nPKxAo/I8Ocoq
N4EOBmcgyhyZndVDGfIlu0qw27reLU5Spv3LndkTuY9l0XhbJnghamTZxo1ThBkFBf4IelsznuYo
QgqAsL4kxUMK6otJA5A0yJAMDbJbDEV+0kmCfPfzfkrxv+Swoa1RvFGDdpzY3h/BzrrH2EsyBjEn
8ohHN4BxafOk3H+DiQvEvr223R42KlH0KkJ3H9YgsgrVgufGfWEkerBtNoLn+xCRfLNeid9F0g6G
pIrqTBwrVzSTo9DzYaTrKFDioaSzJQ4afIthJGa+xdRNpsggj6UG9GijALyimoJPgSsirmLm/Cu0
EbtJ9ZqGL6OpWv81BC7A4+C4monoRIM0N6j5qmH/SzpGVVSFjvwPf0LoOSm/Eq09FGfjPfM0i491
Q7xW1UqzYJEWAG11+XExV0LS28f94h5JJFhKgkFDCxqhq5OL6reOjnvbT0N6v0wKTljX8ZVP9zcB
4nYKQkzhMOfhZaawWsWORWZmz6hkr4AxU/917ndXsVhp3/Tzk5U3lh9VwlSXW2hXbfFlkL5OdzmY
vgNIL0ovLB1uzq2Pwzz+rzeXwxHN2E/apSwykh8FKhgGbY+45Cx/Sf6HLGTt/neDhTFZ5aMoJ+J5
683dYOEg7PIcNFnUP1EE+NXBjQuZ26CaEMNO6oi+rl6UAvgcsuR446bNQnL9y8TiYftGzkQfN7Q0
9qhxnv0ZdsgNuaB5srxdt16tWs3uWrAegFwOpUVnueqD1ML9dkUgxeQm+rY3kmuNetPE2jOj1CS3
FCJ17C9q06ZUYwa554f4LBTuv8elpNrJKcXHEqA1/sk6Ii37HY1AizHeaaGYox4w0ccL/vTCoCSg
y2FzNuYkOqZ7KnQwcvKqe2EylY/RrBtPUIsXlArjzJq+UnrMxl5TJZEymbuHQ6vmAn59Ao96RXC3
Rp/btMaflDx4AV7+a6DkqwZPZsd2V/m8EZ3HllpzkJMUzGhploQ0HPa728yuEX3EXP+sB/RXWQBc
BZLBbaYNFFDJBGo5qmCS3q5n6aEhswHUCS92ejnXx59MD64gdeBNEDeOWr1Pv7RbC7EijQfDLvgU
iB28AdaiDBAj+A+PIHi8+hgHwhUzCV/HPwUatcBo8ZYj4gWZsr1n7Kqy/95VnWf8+xNGdb/BWswS
rxJ5QSuG1++l7BFXyRRJdBmXsacHzrUeIsKytWhvgt/J2oQi6N+hwRBEmg6An9H9QPAw8eXegeZ0
X5s9w6GYa3R/ER191+4PkTgA98NwiuwHWghxzRjWEk8Y0GoGjYe2EOjeUtzyNu1omBEzskJcoVn2
u8TlM3NxFPWimXxpyLuFp+/G0l0LndHKoyI/dMohM3wSLb0AQ13MAFPrM+hb5MVeIUE6e5QTsaJD
Sye4HO8J4RShVq2yQPGvNJNwcZEBShSeJrVAzstTNBz5E2q7B0+IfaLLfSLRxcqFQnmcmIJ/aaov
A0w/qa6kjJfc2i1XISuiAudj+D/aB+QHN6yDN3UITKUtqhxjEBw9dYBbjk7yhurcrv2X9W/5YCHu
qfyH2yCeIXVzx6X6Kw69qt2yKiaxRhM9sXi0XScYjt13DNH2Kp2jkebPx37YMqNjGqbVw9tddU7Q
eNbkHWSXWCxisjxq8e5JcRYOtYu50SQci/K7QFBEZuSKinJvjWFJjIrOS1Ed6jqTLKZ2ylgXNxJ7
4Zh+g4rjb48RBYIFmSwBnf5zioFiNBY5xfgrr4ivqIuWkSP/5TskztVXuBmhDFgWUGTasJ+mjvFV
fwdXN3r3wgkkcwKiWb4cvl+tVyYeUueZwmzopV8wVD74P3pl/DMg1vTtB6XTpGbxmJBzdRL5Rlpg
Vx6umtnWE+4jb//GTuBgVIQEOmHzKkJwlX4jlJh3/m4ZLtyNe6w9a01aBO+iuqXbMFqiFdypMVm9
p0S6TSXArvKWMYkuOVxYNT7L3zoCw/XvfTpeQS7kgGvoT9woqbiD3RFLkRP1Cbtw8duubKiN9VIt
+iorXJ+Ve4ZBdQv2stHc4eDDWaDFVM7NGiY3RCZSyKTtkzqfkSBkMU5KfY23D0cV95wcmarQbjYu
eoH+l96pqqC/3KKkmFaO9jK8NBs27sWzJnZgQglEVVDHBRdfEK9oxQMIFagUKh5rqhiAdImOr0lL
DlSLLpyMKK3dilVB9+eD2woTVPlRxeSyxfhhumOFdBslliLmhbUTqhq8MMs+cU6FbuHrIBliXSz5
PZfA+fh3KTDhMSR4HpLyuqZGQd13KAaxKVxe8ANGMRa/vJIOVq/cIPa3aZ2isqv3qfb9HzC0yPwF
mzkxt3aYl2p4iC2xCBNgd36O+wjQquchzmbMilkaXxuc8lCB/OeeNzji/LU5hjw0Zohi4cLGJSPF
YEUIV0B0WXvGGDyNGhFgvNkYBs9V3B3DGSykXOu0kar3kSZY68FjXGiYuWhc8Urwps5HQ8sDCwLy
8/LEGLQXFejL8WfIqp/1s2JLopjE98QwbYwuoOLSeCeGqS21SYJfNVC1xfsckxqajuyDdYnPBq/j
x0pKkzyFwS2YgXOCvIe5Uvbj8Ls/ZF1ntGxyZL+toW/jdFxPFCZvo5xGvAg/1ykG3FTcyY2PONsT
JGJltCbwDAYg5DlpB1gplVHeq24Q5pTZVu9aMqGqGgZT09hxVPmGymNZRvQELSLkrEI2TYRTj2/n
eJqTUGzLCQyKEgDSiR31bNT1CwobZL7oxfamnYbh4RWLn9GIUeLlmQDZ0xGPpamiLFhvq5vzd5mK
Fzd9HiExcteJB57pYvYLtBlMUZ/2yENqjaNDVUYT8zR+K8JSee51G8//FnodgFUeLOxMfc2elP7K
/RDakgj7tC+0mTPxHpMmfrDhQt0uZTEDWFHYFk+GVciy/PxRwhJr3k/za64LqLwNLKghaHqoWk+J
x/dqtcxJkfFLyy9nccaWvurrNaTCV+/ux8dSRmcNQ+essAh8t5V5BF67mr6PdxRUSUncsPGTJNpO
BRNkRks+eDCAK1s/dI/l6sU4QtKSwu0thXaTKCp2VFmgIlq7LcED0sT1ou2VbTNzK2S4Wk605OyE
d3S2sfduVYRsUQ8V4hPbo8KDLS3pvKf4GP5xqRD/GyTLUTDoetYh82BHzUlZdOzwp8ffY5+/xakS
te9Q0U0E1jEPwRIGqc7XMTVhtCyoJLg+4ON338Lstmlw7nQSfHxsGHPv2g3MJ/tDCK+ctGP/D5ar
6CKK1TQSrO1x5khVQqiKm/FMNcnIirrBfwp9vhhLpIgk2yWJRSNXtv2B4lAf0Pz64NvOcwfS2Lz4
PUaGaAsynvUO2iMdmmqmT5PWwT53TBKq/WaiFqOeTp0U/MLNfdvEU1bul5WZ2BWz2B8LgROqdkpO
uRuUuPJusN2YtdNyFajRcaZzPuvU8e5zJ88Olpo2TKpHsNb3inWIQ5X41clvqC05/y/rlQmy43Vj
XS9FGYPmydiE+CmFK+7GpX/5IhcSTOJVwh4kpVPLtTnt/ZufRi2mGHw+B7KQjUp1G6+NC+nEMsjg
ARK3XEXNlkjReeZ4RrZ1TW7eBChYwG9Z2pazK7nM8rgeLGRgUHZ92wIXey0iLA2LKa6S3z44bDQZ
V8U2K5FciqxhQ0QaUAYiqttxY51RzhOfb8hLFWht2rxSZO65JEWH8NoxAvTdPicBlXFT5Vi38hqa
456j7s1A8JmWhuHxzp0wQAjopatphx2Akz8bOpAiBoIe7PqipqaN+5zZuSTlXRTJq9wwluphlvfo
dcuckaq5xdj/shHlbpVXeZAVgYPOADDgITfVwmYTFMouL38xEIt7Lnxr9XiWWjgi0KEUVTUy5Td2
SUQ7ubbV49NvxVFDbwkO+9mFpIFCfgzIHwweIeu4d6YMKtFl0EsZeWVEd20g9dIsXzTBos5dr6Uk
xc6gks/7w/lYZNz+OKEvwb0zgoyhX4QluOt8eFl5dOST4VkPUPFxXTCn0Ue6YXbo/ljL9EEjaGZC
SGb8clGzJ0z7telbBYSCl3OKpjQJfiN3bSEh5np8xzE82li7kkvaQKka4i5uzLnZxxWl3E70Xg4L
yehzE/pw2oDl9asp++hxITLOe+hFHn3qiuLlSJ6yM8Eoy84mWa5YNN1BH2u95xJjQfXcmCkiEl2Z
/ny3OzUki9oY7fDBtbAV8aTLCBcRs9xZt9DScoTZk5LlouPg7pYW9WwT56DB4O5T7D0066MFy4WG
X5OmIOZgyGWbqI7vhYyW/ifXrYF2RiBRIhAWe/nJo6qnvTPVzdrF5RmdYoBvR2R78aGd2VDS/RoT
BGgEaFUY4sZfl59Tsos0GK53CJAir0Qz+2jHJkdqSgqlnq2gpcTuQJu3FlZUVB/g7R7MeRVx7Ozf
DwgzqWNsEVuurwZIHkJEVzDHFlyjlLcj/Ch7KnyrE8D9OLMyNlcUXxuqvw3IJAXBKbDokyxy8bVA
2OBNoT3KqGZq2MsXkdiHlfWraPH9vOaDIFJw7WgiGieER7yCnjJfqsLQmZyTtIBaQBYPzlPerpei
l2D/ytzOxhQ3Ch+BOuMr24HlaBkc1BEGeONxuyICnCn32KVcq71jjqRpRXEt7JaH53rFNk8w3tWJ
CiKEKm0k7tUJB3vz3v/cmYUpLXHUJvy72V2xi1usDAdegtJ/hNR/2xcOVO64uoMQUyz1v5oRAQaA
5vO/c/HaXMFYh4iFwaDky3cPD5azhPdkFOWdi45V1ykZvpwkwX4TOxbB5iFKBpb2YmDV3plwAN2C
NJC1u/jtjnheI3hFzAaqw7ccQ6Lgkap7eZgz/JWIAQ7e/SCvAO0fuRF4OcUpD+dudi4KXl0eFqQx
JQX30bUgcrepk0SVPtdas/LhUIaBEVsXHxnKR6SJABNQIbCCZJuWrTuExiWTZ2Z4rSOvqj+JzCH7
a4DQ0dyaOFK8YQk7oh1+haJtA+RgA/PvJDO8c9eA01hO59Qb/jcSgxSYkw7GZulBNoiaoYToQbCx
lLjPFw3o2xMdr6C4xubj/cbwnFkReqsGLDjVhGdysBDz30g9lU4l0ohoLD5MM/DFr6GW0ema/VSp
0QmvBbtPKbx7+EttXBYGTZ/AsjL7Ot2G83qW3oZcLufesoOuuIhp1qS78Y5OHtEjf03Hm79/oaQm
4yflHPUsohl7cbs05QEF8vVI6RYpKMPab3QHS8l5uhxzzHVsjiIG5dcH3hh5gzgHU/ZrhB8McQQW
D+tP9p+z+pyObOtvCsLm6KdyBF+vXQO/y8qL3Q1/K4JkWsSHRwuRpwv+e0/+x0QD+VcO7baDLQSe
BzvCqbTsCo+VubVutnAPw95QX1W5sU4CE4cC7xja7ud8L6gu8DncyjWufyhSmzq5nVdAQKzHL65R
3tMNSNOouzed+GJHpXzrkjuYoz19EARFFXt5l63OQdS2WzSsGMrcOJnlHLj6fVw4YtdiLEOEi+K9
058dYyDK2W6CecN2uYHu/5vjgz4KH3ad3dgqUX/bv5Zhdhxt3vC1Ho4axjT7s3Up2dHXkW7sQcR7
BshKiYv0cDUrunPpfRdOXv2yFWE3CN0BcqDVXhQNwoe/RK46H/LN3Fc/hi9bQB743/zM6GY6DPcJ
wm3igdJ9gYofYUiV6OjHLQbcdTyTdhlEjw7GhlRh1Di4zOLSS4x+Dvtzd9bsI5ZROof8c0cqqlld
XQ50DpLxd/lUkE1iN4dXPn3mJTGi4ujfuw5jVv7G8lbdbvE/uY2Z/z3a8ZECakeynZ2GwlvT3Vez
dEF3z9rUpwSEtcHUXHWkg8KIM9X3+gtzBRhnpKLHY1fjKInx+t0cYuym/jIaajsLYFp9RPKRUx6t
ztN5jKkdw7j/2RWRx/Xde2yjZ7KMofmO3oK+L5rJmbl01JO7eXonf65w9YAbNNM3/w/jn4VWl0tA
pd2nYuE46ZuMe2FHAJUEgWPcNHzrcXZefnTKxljZamW55hy8cJz399sRqr+djQRXFF54CttyBE9L
lhbpuSfwsfZV8XG1dtyeEPWq3FW4QmdfC3eoHNt7HYW9/3olvRRB51MvDNrXH1Uztf+SW0at5hYt
ZX+WidHBifQ4+/hqd/+IpKKx1eUmbriliSaQ7IX08NynVwdLWMDwtbjKqS+k8iYFTopw0YXO5ymm
x/iH6vrAFLxw3563bWysiA+X+fWBD8aIZqjZqFTtALRlyzFMJuz9weqrMcG0F8c9UBEobK4oM8JP
Er6XkPRjd83PjeYdMGqRF0/lXSAgep/Sm3yI5FLpCCV+MFwnXfI47KBN7KHZ2tM/L1bDq2SKC+St
mAu/I+NfS7q+uDd+G1rYDMm5O0ps7wnoLBWz/KzYyoBinyaFMJENdEpuM9W+R7TcSH7gEg2OqK+P
CECvhsDWp+7ONhSQxdnRglBPprjnTO+z/6tPCCc9uZmENM/jLZ19I2dRc5fufytBf8c6w6OIzH5x
LWjJqENxM+94HYhQIhuq790wRTNf8PnT0/BtlBidN2lS2leXMf25f1grY6z8cDlCyheHmRq9hACq
VRj3r0FX6FOLxGsdoiYwOJfef3urfUau07p3dEc9H+EmycDfkMdsvkwyBLuzVSJNTXyDqBZyOSIk
I3CXxTUVf+87hCP9NBRBi1E9HBWPja9sD4oE3+TXSLWC7S2nR1YisfFRw1PEjJllbvl35VJaxWoq
DyINLH80oIr8W+8IX0GtE7MhkdzrBC6ljxvRLk0KoO3UNrqX+RJN7MxMGw6wMnLMBqIGLqyOcPZI
5QpBKJG5tH0KRUGtI10GViedEm1cW85SeDm4oI8L6kKTsWz/esfpNpWYKVcDUzPjHy4KhHBk/e6o
qpqn+avvjxHkD2pCkxNxjURjwn4Lw9GBoL/bUG0eDm0HOfgdMx6Lph8F2zCEa/UBr0NbWKgdYpvf
MLQnIAKdLXPp5wBbQFG1qJCAzZDIKWz2RMOKASd3TGwQ+oq0jGPq2hgSgGyu66mjvZgDPuGuqwsu
d5JpRPUlYeMDnlkv3i9Fg70MU31KFn5JIuIAhQM0xvGKnlJbtJeWqbLCQBUarKRZKZUcxy25tQIU
SLAw/jzNnbmt1vUDOxDS5EnCmEvgqWs5T/yedcICz70GwBk512MD05FRTLT2v5d/et9XqZ2vqfvN
KNWUS7E73PdBQaukaEwqhi4W9PeRr0IGLyHsuw57s8xAOyyqpxPulGHBJNpIBfrE4GNCLwvSXPXb
N5AW4nWbidtgd8yFiushd5D5eSTp+y4Y0xEtAiX8HyzT4G9WDLiwgv68yeHXZVETUu+eCxLM1N/A
Qp9DstsKwqIsv9hY0DItZjWFgvlpD6Bil7dYBEyI+zsN3Ls66FmCd1otiiITcKAco5kApIhT9RpW
XDpfDUtpQM5fMrE90NYBUslxz+o1udJ+h6edz2J+q3rpVRI3eoE4clsn69bfpaPJEgS4ZJ5+bhi9
JZag583ISDctF7ERg4+UaLveK4BMrKAqHafOEfchIUM/DYiMY2ZLOYBFd/u7YjwY17JMY9mttJoW
D0JlxzmQrMjMh+N/hCzrbDq+WQuOTRjSHkFn6dhf+hcn1So4JZUJxH7G7fgKUCw5xMIS6CvGcmw2
WV1rM7rO5yqn26ZQzAZ9KCKMFkOwh2kMUas0rDsZlAblA6llrk6mCxsI3B1u9mN9EdADFshV/V5L
2RTvxd2dTyBuRQrmCrhzS8MMTWhXeD7W+d+/6McTg9DnjOY7lZRaxw6GFE56Y+7GhPoFsDOua5UF
jKag0xdilepNYGfvudIxDg8Myt9Us14029wmElJVtRYMqiWkT1GJdlMY3NkeGhsrfOmluC3mYmpo
teYBvOsFHaJkco0wlU+jRqH+Nuk31XPVWziMtFVnVLtWQdfp8w+Lv/rDFI9SMK9DUHKZQlFAippx
R+5+kT1JWQHmtIt/kb2eMDD0tyK9ZsJ/qsxobrry5JfyQIWFMsjpIB/c57mgnK210Qiw6bRrlBfi
3Rcd//cfSU5Yf4WitaUyVqk09UTP0+uykn4o/88GYQ4d/X+SvPeLXbng6kDVfex2tfmtS/slK/UQ
2p0uFdIWNFDlLUvVV+NLvPIehoZa3fu5isBz+cmaprWDhoNzT3hW97GZtSn69bCwYtMKBRil5V/h
rUnzwh9EXRJtQAVou91yB/Pv5leKh09Bn9xJgU0Ui3nbafi/D7sdMTZQchEzGiB+GiADoHruO0tR
uPtJjLMMotxDqm0jxH4n/GHLIHAXbGjw02al20EXZkcgO+dtY2eKPOOohvwcxnHndaQlI4PsxnhL
8kV0vMNB1EQVHU0ENmOcGPX4qs3nHYgf8nFlBADCr2WvDdIEUR0tgKPRK3NIOWSeya6rnarftjU4
qOdCM0BCo7nDJoQkO5ql8ryyNVr6T6D0V4oE77vFPRW5mOjV8FrX/BGXspYx2xIWbJc1XKhWi/2+
V8KtDR8Xth9mQLfgEV26SFrxn0MYd+v007TvybFVe1OfKPBwqVuodprB9GfZu6JTzI1bk6cAjt7k
G5U+5SMjUQO5xzXs/Em1lW7Av6WDZ6lh8Uwwzdp4y2TxHvuQKr0Ygp8ZKW2QLRZqTZCg0WaSIrAP
QgrrM3tN9PCcJnzlhdbK2ESNp+dUqI6PNItf0R4RqAz7b2Od8qY6B90t/s4QlAzvk9ExyWV2kjEu
PCEDNBPEYUzE0sOSgvTZ9GTN9sNI+jkekWRAjF1rfUhvcg5dohi0v2PRz8VuXz0p96SnC6AGiBhE
2Qjh9JAkETWOjax0yID7LimrQL56hAbD0uZJSMyszUSiV/fzOX6Qx7Cy9wqtUhNygv0CoLHLeRhi
x7UaEhPVKxQtGp9vwdptDvmjYtz9k5giC6A5ldX4y0JBNr648WwM7TzHXnBuMFm6VPhm5oj+Wkvy
nwPEvHfaMgYF0XoqPxkfxW8ZH60/QBzEq+zuF/nUUZH9o6JdE49XeBu7M3rr4cypHV43YTypVuSu
HeNYApewCjLHhQEevB5DAUhBA1q1Nb+S3iYCdOQ24MnWcIKDaByURCbxdEOo9dCXY83BGNJgfFt1
s/oBiVXq3nLfqknEl3OREmQdacyUsw7/GHvaAFu8HfBfT5i82dB5gRAbMo5HwfreOB84j5kiiavs
a22zL2spg+JTpyxmFEjyNbA+TnZZhC2b634cRetObJ0Ml1zCRh3BtbPqj68FyPRwrZ6WqtbN6HiC
EBZclD3NlxisVR82DgWsWIltQIt7h2loB6Tx6c3gZErDGYFekMNrofJAl9wjWVlSnkwy5YsIct4q
/kkHj7EWTqluSPNVxkIyLDLANa4W8oBrCgy3d4QbzMZFqyS3w+XRDJDY4ezUXXe3/pN9pSCPjb43
PcKqk7xWp4xjTshL4znOYrQ8ht/w/C763CRtGo3wTbUrot2DkSOSK7xacDUJexMXrk50H2unF1/4
+soIdBOYFbs+1Y8xeg8M40dM52WAbJXMfg75+V/oxEeKe9VlJBEtadrElE6lSmajiqhz6urf6upF
T10HmfHDN0/svbssS7UfudoFVvDtc2tmZYpLpjxuCJXZXCCgwP1ssp/AyCuHJ2D3o164Lh7UTbfX
IwQp9wo8Yo3HvU0VNaGv5gtPegjdcDph7wV9W3eaVS6TlVjHI8Ti1DhMfaEq93tQ4pTi1tQrlz1t
0fOOHtglQC/ltsFkl9soUCcUBT7asnnn64zIwb2pEcf2JZXqw47HoXl2ZI9dL5XH3vojmMn3tzmk
zAuRPUeidB1AZNy2YUxuM59f9A9eU4mJu86fooXXEWZb3HzUyC/RourY+nDgEzGPtSHaOy9A4MpF
Ev0xQ1ZHWplFiOHE9TmpVShBKcLWD4rYg+2I0v+PGnhgs+0l7eG57pNu0HmzgUnSOc01yo4dCof2
1Itq7YdLmOStiVnzD2hJ3OmIIG6dd3KRiw5/FPFRF5rnwM0l7mqo8quUoOheC/NoutOdT/YACs6F
9HCuF2OltcokfOnmPRuwpLBS+2d4VSn6Ve6LWQ/qpCrzoPRVE3H9e7+OlY3XpFSrhxDtiqR+mnub
CTcIVv877EcbmnS/xH5jvMINBElYHd1fe+YScSdzF4EXGEyKbTj0IlCJK+GaTfSPQo8rIksJlqM1
r/V/41m5FDjTo1BfsdxryRFIRLPUuMST5G7e8OXCqQyv8p9O/CLfenB+zsKXKmAE5RHdQ8Rv6Uk+
65jsrjDvFFL8xfU6uUx9m3/EkBLy0/EMAmeg/BD7lTJy2BBsnE8bZHy8mR5b+ztYwlK3ottooyal
R+RRZWzurn/i9ItmA1SIAoD+pW3GrbQWU1nsCocncPXvibnnhuexEpF41fQb1Tg90SVKBN/QTrEU
/YL9eP/SbaPN8M1wjhqiCR3iDNvUTI44q8Lg/7pI/z0IFLz9BYguWITVeHjH8FE/SFILRkZ+O7Gc
tIETrnLLX8WpA4vV3DtvTJ4vvt6/x1RpkROYvXvqZKRw3jRdp8IQrB+CtBq/LTwsXFqxZHz7hh5X
KavafG0qD9Cf/djkkqDuMy2K7nvS+HvSAtiboM1rcfBCgmtFquFCB21vcDIGdf4Qc5v6ekBjTpx2
IpqZM76gLfUOBvcTHNIG2ZYUK7rPAe8qweFkJDxumqqfQP5IiXfvRQi5kd+ob5uKkDL9uBQSJciX
KaANgk4YQLhnBwzflI9piN88nyl/QfHcjaOekM3pLX+HU88LBYHHf1t738gPthGYJ26WNvcMZ83w
rSNlXY3lKnwoSS4FaRLXg5le8bniaEIgkIGXNC3FeCWd1UC1Np+OQ+JnOFGhNRQpLxVwYFqyLzKV
LG2hyUvsqtKpSAnfgc1rPvopQqAfS9AIvN5BjmpqHezQWMoZy/dka5LvHUvrTuYFX5B1X3H2Pov7
+d2KTdPnEUjvp+A3afCED3uNCbsFdECkgt5OyFQRu5c+SYbxWN0EJq9nIJBeOb0Oq2XMAFxw1Bw5
YhOCeYhHHlkqEPRgmxw8tACiM7yXztpIR4mQzLxty6aQ7SWf/pB8pYVuD4rhLpIQKeY7GxTAwMMh
1djcB/zalX/Trgpa0yXdVMuhQfU97aT0QQ29OGIBcDhQoIH6j7mXYfdPXywYGUOsr1Di0eLSgobR
P7QKpgCGGsWG31mOof1dOM4B9HlMBqXuqcNfhIXCbiCCllnuy+cHe4Cq93LRRmRRhiIF6WQjMqjO
fFHEd7/kFIg7gAlC3kzWRa9jJR+QnnADI5htQVOWHKPQiNT2OK0/r5ViRS/vAY+tTKBjzo9EXG03
Ancqa6zCLn+ZUAker06hnxC1cNVMx/gF0aurhKk9ZsEjtt/TnYApD4neIgP57r2erL3Y3qCeWqot
YubMXpjyQVzh0J5lmo/WJXoHd4sXSl8swL95pT7EAVqYMkf10yjPhiHUKC+tQYdvbnkrd/A/DCAA
lZGPXFNmOHAgDkA1Egcbt1z0NyM79tiIzQLOT9ZghMtOGocyDlWyRjUpVdK9KNtGWi90kmAUIqUF
vml25Z5z1K5fqvtHP7X9Bh5PyYbGnxx5vNYfSlwfaqDqx4T36o8AQKGmHtusv65h0BTMHJB/p5DF
jeJqTihhnGvbnMDPuXxv5Dut5/Olc0apTIPuXq8WsUwrXnCkEaChZbnOwOlDkAelgDZzg9NSTtEe
zhVXNd2r1I+kTKB7zuOpM1wHN2avSd215FlPbMCyEx6H+o36x2EOhK0K3EQtysrGEyW0hAn4qaYo
XtoK5L6HpapmgGMirnck7fqi4OXe555EaRvWDeyYaqHc3vf1Ri7IAufC2jlfAkOVQd2Dj9As8pUF
QWlha3BrABnSJJoCB5c05PhcMfcK+ObV1e72sHr/+IUvdjXANhB2AcP6xY5O0BWft2hV76BhcWY3
7EbMBjkQ90lmK6XkhJcabyRVAh561CZStYz9AmRoGUdYlyYYrYbar/TO9q9hWusUezZ9P9s3eEte
y7PHoZvVD5lk0F0M94PH1YSevLU2R6E9WUcfE4BCle2TuYJ97FYdLHqP1DodRdaSFecW5nU9531H
PUOIkDtdgaQph4AMGwF75IkMUuUJMk34N3CMvrtbzgLF9FpiNCl/uRVhj6ukcTW4J4BuU/IpCbz+
IEj21ZTaQ/6N2in8t4r/UrnNVVLtoBpSL+obNkW0bYoRaOV4hCniBJn4DEDyURAnSqNbpwkGmSWR
1na2gjOE7rqQpXnmSIc2OL707Uvrcn2m7Qonzv88rh7caPs2jwFE05YkIjEqp4nFU4WipP1xUbWr
G6WtSMg7/vi/dgeOLT0fWUaVUUiACWQDryRrI2HMcBpuTKLEQcFMkVW6ycH1mZXgv/bAJv5jTnGE
HC+hRSfkzadcmubAq8r8+C0s6+8foXVl+lJuyFip01d0KRmmtcJBfiGuwtLvV3CmkDoFD6auhD0+
vp87gR84gQGXOAEF9TJJUwFgVhDFpbI2jmNiUQcAfjOv9qt5ywcarrdp1QMkaD63hz4bu76D4e2w
eD/mqz9j7V7hiUulpj8vrQ5zRNJcgAOVM/XehlXantcH8TQbl5TA//uATsQkiS9f6JyxTeJT4oqe
FZUnGDCrbGl0VcH/XozA/m3XKNs1YAoEZjXgemQBT7HfdlyL64CO2Q+loR/qTGo2vHfiLkvoBK+X
n2AVN0qBGOnvwoiQCIi7G2vmJyDg75lJM1WiEjrbYnJYqZCdTa9i7Sht+kZjnkOBWYDV27WoOa3C
LEeBa0+NZj5dNjWWbQFhjLGCMwkfVcF/gYoobBBENWJAaozQio91bGsUvTE4BkXnpvj13IQYdqKC
o/MZdhPcEDXM8FUtRikjy5kj4Eccz3kR6iFT80/Z1rS/czdXJCrpXY7lZohJg7EW5JOwMVRgppZl
Z3rJd3xIG5nwQqu3/zPw2q6SEIM9wDR9knbz2zAjHsEDY355ZkazKor+QbQBzLQbWCp9ISiSupiK
3m5RQVzjCMA5rH05W7CdDQE2goGUlW+u8i/6OOtsGijxAln9mklQGf0BF/0QduiBRgYv3cX5dSpp
E66AfmEg3lPzJPlewDjrkUrGuf5b/NDBfWgA3SQJp7VSAynzkTh2ecnvE0nBJ+A6ey4vQyR5vq2O
d2QAvCy26XV8gj9L3cZwGsexcJ2eXniAxO5KH7gtMbiKUOzwJ5vf/aYCBpu8PnVzNZiuhWr/EHTc
yYMfOIZ4Z3KNip1xbTbSjoVZQ0pF9GlZJwpHmmvmToKlDkUTrR4AB/5syPS+qCK9BlogQuz/v+3/
irCEM0Up9Vm8TgeLT+d7zX2UFvTkVX0feSaN65oe1VP32r1gcD4dmjZFwVIeDXYN6MnSfazG45Pk
0oWx+BgHR5xBsASHcWJvU/zlhKDulqX593OyasJJyKLiCBI+OX1LOPImkwptiPlnoqMPsFDHIB6T
PKUaM0oZPWYjI1WKmw+F3LFyEYXTu7WWJhBmdV/L6OgCJ1LqHkxURN2/AcqNEYhkIESOYtM1tUBU
Pd29VTErLM7OjqAkjBD1+mFuLKtU6O3gx+sJIVi67EzfKmd/nwfZWYVC/oxeADoyeh1dG1vP5tHH
xubpIAssxyDMbjmCSIgRMbI3z+PBTPRcKqGpfKPwBWipPNsbVkx+2QBFEOJs1idnkcwhzDidNdLi
Tzlhq2j8Y1EcwZmBwmZhd2DT41FcXFNVutyBg2TfpHE4fV0ajsVwmdHd9wNMSfXffFdr8+OGkIQu
2EWrd1sC7yt9TgHStTOtxlHGNUo06q5fMjvKl2H/PDFZyQ1At13bGWAFkXs4JCL/iCWF8pZ+f55E
qdhaVohZYbQwKfuyfYdXCM27iXW4oVh5SomF2JG6914Avg06cpToa/NcRIqKDledPYtZFjDXcfM5
fhThu8EBkX/nDPLa9hZu9zjnXWZ6aYqK6Vh+ujVPfj6f78XuBQ+how3e+pSBtFysC3F2sa54DQTa
F89YH2RJSqHg1eYI4P4TkJXWB3zCtSgOWzOpp4jaxLHQ8JLKx7bE3QecFNJS03HwKa+0adN50mWz
5GUXdpKH24oWv1oqvkNtP7JploQ00zwVyTW8qF5Q8lu6UqpgYEPvKIRgBZ9Z4ixrXUsvRvxsBVI3
vbMo7CvIcgMcoJkFMEpf7SEFhcccCQl1UwPz4/+A9R05Pqy+cQVDL9Q1/JiSG33F/dOatn1AE1+f
/s5MlH7gG1KN4jNmFsZV8jk5+PKJCZkihuj0hTcyM6q/ISh832CPuQUGV1LbBIg/fhtzywEWjS8x
R16EbUndVwGenj309Q4s6CCa2s2wJZ/w0DU9S73iiTaQb6HPA0uS+cDaPlikYVNAv4JlaKgzS7xR
Ltu2uO7taBuCLK1yAUZI40fng+qPkpexiSoIenA+mHq7QLk7vait/pDvqft2qp8mBjmfyijC5REV
cg6mV9tHxTwnl54R17jlAzCijXV2DipjeLFku6QU5Tnd1yShUFBaZlizKYa9Lq+ZdBtJfchGSn6i
VCKuG6pz/5Man09R47kv71Dd7/xV3MaDgwRspsgb4xISX0+22XHiOF1/weYE0dSxOQv9EZXDvErK
vjIQTGVm36hw9dlwe6fk/Gx1SIBnxsp1aQrQwQV7JCVJLx2WxrHY/x4rYMSsVFzmiG/oLjhkLWm+
2EcUkZMcboctLdGgGYWZtbqjt4HhMlGewnUgjZaFoHQ1uvJoCUWIP+GwIeettY+7y83jKxZMwqIJ
XARDesv3e7vYNzZs0EgfE9QWEXNXfhr+Hm7MLpZSVr9inlAdq5UeWsc39oA18u4MTM46Gyz3Fhf9
EkXVt+2HLw0hIuM/vKhhydEED5GH/LyTEJQvgzau8EuP0nkF/mY9g6VjVEdWJLcn6ZqFm9xqGbuw
bF9ugNWLmsud5fWR8XHEoon0fuua9DCZPmD3uUlFEMNTPFSPROPYXHFkcOKJYXxLAOqBwiHgX7aG
FcwpEutslSuTFhaQWWyhaHt2Jdr409DnKXXSQYpKIeHiEe+RmsFynQ5WAf/xklwDj/dcp1G3AVCJ
EStVFQVwyAZWE1Ssgepu9LXN2OxkdKsrswY7Xn03MVZ+LLieQzpfynRLcjYKjWE1gRdzx8cwbxgb
PFEK4IaE12tHkidyfKvA9ZLbRK57SXgk9jjTI4OGIjDBb0PWubhVoybzE+OWCrkjpAOwrcIJ8hz6
JBCXMNt1DsEAs/iLlqrMgvP7530BuAODAk5Pkl2TKA1KRQk9ehgryfWxmG3oBEQN1thbTqKiMbQL
h8AMq0/UYJq8PXo1+ju5v81ZHnCDcvdbe7TYqt0oh4ogOTl4LUYc0pNaz9zI2Pst137lWyN38/cv
AJNM5eI2YVzNNAfzDAnGelTAGmpXvb4a1BTdhtaGWxiBVvqQb+AbpfK4UpSA0GNSKnYQt3krWXHC
p9uWg+OpYxx/ECbR5rzzMnSZTKDPiEjGxJ9aXOzD7KmKgACf+MJueB4tlgc5NIv29aDzLMSJgi5a
FsfHqM8vbUr00LM005UvohRkz5R6raZRE7362iSGRkZscBPcjMFYJ41ppCMgOk3sIXB8w4Z/Qr80
6mfick0IUSlYxvl5ejcYoF8hFRm4W4TJ+KVZDZYIuoA5lrvbiI7ReHAtvHCW+9oO9pzO4Q/xAyJ2
fDu+fGzowxebHgo7Bth24g0lWS6EAHcUzbXhroMk5YE/AiynMH5h1BVEqHGt4xpH5bJMpgdMNH0n
WCos4mKCUPEzAlD6WR4reJPMDI37/co4e75UnYE8MIUjOhF63ZK4ClC7DM6l283rr2dWr09PMhaA
06CiQaN098s8DUA/0+i9BK9SNaSKvfn5A9NrVWEApS/WChb8VQFIN7zJuUrhL5emYlhts0b7e6TT
mvDLQVVUKfKhG8KhXNXrFMULCT4ZvoUbbNkI0DO+dVzrrFn33zMIHnfiltSoBl1MYGffxvKU92vN
3htyPyBk0oKi5cYbual0ZcU2GkNYwvtQPcseVplXZd3RRDB73htKUt/cdPzcqAawEP6iibQCMDWJ
DGhKIwG5F3vPA1C0v7+076ZSE9aeEopiTOsg9mjbSYWvn6HwX18xghk6zI6Pk1qEA3XnTYfpegHP
q313fLuhCCPeIbcH8fKmvmi6oRtj8/w7PWvC0t5vUc+LBWknVRfu9PWEFJyxley7oaRlFiI23lxk
IqsXe3DaGyamUUUfsWIZ+UaDW3oaQ3r3Nf8Ad8JX1cmVuhxxKGB4n3UnFCk14+7CIyBXhCS/EXM5
5FwamXXwKkR9nPbz/FQqbWmIhK7AmfQbUDob39bjk0unhZmIXmI/JT++c3QNhkFpUrK8FZSGTTBL
pCVwyIcdRn7Z9isc/fTY46dqzwHxm8O0VFW9RL3IeUiw/aMV+4o9lGecn4AcuWtvzumM/soGP+H1
cvSzSZebexEum78SLaTGzw7+IGeGW1n8lTnfUk9FfDE6tDugr/TSClDk9/vAqj0rZzOC1wqprKnm
Om+I+cFuqJoH8dtnFeU+WxlDePzeO0DPScIFDUQCqWl/DU4Ct8UcdMDJ2wJvKNJHygOKSzzJEmry
4WAnhgRuXExDNJSocmE4fYxrGrUuBTdRGeB38Fvdru7+43e2bHzJ8RWjFMGRP9jMZ8xuuc7SKPZ7
/EXXyCvJHHjfmYJUSoMXMargtNHcDQwkBh6BGdOXvOYynX5dcw5mcHiSmIkSxisP5uVGHicagesh
qo0D53iH2uNTJaFk6Lgl58d6bzHnQVBaYy7NRf3O2eVocwlwUA/bci3Zb9h2tBl92lCEn0qWaDS1
1WUqKOEy53J8rQwMXrFXYwbHyiA3WR3HYDbu2anMBa8YX9yrPzZByX1VKrj60v+qXAFNtt7s1Nnv
COha5poiyWlj805gDJDOM0JMIEBceNvy+8kOsNbVuFoh+8+Wd2DSZxsLPvD+VQMHyGcH82lpzqFG
rkf95j4sujE2mIUbyxSjq0lVwCmqgUU9lLjtGDsU+XkWptW+1CbUlrOxlPcU/HlzYEJkcWTCCoHV
MaJ8mfL0cOH6sBhf7NswW+VrYR398ukI/ekAvXiAvDrlvGO5KADg9N3EWt76MBKIY00IiyRxvrdn
Rj9Cla2umA/ojE9Wu9DyGZyvK2qX6ckj1T8K6dG0F1ASUT4wltV2ebg9y3TBLE7GbP46HtO+pL6c
HGpxEHQv+UqKoSvkCsJfYWCLdkOXv5TOwbF0SjQLry+APEiNUZujlpH7yxHQt7g0iah4n7z2KDJa
v4CdMd3a+XcCzV6hy0W5PsucF1ZJKnojIYRjyJ5KQysenBi2CJ8U/G0affJPGid3OVNgj2HDYwfY
ApsIXUjmuhbeF4oJ+872gfQWhQuew/sRH7H2EKPRbt5sxilQ4jchtLCuYPMRVyuC8z/y8a8UpiwO
8OBmmQrm0BpYo20ESpI/vVF+du9trnatEADxs3DiNkgf/U4WTPr5QBmftUAmjUD7C00PcABLFy2G
BTGQ0Ea8H48WV67R+mlxBu3Hx5ueWYXlydjPDwdjP/fVj5+K7ILPCxc9844yKcxJQovYMstzPHgK
xyWZ6yEBd58jw0/FxN2Z48iEFcL/a7hpH2bXirjahRJUBht8mq3rQEsqglqVolilnbYuH170waBB
1WJWn+GOzHOM4AO95PREcPwpnPkRG2b5FlWIHDTlQ8F2eToBVg/Ckfq+PFuglPlRvUfsJoecb8mq
ir7MeM5lJQvGlpN3Rro1iUgp9/VdNCk9yzfZ/BoTAgKDQl8+Rb5VCAvsU/aAkrdD4xtPyqjGsluw
Kz7MDIgMSaCj5u303HBIJaBPr5MyGSz2Eq0t2+YR/rFpyZNRgEYv3w5i8Uq8lOCweGqL4U/jqfA3
KcwyYkPcYLrPQyIA1NG896vKajd9K36YUobFCvjIRVIB/BZp7xOaCiMfuJ59NdwV4hj4OT5wrjF2
szVpE+0bIkIIo30W/O7+utmizRb7qvWfyiivrAknAUL82jKsm2AY/piRTC5lAsdyAHxhMEEzr5rw
kh6NWkR0+wERMHDLWOyqKzIOFkp9EoSmneDBQ/Gr7U5nhBOA1FouSCZ87dw+NobzTYHCDSh4HKoL
y6Zz4mYURzbTnQnhTN424wnknOhx4RoW/gybkPBFjkzgw0SqNU1if1Kc8/W16TkU7/R8rEHEDb3e
0/KY+Yf2O5BYMvRr+FDYLjWp8vXjF/ND6BamqGUi4EkC7DbQMvPXhoM/LKnsDiqypMr+9Eki/JAQ
KuFqKeme+O6JLRssr96LgW2viubgKHHVRzNJ33sB9/aNfOZXDcvaK8qCKBMFR+WiIxdJ7HD2Y8fr
H1XF5WDS/SCzeBDooTQRRnhmW36VDnHA/4N8XEq0dTcOcwexSDI7GE9m0XnTz21xs+YBRP6Ocn7P
R7z9i/LgG4asM4zMXdmEwuHvFuUFQ9bo+YIElBZT2I2X+l5f3X/tfnDce2jBNJ9V9jQVdCo1tchK
yjL6zcmWkJw1qkD1LTXrQttBaMIezdLGcMDuSU8pWFUFEE6wu/4Zqymit2EYU98c4005zbDUbP5i
ef/eI+FT41w/rJkRi5o7QLBFgw8i4CC/N0vXra/m8JLdwPTK7l+RTmAb9wyhfQQS2m17lW6jKyFF
1n6mpIafBh9H4SAlf4PaIwIK+IF/1g3EPXB6dnGg4cG1M37PceR7Czk8yTWSBoCjIEFk9fZbR+uD
GvfFIgjwGddM/eq2k116RSaMcLfn2RKRjDiFjUyjKWnG9t2RkI3Q5pY0glHA/06w89dnMSP3PULQ
u51WDRbMqV9m0gRSO1drIUwEqb/eotZBxRnMZtwMP53H7a44bOSsEgcb3Vy65aGaXedhZ1bBzggy
/wcEhJTKV6z8uRpmNcN0KSwyqgeuj9yTAUOAe/xRf7QSwkUmprwbLbNNzkAJPLR9JXAHmATvfQWK
H/L2lUPoOFYjfEbXm8n3S4EIGXBXBTY8/eR9sfItvcX+qLKG7thRMobrcSNZZZs8w48en8+ygpAF
7qwGZQgwwqUD/OlRRuLtc8cv9DG+tuv0RAQxguCgEym/ocFhTQGLsV5+epG+TJF9TaKYEuJoRoCl
hwwFR2ZHRNnT8W5ZtGqW/WiYaglxO2cdSLkkqFthF6GQkeNBagHYX+gumV0TAMQ3NsbT9DyNSHww
VZ7bwhFSl0lXlCY7PLDP3FZLi5NRqdiPU2X8nrnaepURYOl8BBoRFcrZ39+5kT+do7TSjKBK8kmg
Khfg9SyfktX/kT4fTYK7ou9uePtKCh/6PGelzoNqlv7nVt/ea/YphXwDxIJXPleBwRJ4iL2BN97R
wfA87uCxeYjcaL0niiloQ2BiW+ftH0Gs68QcttRPcSO5Nrs0KDv8RKgSm0pFQ4Q0gCaE4uDb/bDp
XY2/UTdtdKt0m4K4P1B0xgpuWaGVqBer9bO9zl4oNi4+clKpOn3Hoar1+RVrig/Zltke4uClGqL5
AKhqZXhJbW4yILZUN2TUe4PR/sy0OMfbGbIxd2UkWPtVnQrZmfdlL45F8fqG1IABUqXukwOg86Id
vZe8Il71H4y4aY3Wvz3va97c3P0cL/SVFufMroUwtgv50q2KE80+NIVJRFdsvKWMNZh1d8LLlBwf
GhvvywrWsb48Po7zBgMoO5kBa03HOWXnR9WMzICjifpY/VY7zWjD62onj74jASAsAUnb2OTL9l98
+LUIhy9WoW38jjE7OnlYhVoTYna2+GOByXPWYNygzqPbMl1FjwxxRNR3iilLZ53HMgQq5NWUjyJ2
bIMsOHvW7nvPK3uSh+Y7LjoJ7Zq/5nH4jST3Rb3BV5+gcYanEJfdtTDrkrcaD2YXbYtqIzbg4l9J
P17f+wDzSR47IIyxhnsc2aNJgU8/mjdSJO3WrnLkeeDZekDPtilDZGfwI9p35CVYT6YjzLEyIMpJ
/6o80zV2VpWvlUFNdFLCCl6tb78ZGVfziFWGXWmBqCJPskz97hq95FIot1TExrybOShCgACHPUcS
+K6p2Besuc9TXIBpZKGXeFP9jOw64p2yhLoPYVbWWglGWmp4ExA9ctvt+ys0iJ/y959JF7j3lHke
VqziEpTJBXAp9v6MABoDoqJ/s4k9+xRdTj5YOC4Zasi29PklVYrlWx6u7vPi76VE0YO5+OM0GyeD
+Qr6IYTG758aIl+KFfzoRymRgFSNDL+0caOvWiNOehy5bisSh799X3jQOBuEKpHPCr5Q8RHXlOB/
e5yWLV4U+qG6akl0tABmcrQtZfYD9F4miwwqT7S0XkGGrVnsp8C/wcfNVNEGKrUCghV/YL++sVmW
RsDqO3fe0BcfK+el/b18ZArgn4ocf09KhBZB3r2HP9qA/695x9APOcktRppp6J27h9oXUc8Z2jdF
49ShKF2eYY9wCUDt87QZYX3I3GPcFq8xZivtzaOXjoMWN6NfemnqLHFMGw54+Rc+Do7SmWpFqAVC
cLaodwaP9TuU3QescRutG1oqXy6LI7RTK4qgNpiifjGrfvhOXs7uRZ/lAP1edEB7zwhHQtNIRvaG
pHWYD3ecGWdV6jyhstrnHYdMfG1xTTmMG3+OwZVGhBmkb5Wj8hgcHfr/to9NoQBQjTWcF0rkptBV
5tI21JSCKsKwqpw/zlmnMbPvD6Ckev9ZGoXYe2yHu3YSm4l1VpRQGj7VHErw02t1P2A8D2KpQ61E
znxMky+AYkt9ZT2KTWFMXCujIh4OEYQP88JfRDI5AN+jQdixWZGUI104K1rMiAf0Z/hTESD53fRA
4UzrT3tMHcoWA6kOTW9mpIWY9NOJ3M0I26YBfb5FhCLdnc3lyyQ5ett3Z3hz1hY9rMvcBo+L1OrF
I0l4doj1nYMbStOBUphzyt+VVBSI8dT2VMCzaW5kRwocXCbQa4w7Bbz7WAwjWT5NhJqxVDVuKpxm
1Z5w3KDKGYtQQMXcVIxh+Tqm22P0wbbp0nR93wD5/4E8ed8dNfL2K6dbl+8CgbWmZt8U/+iCAhJw
DsPtlGawDTTPrt3E5kQX6oJBSoZClL+BhFAsvtoj133LOTVX3tX8qNrfGjYwgeE+6o5FO/J4TSOr
HsWRDapUmOjO27dCGTt/eaaNEMVjnfO0u8L3gaAUbgaylNqqG4OXjTm2NneVnzI6DDf7IgV7fe+q
Sx5QOFk0WtUMn3ZhwUuST7KImh2egOX4QTT0MdYkOBKsGjqysF3P33/BL+6n4oUhpQs2SWee/mg2
IvpVcE1qVgiiytWrFMQM+gATTAMkIMGMyf0QqTjI+5Vem9T6f/ya5XG9oPZd6T6qmhnsqyRm4sOS
8QHZRJfdE/ycnzC5jzREBnC5MuDSnSFBIJm4TLgpMLhuzHNqmye9o8raqkYSIFhJiYlFBX7IZdj6
y7FpvVwWdYmtee6wtlsONZZyss5n1grsY5hgGk61WymlEA+j1/K6Ztc7dNhR/CsF1wfXAqgSzj9X
N1EhViMUAhduliTNRkK06kbLQByJfbP9zqrhxzKPivUaaNjkUos8ADB7475+MY/Q4aiSdfFmKWib
oNVmckegz2jA6YbErfZBnreLTbIUOvOXQVaaK0hd1NaItNxe7V8k9VS1VKJKVwqUqhBxOaDiBxJ8
OICy/S4wvGzJs3HTmfiBQfhWeV9Qrx89d9XY6c1VhTnIRX/u02vc5awlnUsDYD6zuuM6I9E+XsxH
tDqixnO9FMbI3XBxa8RLDk88sR7DzeTpxGkerZsoPoKoeIFHTS1IrWZR77iQg8zHdiK1Z7P815Zy
NG4YQT7uOOIRdmV4vdxKTQiQPc8Ju5YnRg3KVULnmtHQ52tDH3QVoPAivngp7kC5yd6HdbD5LYyG
I0A2Dk7oY/gWS63/S34AiPYklKhTajCrtytNebVFfdrHUzIuisFzuJsFUTmhCUWbXz1e1O8DOSUe
XJAPGnYeICKnp8G9Ufhppclq7taLhLrGY0qfOTQH/K0Ef7Q8DsvGWWRRv88f1mvNV7aje8Az/JZo
rZRB56hMPmsm6Reb5t5vnoRWynMlm9EFKTGqFWnV23F0J2m829fgmKZzj8jpjAjxvCKd7+Anu9iO
i/CS4s0Im2JfSHb/DdpCE/M/P9/rU8sQQq9/SUJg26suYPM1rCK01ZfQcAf8mpPhTUCimvbdNEQj
JmvqT0PVlPbVP6KFDhr6Z+eJQU762uoUED16ICdu9Vg0tWrGkDGchbpq19TpKAmCTHr7FehlS0FN
RjZkY/imtaxeYCnXle1lj8bt8TvTBggZeVaAMCftz2OLFCYNL+rp14GP3cjGouvjlSYueGKnrsks
Ucwt1J1ZFV94lw/eGTLl5pBwXt6241AAjmknL0FYQUqNVClKZ3ZgvDfneApYz0FZxq8k/0nFybJb
Ky+NkW/JQsqSn54rHSUy+beVKINVHeDKfOfTZqVjeGcE2rHgGi+f+5wFKm1kmjIVHBO5K6Rdd9qN
awYK8yoF16gjv0sNo9gtqJU0Hgh17lVck6IQOIVLLstg1koAyEcA9IkmnLO7HqwhSLlRsvYyRLF7
9ttxA70x7lBgcVFdJXf+XVGlCJTcsGropV6UP8atVEGd4h29OFjf3u7yt5Ap/2y9bHpSWZfy2ndU
t13A33TJlqE5u20SsgdCqnxI4NGRnBUpZ+Y+mYcNZdDuRrS0lg/u8wVvPA+vmx5hEBwb+anP6SNR
BQdGnp/2t/gJbOp/BcnmMVOcFQIzjVWsjtK95HEcOPf4CNm3wwE9UlKGKHpc/15axn78Y3xPM4Kq
8lP4mx13AfGDnmJTR+bbM9OCz9av8IUFqZVGSrnCS/XIxwdMz1dtjobTco52FtGXuGbsnmVfgp42
XpJXM8+yCHTac6PasTxgmerpvmdSuHDJM3H3Ytb/AcLv8pVg1SfvgW2ucbPZIplwuyL0Ozk74Xo1
gblKpLRIHlZ5OULbP0JvWHtfzCIxzZs6eZDd9BrZOJF+O4mD8ftA/i5vPOBOgOKzxge1EJkVS9EY
ey08dk2Spa9UnrGd2sjpabKtQ6AFTUg7FwPzKb3lU//TXOZayQdqVkTNw3zs/an+CbNt/v/CQpEw
FDNpdFJX2jlSrO1upknSIqtekWygwTBO9DKh3ziYHJf3HMwJwA/1QKWG2pDzZsPDoi0lp8c/YG7b
0I0RarA+/F3SNFl7QGBd2HWdNpsuyLfbyqNCgkx9VQi2GelNW6o8fUSBGvnINxn2wJnCxLwj2Vv8
YQpEqkAUzoneUNChDWiYQFdH53LCWpiYR3EwCrsz4lEBD7k8b1lsJ8Mgyy0orCmSJvqw7YjpeiYJ
uJ/2lQXrqCD9SRAVh2zelGMONr8ly97s11P97yAd2m+GybWwXZS9EyiO6SToz51tVaG3joi2Lkq4
IhQlKeAHLCGs4SVRFXRP+0Dt3+5InZ9YavO4Zl7c0ctNJZem6pbtiv8i/N+6xhuxWC3sfEYdXbzL
zi0eROGS+cwArLiDCzuAy60//ufKLz2/SWij88P2uwj64O2VxvxcpvAl9d0aV2HocB9JPkM87iCS
br9H9Jdnb8xG9TVjqBEVkVe+ys1fW1SPnhTNgd35t2J5BEZ75HKIg16O2h5Jir8umwA4omXRmCXe
gIYhPj8F9pAefkISvvjxNkvF6+40MkeP6AquTFGSOn/2NiLWx1Xs4E9xphvgZNHmpFy6HnqFtgba
j4gfpc2atH3dhN8cfVk5A+QFVfiLvH7IKxb++9qmn0LpZzpFUCwxMotVlCdMeK4EIzhX6aOJUqnV
/1KcluQtx0VBEiZYEDRfMTMOxnWHeN0Rx+f8kmnht2vfrffiKm1KOmLTrJ1QX++aH82xX85HgLj0
CMjRcKVDknLFQmL8Tt15i9dh5KpxtOM4mU/lg868eyMzfqqdiE8Jifm4Fi6cZr0gWyqhFXxOzWHK
I9FywXU4ZfWrE2pVeYn07z1iaDlVHeO8xl21dq+u7YIxMk1vZNpsarh0mokVMuEotYBOpyd1OV4f
wnHeOVjDt0oHnzZRAMo05znfxYpC8H1y5ICwdMlFARzRtAETgIgN0NgwFDv5OkMMUDLc8YYFXHdt
e8xOLbLhi4WsYxdRKIhKIZDJgizDoBcx3Srq6cTXMJPMjzsS8ugNbfPhOo1YNLZAYmyNBiMfAUMd
LRWegjmeG7bUl3sYvRtjmT2x9tJlxkVSlxkDRon4IvMRZJjThHBMUb0LH/eqoJD2dRE8bB+w5f6O
LPb4ZtVQk+rGeb6DD2KjL6+ofZI2A0HZYgePV/wh3ygLR6ETYVuokeJSH7ULnDZSu0oPI8zJnIAz
VTOevYvnef/2RAcQLzQvZrPTuX+9pjlE4heYsyFbgELIUItqzfvCtS/8OhVGDGTfXsoloexKeQRg
hblMyBEOI3sGtmkJUlPhUHeaAVb2LV/nG6vD4C+IPdAfY04uFau15vzbXBgmMJBFdjpLxmk9FFra
DFqM0qGNyUP8Yr54M/RZOxCb9H3irXGx1VkOqTJv3zC2RuECmouvZv6dTBvhSTm6o/Nlywpq5HAo
rpkanfp3ZK25St5xmJKB62qzyPHJrfoBvaayD2yOKHDsl+bm/ZxOEmZgpl+C0lIFDJ5t2P7NqI8r
y2iozb/J1lmCkRd++iWJTB/ffA+uQEtmgcANnwD0IMG8Sn9iNR9Wn7Kk4X7EmmBkGmavtDujPliR
AaN46hDHm9XXOepv4/rOWTX7swgfWuWcpyUhiV9z7xLwQZoaDWUEMxQFP6t5mwqIWjjou9m0fwZD
BQ/6nCEJw6/kIl6AIJMsslZUXGPNINTwogccgVZCeqfNGsDap8as9VEo+/Q5buHL+6Yonbvs1VoE
2+hPBfkiUAMjws8Qi+9Dyi7ufoq50XfZLIzxYpMKYVAK6YJTMFz9R4wfo0+li2C3nKfvMhOYIpWK
Lux2OT0VXTr3GMieaPTcydY3boeYRtoBHP6OeZDZrr1iS2wfTaHvynXuxIEcpOK67aQTY1RrytLz
ZPndBYTpRUKTcI+/IACXL4bMF5DU5bl3wI/WbQizpmjPAXcaByLsuqBUwBhCJTEqMk8dCgLmOXpA
6ci0dnGTyOMF6GbYl8LEGc6bzLvrDnjo7DU+MR/mcxVtQ8c3w2pLNHYiipuLdHNWvrBbUQzMoN5K
qltAb9etZodW3UsuEIvjIkNt/LtAvMamfroUYRTB4xUQTz2zAbtsb/yqvHEafR8QuYLPxrak5vpE
PrMCch/8nVm23YgPHnTTNvYma3S0gha4qZCwLsHwgmDQ/XTBLIjYBollV19qZeGU2+BacEwhOota
chNZNaV5Oq/D63Ta59/MLXDxTkz8IXBi6MQsFBRSS5ZrV+OJ1pYLp4M4GkcR25E+rbB1xpwFCVi0
Tx1lEPxV3A0OJzb1lRd3nq2m/9fmtoL1NIMcc1yuQLEsYPrZO1ZCclleTsnQTNVE+7p8cU4t0RKF
EVvM+U0mB2Q9LRe1LfMbWIyz9qkILcGKv6Ii/ddmZigOqprzlLcgOiQ3qzlIgTrlth7PD67OMxXb
77Kl66PMOrbVLhVMYOH59soMz848T9MyZjFk3nd6ryWzRns7TPeHQTcInG1uFqU7turTSePNDqmD
Vo9r/My1pUiwtzpEA8WmGaC0aXf4QD9KdKvgBZ7aLtrgulmhZ+sEH8KevXOmyx02zqH+NtL4EpCo
1LEjmIAOMeSAtVWxmIoQb85Fh9kT/te80k+1678XnB4LML7D+rhb5OU1ejk5z+HVVbTKccS37rti
Mtnkj6AnhGUxhij/amq0HJIfdGavFvKR97gm891sAh55mZcriyzD9FbdiFdvaNZoNQdtrcRHgJml
GAxuiwdBW4SMtRFZaLt+LuyRCFWQfXfv5aCMeXkqBz0WLc747rvQKX6VIvbrIg7bICgKD7nlUhP7
wY0vn1nkIK7oKZCk24wzPSTPBPb5iDHPASdvY33VIzCm+nd77DCNpq7A9/3FeqdsBxQoisXZP1eQ
vw7mfSSDNNOZpvZhSwg2mz1Y4Wgi6pq7Urp8KYp3Qlpo1dWcO3AErS3BWcGv3ZLiuNUVdrEUqkGv
OAFaKugD6wRSONnqrfvIG2Hr/JeOFgxXp/k9lUjhYwEQA9b7o3HO+P23NvnJ/XeV/8OfZcxuxzyV
yfSUXWZsZsQyJkpjwiBpfNc4vBWRQqKmuTIWcpG0glNSKkUVwMG11CV/QZGmmU7lbu8ncMYVSUv6
viahXemucYMBqATUhIn8139PU0l3B0wSlK2ORxtn/ZXM/oSYV4sdDSYCqEyKierP6KyHPD50mArc
TIGkXjfe37B8B/gnR9Dg9sXeqosGgpLFp8jQu03LebRADGgeufeyYUAHD4IZyHrKTmesXem0x4Vd
IOLwM7CBMwnxRRgt14Ro+qPxaXtUnxu5FbX3UCsfG0a3Q7hqAr2dIwaN9hF8WktgCJGgyU7jnHnS
552YjwmJ6ZnlFeFVKskTe7DJjAbe+J7A7W1qRWis33qzSurWSymfdftONDNUIgtN0UXVUvkhE3Or
MG2QXrGO0tCJly4WiX5C8CHKQ9YUOPqzVBLJCGcgUhf56I4/F0wsduKkDqzDZ4OkJZcY0fwM43Mg
FpzFURU0d02pCN/eqMYc0G3RrYYRZmqbpPUi6MGM8cWxc6Qf97TViwUo8/zRb4X0fE9gPgnRI541
ZXbHzh8o6yPZLnL04Tx2T+9MNsuxjETG0Kq0Q4yFomEpRfAodBFWDQk/icZ8hrt9HzAA1GMZvGEk
ToEcJH4pZePrVI3+8xHAUy3L5NMi9AtJsua7f+ccV/aPZ1ttGhN71EEBdXMGm/fUkE/LmOPQx6EJ
P1oXd+BNIn/EYloXOjNgH4d7PMlRK96cOSV0oXvvufCGYfMpBkS5dITgx0PM3PzaOzMK17/+Ast7
q8/hY1gwyQW/LNAgOIuO2XUD3oI3AAj65queX/4DCvq1if6PG8JE8WvqZtGxIzpnQkkyZUgWzezD
QWgWR2T7YDX9pEjdJ4NM5TNLiLk1mITgWWLpMZLjzXNL4Pe1KLw2gT/5BP8rbBe9Z4cv2UCLJcwx
7C0n8fLpi80cgqYNxPuXbYyWZo4jP1/qn2xWPvRkEZPYkfP8y0Jw0rZabv9mrdNk3mF9rKOYRMq3
kahoWRJW5QQZVqds6oJbQMmWSiMGNNdq5KRxg3C5sXHHTTjho6dFgsfjH9CqsuVtkpfOwgHob5Si
KUcMmYwLaebYwhtNLbnNFxru6g1kZ4eT1fQR5e17lExW1rpOPKx8Cjgd917UNX6yK67SHQKafNme
3tog8Dk8w0B+8t/DAU6YUQ2LVby30iPav7K5kFTPr5X0lFhck1SF76Db4Sl4w3oX7pNITWZDrux0
iU8Vx2oG5MAWU7dHOOvsR1/xf819lsP+kdvevvE2/v1pKXHlUdf02HZMiKBajkl7nxmxor623/nr
wIj7hx6cfZbD2pkHacLDKqKE2BJGpVw4imA6NyKZfg4pviC0qkaDdDOups15Cf22LNHZTw/If4t9
uL06pk0vIlF9YY2ZNC3oKo8wYVxalaTC8LGFsnIDulEmEW23mnu2g0QZ4PQjaTS8TQ8U0rdRlJJ6
5P+E9FA+lJqH4Bq8VrOmYd6OnBTVhkZTL8xuc86EWTH3zNkaKb1X6f6mjKRTCeWNAN1CbYsAcrk9
WouEn66tqe8Rzmx+tSNqT52Xdc5uNSnv8wJ5aMgeEGlww/Y/2VYbPRVIDmngorvWlcWRg9rm1FMp
YZli3KwC3rsk0WRhE749DXqQ8HzQWKjGA1xNQuTwli3ZDhIy9n/D0bwamz8NkBykFpbLEXDNTaTm
d1EK2azcvFqXxRAkiNYEZPW1b6//dCzrSsj3ayrWU1hw/MTiKtp3ujLzJFayWp6vyeQIneGuKTnZ
lMacbs9vG/E7GrV3NsaKQ6QH5pxau0DPslfq9cpmYuwvB7eeTKf93u2u8Yqll2Y6+iIrfRFC2ttj
xOFXkfr1uNG/mL5UU6lF/9yyu9Al5n2ScXrq08FKAT3cotRPoGiBc+Fctnnxlw3N9xG6V7gPViYi
yLC78SiQnjOsA6KqP/7woGkrodL37E8rbc9LJR+/Kt0fwNQc47qZGzgdEwra3584HPnXWA0L471n
TmfR48YvLdRZabzyA3l/tLyFk7JBgH3GBF54CjSagPxr3JipOItdwikCUlj0V83K5tAiqxSk9iOG
BVZWzQrAKgPaDMidonJcnfB6+Mtcc+WnMWm2KvhqmWf4YSiOggDXc8Ih9xM0BfDy9HJb0fhUGd6s
Uy70o2V+0eNBQnbxG49y7Mw+EmoFxlk7yk0oyiDMsx5GcR3jjIpunee5zzPOLUiuv/KImSw67n69
0OvBM8JMlN4Cc3Zyd4F+W7xgmmZAtooufagT3a06FJ8eNUXalGw9LaFTqzoluYsQpChuDfMdNX4O
qh1vDNLxrlBDZqXuKl8Oamcoe/MF2j8A4QHFKan+X/Tvf3MJ529RZrz0U9eKz1ziXr+qV2764M13
zq4VZSFYVljKjBZC93OZKiGUiE1HrGFLt2pszV5XlgsD0Iq9Oic06KhAsGl/D6Gs1MxgPbv0PLwB
HRS+geDgftdKCXhk+V1WaubbawXtRZaWL+MKysQCxylnVra9z8LbeZmW8mGkf0xJy0VhUDVT6Rj7
sSQ3L9PWz9VP3k0QOL9WxnVHgTT1TfSsPD62+rBlqLWFN7hDpJUy4gfZ7CmsyUPG0GGxjId4a0Y4
yXjfo6lpNFm77gI7bAbvbBOpVAIBpc/7c0PtpXpc8pGvBBgqEiRX4pqhDLB+c+fyIPELT5dqAape
C9zsly5tDj9y4LMqMvfkyVgDjUyBcb4ohUud2+StWFQEBhEUPnrNtNjiVJjY9XOaAErl21Q6xQtw
VTS7IbAC4Nxcowoath7TPIbAwOwG4zgkS07CFRAHhUb2t2GDvz3vX0LtPOWljakMuj76teEYtTrE
76eJm8rCX3eDHIiOhvU2Zi/Ys3bEnfl/99eYOKmCGPKmxylKcVmXvTOGOpPjIG4yzs3w9dbsqgzy
GVjKumc7A3JJjex8To3t/j8g4032TYhiLBNyd2qvLPi27xHEfer7JbULoWMBjfuq6okr6JfCipVc
juZLiCvVL4t+1j6nGRC8PLvV10eGu1aEyRQZX9TwHcMUXrhWB7hd6h0/nNqRmA9fvYjExRoz3m8L
ZrjhoITj7r46CO/AQYzISkatMBnl6lfgq6dfEVIT5aOuRm2hegBtAyri53Vt40YqCOCM1eyWP/7a
WyK/VqytP3YY8vLoBedIEIpP/Er5h8fkSHzbHd+G1/9MTFM7p0v/FCmrbhRAyCLAeK380mqNNopd
sqoVQLwGgX5IBtgTdX25p9Ox+PmXt2IorlGRpaHzslXMEu/LHTbUqjL6It/xY3FYfLUFJZnkXuwO
UkW9pv4SNsGT06uSbbBdOKVJIPeFDBETaFbTndg0NI1/Q2P0eTkNBlXzcFTdVLTPClk4MOSQiUHw
ZVP3dS0bFAr4+qgJlMUgO/CRVFSk/W5j/D1S0nzeK5x0tmaMI7e+EAukhmcUGQ5TMDo5qmtgkAMY
ypWVh7cXjs6UbhPXO1W11PuY/rPH2WruGZOzD/GJWgso06mN2bofxuyrsiBHAwG3Tu77iAxk8oFK
oNevTgIFZZtoRE8SKyDos3WAL1jhVwIydGah89W8cuqfdJerqDb6+7UhMSp5oc/9wT/xacXVWDHf
PHKWemkY4rWOaRq2kmH/7l24rsoN1tmMVH6AprGVuVp90n+nxVFSU5B3ZQvEzaZnOrobhL5E/08r
7z1ZkUjN9fbsdYb87hebqDqVSegFqi0H/frcaNFhDGttvKzGkD+4y23CcNdUeapaMwrkcC9x0i/d
YXbV7C/WkBesjM5ULyLJRZX3hf6NwkQ1vIhx//YRTwT0oABepPCPU4EdYla7ZoxyZcS7cECvFE0r
h4DyqaceYmQFNy/o0Bl9b7V4i74mn6pbIFAMBRV2XE7cTpmv+ljYhHM1DGJ3tSLm+Uusk7cXtLex
rKxlbmRwC/2k0TdEwrAHThiBpAR9rtynPUifBv7EvJJ5f7BwcHfc6Qr3XMnMXs1ZJj1Kmo3/2++v
oM+G5icXun9kOXw+i9UtGDaDNz8+rMi5FeZLV1YW4lcoygLRPFTWFSHwsoxXuZN/nBLMrB/7UART
joaVAQkbBP8Pap7c6I8Xl82ZWA69YLisxXohhBKg+vSwdt7MHSLSAAL+kKK3/mudoQ4b+ubnVjGs
Q03Eu3c72gKEtNF1XZyrBYXhW2gyM+qDWAja5EIbNAKFxtlY7iE9a5zCnW71SDvJ0yOUJ4rciEIK
EbFe9cZCQlgQqKpW/1eFscV1Iks6J130Hlj/JDTHpVlE6D0yqEr9puFfa3ofwjeMqBMuyXOSVwzz
Puc9Blfe17k98zaeIz3ZUxgJZsvz+YL5eziZaUweOaN/2JjQ7dlEWDl2hqtEeQCS51DJNpj4dqcs
CPR5KPZgU5565hR0SOEMjh3iSjdYu0ax243SzD4Z9zOt7/rzbhvMJxRaX8INUtuNbgLYIf89A7WC
zh+Gn0ciZYlu6TXww1T87LxgSyzs/Mdm4NoKFLVkpHfZNgRXEYZruG8lcVTPp0CIguo4ehY8Ltor
D+qjiqZaRvhxgTMNy5lgzaO6JqVhd6HzuDFfIGCr1L6v+UC30nJss1e3p2s6Yj90O8jgXSdKfmYT
xqK7GaijCh8IiE5/GJ+6XufTWdBnG9lMbM2UIw272N6AiFfTJ/g0lU1echCBO87prFI0ZLLAow+i
C/rRLIPzJTE5wZuHGz+rhTBF+2rEOGi5GGb5ZorfKpPLXS1zovQ31AAHIhjyhxLiujcMZ0VAqgoX
DNkI6Cmlpat+Ll+dFIhjBhVDjzcf889jtlGhjq1FhsAHg+1ftxvMPweL54YT//NNir63R7Wj62+C
Gz6T+1/Eo13IM0jn+NVb/4vSbtNIKM2tyuZXlBK54Dx7ZRnHmKb5+B/qWz2E6Xa0sUdIIr2lQrEQ
PJ4vD2aDgMJ61ihS269faC+YbG0KpvVs/f1t7gI5NzV+fisTP/0H2kn7a4lEjNyJdnDuXQxrjq5Q
zBqk116P0KYwYv0CADCXM0JuqPALIrLZRRAcUK+lZ59liRY3tR2ZoM4XNzFUYjTGewllVKSOhpDR
/XayRsmLm1koBc9+cJSPi5fvE/U8xHaIE61FhF+/AKPOuAKBCF1GPcsPQAbdzT7zVDWcUaxsDxJf
BhVNNvU368DnMvSw5kpKKSsGiMtY7e6CU/pz8sSHa9pAOiXX9iRF1ba21upsJLN80DrGvfA+JLc3
E/bSSxqHphB+qU4+FeZAybedT9YVUM6YcaKL3Y1bGHlryyfwtjrZGPLP5P2jCcwjeW+RMOn5uKDd
jh7AZbU/7PciH/eZtmwaVqYzd5m/kCLKzctsZa94cOnl11VsKJlRf2orZM055VljZUmPJP6GTjHx
kcHxWbiKXHbS780D+5gc+se7TAk2l+UPdrUImrYLsH9oOjGAcAmzIFmgOQ4qZZtbFAN1mjfz3aOT
WRUL/bqiuthAAYWh/F0KR13IJdJb4sMQiJDFhyOzR+dpikl4+sGRBa5h9pzToY6v9BApJcvYb2xX
VYE8SAmp6gMAtcXl6IAVgf+8qR8+gHA6cDz/PeO5eKUATTfe5gGH4Nn2Mtd6djEFqLQXiVMciTmz
6QfxoJcr7AYToRTIEl+EjAwZ5T3KxfMeNl1Htxk1vKtPx8BgLGfRP4upm3pmYS7LiSAQAYExTwUG
jeyPKbe/dtuMEplUwG85svoY9hZX66iXNOZw8JxVhj5RZdTnMiQAIPpryYyADaL3/YN/dQBy3phv
8pWOot2qr19onOvuTaEjuGZq780MELN9iwnmWmYFwjkHgge2kyEfH+Ar4N4SpcqjepvmgebxnfxE
EdQlopzunrJrbX1RJagDKlnu0TRNLzyqo/8+KDWlZPXyyhhq9b1sJLyXAshmIPmj9joxoS8NPy3m
Ey4mT8CuMeCAWsEy9/+E8Qu/CeBKH+omMKtyZWoT7ChR+vRTKA/nE02YXyDWLq8xeQgLFYNSDmSd
tz7IN9V54r4VQN2hxtiuWeatSIuy2NZx1LQM1GvHgIk7P8pAm7hCzwopKBQ4CHX5xrdIfGFUhG9v
7MsNmLQgtzTwZxw5l5dFknEFSggm5QktfbesdsmD+CS+05/jwNym+f416xs2WgeJf7obW0XMKopy
TyaFmTxod+4fPLiR9vKsoV7jMZlT/slDRfVk1hC7d7ZztFTy+fuebTCBgdwnIilJ3uvBPRAZ4MVk
N+g0FPlNN+5dm8Mavke0+M6ei87BEMql1QB6whB5JccyKlW4CutjRurApdyuKX4pvq+o+9DcVocZ
k6lCACshfS4LFWwd0/7GvcOXo+GU/T/SwWCM7UOnRJ1QXNPQ6C5PKLQyFmvzUJSwAsDZWp9Bi40s
Joybuaelb83EThlX2ZPax5BvxwDuepER1xYetfKfXQ849m4I/gEmwgzJwwNSC0pBdqfgMnF5KS1x
li7MFmovop39OfNa45GAR6a2BPlyfCgFfPRLL/LMie8HC6VtxnON/VHS/D3QabaHtu8EWMmbSO5m
kX7HI1dXPTDSo8yhPL+wDRFcJonfI0MlDxp6ErPHnPTs6BrIreDVNaOmAoWfpyxRg07mLh1kS70m
9CtufqhYowLpIX8CQOheJL2eP3H+y6dAnXrl0N4nol9db1oO1VD5x3VNzhiIKdPjx1Rl3u4Y40gB
tQ9oWdTHMHIzLnuKwSro1/xsMeLBkZvBulPVaj3MBQQw8f5JS/oXCfeY3zdp7soJEExkW4Vptjix
eKjDn/Fsq3AuwtLYoto+UVZLE3Kmdxli7Z4MCv9H0+WP+KHC2HzIm41Zd2u8WAZ+1JUZAW7/zMcy
G6rTZVQU3Osin0B7WK5hEGTpVNtml2kLHco983J60Roe6kXKt40ieSf8DUdCewlFCxEAVNNc4YWK
gLJI7v3LF0w8S7VT+09FTAxpp/Svcdn5BaceG0a/2jqUV1vKiccrA/d/iBg5TiUyp99qThyXQyRJ
wixjFsP/Dxcu0COKmRT6rKCb3Du6ZhEVoDUjGZjrbYaCflRaEsZtAkv7Usr+p1lNAKTsSTsKr7A6
cdiWkSO25S2AsvgWFqYRwVKPsSiP0TUEfvEayKmhIcCvs6imL3QECQItHiZ8BMSjG3hgwVTk9a22
vmnjKjdwGqT7qK7Mlwtnz3/eEmGU4bgk5IJPtDkepkYbnB9AZVNYTwTSwlADEcD8+Lc1UXMkVAd3
e65qJeNkBnfiMIVLhKnmiZCcOc1im254Q7lCOjqRPwuEC3wE3D3ilbRJnea3reTNA9qWruLayloI
KM47Y20WE70OITmArXj51ojg4x9jlkavBdQbUjDYfbQL6HMuPgd3fvQH/OjjlGVCNeGITzhxvTAC
eLq0QtQ8Q9u5pEPnc+QcAWopt+r+DDXXbZB0s9zlZGePv9+Gzpd8dylzJ2Jf8Pk3v9gXVc9bXh/w
k1BfdMyv2+GTDZZ2uwdJA+28SVN5sOI0vWJUVzTQNlqqPzsB2SRIvJxNY99vK1Y1fsYkQY6eOfI4
J9cMonU+nfG1+Qpjic3xc4du6IHjcGzX7LVH3mIzWyjOle6+kjJ2TrNciWHkgdS5/ACe7PzU4mCJ
VpJ6um2d0nf07zuqLt/nlLKN+x3C8M9ExuX/qCNwoinycoGyGeDoH+qyhULpiZtjZ6/8g2nZf7Ma
1yK0CvqWe2sXg2wFsQps4yrpS0NP517lNLZlgGL7+s3J8qWgpOORyAU1y/b3VZKFqLVwMVAmb4Aw
hi1G3igVWhVfiZsNwFEBWE1pWjQLnuuxHH9SdvdaPFyCGevwDQWIUmzKu9Fd5k5ZNdUpWsEv5Oz0
szM26G0nztcGqQL+UmX/lW+aDWfGGQKCReRnZTMevTZFz5oDJp5QPENXccwkHkFJFrVLP4yGGw4Z
onlxY53niEQUBEzwZcS4YIgkiKwm6KYn0uL4a+L5+ONiu3N+FpI6MP2Pk9BZ/Zd4w5RPzM2gxAXE
l6VYZtS8+UtOkwxEny0SEvfcf0YsNOyc154lfIuH+gywYc8Gi8SkE3HqtcY4N+uQjlNHsZlvywKq
dMEO7k8FCeJIAvnjj2Bx+lBOeCkVfltZTg0PYrYXnOD6d5oqL7RzL5oE86993BfNC2J0PpOQSKZv
hcXvOxji2Astg2wHiUHqFaybTJ7moDpQcGipOeLLM3qqSaARGHubF7vpRr7sRiglCU9pyIgjvqmU
JmR3MioJT7rggdlbF8Z5o7xVtaI93CTTTBzDcH+Frq+LuaqcWmftDq6HGTYQ59UvEl0+GgNRpWXd
64j9vZ79QsCKjDMtdgh8QAwlSj+0AHjIatGVW7nlV7gCzL0FN1D2zOXz6aeJDJBlLZRrAn3VX9y2
hHGm35jZMEjlrdmjpioxybMAMJn+4dqyAebGfTZHPM4q0u7RSQCiU84IxJhMI2RsDe4u+s1sJ6AR
2zEno5Gwv1Q9GDYFh0BUrpcBqoBFf+F3IQQ5fLecDqu7rlI/JiPxk1K26n3uocYXwVFYVt9c00AY
f0Wt9cxs2FqXvL8VotX+jvU87bjYdxfDDXRiKis0Tq5+v+mO81hmyeudJEGUsgHe2lzqNpq6NXG3
NzZsKDwhQ9tXkfXkYyv7cVSjEElSCVXyvU4cMfwOxWEskexVxJYp2kLkprhU0AyV9riU5vBok8+K
2fpEifJJujHiFBu1Ug7xdNFc7UxL+fw8/KNFHKhG3NMnjMY+JlIEcw8VLfNbVotVb270Oxi/Y7E4
j5CBXyxz/mweCp44PZhVgQIdF++6V0dSDwt3foRVcy4+dOpe6Zv/TrIxl7Wr2pQNgOCcr7D6CLsZ
RqW66nkVm2Vemvg1DwXePKTJ8qt/Aq18WU4gDqYiR2AmSKDtoEytdA9uz5hGw7YU/StCB6DBPbrC
rQfPtLjvkptp+8TXbEpU+OvLrb74ACRtXBk3Q06DZ+1YS1OdWbEMFqxzgp4lHXGQk09ggJpm0HMP
zHIEHVo3l6fSIMOoBtnbXPL8FDzlrC8WrUrZKweGdLEan6cNaXYOXA+5E7JRCzEX20GGYpM3BwaQ
ipWKvmkoLQ9SZ1ByX6pPIYQ2OhmBvtCs5sS+Nr/vtsSIQJyTAwvkjYxCQxfykNcfLqTiwBmrca5U
COvacVuQIX5txQClXPwwX4MbKmwyt0TnJ8ALCl7N1rW97Afj4Wgj0pC++oM5c0XYcu6LGBdfTPmE
zUun3imRHfaTb45SEuyF3bvSLiOv1phsJJwnSXB06dyJraCRCaUXUSVtVQDtrN60crgWvOfw2kRx
M0H22TBFja9+yj6dQPyuSQaChLal5VnM6bzf0YEwyyCy/jtLLj8aePQJdWpznbjY8GOQVpWclxfz
VzXZToSYYUeFixuKU0+sfLFdP4IMeTe+G2M4Aap/vbokCL3UKPpM9ZiTMqCCqSRbmGhZGOT9lFY0
9hoMzbz9QtNbAEoznuwuFJjv8QiNDQ/e+h8z2rGc9fsA7XpKPj09KqYYQH9cwMlUVmzz3DAW2KMz
UklN5Lky6BmsbSNxgpe+TPJ/+VIhVvvWBPwoS4DjaSKRL3+X5UCbNL8ANZg6HnILdrPR9Qubb3iZ
syt4csqTnnSWL5kxHiGVDI9lnFWrRfZw0n5UT6lwYbfFrewUki7pVBFkrcH7HyGsCqyPHStP+Vnp
LMwixR5+/2lKNcfuBCd1JNi+jsu+qBup2Pn3Nw408Xyh25vz8U2ZqHNrd5eBBGbPx2lixVsssTN2
TA3kDfM0La4hqVye0ha04lWRiQWs1EPjeY1CJorspDMlLMpLzuEFu1g4fWVuFKgV+WsreeEMlOZj
KYFv0/n01nOFnIlWbUqHLlHt1zk8ar7PFNy5Ovr29v6QBy+xornfzs9aaZC3x8MaRLF8Td4ZwolJ
6zFRqZuBBtwUb/PTW09JSDGX51LBmVGMVH7ejJHBKW9oujbgXCfsG1uluz6XBCXank7LAbokpfD1
I3raPZh1Ty3VD/GdYgB4MgKOgSawqRkR00J6va+GvYbpLSzsZXCkGkINpfDnYeXCPuFB1k4vSA92
UrEVQ8alDTGPqCHC0qCH1gS/vDiK1Lomc0yEiFyzwqvtkK6H3I2Aho197wLuGzHSEV5xN1WGnAW3
1h0g+gn8AfNUXi95ZRefrOwOUNu5GsVAW64l3mTeBEaCUNZ87q0gGIiu1RJwkRDIr2BdtRchxVvT
aD/vF1MnEPCwqiTv9ki260WwdfA+rvmVfrvrKqhlsZRiDT6BD3x31YMOzr3Qcpri75vrsntd+8ZH
5zIOGgWBZrf467gZRbXsDzAN5kqLSUr/Ryj6ycdB4XGQIoumMTxYlMtWvO18y3p/SyilYKTIEAHx
c4odFb1+guRs6gFXR9NNgw0CEjHzG8Lq92V7BRJUbKn83fc0jZKXXidScJ53feHceCD5YY0ijaxU
C173yCClEA0rEY/Hv2yE1uKgMbZ6lUUkTPudl6x1X194k4ChDxq/FgxYmLNKOmT6zPfm+OYL6OGq
VQfM4MkF4e2lZeRYH9iV8mmz43jJyGG9F9pbsJt81jf08HxrfUI0iCyD8ozUud5JVTO7sCWxVHSp
d0iS/YdvfNV/ZGHycI7LpiJpyCBLNFruhmGv2D67B9zSZuy/FHJGyqQKDdW4xO8/txQQA/aQqDb7
wqUXflmhnWfFrEDvM5+Ri+5FRB0sR75pr1QvIh36YUHkZuFzpxEum6LKrpifSpoa7sh687aa42Ix
blVgK5aMgHQRnFHsSyljaFOMckozgQTpiYf+3Nte739On21IBd2pZvADv/59jjknC0ZUhkHwvluR
uqn2Em0AhJxQupA0aBR9wx2dXaJeo5bTQcCMNlB9my23upt+Q6W1+8zB8ABxEWImt4BQXZ43qH+q
Jwn92LeF/5F/FzoikyPX8rkNmS0ab16YR5eS2rcMK+UhNaPQvp8rsD4PbJzKhzJE4Ip9fO8AqV1w
k1kNdpC+RabXX5nRYxtNXrc0Foah5D6N7P/9KZDHHNXOLkNikm/jCLYppJ8+LIvErH2zaFPcZFmI
8gkejVvxjZxtZ33zOexsCoHRYQ0Mzp9NDWc/gqvsJgXpJRK5/210qNfBk/DyCO9HCbwEelkqEjKz
ev5pGhYhFnkhlIaH//oab/rfCdd0t+NJEwR2H5A4BtahYlgApv49Ow9ggqHoBGArc9Np8AVtm0Y5
kKeWHQw5Tbkz9lwoBrtY54TN3J1a7N3+ijQICs9d/RZfw+HkkomXOeRu/QakE/n+N2xTt/wbt2/z
ibrdOYv/89djYube/q72US74+FpUjVqfKo77BkDA5Cy5UmXLTGJ1DOyc77v8eVQY0KSnwe3QV4A6
1Vapy+0hq1i/QMJJ+dQ0zjiRW4v2SxDJsz6jsm6lZ5BpMKMaOg5EVWbWkbb/i/Y5KCac1Z9kTIib
TznlBHG73c5cfq7MCc7Ewh76EMH6svuWWXSyhrgL8b6d9qS0QjfMATxYeovMBdmNL3vw4CF0IT28
R6LFGlnVPhweDsVndMoZINVSS57szGmtvR9vY3mj1rNOZaqHxfiiiH/W/A75yTy3ycvPmLwLRKVH
Q2AVaJZKXT4ht/jm5LHwUPPv+/NTg75I/DnlsSmlyCCT0Hvv6sSRFM0lKhD7P0JT60MJ26fy1ET9
24a32+fF7e8JqKY+6EE0E/Y0wej9WWtvmtlxqUMKNzcLkdQl90cUIDq+IsAzy2Xs051Ed/+SEout
hHcgT1ewuKWfH8oh3wTUH0wzH99VwWNo2HboFKLL8sMs64AtBKJxP6jyzi0cIaRMjMbjv6cheC6o
KjJJcUeCMNf52G7kL1lANoGNHYlMA4rEDpqQEUd+fVAsM/Cj+8eW2OWicDKWoKdIYmHgfETbdey8
vwqiqih7PLe9lzO2hg+iSpngRd1TtoOOu/9gE2cdQP9qaIkIaHfyEiEH1qkX70oAlj7DREOTYJDw
Tv//dXfpprAAGZnnY9N+GtaY5mw1LVwDxXmmvmhOMs/rr78WjjAk0EzDBG8EcRio7yMoyYDLSxuB
UeYmeav+NuC2trV/kgrjbBRK4IOVHuMiTcCELHPAeapYkvZeLwS69H3tLQeklvHaSkMlneF2vN5r
5XempZGg4PRKoiUBtpe6IlAJg8zYTWhF+/9JgkZzQx/IiNvf/iR+Wt4UwF9Tr5Cpvf519KEM938R
MJk9KRRhZEb9UrzPDzD649L450BKQwMDm1Q2IwDuGZp/f0NrPNyPPBwwl4tNh/50quW3p5pBp6d4
7W98nbJIyiRsjRxSr5ZhzMYajXIizLX9w3IxoDWhmhhX73llGH+7KZdJUAJbaJxrbJGpzdb71hl4
4s2sUh8X7JoSPQ83dMBNYkIu0ljTpyeN+nYae9twzbFzFTag4iS8mtXMicntgAEwN8vzQ0lQHyNE
bBPpYVvTLPzcrtavOE1G4up5nuXI0+IjEYKNXHPu6TJH8dvD9A0vSD+aGXXkrhm0tTyKqJTfMMz9
VUPwdH1CDkANpJ79/Gh57XEPFF4PIGIOopow6Nv9Tymw7jJs28D0rxr70CBpoNa2Ytq20JUAYXd9
GYFHk2IAkySmSBevBfjeUarm2Aw0q4+ccMB9i1a1yBcOx55PFB5S+8OKLMV+754RBymJRfJKSCM4
RYrVRqqoDMu0AVay+mIQsklSd47yUF8lV8KdxyLjPcxKlKHG68w0cEoQUZHGFbFmbsb7IDYvznnt
Ja3DECqmmynio6Wktmo+5zqSbrcvAIM9sOd5hd8O8fN5YPa1U4snYUvQBlGLtrGnbTEtY35DqNIQ
YyEQ4CYSyMiQddxCjV/79hCULdYeo1pO/naay2WPuUjx6H27QX5WsXGNorpG6dpF9yIBtyRKlE50
Gasl9NFWZ8TgGlGktJKK7Y0olZycPfDQyQCbimS+dvM9lCD26Xs79jC2EC0zCNBiaGKGwn6yX0sI
PaZTC8fcWuvjMkiFKFvBhbJZkEw54M2Xtx0iBD2hctPHiMsMwxUwytKnmve8425sjTyyRAYZyazD
/71mD80aThse8RbTl1v2ez1sVUuqHlFvSB2I00Va5pLm0qHR8FsrGPqHdKooqc5s9QMtg0+9xX/z
cFj+SLvCEthHdxd3Y0Tt6fNHPVaqTbbgc7f1vZaH+/42SviNZfiyFB1Y6ImIJqWH0duhjukwlKLc
k5McqNBBbXALSBkc6ECfeurXUUYoqYwdrIv0nVBOkXHc8ZkUPFnIspRqQPY+e9cyFK/Jsdq0fKtL
iFv+MiEs8dg9uf4T5XtYW/LYQX2+IqKeKilRyEKFG+wxApuOUCh/mx0xWVDjjPJX+apNszCdarrH
/kjHCJMQSCBNNGME3kd7VQNTZ6g9SklNcdtQZcLe5eckqBnMemMSn3Vx0vKC/ONWn+AcnZsGw89f
8v7xU2yRmw74FhtCMUNBXCXWuQ+hw21GGBKSBK3WVVF8tBsuxwHln7X0Z/ygfSQajemf6K2LYRWH
ao2Xa2h11hyVHJX3AOCBthD/T7HpCdED8FoljbfgUZ24WsMjMfcctu3XW4TURR9gLbt4D30HGnkw
BVBXHzR5NxcxRFGW+AS19HyTm+VXDZEfidQr1kIG0OG8/bheIPChfSF8gwqQ0+pO0Ey0hTK5COBW
Dc76wgrRouzwAOhIzNPtW3AGZbbOg1fUVdgU9lVuPPXYxMKQNns0i/qKseF0029vidMPsAhd5VAi
t5MWRfGQJSS78JtI+MwAc1jG83eaafCqknQfLg1EPOvJRTiwGqYZ2Y6/HdYmm//ZMc8Yb4NLmLx5
FqtW7cXZiou5JFFjPbnfpfR37a64CWSdXDsWgagccczfxxb9BRKsQjfnP2Erxn8SkfmQDcifDi9O
Va58B6bxIugR5h4kz6VMcTJ76dh/jsXzQ6ZkdCeezXeZYaEmT398KgOVRJo4qSItsIQiMyVvGKTD
6OP/9UoG+T8yqj7UTls5z6wvr1IRoKxMKtglFeQnmr9lKBxRsE++NfyQKQ9BOM6TXbYVk/BzXcUq
vY6avohsR/TiMQQ4ejOiTEYu6hsb1ybs18iFAdIrdq0P4ssGyWgZLKbfbBbrgUexRPZ9CIx3DnrX
hVkKKnzyz6wIUi7KmP6/xFUC6kRMCemYm/xiYntgZVGyNy8NlOu+ONIzbpIYL1u+O4gO6ZDePAKc
haFSQOGaZVytElrV6h7woP2b6lVOTA4uFu6YExbM/Z54gm0SX5edaMOMSFsMtUIip2UUAh7wln53
VLQgfApmdQqQ0jQ3oKeeyp5yB64SteTrbBxfzZBZOlwIwuZPjjTqQ9uoB5KgVfTQBllcVs4rUwKN
Zw4H5CC+UpIG3Xm1Hgjv4cFbC7ziGWCb5JgqK5sQtCTLjRsmNMNoiGV9vnSo5nnPvHnA9p/nym/5
YWtpueF0zjSM89xg2XuuAnqBO9x1BUM8CT8tz9rXNaQ1HVKyFyQjcTG/6bmVChhYv1OlQIPy+APn
w+Gi9ZY5c3/UimAIDC2KaMyTzXbLSnxVe1Kl5M/tCTQgqb4fbHAL5NKEjC04GWr/K3PY1pw7V3Yz
WzAGwkgj4b7zrFIV19cRMmDb1YJytf5baemNezfH+WRKvKZyJOH3ZPQyucXSDJyrpR3XdGKqLEht
o/UwG3/nMwjn4ZoeZdy2FSGXH9ZzgR66BEzN+J8ipe8dmodc40KLMGh5T7ydJfxVOlI1lFHS1UJ4
D4VIgAHZRBNw/5x0oUOaE19gR08nHRMQ0eqz7w/oaD0csA+rKHiciy8dotSN2SW82cXwYTHbmcjm
A941HjAvSb38TxK/jwiv4TQR6GFleZ/RIivUkWiWQFMbTKJCm4tzmjPG7LmRDyWMmXwXet3+jL9t
5VjIzWagt2RfIRHbHYZRjlCAW6ozWPmtCfv02wnGfvt2ufcAMey3m0GqrojwYaX+5IJGG83vmdIV
bGIaXGrdBc+i0TNviQjga47DAeXf+K8pxxAxytvvmixOcjenGuL6xDKwtUQLlFpQW+uEr6rJwCwA
q8NznocX8sD4Ix0/NciBKyJuMaKS+aZ6H7IK3DvQk2tTM7l88uIj//4r5zfKHrCLgpKaTJ1NNolk
I4o69IgVL7dx1hYZYvHxK6IZzo6wocNdY2ScAe+Wav7wPd+qoa42Hy5ss1wVTMoVGpU2lYKrRDPs
JOA8QaDw2QY419E0w5FiQDdRO3Ph7t8iYH1Uewg9XCM9ZMc+YHNYD9qnsOK23fkF1EO4lg65hiFa
CuPTbFtmPTujRkp6VKZQ5fVrEQpSBe1rbSRq9ST+TirzB/uACVJB+jV42TQhIyOgC2vV1QCAtVWY
C+u2tVLbK/jl/sgja4MegNfEhetCKfXtiQmAMAzAOnHl82r8/2cT5+DqALv7GRYXgWNr5D+7xzFu
MWS8j2pxFBWdRfNQ+T9RocyiFl+HP6b+S3oBpBlyIItQICs8qHW8mKU+AxZoN79ST5PncCfp1Rpo
xYkgxJNqT4G98cWbYjcu7iLgz54mWqGWg4h8tSLdImNaIR9HCU//sdJ0AlRmlq4/pgiqwoxe7R63
AezPmW/KwGM/s2b5VdkyMFoEZ0XuD6Aqc8vQMsX6e0GEi/nTrRHEW3F5GFf4Nj974wrOtfdfADn1
dgvH1nthF97xxCjyepq90035TXco7DAQZi/uGLhpvA1Vfp2WgtnqMyWH768cGSOY79Q2DpAFkWyD
spP0Kbe94VktYanalHUr7oZOzxAEjHHdG1qIdbhV50w5gv1eRUDtDY72g/u4+NdkiW2x0221Bl8d
IjAgh9eauVbBbBeJFcxTLNbwmra+NpjnnF3sLs6HLRCROfaDLhO5Z494bsBaoBEf3E/o7O2N+Kce
s1nqCxwMUrPWw5E3DCHffhY8x0BzYIZw2Hhyd1HvtMv5xl6YQa40kwJci7mMhboE4HVffZAaucZS
A2J00+rIRfZ5VbqJVU2mt3/XkUoAZTMiaX954Xmc8q5ZtZzTyXv7NjPENwUvWu4thJBe7lcB/GIW
N4hWzIjytMJf9iShQKliXI9ARo/wvJv0cz5++Wan1J8wKdFUjsMgBAT/J6PckIu+Nu0naDUWFKvR
0TBNgzHHlKY6r/c27xLRCy/n7Oe9nFcQ0eqXSj5vdGSn8A2KwYRwm5FfgORcql6HEbzIvEeWIyUy
ScG23YvHEYiFp5oZRW9U0QGA6DAi4TNfQulvM3C5c340F1kLQKeyG05/4b7JdbVSkb5FtbbhgBab
SJ+PZiB4W5j/5vN5l3QtP13lfNZVW3d32/+Fj/6mdcO1+z2UrqRSeNDICwvidNSN+Jh3ngcljWtx
pyuOfgrqIkhOZVu2XHfycOR5VgnlB+II0FU/hcjhw7szu6UnRgm6t/Tcfkwu6msyxoeoPrcbCm2L
VOcgUvJQpnyDBIyIUq02Hw3d8ECk9UhR4gBmkF0UeYY/eQtlLV1gZenS/icZRUrM8aIq1SnSb3V4
2zKs3/ngDc0bZfeOX+ch7TEU9UiyTT4ZZZQ/gBWvV8JGV6+Ot3Fhbo8Bh3WYROtT4E2M5Xl3IMZF
MnG9db1/spfkBOZIyB3YY5sQ+RjXgGsaTXn1PolQ2VrmYlOWeG37owJOrdR8mTwKI9OSbPUKlDbG
+qwln2uegSTI6hZ8LC7ggytqasjYW9wfHkgKgqTjKl02X9RjISYcVWnps/m33sQDdzS4I1T4YJTw
gdGlXeeTrxG1Yr8Up/uRtFei3MQHFLXMBdoIqJD/leZDN5i6h8wFJHGvmxmQFY0DYclayHqCqJS/
mCF8/e3dRmstPdy7a0cd1Jdmm4TsYwjGYVFT2mbyey4Hwe83rueeh4SKMrsZgotS0+Z5sNA/D46r
XvwvU4b4DEqKkTSMMHDNnG1Fxocztr5ZaYp7AqSbNxeq9usFv1zVN6zR8xo9SEqEWtGtcsoFLGNg
wY3TVjAuQFT7IQyvuFbzGkUuuKM0earwAeAPyEp3Gc5cRHCuKcrm0OH66TvkzOW8C27lcFY1+ikw
wb96O9UWlTdakmKQKCTcGds7Isb1lqQfxuBDKUUg6F6Zw/aABpJMqz07gBrtVIXlvNDmHW2ATx8m
sIUH7H0C+3P3jXzPygJpHVQOyuRrwTfCj1Bgf1ha2T0wkRb5E82Q2DCubpInwk9UmTG5GSFHNu1M
FeA/dALoEtIwjSJFXKHFFJDx5pxGtV1On6XTGoXKMAiV7WoSg2n++uFhk0bqNGgtov0bxVx03DhT
IB6ix6ekiQl6ozG9ubk4xeSxZksqeEw/ruSOVoY8yIM6idFMSISsFG9IMDCnW9bDm3JZZlwuqJCY
zBSh4anEoxjMhMDzrYWgS5YW0nkWld7rJ7iB9H0HpDenSx+YvIY+ccg1rseC49SDu+ukmeVugpuL
W9DNvnWTuKILio5oZf1UKSLmWkYtPzoWf+jl+q4ZCgMMQ/EwJd2zYoiaY0sI87W1QH15bCe3ed9r
ADKyfPoJ8lg7XDP1YTUID/JhDsLUWGK1DCiX16cO2d/+XZMeeKwCbKwxEn8hPA4OyKqfp43Ml8fd
FCJz7un8vKy2w+5R5Sw7NFhOMzepvS5xCk0ISSYpMqkCFvWrQzllSRNqJD664G6w/itAQhBYq3XU
UofKKhFSIOPJJBealIgSQKF3FxlnJYm+IaLYwy4xGV80xSWr+uLZuD0WHSm8sKNY8S/+zU86nGZD
Vl0I5ciYsiRQNXZa5ibvbGChms+I6NzvfUnddmz1XKauBg4A17DxUPqF4nkxR7fXiXxvzspi8MAM
xnI4Vphljgxqk1uNHyRHB8HmHXRz+6kdMAtJssW63tmZp9wEQ/a2YNp6iku+ETZoN9NM/vrbHmXL
6MZULfoRi9eUkDnRbBnT+w5RyEIRLrn5VBQsKm8XfglAYIwPHrbwUvMg56irhO3IEbSMAWrqx8Aw
kc0JT5Q5mq8H9bTLwFrEjW+rQkOC80s8PUf+wDykSkLqJJhSZMtYglgRT0YCrVvi8n3gTrbRPM53
QLvsG0npLzL3DwctIXg4E3+u1oCFlJpzs5I836nlORtG844bhEeJi+aV1Az+m/sDcOt7lpEzy1t3
c3a9x0L9SJXh+LtwxrhVjYuacPrutdjn1xuaLXYYZrM3fEF6L3I4lrhWCkJGZwh5dIHOf8/VnW9O
EdlsSTSyreR0VOP4ptKcX2jJ11VASb1vug06GM66RWgERb4uaS/9FY4fJrjyDkEpgnz+6xv3mbsH
jYdK0REdxVgkbc19LGjkHRVn29SJpCvvpNe08G92Rrs131dSmGt2Oxi9jB16vuaPcAG6z9AkyBvO
dU7ZvX7see1GKRocQMS6ZMYoVOFvofL0souCtMop6GdQjVAxt2F9rHVa4MF3JHeiiNYhSvjN/La3
5/Z/AkTA5PkZLVAwDQxg3fjiKjRfvS4d5VXw6trcIbpctLuI5mIzwMy6G3tkTFNJzeG8Uz5wVdh0
wCl8Xz8kHnoNwDtnvo+kjAoJ/sPDIArRh3mmWRUE02rbu2hFWoGJJn5VdD106b32IJPqMuOsHrb/
nAjicGMtZxlT2/vmyRAbSQG21xGcQcgFZURcygkpxRf0H4j/cfmuRO4scUzKYTG15hQ1DhFxmMDS
Ylkxsbjas5aReGbM7+ySoj6DCvtsP7FZt7AcaBgs0RXatcpifUcdh2rQfLxYT0U5Z2VoonviDcrc
XFV4KOm3euShYRI7wF+LqBbQkK3SFoapmTsNCjFCJpRz6+9X5WTF27073+7aSCxPa04Z/DobUxar
+wm2aYZzcv0vWHCMu0bpI3vZup90oTvu5oD2JQbPpIfOOzTUMfaumeX2aXHB7poC+nx+Mq/FzvmO
noexHUpJQ8OqOKWMyYaG69shtxVYLSoLffERPtz8JcBhqrDtn8PBvmpLE2E9NX1dE5J+2GmhSomH
jTM6jqdO3XFaGrvnSGFbakd9JnBdhBfeOOrWAbyj+k5qOSvLEH3x0N9tsKLa1kByhPZzJ4sSVToE
BC63sxK+WopYnTPPjSsZHAgKVP+msde6dZAa7zvgxXrQR3/rO/Lg8vn2+ieGKGeaSIvLceUzrfyr
VNYJ5M7Lo/VcXGpACkALFUtPSEgZr3Bg3WCBPKDGdpQdPszm3C8tmNnRa/FoWiu3OONz9Hs5CbnP
yc7k4pJ1pIaFs818E8agAEVSMJGeVt7SGpUXmsDqG14ncthQqivFFQ8/CaWKn641ANiqVmelmy22
WXu2U7oUFEIF1QMmeauuZStII0McMZA4UIMQ1MRO+jTiLaQArMEe9i2KOL/sn5uf4MEWulahW01D
3w78trC7e73a0zRI1K8CVmwa1XoontUbGMwFZ4WLl6bQtxvetGa6KLJlDyTtP77gKyTkdZYw3eAJ
3AJ1iztm7SfHu5POFl0fzdmpQ2ZwEzXeX5xOd4lWqbyzpPUfD2U3A0rZpE5hJ1hXG+EJ+fZcTonZ
FnMsjzW80LpOwcS4gzdY5Dj6vvf2XuUpuUyN6ffGH9Kd0VHSQ0VZFyVamum8B7GSgn63B3PVIYCK
7FmgAmqAgiX8rHvNxiPfeD3EfZezEPMMbrUFW3wkQaIsimL1Z/7G9tZZK2hzu5V8CrqGYzOEpT0X
NOi5+XJ/zBaCn/tR0rcg0L6oXcYHPUJjMkrFBGtXXyCWVw6qxHvVqG0hh+JUnDWWqZrA+aFaZHzV
XwKZ0ncUaNk+8s5UqM0IqE06wZ+JZZ2KjwAXGrAggMOBJLpcKxsO2aY5qeAAHdmBQ7Mo3656HYzD
SgwA4lc7BuVGZhprlwCCh+Ml2U76JesVxANMO7uld/DCCjXU4UTaEfe7o9qb9znr8VsCERoC7RvG
Gb7g0/nyDTjfF5sdWzaEsbVNLW57jHwCRsW3H4UiYH31iTEN1G28kDq40dihCXECGAr8CNIoev6y
s+NqEESemArE5YMXgouyX+RCO6AAnFTPY92aXGZqMAWh2cXZHURUQhljvi29cY2MdXR1V9PFU+qz
sGr+bpd3FejzpTskcymyv/KBG3Lx+jjz515EEUnz9sRMQXmFoeKxqQe9FGqx1HABGZ66Cm2w3Emq
9L/uXUr7taW9/x7qPq8Ca8xybX8ahGSs9uFpxg1gIBj27ETW5bqcWz91NqUV50DMLongCgOCmmmP
d+IiWL/XKHGvH4Oz+yWuYFzBEXCDIgPEcmUZqgNihgGZdK0zo8vo0jLmv7yTTcJ535QIlE6yhlRN
3+01OJtdBNRxkcs/o8jjcL+QnFG1zUEauTl1ECkWAvPZy5o5QRH7bnep/ZxeOSUlrtmZMsj8SVpT
a55YOCkSugnmgxdGtdaxCjAk/610dEnkWPDflHyl/KYjkQa/ozXCifQKqNFNQi4YAx3zXMrR8Qg/
uExYWh7lIqOO2EJabppzs9S9xOzJgXPwlrEOEJ2gxS/wgZsYbk46hFfM2/B0AbfwMaKpy4jEqLo8
YYhOAmo7q1rlMLdlgc+pnuGCgQTGvdBVtGr0p75LxXNDAu7mfBrHI1WFx83Pnx7sQLPcEywv7MHI
SUWzdquEJrQADQbK5UHUqKvdRnP4GVBW5g+95DhhUUltw4uLYrFRikFh+kgTG0v58KxQNmui0Agj
hHNSP3WCZQLYxr9G/89N4dlNttCuZI5GWnKYGh0RLhVs+EgSTMqDQbmyEjrMbGeb0+G4WvaUvy93
QOcquMmy8cfxGTj8mpoGCVAD9ZnZHFoZr/HdGwE5TjcbHPccDkIUsiyfGKocq17vRmKlTrFxx0yx
cE1mdRCS/qdX9jF75VcwoX7U0wWdB78ca2NcEaKU33dZ7GOreHSWV4isLSJSHIqxlrT6+LOQSACs
vVyfHN7dQyfoZw3T2rbjxS9lC4n1Pip5nxhz81WNBqKdIWEjRKKrwZP+cB5R8aNybfd2IeFUyXU5
e3R9cARGeo++8XBlHweFI0w1ecp2fnS9yHMKPZFcSs1e0rUFoclVZ/MeWCSThBqotQwID8qGPYb6
t1sVmWerQjZbiikXjr1jpYzEKKuckJueIQFxCNXs20G5eoXKWuNW59fDHTn0xeg6wZMe6m9ZVy3N
MrlM0RyQGXtdMH8DoGfv/HtXF4Haa1hbedqw740Lk8K7l1dYQYtHiBIbfhltRFhM72oGplL9DM6Z
FFj4eH9IBe4HAtaQrXrFJVEH9vsCqmzmPtj7tsUQL67bwyYVy8K8WB8esY7rd454c+KRB8z95yNC
CyjLqX2MiY79TqgP9hu+kd03Y7+NJim/tHHodU2u8Yro2oM3Nq82dPZIMHbH+fSIvzD6FhNzTA+4
S58L1whQKM6jPPKkrqMyAs9wHIbtZOQA3NiihG1hP5vrmcznP+ZXU3R18C51TcTV3E02sLdgvFdc
gBh7UVIYT7QEDw9eoTMmGvALoRagi5URsYx/UQB6ojY0RFnXlFGFaa4psCPmg83tKhIxiaz8R7rr
PYR6DiLJP5M8rkIkIZzAjBZl5IqT1JosAdRn3V6SrNkCmES9DWu6aNH/N2FVT0GLH22ec4f3s17q
4S5Vh/SDnEUC3dWJbt1dUxxU+WdnbFSmFpwKWf3C/89moeSFjj80JwdsFy18dzLDDG6XMWnjJPuP
FguwqKiDsl3xuhpPGKyhTbhuD/s4E++wXsxTVM9NBc57QSAhEcEKrz/gKlrozPo+dggIKrQt0WOB
ikUtst8DCZigXQjqE629oFyNu4syD6L02JMp7VMbSgadsxthX1U14DiBgX4RMzqBZ8mESLdV8NV9
Tx7NrerWFM3cF3lCzAA6FnGnm9c3Z6in19FLiY3SLBhgNjdgiRBX4ukiIqJo8UgOzS5htUNYW7i4
8Wwb/bl/BFeHvERa2PvJWI5j2UhreGpWz+N30zXN/tFHp9rDjkBTZ6DT7SlmbYVXAhEtoC013n88
bEDJOctT1E+6TCwa7sOgTjCZdnefKGU3EEH7CE1n0E9I8tB/HUyza95ZzofhokBj2IzyW7ZM54+h
0YgyHgT0RyN7HQADSAcQ1MKHCpY7GpbnxhKt6uG/BdgrVyYcE5faBQrm48VtmFXYpKcM1choE5qG
jHFm8s59eXdheHvRcb3sBof89BbiUlv8g9G3HiVDmG7DKKeVanJWhcdwXK4lGkyO0/0OWi5GlqY9
hXwLi27mZFoVSjsUHg4up4ndWNyKbwo+tIO+uIjT0YfdIBzR3Pf9Ehk+QDHU8lwxoykXNqolOceN
lb1Ar2+hthu/Oc69BfiPXJGNwRThBUzwJTJQdUWKti0HP9sKFW/YoC/VRMh0KTgcHlAIT6n5+1uM
Km+okYFzs76ossC69z3zVY+51Y4NB0JBoOfSOLgFCIKJguzYGgNkpAOwZmTZ4VTcdCExbz5RYTWf
J+9/akmnIZ9AAUCJSE6FE97u/sGt/YJT3JQVnI2yO/i7MQwsaJh3iR7qg7gETqv6jaP1v8fUhel0
fXdXE+k46bqzPS7CDeGBoVTAjRA9KcwqpOR3cTEJO1CdRsVzTUyAu1/dY1pDDRdv55J5QXzx1FRI
UuSF6OtTxmxrnqfUdw84DWQOyfEG75UtbB0K646xfjlNx2d4+vfOLbz6MTJOATXyElFoeE7dwwhT
/w6ejHuwHbLdgN30fA9rg4OCoMEaUt/Qh/2lfCo2nAQuJ1l0JRKmlf/Ofy3LQmUK16zjwMWLAh/Q
5ezQtmvWjISNf4BQCY4iSA7q9Bavrf2xsmXOfCxhExYc1AMdmtW6y4hiyLKMhT4dxfViCRJPSsl2
sp7qDBVxJwxcKw7cwSAuRxKKwUlajQQPpzu4CO3oS/EIfCGitk1G4iYh6qNiam9UZ5yluoB6AcpI
LqIPJp9gx+uJQ41vh0Vp8rPFkV7lIvqo+6nwItRVJq55BxQ0zS76xxVOEvoMRrU2DYUkEJLS6812
cc2ghRKPP0cwYJ5s8Bp1sCgiZX6wxYA4wOghb8hXEwpHdz9bqzAJ+uBhDbnZETk+RVSXygwpTlBz
IkgC/vAgxyzPR+IUBou+6dfIOYn58uQjX+dNCMk1aCaDeyqptAP4RFLFIIZJlmd8qmideiKu/zg1
5C5PAmFRS6IaDELgAgmFBS/rkyMLR2L0BbbkjaBw+l1XI7jgf9L9tLNsehDaAfmaty3+IGW5EmcE
/TASPyyP85L2imHcFdAtsw2y1KTn1lXJNSNtV9av7/6PuTCP+OVUfe6NjaYLPuQJlGeJ9dy/Ir7O
KH6BryuoG0QN6jtQ+6YHD//0IcG2xbBveKL0GINXTzRG47kTZN/zWZzmlFBFOcEdaemqGv1/5/qh
sQqcZq7r0XEDYAeiMl6LsUCgvgxpBHalK5oCO5/HMfV+DZAW4ZQ9HsIYxxYeDrnR6h4p20FHlpNj
ihUu/9zddiyJNrFbKW2euOQh8r5FHGx6n8uNiu4kX6hmY/MJrmaYorgm1NSoMfCcze9Q2CZ6smAi
sWeSY5a+5pXhcxQRYxdXQdWyQn8tH7PkK7fSpzvsH57vhPrHQIoDNSkIqaSfLzsVu9Zke0ujy3A/
jENfgZixW5XVE+HgqrZo1TdImuWwTG2/Qve9MzW1yU/LutCJ+GZv0J4HMrmtTDtYsgEvd7eVcZEm
N3dO06dIprN0t1xJD0WDIW6Fgx3zNXbkXZnlV2WlWmkJ6Lt9UUtilC/W51GfSLPdA0PYi/zwLHiC
EE7yLI+iNu7I8bRbYbU9ThiNgzk3fZrBb9vhw65yyddnGVF+RZj4hrOmRiWmT8Fws69Hfz5trPXj
rFFYY+/vsdhPF6hYven/X8SYoPltIqa+pjxAY3HFj7OQfugH3u9NdW57tEmGjfMwHb3efHNLBD0q
6JPpc2Pic4fFwdVvkVFdfycMLR3da99cK8yoQcaZbQZRWbVnhmpjqlurnEExhCTwCnZp57rGkzDY
g2R01yFseYvH/zSL8XPoJlr5quBpkFMBEdylyQTrpkAXESXBVcvErHqnGzSYbfFePri02ROToKGx
hQic7cuuxhbCJi3rarhyW+2lJR1eubyvyNlS//hyeA7IBrv6lyxbOIVc37NLLMIrepPPVmIpT80h
qWDt9NO9iCGihMYg5AMIuxIvUtvJEmt/jUuZ6WkzGWc4PNSfwicnihjTogxJhmv5jTpRCr+l+K2y
NVh32kqgu9AzoIKxPwH5Nvdutniol/GSN4cut4tJU82X4bnh13zkWVPEtKLAnoJgPn8p5D+RK6yS
8GXmNgiTupVpY6993lPeqdq0JpqA5htnaU3f6a4179r9GmDPw+WlX91BQXjYbONOBwKmgqqy/0DD
g6M1PAhKUB2YC7b0M9M4GHO45CWvTXmpr1pDcVFuMsFVge5HipqJp0I06As80nvStVYnwdb+51e5
4QVCvKcweMm8RKg7zsjvVZG7hFOIb3jQyehJYeJb7KQUkBO/N53bEm3X2wqF170KJzaLw9EJw4RI
0WU+N6NRyeEEgpV9/HX3ekJDyAtl5gesWaTZ0f2O4h0/ANjgAvI5g6it3OOVgZkYoI80sn3RMO5i
Vg60AMcmNfYjyw8Ky2qyYe/MAGFmYlnCi77rGkCT/lEdN2ankBQZk1ljEv/towlYpbgS5amOf0VI
zh7LBLChZT9rOPEKVs6H0ZoVBZtyOqdCoHT+tiU2Zfts39i3/8h5/A5hjplcYe8oD++vkFTSMHA/
bjm7pEhbiZxIIc6tI0PdHrxoPCh2iyM60yfidoeuUBSTPtjOhjbuI69ZMrqqe9Tod7ny5F50I+OB
Fk4ZwVGkJ2sa/R+4mBWkfxhkNN9TFu2AdGow0yKINOhKqj9Pesp0wDONL55v69jb0CJvmDyJN1jt
aS+m6KPXEtq+ICs+A+xsmsnRRJYaYalEE+vug/DrMGVhiPCA14PnN40qwnYLpMb1tv2peKN0/dOX
XxfYFXV3w21ylIiwZGYBepj6AUnA3lPrBWomPGWICE7OB8pmtf5VNCSNKcadxSRf5tl80gc5Yk9j
2aSptjcVe2y9GEcholPS9hrlB97rLvW7d+8H/Xy7yFfQxY+ZDDdOm6d/FTciJAy0UBfUnktB7152
Y2a3b9RQ+dbrjmcw8HNFn1M67t8IgitOqGLniRZSqS5C3n1It04QdTVHQI8w+y8I3wPoQ3xwNZAg
xDwnKapGPFvHT0xM3StYY1t+V6wb81FbpmsFmu20kI886ulTNmdfQw/HvpBnBMusOvkWBjH/ecDB
j0BuFxB/y02G2nFTN3/b1btb0ECzfK6Ljx3qN7kbBqy0gU4fU5wo4n3vm6Nu/+FVNGDc0HkJnhg1
c9O6lCkoLGVd/2aMTwczuyPG0LFGsrIxinNHt6y56L68koIjrjvxcLQ2Q4IAkFRW54y5oypNcZaL
i3DIXiPPcpUXSMzv/KalvtlsVhD9tOsCcAHipXgKhwUVPmBAgdlCLIRDnTnTxsMykOpyYVHLLoyt
ulGJA6+l3xRnVRHUHrsFjyM0zn2IiB+Io52SmvEoS46b8Wzcfi3NZJI+6PHwVPNNNdDuKh1ZEMxb
ZO0HfDuXqxcUOdeFb80Y1/VwZ6qJDSIriEhUjfvbWQ7dAPakIryEWadC+NChIMQHYfsXq0NoVZH6
lnDLfF+TRAj3pQUvIHEe7BmHr5NOCfGfCtaDm2JVUXaBc/Ogv3W9f2Ns3uZwdKch/ZvOQ9MqGY3Q
V8lZdWp7/qfpuzR3CsAlTHSQAgZW4FjsykLXnFmHlSZinhacK+Piz9860JcSbbg4AG3GbEstzk0b
mnBzQmrqNqBiYkoCAm6GEaECBxOcyKfWaHH1QNkjyTk4h1Pl78HmAKz9EHqlsb4epV94x08RBRRt
Q7ghh8oWHhDbyNUOQb0piM/ueqMQY8Cm7Ph8lIvca07ciThFiMobbAk1K9togUUi3UhtuzoD5uUM
C0tBRRO3cux4BzIbdBRysrnicvBlYXhg6brnTXqIbW/4Wc7ctmWxu+I858LIrIdDzhF7yfI3QawF
l/V2/f0eU2YhzmL7krVWbN8YIo9dos4RR9loYVDgr3RTNHUkl2cA3GfyDqyHdrzcjJ0ALDq5reGI
TpsEQZ0acu3h1jndx1R7VN07HJ77KtVN02PTX5TNGbqPrOEHAVls/DtmevtvR8dQqdta+Y2mQ1Fx
r56Sap7g1Lx+RWAxMmXpUPtS10u1NJTLNIIzR79TzuuU+xGaH/Uf2XH/QA6JqMdxip/gIFsOQzZ5
aCRBevsUxIqyAtAroOWKmuno1f0O9xLH2jnUU/L9ISnDiRBItGutkJquCH0KuyAD56cPRETKk6Ub
Xub1Ctq1MOnLnVFpslOh7kqMH1+5cJfu5hGFvpJWTgOCMXTNhJNj6uou28MhId/oEMYttVnw4R0z
RStWgWac9aBuGcj53Jn1EUzCpK+qsyJxPe0fawxQKijswcbkrmWBoBB05rbblXFPTMnmvjWfln3z
J5TxDhQWM5h8DuTbAWsqy3t6Giyw0LIAUhtmjOfqTZo7hBG9xYENV4JZ1LnAa866yBELWWObZj+T
+I3spAHZ0usSbN+rlalmr4yPG9YQm7eIFoUQgI9zV5lbgbytmWvut7MTziLBbKkKloZ3oaGp1c4M
MXZFCZu0n6ohw2QZpQBTwdDVS35Z0xhAyZmuEStNWfA2TaZPRfbOL+bQSxxgjgbGbRn5IjSZSRkx
7sa0ltX16hmIbBtZeo6kumJwaz8bfhARaoTUEomJ2HH8lHCylI0DTcax4JrjaOTo/O2V2vH3JIaM
78o5rmD+fDKvBKmYGCphrfxSFNJQxH/65nQT61QwXJiTivQ4l+ONSHNWYfQl2ErSUPq1s34sM9yK
9YSvuWi93vz/1ySjoK+u5GaFrmYYPRMqr3VZ9FXOMFhUWnchrEYDLypsvhPEdBxW/1P4i6lPW57I
YCG/ol6phHoQlvjHWXoIjhfQjS1ltwYXrjEvUiVXQwqdiHHwCQsS40yL7xdKV6bFswCC2ZM3CtV6
lgEFQWOpvdIAK2o09cd1TchhQC7U6VEVHmyceLxWHpjnbGpl06XRa0fNoDc/JpQl1FpRrdg3tQHQ
yZDUIkubDtF2DtTJ15NbyrQdUALVGw26IVloeEl/f9cqRn4i1HAlPxm5mfbq43JSM/i724+5e27j
ZApEuttwZdUHASDxuz8bkxOZ21gCTSaDfZSXd0hNVN7smD+b/+5DZnIDOrcoP7InqKiKDDIv53Yp
6addJ8CPh35wJktM0iiNJaumg5x2f+DwvxXWRu2clNyIreYBthecmmGJNosIJlurK/hly8PKpNed
xUVygHf2sMWljyLkQ6bamq+udZPe0HqbZyQO6DTdLA10yMMwrdei3AZKgFi/iQB9Zc25kFeYFxV/
ZyTCHSI5zoSIRnm5cwIFqRklYKV69fX+/gsB1Oig9d9Aci1joJ/47NB35+hrCfWQAGkUOH+wmxVa
s+iMITbKk/lqZHMyvY+L1Ac+OcFV4bsdEb9kgncrLrXk1LIFBuplv9JoEdM9h2Rz+gFUC7YnUmGH
2wBHchTVbo1evr6ztdTrbOqxQsCtax3SNIZ1stIh/r8w/mHhW994N/j0Mzsmq7tOZO4ok8otdEsH
II8ke20vXdzQ4+8cTHmRbvv3G4c/j7Ylp25CrJKaakaIfXYziQsfxxn2zFrmGs/1r5YPRyEn9muE
uR6/lRhgveo6oa///nvLrA1ZnOul6CsPyo2Z7SsKYN41I9lWXOxPGUfGGAZcpV2gpPLYZiJnfwlu
gk/GrQyRX5oL7glJzIVhQ2DuQBhDjBv1BKv3QO0Kez40/m264PvKjdLBQ+RK99BPM7PEmurHEEn4
yRDaoT9evDV6urux7odHVAetOkxoOf1pTz1BpQJjP/HJtVDJ4cqcqpxC0h4CFaWOlW/6OEM4O8LF
i+ludBckNIOlJ39nJcaqRuVh85HYAeWYYqVGAHyNi1xhwkR8lF3xSP4/YKyrI0if4NXB1ujg+nC8
TL779lVb6L8Owu6KCL34ImlRsQeoTAPc+TMqzN+QQS90NAUV2ZiOLKTm8ewqJgbzqiW0c7BewNHb
WTfmytbREFxM3wDDZshKWlWuQHnn6Kh36OHHhZAodIsj35ejMy1p0uKNcZmJjEHhlRR/q/e9MABK
Maj6K9L40U8lCkdu3mX77NydxQvOnr1yHxQZUhn5uilhwGStBHo3DrI1md+P72SXKzy7FrCWqHav
7w+2HWtDEphEKNTLDVUTCGZmUkZ95gjY0MhJoHvFHIc4qjBfXlxlZj9s+y1zJB5d7ZFjdiJp3Y9S
uUvVfw6aAq6+nOJOSfs4fPHsDn3XxmR5NZ5KNT5lIEFaDeYKwSq++pUolGpxqHX7+mHIBBY5Kxde
GwZB7jpG1kxWDYurDylvSd+jRBfBEb3wrCvSUxa4Cd9n+MRActHciNI+n+YxQhBQ5ga8kqK+WM5T
AUCZblB47l62R7CKtKgb+nJVRsqG4EClmGCsNGYs+q/dPmwQHPIrn5LGsU/Iw5ckppPVIb/eXHZy
ZB6nPwMTfXb++epcIbyzxpbsKqqSLxPTlB2lJ17NrDX4ltf1gqIJwj8f9GVPib9+M70oQDw+e00w
tWgzMdAv4QGuTbgKKIqQrB7YhsUsNmN4uErSY9pwHsOidj319dEADt2ppoQznavVuz2TZygIaMNf
yTxCG55aXdAi6juEJASdpMuEDoJDpqgjLtu8miWO6KrgCAzjUeM1RenGb9m7W8DarxhL2mhJ7sg3
gXH9belFL8pMW+/oSpSJiCo2Xo5Ml/1raC79E2hJVNI3up+vV577pO7XR7fR1U+egHmdVZkN0i98
GIjEdhUMHvgcg/sLGKqc6XG7W9OKwgiSyoBYlocbNzbaKRA9yUV63aDNFBwWiwdXI7ah/Rz/j+3A
BIXjBZeakmQ8a4nLVlimGlEpjdxPZqqHiIyGIe25yiPBIDSzUlKPpQk/OqgE92AoBFL3GDirBOm3
BDPNzdI1CEPwCAhaytbyKjUS5MN9JRYelqfVM9hYHJkOuA9rBzGjRQraaCvTExVtvFVTyvOoDLGm
eDOSRtfdnUfE2r0EfuP87veZbCfq3uNzAUKWoV3jc9cNzeH0FqyDGqHSjbLywrkxpNFENuPS8iVE
Hn16B/A/Kzr+CXcCIHzO2wP0Wvmak3/KmrCbXdnPEPnIFWPam/txVswdeh5cxZeIRt7KPM0Obeav
6xgjXOFyHSKpw3QIvPwTjOhxd3/fqjKaGwDvZDme5RosbxwGCR4uc8RW2j9VEOVwfirz3jYYK4q2
mGS2XAz2FKrKsyJ0ZBO+35EO8Rf2BvQ/cuVn0/6Sp7h/vkEvwa1FUQpHTZYtLHb8ycYu61opVRY7
Nzk3ZCvZ+saGGb+ECo9SGjYOi7Ey8cwB10XlPpUBtY7PfemulYtEe1WbExKUXMu6OOiTWLcdb3jF
eXo8M00xR8a/6qsDXo/PMjRw3QJinakmzASHx7aVlHBvlVncIR/iNPq5vPQL1w+IAz3s9hMH6wW2
M8ctnhLLAymEJREkzfq4iNVTcoK64XDBnPsPtrOMrRta8FlHiero3OpxY5h51bLbtJ2JJ95AQDZZ
ndn+whEuTXervmPwaVR2hDJeFloRycuYLWwMkthVPaGE1dJY9kKOEmN63WqKzTaoU8L7mCEJGBlP
M6RmxKRcAVJo5i/XjYFDoM2SkHqI6JR61LM4Zlg0gvyvIs1WkaaTg2Mcpyj1MKo4vFcrn68MWU/Z
kbefszmI8eM0XyVHptAVpXdGKS2DJ9p+T6MzzlDhxbiDJHYykp8JRByktm93s1/DKnpACqYst1It
p0CJttwIVdAbYYWCBlhAxJuKRDQcgDjRb0KgtxRhAYDjkB1ufLyWIwyMHHnWmP5tHZAm7z/cdEeX
Su8cB/kMr4Ch9OfhoohY9UvcEaptBIvk8pZCghpDtiWqXYpG2ZxWhdHB8MX0SergJBBgTaozgq4U
VvErSqPdfU8CKHA8x6WLfbhe7+k6LneCDVqXvjNswKHD9gYbobVl6XYzbY35vQYkX8Fupt/eKbQy
xHuhDOzFa6YKbY4uu4hOmXQu3Smoztvwx/HDhbiFLV8gl2NgkByhEG49dUxrG1qFQT6O5msYNdU5
aHovQkahoAuzipzoKjNJyxZisXtrwuDr2kjC+7LwwStw95H4iRZRbkn7dGGWpEGsVhP/DQpum1Jv
uM6a9gj9E6B1Xa2QV3RY1IigtUSRv2y52fAEHPVw/ReKA8EXbKCDRYy6JQNcZjNcFqH+yZNxsd9A
u4FxY5zogyu/rcZVsMOucfkY7LRBJ15QjQHySZxfb+PWkamXIytjhZCIxVXXFURsPujCo0kr8I7M
KQzRzai1W3Rr2jukJhxJRJ+KNlWD4rTlyfymIU17nimHjQIfddYXXIimFUnykAtCR8m8BqoDTc5s
ok/btv62SUAve+SVLRuS1uPGVcgHKye22eARnNYQARgmkd1SjnI6F192bJhQ7w4pZJ1O5qWQoqPT
SCAmQwx7g2pz4wSIPoi0pM8eci0q1ldtkmHX/KBZ645lzo4+MR7urjg1RsK1IUndMYKbIkJ4FSe3
D+DSFBYGPhPKWEWku+x5amUJnAvCGLHnwgx/aRbqAHAjGuu++cys9G9xGVG+TWDeWgV6ezIiMywG
Yr9hbIgOEWOkbG8Fpsvoh0NFMjUOpM5JqIq5jorBrAZ12qrYHHGYEMm9MUjXkBs5yy+vKxzn88CW
3+r4FDrVaJffAr688nS4nrSyTFY928w4wZPVqqxLmRuzJ/XgT3Ym8Nf6iOIbmmj3F3gGAmvLPw2j
Do4lbmNhvilNWq2iO8E+QjxSerjq+A1+SULL/ooPelQLCKBx6DEdzrMsVLmIJFlnC7YU5Odg3y+Z
boWbb3HtAW648wc94Xs+UJWXk5LGo4FYD1y4AUqeViusER98tLl/OL1NvWliysfB2O2K6niD7gN6
FpZz2zwnJH6LMGbuWVljO/jmW4BvdJZhDn0YFKqJCjWU6SAG8s2UU+Zuw+ZE1Xe3meIwVp0IAfaB
AWJOgVnehSxxAevgDaTAMSOQhmL5W9TWw2q+qq+Cm8SNu/4q9jKkZDBgybAyUPfQOjPiMa7mdf+o
UIKjDu6CawUfhz1hGfn9oCKPNI3+1EZZHdpnZ6X3bvfyGEMf7OeiSwPFu5FE1YgqsO5FWVE0xRS4
bIZ5Gj+vQiDwytb/UPCwVuNNXkOOI0o3aG2L0IOyaVUbYKp6+JGb0MnDk09fY5tyFNAUVOZ5g+c5
w/Ub/ZbM4vY3RWx13JnPcnffChQXxPE3YBS/PrS4n5cmVN5FbMo/iijmZLdKaQULuv/yW3Q1FvOB
QwFoNxNrp+9LiWMFzYdo02efxXoMAh1h9/Nl0bPvIgQFQEfgbnMwhwf22wqON0LiLd7d6c5gqZbC
VhtwHEB9vmc93Ztmy9X58Ixiqr5ncLIC+o4mtCdIcrNptAs0x9X0ZQpTCEtDi3/Y+g1Kbaof4qq8
3bGs5UQK9Jj0bKHmhuuYlejBUu9PhGLzUf8zidaseXrlH+kf+LZKr/pfmVenyhqmLXGz8i1HJq1s
/nC6I5YZ5+kOaKTjBelu1Zzn2cxQ42fJIdiA3lavp3khdgXtoGunal8whYhky+8uih7ReGFt4fUA
0mYfBEWQ+pYY6XSONDlgNOi2PNomzHIk/vEcN6fNxG7fKbhh/hnNzx68Pp8E9JqJ3zEMJXVSeGoo
sHF88FJWCkitLf9yqV1jxhiJT62lsqY47arLmLAY7maYXwCSO5vAI6EZe8Y/jV7+ffjHuxUMqOS8
to/UKyfWzi2tZFhHBUEdZw13CkKdChURbGRCL2KKgbGUgd93wzkxa+JQ3hZUdoyuFi66YhiEaN39
V/CfLKEO2rNZCyBwahG/qCvnSRsgy7OAxgezL0DpqIr0UcfV6ZIfebVC2kMpw8Ldrt5PB658IGnN
PytyGWCGGLdBJ1GGHIfj/CafY9Q3KiAthQLCJAcShU5307TI+4K+QL0VZIt3F1UWHQEbWecy4e/6
zHVC88c5WWvl5bnpDHcpIgmDR6rmr2+S3i0XVpQ13nSo9o8A6LBUzwRGVaguSgrRMGjypbJ5bOiH
Is4TX7vbpz15pEySZgHrPdqBXxTOh8S3MiSpQ2myRyk22QxHiXgMWAhIluZKARJnb+NyVZeajm0S
O15x6aQwL0xBZz4D68oYuz4ukWiBeeq9LMh0ZBRe3zRTFcnm94oXgns5pblhd/J+XzZ6fC4Xgypb
w+sfhWE3KEzkWjbyyb5oqYgVgjAnvVjLTnxynNK7U/eO2H/XRj1ZBbY6IbVvDPgvcfUEzSbnoHKe
7KbOkMhRQ63stkynnVODufJ7u4bg3HG0RcQ2C5cXCxY0Sw2e0hPwIYEssn572dYk7JHFQhdYEldv
VaHc/H7enygMsaeGiUeEWLS+hA59/lH2GtGDXPWpJ/pK1BGEWSRBMb2wfhJRsHPCk18wxKSvu/yF
7/YrMxHjFOvtlHho9X3wlotub1JPeRYAJfFATS+nsrTQ2/Ya9i3EsHqwrFsz5cOYZbkWc1EmNM1g
641KTYkcT/jFinKQ46ahJ63QJbjBlGJfX1qtiWnmxIyRFvZA+uYzIoOr2z2hXr9FIFwj/cArjb1z
OG9dObiC7EAV401ky1quWwi5L149/uQAY4SRy3QT88y7U0lVcOk8AjKWkZwOAp8sLxz09hbb/Tu3
uekhqftkZCUjcvzjTPMwPiSNSTd+f4VuJe13W74teZMGFi70RlrW5ZBPC89HphARwcy1L7/9ssun
tHNmliZIk2LCwUlfQFVQYfA/CMB6ll/5xY0AHg5CQPYLCWXPHXEZpuL87kcMFkwL/x2mlT98yGkw
kcBWf2120sU7vyraT3YKtb3SCSthyq8i1MLKbJNn0jiMrO0c7z4eGKaVtC9Xs4OVyHY8M8xefH+F
FDBonzNeaA2Cv8hEdtZY/KFlIb9nIXIasqKi5pZTi4m7wKSKRN+C+QiBTjdESJV9BhfP2XNzWr5i
9rC+3UO/yYmFxR5Czzl0QSz9uNqHx7iXsWbStT6fti+TLkwvo1ZUxUTUEuaz6qzNczp3abalOgd9
ljtVxO4EgIS1f890JS/QHUuZYCP2cYRHWFZqsfS4scEE4oCsCvsNjEvQzvR/0EAkAXavtutbca/n
9/xH1J/OLfBA24c/ItVI5pRLJ3LPvmCVtegcVqZ9fjhF1Y5BHZQD8yvHEj8Z1IwFV5SFrlpXKrwA
sRvpPhRaownvXy0QBCjYjHeZyDdWnYxjL7/DJZnmybu11cZYACnxJrYKf/FF0LEG1L/wJkQyssGp
TrSPDwLuV4A7N02WOiL0J5asgzvXhDizYwBQYTdKnXIFTE9zneXVb1VXOHWz1nU1d4pBFMIPNXpK
IcIzpvOhQv1AJzkSthzzgf9hs1Vmy9TDjjs6Y3k3A9IfS1KsrVQosLLhysmNrUqahVJJFh3LDY3t
MEb8gRf2OOBtDTYrlR4fZN50Ue704zQ4aSCq+FS3cHn7LWdC9Yh6SJGtJenh2E37moan15r174aY
dl13C2Btjb9AQeLGC6f5sONkAnOI3+rJAPvytEv0/0juY6GOqy8Ts9b6KaETOUv7mdDvD4JgAro2
uKzO31EwzKN+wkyTlJwOZl3Fcgek1ryR3LK9dVSiErMyva38GkIGjZ/W1+v/ofXLudMbYs03GUfU
Ro+ehvCMR24a7XZ3/jhUuLu0wcb14P1beW1/OrOaCizixz9jZ1GPh0gY72UyZbi5UchhS01PS78w
IzoTV5zZKxTvEnbuz1EhuV75B/QVC0G5TPAkJX1D6aFSIdzqy0Fb0Xg/+BiuSCI5dinoLez1xc6/
umzrJGXQ2eMabNK06D7TNrfafUY5sIWEEKxxpmgn2c/jXd7KLmU8JzVfr2qCv1M8SEXbi/XxYpRc
GLp8uoyNyYxPN4xZ7uf9IQuGfrvdwmX6S/LlqADF5pfxBdO8rFOa8cWnAVziT10Se5k6QMnMFOdg
1ZqjsdEyTgNOzlUYD4Gs8zC7ih9yPSdE9vYmzMzyr1+JnXj4G87rRHAfkD1CqrzYOWzbX/KsJgCA
iRhB9x+oE75j+JB9J+czkTR/Y+IvTdMJBXPEqGtRNKhGSUq84MNI1hBEXK41dJMlKX/D1WuWPbd6
jXSSjRMPXfoEYoN18a2ju+SNi90QA6y2yQhrTlqR8rmy6OAqk/pHfp9LgxQeHyMqXGAsmJlkQ/dA
tDeeURzrMWvy/pb0mL63+cGHKk84PZEBZfat02EeJ7wHo7JPEQ8eLyO4zC9tzaWcrBNLE+FxL6L6
Aj4+6LDViNqoVrayDukB0mleo2f2ERKNIJYdGGWkt62EJq3HcQFY4oYgQJ+ThdIMSBpinXvA7ZIQ
NCNuzrqs6Qr4uruOFx9ZuEN0+Z6dJeOx4sRQzSeWELARg7DQpn73ylR15UxwFUS0lIEh1PatDJe+
zfjq8ZNROBwuVqruZ1Qp1OC/nhPYl3ZbInTSqk9TxhkzvjGP/f74fnk7P2qUKS5VTGQKfP6JN4DB
mJzlPfEpqKE5VZWl/rW7DwodWvIVO0O+mxt3Xr85LhE5Y3xkPTnvveHAnYdP9GhcRmeCxX8TWWw4
pFVmvUczbtKhzj3dcix4N4y1i9G2qaY5N9FLOBWs49dXi0fiu8qbIXgevzZZDVk4xrjskd1MTLdR
PLeS6JFBlEnM3hwZvrLYnp6IX0PbyZ5L6Kix+xxkvJBDK513WWajR4iEW+o9LaRmilCQhUXHn0xh
j7gcH7ICIECOmYduk6tKWfJkU5yytr/n0JSjtHEwPYh+dKGhWcVqt0M80olP2k16nCx5Q8JmsVNe
te9e7OvwKwhT5y32HvDQfYnP7Cp7tLxJSYZQoIVcdlhnx76dASEgtx5jEbF22igoCoiNOZtA2YSP
Tyu7hUlhuupb9rRIfOpu+hYj3Rkr7dndIL/meWZhXko9xMv5G68Cs7Z3InpzrWUxJh8MYIEqdlsh
/12rGtnVL0SdVfzdsFD2b5VqMhIZKI+oC2oUIzZVYyVvNNybPfOS4e842x5rkClrz8j+cF9/EvWf
APqlBpz80qNr9qTclYONoEShwyxhdx0BUAEJ3RbM1IXGn9/x74SJ1Qnc3tOvgU5qsokCbDJHULM6
OIeWQdOHQlThi+VilDo9vigr1DH5V5EenBAvLPY22z0ytKkV291jgyNfYJxbIBdMt3K/2EJJuUxk
mgCKUHOpMq11hguew05awtQXzq3JjApot32WkDqPzQJqtSqkSY2pkFA0S5IEMUxecyWJ0VrkmHEb
9pwRILNFBmI3r4wAhRdjuOSVg9BsF6SrpNM/NLQu3EVJArjN9NHHsbMHOgC3RRlmRsfzOS/DXx89
7+bHB58QM/pai9QeD6e5OeY4d2872dlsU3+23Icq6zdqjIb025AfGAKLS2YKsI/Dt3CdWl7n5Ba2
W+kWmTdAs98qKU8cZ3XNqOQ92UxERTWIz9lhBgjCaalz5L5FW3CgrRj7DPNV4/0GHZ5lST3YIt4A
DVLzESRQFqbu0+EM7+tU258EktPbKxihTb/g83DAnaT2gYPsbHvnVEW+zf7WdnmfgZOejO+gEDqr
sAQs00HrxSvTD6eqF9kBWBmgZ88p7n30zwVhRDS6DpYpcSnE7AEBvgCs/L52FvORAiNmulbtlk6l
GG4fKZSMKq40c1oMM2grfixVcaISbiDwHjbZEIQ+UVGBf4neHjc98ktRrUB+b/cC90GkqVZIimhS
L5Y0GD5WQ+oipqxx7p+DhtKZYINRV62cozjDJsizo4NyxBJCi4wMeoyUsQVoPK+nAbpKI+syTQT2
+uA0uLzEd8NhO7Cy43CDXHFWRtaTy6cooELbDE0JGEM1l9h5TxEImdDQRj5h4txFflnf7WzkEwuN
7FIdMEAKkCsWucoxpYHmva13OZ5ZwwWBDgThXpvWxwKC8URrz/Bi130txY+S2iDMcI6GqLp+nTqP
EFxML/N2dvmnJuM8cdAMdXkifUAo+LM+DDS0nUnYSKvDi6NCu1r6HCW1UThUlHpWifm+GSk5iF1g
VUO9KOwXDLVlLPoQ/Ml5ZcC6U7qtfGx6/Vy/3w/UiA5NgmKcPY43IJtBFz0khcuxebNp676zceqX
raEUBRCmYxqaUmCWAwJWtgrF1nI4LRqf829gC5UfBJwwECo/V8OcQ9tqEqKzGkS4r0puVN8F+MAm
zJiQhyK5+FGHu9fmay+KNLf+1j/eJNTbKbL81q+nKn/Jo2g82FLpljS15EMQ9f++9Y2vGY/OPkOL
CD56+XeBWg3CxTraHtvu0vGiDhDA1H/Ss2b8V4552R0QcqDjuUyG7vPAZF4nz5WiZwfRA1ERfixq
MSdieD87GndBm+GbsT4Bnt7F3exmBNrRN1cYtHMg25xvd6pjos3HbOuvTVR0mn7FXL5HFMGEKwQY
KMqdPdch3YrMjwcWfncZJrqydA8fOtF/JNQP9R7HVhixCv+EVrvmmrGDe8ntxHXd8J6ZSEX8bPZx
ucvdLolGQnWIDI/6QNzRXJP9HKp+a8D/0SP4EN+BIFj99Bt0qiYVS9LZHc/eTgTOwv3aqhwAsWnC
JrUfCQ+PZoTfUnjx/FGt/Kcgnv8xc3B5v/jHlXL3olpEoQjlou24eWysVPGI7pn2WXv2xlFUDOKF
rYKhq2Cr882PDBFZ4NEBTof85l7MZcKZC81JOIk6XTCZ7WTixjkzNfrhiYWdVAZI8xCG83+ZzrPH
MziE1DMirLwBX6xsBYpiaC/806F4KI0zYgQEF/cD5e5z2fugsjgzlSaIa+jzPE+C7meIQim1LbPK
/3yOTb1MP38C6D1w6YZZUrqOC6VK5NXYFtirbVlR6tHTB4y1qxfIhdapx45P7FaBT6QnCHzsX2pq
KyDNNBaY12c1RyfMiMDWKJZ/osbG3PztfBg32xDUBhvhL0gLpDBpi5GuSna/aQ+VAjGv77h87gAg
Xm0pk7S0yvn9+ro3kg6NhT0xm6oGDJTbaY1D8oWEsGqmuyEPOVO+XPnOotYvbGaBgvDteyNwaueX
iFLadjvCu+tQrITjRmDlTNVm5LWqEwv4bgVQeBybjjSCZxe5HMv5yXerXn0O4LWNtvwAUqxddNtA
aP6H9E4FM1GcULVGKc5QfCAkxGLVs3R71cEilId+qTliAuzJ/75/a1a7eAhB9vsNDqn6uUcFXY6M
mgeGgw+NkJvP2FC9YWFJkOI3ZiiJlszH3npQQaAkE4XqDiZk4tNZBsUuNdcztCngQ1YeoVdCmWTZ
dMMmnYF+mBmo1ysP2Iji8JRj57Bb8ZxpdjvP33mDSVzCISuMxTRaMvoSrx0goyvEkjXwrssIp+P5
oP9ujpdyJnmjK2Iu/Woubc6btGoU7Vn0oyLyKCDN0iTHmLv5UERZaEN0LFcyJaPgPAlYx6K4NRN5
1CGoLDheisWo64MVyxRZUm+HX+hZGpiuX3HCGfV9j1Ulp9aOyaQHCvrjcVjplcd4rOKqR5lNHOgr
BRZzWGqhXN/K26xadGKUM2s/jOBQJC6ViAsWDJWQ5kUPNZLnl1iAc+1kuFu7dz7+Z6NJTlGNcKJq
oQ+o1rGq2r+h1oKqhThzDdPXWa2/IfPXCubTMZD9mpscd80G1v6sZdTd/tgkN/3Fe7qklOiwRRyX
UG+G2TMDpmWoEsLCTut0Y91Rv7/T+J946yNikdpqRJF2f7DQqheM6N0UzbPDV1XAICR7+yQZyMQU
BVZ0agPWW3fFPvY0mrkiIplS9KrhOqgOrF2RRDDKQM0Jtja9do7tmLNwYjgN1EmmeRdVHiqZznyR
sjn+pG0zHouKHf33Yj3Q03dsUQ7MASa28gpEBDb/jc34jRQrZGX6ORTQo0OfWOWO52fiLMB98PY8
4QGVd5xo3BIeeCb3MrMgT51K45UBB2RPRk0rMiDrRcUYteUZzXSiUAXMtWlXWgQ/3EPH0QlRUc5B
rQXGxoUs5sJwG14kFjF7a7tSDuaVHQuv6oE9G5PBSp0cDTtlX8u0DlECQJs9BwxJ1NSTf+hMfFHU
DD7zHjyac12YQsympL27wGyRHVbhRzHxImqVWsMkFRCBmE/6pFCU7yX503Bkkg/Zb9BKVVTD4Lis
LYhZC6upj8gtBj1ZpSwNVX2pU3Bt8m2+i/Yb2Asqs1zXFPiS078tf1HHmALLHIv0q8tyAQ8TvfVX
krfZEH8SRS7QY4J+EI6G4+kEZ3lAHVCf9zwcWOvKykiCv3XrWXKNUS1weaV52Da5WEQkxLPgn1uY
x5wV7RLQ7+OFOURK7rjpWBCjOBSBfzOaqRC9a3uDJHfW730h9lu6CQxsuFPhx9UeGsoE4EFze41K
6VzaaqGtsLuVQEGVLurf4fAVDKBDN9RAvMWCdLSLtkyTwGy7xPLgGuDNsHOjXCVEVcJt9F/CqRz4
A8YNNTUaTqCLvJnNOF6dy5GONKEUPNjCxo1pplgHovPOmFti0umOvYKXrhk9c/q8NBYXbElzM0Ao
6hd5MtvokSz4BRzpvVx+gNcLmhiXsoj2ymwYUMR3Zx9iJ/Gnwl4BU9ySRRZI2IpSSjj4wH/JNK6x
tTdUe8vA/wQ/wU+pHBaXTv4rKwdPYj0Dw3Hw0fCtO+XBOVm1UrXxY4ik60sG5Zg6VvVIxkwGsFv+
phsoi6sBqf/tQTm02Zg2Zm0yHI+eZOF9d4XhsQJNPvIY6AB6nC7HYkRsaXgENufLvJ+yiqUH7Rat
wDEonL/p0UKLKynfRx3HYmtNPbPakVrS9NBNYs96SC5HEYWzfQrBlssqdr7DI8qrPsLTvxO2h8Dd
dR0UzCpu8WCkX4s925R51ZdOKU7V3lLPRw7KG/ORcXelNUWRGRo9OwcmyvnKaNND7wVGCpIybeJl
QDaILGdi46z9qfgnKICHkfw0NCE2GHJUtPF+wFqKg0l4fskkltS1N84SMxSgEg5Hh0rv4sJhZ9YJ
mRhPj+NpnvpOOZGBlpCzbNcTk4KbKYvJtZnWzfabjUbqnE4W63lbgRJ384zYlzeFbJbsXzGDKY0y
ycJDobTSI6g7GQMesbcid8QvdvvXFqLYoir8EooZCbdmN3LFZgASLO/5D53A3mUAoSktyoLdajf3
Hntc/k9d8K6UeagJcZFBSNw77Evwc9eS12Q/7jVkQpb38q2cDAjEfX39BaZG1ei9vyBCdieWgKaO
k3Z/7HsE8Fm5udL/Psvu4edjKkJoxAs3+7I9Qa5pwTyuOBEIftDH5yrHlXeNMrc683e10ndRU3D3
aM7jAQlQjOC1aC7FNwPOW+UJhI7v4WphM/V9OMpmnwYpzUQvYAN+pBkcx9+o7ALrvQqH3clFjPUB
Fll1p7aIHO0mkUpUveMlVBBEHEx+/eq2KWqrTLtqS6TEIRDYihFKfuQm0gErEx+WRAqG5VPljAHK
UxRazzFEwq4MprLGwZeg9JM21jlyX/YJyGmvYPzGKQpLN/d5Vut6lDwNeobsddaEIkXRDS1sCKi/
Pa2xslp3VNMgiEYgJDXORNvUww6wH3hwHs8GPJZ5vO0Irt64A2XN2rbYneDAZMjkOvBRfiztwucq
A041BkSR5gCo+PHDEdEDwf1iXTBv1bT5oUu8aQbSoW3YoqvrCyzzMwf0duiifT9iMhrva4w7xa3/
SEPI8oY78sZ7I2z2OISU7tG2LuB4EugIecEFlFuQZbkaUCdwNucXVdiHLrqqTyopzu52RxZ5x6XO
bk65+2LP2mD+IhQCCypMjN9VSI2YYrIKulqMuQgJTyTvydmBq6oKEJkU/6Q3zoxek/GocH/CZ1a/
QCdB7pShdK7Buq7MFg+cLz8SNd12vcEAxewl22iwCQoy19ood9Lz9qMFp7LQbzJsGt/LdSQ+jLk7
ENO7sKo/EW2S4nmeygBRoq7pZSgH7L6rzGCiUDJArT4J2exPh0RAOXNr20pb6nb1ZO9LRaH2Fwcf
pLUyecuANoxapHOaK1agT+wLVn0GY0IDi4+7QbbKwhCGd7eu6vm/ep9zjakeMKckmKRT7NykUOKX
JJmHh2kLaUNPRJ5RIVa7pxsDuSjWsvbavH4k9V8ClFtNnag5p2Mtr0ooWT1ARHVfDSj83G8a2ZBL
98TJeBY8zfXmJZHPSWDc4iMyw3dIS523gMCkZsq7AZ2IA2RjXxEGXwDlssvat07NeWgG2v3srIyf
XRDxSSBzdaJdlbrccFXK+jDn/O03Pgcy92InLbSVtdY7C1LpjA+itawoCX38lqMlNqwbarNX7+kq
Au+yBfvigpk8EEPCBeXdlsNYRjMUF5Z19cVGSpU0Uhz3Nay21Qkr98yB6m+DBDoE9wAY04PJBTwR
M/kuZPVH6O+PZsOU2RydqSvq012ul/ykrxDd9S7IAxz+osDB7Qv4BV1ssyPjkPYIvh3F43G5GYfx
uAjqOVHOKVYQJPE1TRvfi4rXfzSvmLx9bdvfNGqVlYpPOohnIf53ZepeCvzOadOVf70A1/2yWlN1
HHLoHbugm7joGbNS+7TBuq30weCdYlEGhnNo8R7g9qxhThjUauU93mRPFkiYZkn25J4Z/hAnzFlU
07L6ZkTR7DkvtwaVZ5C+quDpTIZlyADs0isvvSbrZTPJcUa/CNeTgyeTbQOio1ht6eyC7wjQoPZR
cWYn9Nuid5Smomsda98jCVdEp4mxCSUckw99J7Njl6MdddlbV3KKPHv2knKErgg/RiGVOGyxunUN
vvoqHlHdxfs71EX4xfvJuH1efpOYn2ATKkNpj4RMe87H9hnBvvDx9xy+Dx1MIL6kYbRGQj5lWuLh
mlrXlI8xumIvqIHCE1hUE4pT+KqPnnDKkf817eA51w+PqTe9tKvvo0vba4oWEXaVqydjbCd0SEPX
Mo42kSuJS9JTg/1ck9voI7NflHeBSRBMs85aAa2g7JIs0mt1bqsiqjLn3bmEvTp4nRea4jy0i7uU
jHVlkcCNQBiAHvGj/6//pdZUXhQNF7cyuWHt6AAkBLMRNtQzU/Bt/VfqhJD0dVew2/haru3r9W1C
ngST/s/R9i7v2NX2BXheUwTciodY3QZXNUR/xjapDoUENk4+lU/7x/u/Qbe4W0UcyfrUNutm365L
NTY9Z9xBuEdwEj5HUj+t2ZBwAUS6pkV365cam0mJ7N5nUJzka+cYsRKeT9z0u29/M0oNQIulQFQc
CgPm1jR6dQBVbRKs0d2PY/mg8diAsMCpHDa4aTRZMaGXa8/2LXu95f7aNeVos1z+bFgoVFfruEth
w+4emoqAS+QjcT3RAa4PPdX5RGJYzocFxUzQIkM+nyJLGaaAXnOuxXrnVfjtUYjm6Mn3t86xDqVD
gVt2A5SQbIJbS2VpKwKyPsaO8wFuIHJDw9mQcVTb8zQ5fUhFPYgcbFjaj6jlzlTH9VCH3xvaDdO8
7bsaJYiH9hwMEuRxPtaVXhEeaT3/T8F6Th3L7qOMQBVXOlMb/GrykGWzglRXZpAe/HAADrF+v8uP
0m9DgFijHYk4HhTQy60RMQKS7HE9s/X+B7EdKi0VC7g2g7aWLCNbrP+l25v4lftEhEwHQLPk3ep9
2/cyq7xpoUT3/Avst6PE97EwHKJ6iddxB+492OCNTS9SZb53VCiLFDGGAEQSss5mtaTAiDNJJvRI
A0q3ntV330LLyVbhBs79zjKMaEmfNe3AnoLFCzyTATwY3HuAtZqSNd13qCP1+krsDLwJhe/ojq/a
oCILPNKO++b390wuHOqMph/Vbi0IUcGKA18pj88K+twQ//0hTMD+teilKkm3Jmn4pTIbabJiWC3o
oW5H5eLWxM/l8f3WOcVcR8LlCaZq9GAoIhI9GMgEu45n4pK3JvkrQlBjkvxUWzBb8wV+MJcGr6HO
uOc9V1jULOCK81l3NaIKm6hfkALqxG3eN3fEbr7UMGwsGyR4iuc4/EzkKcPkrAJ5H3qDWZjfkVHE
Om85nVX/fzRa0BYfI5NOf89UhAmgQzPQktEvFlJr/1Pte5TRtrf+7Ps8Ba9/xiM4xdfUwAaqOz0g
xIVJXgIrQD1DeRNpUmNQcyEedXIYC9idhq+ALmXw+cGX3DcFPGCXBKmi+H+qUslRuqQIj2YU6PZ9
W29GoFcjBpeYFXqcBSBPOzXCUC/r+VMwbdfm126ZIjGS5sL7HiNJ/Orj2+mD0ILn5X1awrhJ038C
j14z0+u0Y0Y91W0r8bRVG4ldCIkA5v6QayXq/TjfkmldTA29Jt5kW1Lut7dQP/tyw3uSen6DdeCB
y6GxmyfrZ25kvE/y1R2cWstNl4M40uyO5Vc9VJ7CqXMkNa/osyzAYPKhAVm5nEb4jI2b6cxqE06z
lpbox9T/YDAdY7E21TSlPGcWDKXL9A/O690FPcsdailf9WceBZ8vP3TKLebbWSZwUwDzMiW9AfKx
DvoPIG+7xpEbvBnNxC0JEd+vvY+cFKCtfd/6fLEuIBD9Yvcyuugd3WVUr7YUz2QB+M+EoQrVRf+p
mbbzqq3b+Y7wZciUbhYk0ugQWSdWlPdoJc4MI1YWL6NXhAVDMouBK4dOkIZPjQU7UPPpE62gMwKn
ic4KbsLD0aREr9ldP54JhwbMv5jgXDqZLEk7k6FZm7yhCGPsXdIhy1Vi+NI+RMDC/6rdCVC6Yxi4
V/DQf1a1A5oajsf6HaahPMbX8K96T+vnc9tHiyMAqzVfTsHnBUy7QwFb+CWxGBqSH3jiqu+jMBem
Km+e/5ZcPzMQlkwsQ1iLPEGXezT/DgvFTDGmg3V1yUghOmR1KYOblevS0NqBwjKz1l0ttzvqX9TF
CyhJJ+VhEGTvift4JjRJcpLYnZSMJMS4cC2CeG4ucuQre7FWdkKYwk3KMTm8LW62rcB7+UrADSrd
eRbFkYGcFthFYmzR0ki8ISRGjFUlgmJYjAJHI5VZ3Z39BJuiH3SDi6iC94a7SNu8rCJCB0yQ30Uv
zUQHCxjPwKUOnjWDDB2Yyohs8n+QOnOuaGmQo3HqcasMu2edTHI68GXfAJWOHtYlgrVXkdtIVMKV
13MlbH6/4PBJODsHxD58OmSv78Uw53YIt/TJfAoh++pI2H0iRp+pjEVgGNeRt8rbTmgy8zYrvRCp
pn/vPtCrMnx/U5sNvfMZzKiX6bEj1R3BWP0jiVkBzM55ZRetHfFDl1Q73i9DHXL6U4vWJMpWX2b/
khBz7LTROXFeFLyu8mlMvkSxQopO5niC1rMaXkyovwxI21bH2cuUI8A+M6+ysgBXHFg7obi3e4R7
KogQSwC1H+W94BJFyMNn34zsKNc/k5sN/8d1dSsI40yJD9GegqIsPR2WPJy27vj2ILc4GG0+6hVj
fSy9k5O78Qdi3utYRzdS8HqZ6v17M/k4jYY1DHR+wAsJP3oJxlz5FpizqqmZ7ROWnNAYN+e/L8iG
ez3pZ5BGhq1PfePCjzT/kz4X85q37iaDcUtoFp/fg7r0mPUgVHfABLl/zDV2IamTyMz0absaF8Ya
n+lQr+oR0iSoHPWUeDhgjQwYjxu7iYNzqSq6FJLx6ehgD/3dP+yoI/kzSHYUizSJIp/SIK95SuxW
r+xhwvwI+kkUMe75MAx4oyskV79+yRjNn7Z/pGsnC0u+h+pBwDocjd8IjqV5VL4wcT2LeM8G/L+N
DRCdS+yvPf9KNxAdBCco6MDCUKc4+GLuN+UXt77ab69J0ioLbiYrQPcqK4hmtA57EsPG0bfGSpfL
RPWDNDq5nscAw1ThQjGWLng12pjygTzEAAZq4QPj7z5brYVBkbP/c4iYeT3h8ju9i8C18i2cvNF2
XR0iHjAezCeWM+tJ6L6QJ7PUzaGCVrJV6Uo/yORcfXxGBapn0N3+cNqL/3oNMjjXNvC9250a4hUq
GRKvjEq7tZSQqVxUVfaKmt1TSf2KEyH8vpDxfhm6cR6f5UIcDBATKvcE5Gqoy8YtpZrTPjwwGeGZ
Ua5bSn2bfQtOeLDw5Jw7k20zHsXaYIZRtLDQfdn/t6OuL16EithCXtY8UodjnE+ShdvRzArBCAtY
nNtBv0G1lqcwHS/eFP08hHf4Ov3sRHGqKbGhM88czPSB7HYQONJKIBZmBaWDDY9Uqbv00k3ocxTh
sr8rI6Bm77qIpyUdTJ1IhWB4R5oaZPQpMsxwdiUBA1W5Tmkxxi8o36oGEvQmcmmMpo33GDJvdD6X
sDa2FtfyOcVsBsz5u+AniOoWX3JIdPvE5lm0EqEgG4Rn5leQ0AoVGjip5mduVbEHwzPnt/NIUSZz
89AEWSgah3mIUle0azMNfBDIBb+D1mtaKrn7damHchbViSpilkpIYkKjgLgK7kQbnfrQQKH8WsPc
+HYtB2FvUYRDjGlJZaGI7QCU0ldFQ0zs4vj8x7Yo0atYxekyPYzl/3ZFB0x3ORFxs3e0TGq0UTsy
ZG7gmTcjLanvAWgHtp9kK/1HSed2uXs9SClo5FoL6sr5N9AXJyVJhCh6ZKuqNECBDEl3Eg2WcWkj
iXo8sOKevT8Kz7Q4KwBj9hFbwJNgH+YWOkjrnBXYnM/2y4hTu1nS2zdzz6kyNk1oock7hb4qd12m
8U3Ljl+DwEbYBRKIRRwkoiFjWITtzlqvAa27IWEXkjKStxzyuNf/Vf4UQy8n6suIga2I+bOyq9hn
OmYozE1Od4lg8FLSY10gz3dEUjKeuTMhVTl5/7V1ivnZHg/Q9BFNf8kxeYmhmpfSykf6tc//+qXQ
G/83Xx44p67mu+Q+ZyvntBr7cTjtG4l5086vReNycrW+DoruLfsoCovEeOmvEg8fXWeUUX6jdQHE
osj/hO6FedRX4plEyA4vPRdnu7eZeghJs7Illv6TLacg0YcqZhfcFM62Asskz93Dm0+ednct9UHH
NEKqwVxXXQMGZy5V6YC/3QfFyWc4yBIW53KQw9e0v6sDvadJZ/q7FBmLs1O46aZPljoC+hETPmUl
NJtD/oNHSP6OMuLCXXwyfd+nK9E7BLY31G8rUUGVnIQBznk0meWzMWrtp7xNPbbShJgoj7MbLYjC
nHVr6gUtXCSFud8+HH34i8WeNSYEDd7AT5V17em01PkuR07zCL+/BXxUkpPv5NCZjflwvy0MzN+J
erxLGyNLvmkhDoZhwIiJOKmj4hlCIvzB0eKAGcFiWdRcscJGnfeB7KD4r7NC5jKD++VWYc52IJ3H
ldSf4qKCB/GyIxg0YF2TlDBkLQhHPUQJG98r1K++M2x+IuHnbRcK4kZttiJLe6+xV7qno0qPmLhV
GvmfXFP0yAqL3s6bUBXNdT1wKUpI6v4h1ij84xEDbZqJyqeYou9s5NNgu53kLzLbPCZ+W9YkX0nc
PtDY4TiKXx2jckYmNd3ze8/x5/n6YI0EAJPaouL3XO3cgYeSQ++kktgLg75trIXMdrx278MfF5iK
ZACjBPe65agy1872pvyGfmcF52RxJy5VvyVSsjGFaFBWsNrAicBd+0mvDnQq1SdVoTlJ9zg6e3z6
IqM1jB4qX9ddAivHRYo4El4IzIe514+Uqi65aeS2o+Ej8GqBbuw0R1IbjSQZvvS2KW/rDWiwBKKy
UF8Zp50R+91JSW4OdATikLdFBTVjXtBuFHOkrBMmxp1Zg+J5lOuWOX1SD0tz2uvqFsEYgtEf8Hz6
l+2w0J4SNhM/uQI3iH/tuv8yiGcxkalb0wyyc+P4Iahp21eOA5Ki6KM4WLVuu11XQ05KGZmnMXcE
umZAR+JrkxUVrbkdyXTUA6mfJZOrhS1baN0Xs1ySYsESve5TAHiCIuNhtz69dNEO5qyNN8r453rH
RG8j3AspVx2T0iFxMGr1h1+JL9S7oiQQ13TFa/AeIBwH7eS7tfRs0vDAyqRLLWu5uskkCjxbt3fJ
OS+NC565HR3mqpdIUZnPp2Uer3g7YzbMLT2KJUSnBciZKfLKQEeEJIj1KJmCzQtmLLiT6FAhyrPd
g/DWMYzPGlW3CWcRCFiiymyz0nQlnCAw8dOHnviRb/6zgFeze6szeEUVIV9kJs9zv9PFKANAtLon
tkkEgi4P7tzV9LHJ7bw/WHUfrACJGaQy2lI6uGETS+Twf3CMkoCzK7PMRn38zmoCfs1h0xTd04ha
4WMdw6yJ1c/2ZbpA9MpTnAe35uoO27MnBRlQB+V50ySCwS+X73tlpzJBoLNUO7ufOY/LR9KZOqOG
/2BujvYtvxK+16xEZpa4yzj3IdCt1wMZIv4ooCxBD8Vximdkb2FUr/lKd44V9gIpBKbM/UETTGEW
qt9qihN1kzFk83PHQjUbm7D4QMjUFUg2/+Y9afb394I+X99zdKPlgdVGw/aVeK5IIRQmGDWiH4Gb
UwRmtIfObdet0lSHNacArS3ckkcJGtvlNBlZE95LsnbcPBGnyD1Pa86JdkeJ2qSplE30xAc50Okw
FosYxHV2WB4lxTRa/0LzKS/wcoGmf/X8zSd0s3m0L8lDzeU+KJI6ItNZ4ReW9kZPAj6Qqd/0OfbL
74ZaozPzqI41oKlSjH1jaUnkHZ2VoiPVvrvGUbc7NdoNf8FquDINXiX4cumF2ky0w7YvThaGLExN
yUoScZDPZwJTBGUkyG9vWqQ4/q2FayDpZ/XInysYo4d5uCMH8Sef5UMoCQuVMBINaqCrsIb8Ep6p
iVngDsfzXQzHre+mm+KHZkc1B3c0WkX8sgD9i6UJ9j23scmT45YIQGT4Pchr1x3ZRoRT+yFUVveU
vWEuctdASk3VJZAbQEnvDyKkB4nLDG7HcH2JHyuKwCsvUiezUaIVIZOPFxV02PInQcWCOkFaU3/e
oBhUsFgC3l51erD9t5rafcUj1NEM9Hb4kvpISoookrnjrJP3UfZI+q19FKUbuUMWTBEx+SCq/n+a
Bc1/X0bpQySu6KOn1rgLOejii1vUPYWR8JVZnjZ+TySE5FecFOgQNEFRilltt737imN8MOZjYOgk
LsSS72/YvRA2v8FbOSFb1/oH06YnX4nD5wVi3YhfJmDK1SWkoBF+9vLvzH6XalSQ7VjV+ENzBHqO
NaAATglFWAWdCz/TMsvDsSTSS6zCeSuy8MF97owoiVF4XREw67EbdvpGhevKqUTzLRpZTnSe3HOI
4Y9XuA6tcXYIJJzAxAlf4MBatUdM+GnlnVkIekBJ42KQ4L6B2Ye01u90IVeaKg9iUA0ch3H+Yx0b
kghjrVa9gqzN9lhuzhv7qhv8g2C9IEoBsd4i5TU5M3siD0KehqNfjBqrFc7N+97DrkMZXMsXOBiY
IXbcNtVKbF6nYDWBXu3jBTw4S2lx5Qt07cd4kf3AVy0dPf8v66C56uMGbQbEoUmMaS9zhHIpzob2
Q5vbf473eA6Oa95PGgclQNXNRyKgX/XltAy/UKDkEQpSrXRqSkDl8zpkTRlLJHP9ySBNnaGGXNiB
6jXnTIw0s+/WACeSh0NyAziFBVCeoivTblyWse1/Uaov31g1q7NY3DG9SecItwpZQ1DV9FPpS6J3
pQms2t79QEEqogNuA9Udcs3Vem9eQEJTaKRhQizJV6bO2H4cCV+1CyMw4dpeYOfNcfQ1QftS6n4d
zavCQET+71gVQeUAljU9EhMIlyyOoV28kzAxNM154e7vCeEn37qyIKf/5nnGfwYgp74fH5Nxdwja
Ge4FrxcoAMczPDPs4Qhdx8Clulo+14Sla1Oo9VQj7nxSaYYfSCdfJhbTx3iItNg6Z+Jy4Uaf9jTh
JLKagm/MlbcTUjw2zGw8WrppsPmTXpbH9Kr0HVA9wrDwiXTnM8BkxeRSekH2V+r7iSVneBHpj8KN
IVNA8C9vJ1WjfWW3QLHtdLRx7ck+kbn2KA+417uBlVTsvV0pVVoJmg8b3E7A4yphzbK3wOWFYvK/
tkEGRFQb09au+hH/9SwFUI/s6zRYgrnVq0GJEqTBK3q7ubj24mJys3PMwzMi6hchKBwZU5vZnxOh
KlKEV9ufFMZw0CMiw3+8Jze+sWyJTd6mo1HVZJ0REbs5Ah4nfIDDOmMPzgz2fcVZrjv1FZJ25BiM
LUH2fCDOyYfUEFmD3uwP4t/Q5vmBVRmO8rHIaaxd8ifUoAamB6RcKcsKtIGje3iPSiKkurTqDkU8
Y4FgJwypj7kNuTs0L9GrGeznIn5rXibkfRKAPybTt0ii0sqWohyJbyW5QCtaSD2P9jDzGUNpr5Je
K6Cnt+Ajnmu4FP7T862SE9U5+TROTU3CBgcibBtoYJOOfrc7UmLRr0tA0R00UQXF4zC4ygDnPtIu
ljsKUoctpQ+7Idp9K3s5Uh1VX3ECIP4UT/dHbPymxKtUP9NaWoUlFT5R4TdDgyy9Zf7fxr9y8Yb9
pZ17iVJOrUnE7rlFFCPKYCA24h8TlENRWu4V4o6tU3S7VOBXs62t0NHWZNj4TVSCrxLpQ+ZYNbox
abULZneFBZBsWXCz6RIS2advZzO38ifPXnmc6up6i8HRf3PR8+1O5bWn22AcLzTmCExUlNW5/l1x
GQGk9HKdI7UaVIyP/+lYYKCL2H8hNMg58fzuJuz6KqGP9ISvRl1Tx3fqDA0j0sEEXpDf2IbMvtnA
5P6sAZgYiZ2icW66nw79YRPEFrSM6uwv1duhiEh1+vIFfbgiakhXxB1FCzdSMfre0S3RhESzbN39
/yzMsgv5mlrX2gMI3Dc4GnEFW+K335JDEf2al5tuLpBKdvDWIZgeXyTC2F+Lklqfy9ARCDhY8Rn0
xEkZq7FpSpIH9BlbmM0YFe//G/aeBHXVasQN1bItA30SbtMpWEidszt6wvTvcfovhH6NHy8ePMqJ
QMLHJqS7hwI3O1c3yQbERT6mUVLRZErPxy68hhorrcYb5cxi8PjH4QJx+o10VegvjbqA4nV3mCOF
aBnAievKzM/gQ83oHYIizmeN1BsIo5xscBkHANRJ9OmopmtBd3tRO2AifIaunOeP60YVN44AJHrY
3Wwfm0K6jAN9Arsnjviwif0uGSbHLvKZmuzlqXVx7oO21ZQiPiXX8P3Vkl8Y52xOQjB9ZJhlCptJ
YWL6/g7WuJi6fE8bwOho0UvzbXLXYHJB4wtVjw8mQ4mGAI9tYRJZs3BZCHprLI3u95i3a2xecxdr
pQY+tskfCJINVF9gjmDuCelOxBaMFQFbprDhjUiurqNUxqgiQLsAsqEsSAKJ7jxrmyGrbVZNFvxb
DA7vA7XaUetbr9FnNeGdMvQIJFJBET6QqC8IwXRRdJcyD/1nCOJdLAHUSAoS/ACxpbWUWU2qPhig
fbB0mYZDL+a8Xjkc+9SnYgdNmdL34D0OzNUXrAZNLMKw8QR1YJOZCesh6UbW+QHxdz8vEZkSefSA
rp9z6QM7eedyTfyGVe0Ndc54tifU+DFJXYusHKfwZM1Fa/s5uEScQH6F+9SE9tLswKvaqr8pFyTm
wJ3rFgK3ko+pAC5Ens+BkHVBDLskLCEgc4+KiBcbspYk7oipNThuyebGHPGZcMUJyj1oCX/keMox
vfb9BWIvwUeykrRSMvs7jH+uaXOFr0LQJ6ERTVmmLb6DvAvWNeHQfyZtRMWOzeZv+zjPq+QsKV2v
SimR2labCMlJ0AV9DlexTSLtc+QLUOuajpZ8XNltFooWUyyfMXZG6e4Czj+jd6phaTyfFVh6nnKe
gM3wtDKv42KQg9acq8CYROsJKamYKWbOwKg90YNz7/rIQJnLibniakJaw2q6oeGHztPPXZse00Bd
zSZ/yqXRFwmk8Lj+DlHtoQ0plZHCB6ZHq9xq04AF1tyqQ9+lz+jcm27f9wmGVdyYqFPp+YXlhwIa
G2gUxzJvU5C6Vo03HWM8KivfVrVb6qFBCICP4gkdeXCQXVD1dVrzHYnUpxIj0pDDFNSUbos92Yj/
lre0OKOG/XqZfdWuIDrHOHVMW67zme0yhiKrU7x1erxjJzCRiYKz6GFs11cUZx3r2tFyf23TQRxo
x5J5p37f7sh5GrqHkgc4Zy50McbAAKo5OYBtb0vlJk8Wfa/Z1OLDxFSuUed4IE5KWcK5ZfXvddwk
q2VCweTnnvCqtLcQ8X9ETJhrXOMnU+br+xXjz4GJTu+albcJ2lnM7Uz7ee8VuVlc61Cr0LrqP2/8
OWmsyFw746j9eq2uuS9Eq4p4/R7nZNtcCFntPmJX4wMokHA0ne7jaa5XtXAY95XQbVjH5VB1QgKR
urKZHM7P1CpNEzKJhLIxBiaDE7AD2SU2TV39J6nJuZjv6CG0JOrhAwja+ev2TWBu3zc9+eQKOib6
rr/w5cGBIN0SiUYZle27AswEAxKqBTSB6eaf7RgPftt87TbJBRo5oJlxw3DJmEtEggQXLiBeUDbz
3J6BHWjwJi4xe7XZjqOWb42vUx6+2sQBqWpMNVASC1a5MIiIJ5ik0XW+ZLJtvsWKEllGfZxpDhCY
ErR/rWf+O4zHQ+AqAp9vABsx+35gaHYAO4KmmSDzCXT+q/uKDExli+zySqZ9tYbpOLreBzSpf8IT
M+TCCW79Z3+3ulElz0UBgC/4qtbGrUbv7vAANzRUopaZE02vlAOKsnQqvDJk5Xcbs6HaDktywhCb
+5nYDw6yxafNnQDAm3s78weQF6YPz5YrZYUXS2Mrzh/0lUlz7Har10bTRI3hqrrRcUsnpQxpnhGB
T+kKe3spAXauLWZgH4cEhwpKt2VzJB1dP8GYU15Wr3zfmbEPDq+ZURT0GMwoUPbs88HJGcsUfAOW
cnwudJLcvZH+3dGxeUVX2AnOq08+qu9YqBTbiqa6wgqjS7gF5R7qvQHYrzcF1U7dixcOLfRX8deI
3z2tbyBdf4jg/Q3ImsG3GyPqeudElZfSomEavTw+uYWvVtzf4VabEczafjgrvvCorJngEmbBQ7YC
A7OhmHWSTJpuWPLpZDSaNyTCAWUzKkEa0J5T+HL2B0vwi/5/34v7USQEbiZ3ulsyg77UoYlYiMjM
mXVD0vVRJv26CbFZdPPbBlsuBqyX0nevSYmRtirEOFCvMHWBmm2nTshBbC/4AdiulZe6RG4jd2Gs
cuJz12bfavEJRff4NZnd0WmshKIrYhVCvC+jk4LHHt5zU9vD5Yom13soPutq5EK/Dxh8TQhk/oTU
kdR6GBFXHdIQMDuag8SK+Poy+AMYfus/syrdP4DMdKRBs+2kuiBCTWnZXoUq+BlPmuRJYUxDczjq
ktph+f1DdZVrRGT2P84poI8T7SlN0Scgb1v8li8cZvCkdl37wx4VtFNeLyqLvINuuT8lJWTJJUJv
fqk/V0q+NJEg7qnrLUZQ1L/zcnWM+9OqNfBekDtcyyikt8CChSPg8d6voMRfOPOlc2XBTw9nN5/C
Cb26JFL70+JS6npSPd+PNdSHMeF4EuxaSP8oBN2ESu9oz32ubV8VvZEeuttxkhNJR6lqa8FginM/
msxKNiUJCWCM5gwpGXp1rVmIo/9WVaBi2t/+yyMjYSr0B0ZSfmTZFHF7/SNZhns6V3ZpEqeS0Eqd
OjRvhufRMB80NcNHbCqyFE5bWbzA3lWjlDDLhMaFBDRvUtXbdYv249mqJLLrjA5nYgBHmtsjf4n9
209p9g6DDbdrp9DQp5w8IOrPK7TcPOpiSk2HZyDS0smP1IKiL/FFCzT8S0Aed436QA17h1sRHAcU
+agIvyjDTq4oVaYTJSnMFB7FPLBqEiwpCG4Oku2d+IqFmRSdjoJnv40XugP9Fqlef9422gL2Wuo5
Byxz6CkZHZa4Nqg3Iuj5geJVdg7EAAO5xjxELa9zQ4pz+9dBa+dmEQP9GJxcVqSmWvsX0Z5ykOH5
1U0blxSIRXvCtKxkw9sc0168+wTtewCF5cMFopx9r3+ZxFMIsHpJ15FglFhIZUy1brnKHlIZP05H
LY0yXiXqn2xzLFoC1LoKAvlDcuG9sGM465z377JiupnOxEJ+WIEM9cQKEAYOtm5HKfCg2M0vsymy
iM2bbHLXgKyIni9sPf9gWdUI8uT8FzE9sS8LtIr5Xh/PmyVACN8waBk70JXrM2D8PKfgiqtmsMBQ
vGjplJr0m00BAM7RFHB9tEDKLOpjtvDonjPoz8xrOIZuRaS77kspc5BbVvTENHlYX4/dBFoeSo6G
3eiJCXHOp/pqvrDDLBz7O+li4y0jqZGf/lJb7I3anvD5103FKEVMrEyR3uU4Y2PisdSZRI3357LY
pGEe5WewJMbiKNfZdkN95yhzPFsv66doVwZtP4/zPJvrUH3rRHmCevKZMHOSPaT4Hyy9MIozdtAX
/sNba7NV0k8Qfi3ruZ/ZIbbJFvo/DEH0Kkgl+xYPWJt/xDexbjGBJ8o5sfANo2OB/NzunImLmu7b
dAS3x2th6ix+dNp/tkA5Pnvnwi7xAb/Q+WNXYbmsvYXkG1MK/iK464abO90rDMqzJbZjHsT5gWn1
bIZ27geORl9kvZVbCB4r6MMBVn8j82d1crEdNTQPSbn76ozlXSwJ+Rc2aIrsonbShtrFayOht9Ho
95oN82QMY7HsW/bGxHG4LzSijbE+ka8GGAjuhHvMkjrVrSrD9s5FLHfxdhNT3Lr4j9PZLE1uS+By
CIdgRSaV4egQ8txZ0sLMBQIg/Wqqb6Kd41l03d4VRc+aFb3ioqXgeS9eGhGbRZ1tRdXRRBO4ZUGc
E/Vg/KxFypxl2zS5BYjSDlPBBu+/Tm+qKh78SYfbqy7gpNMdM/StOmv/nSAM2M83jN4qX46CYJq7
bcyM3r0NE+877gOvm9MRrK5tzRUWF1bY+4BgwWeCC3c5eB2bx3ynf5AiLUdnH3ILfnn86u8lQ/a5
hb3RudhV07tvd/pa81UVhA69AdimDmjxP0bw600iM3Qp/yg1paahWjwxfWGJAYsilclxfjmNKw8u
6PonGHG88skW7i2cKmMYkPq6q3drrXUom91RI8GtPlJ6ISZavkjn+c6SszsW+gUXcudUz7naKwJY
c6YI2VdPudW36PPMTpdthEZj+bPMaKf//uwS4o0W2b+tfaODx2bG3boGG7YU9hiK8v91Q+OmlVK/
O9Ky7pgz8UzaD8ZUg1ixbV12kDLldWPF4VCpGJD6UeJMebQgUu+psHLFXf8WI9nKlQeY2s0GFCxE
r4NyErWUzMmQ3XooULiHVIWq668Rcni5wqpEQvBM6H60d+f4lJuTxFV5ncTlwgTG9KMIan+o6ZCk
N6hnUZNpKJFUnvviscU76m70x0XNm42dPestM6Gcj4KM0I1Yu5DrfF+wnOTWhIXKZbNimHuk3PSZ
xjb9GDKdN+WOmtJhQgYDJboMmobv5SrL3uFeXnmgl4eeFPwc/1H1FTWsrDMOQN+FydL0SrhCUjtp
z4MoCWrvpi02ai1Qroauq9XHhRLYVJQ25bzPdvz35nSUVkoFIts9lG7iDr8w6a9VRVdX4ZVmu/PQ
MzettXU0TkNQb56/z4QkyrDD7DvHBGKXcOMdYZDefCDy3pw1JtzFVmf46PstI74T3k8kRn+6ZBd8
R/CNH82V2Ex5yojD+MGSQS3FM4zgBhdYnUOMdu3rzbcLJU1Rs5E58eVCJL5OAOUck6YBxzeZtdZM
dZ6wxpozbd3zAw4JxVgoEcpiMEdHI25FuSVrQ1szmNZkaltG39seWJMrVdxjqehI3z8g6y/D1leY
NWBZQkLUOhM9Qmc8zte7PpTUBrEU3h1sI1oRefor9pa+kG6LtDucFC0R72tbTxC6GxkCD+AhMx1Q
xfZoL2F9WVYdU4ouTdxdsCAn3ijc1JOKIez7ify0wo0y2eQOBGlhbjsUNrW3SoG+4DsFDOqU+5me
Qm26XQKfxbcvduSMUgJVDGhvVkM0fI9l7V/3Dn61Hzc3HhDzlo+o1SNW/0d1cu5TKbRTy2z8ax+5
r+gDzNcNrSLGQDbvLlIl4fUUJSApn6iDOVW50Nz7rKDySJPYMGcMawv80iLn690o0eN8Qz9fnKAR
2z1Q6tnI5pJuQrwwJTACLwp49nYrGu+ANCsLhSvtrRCNvdbW3pO6C6CdK+5GcAy2Oaz3qPbvw17O
F4SEoRJozw6IOfa3Gu+UWUwsDlunNUYCertdxkatX86xIx4g9H5We80wPgd183DuhjXowcCBrMVs
S0VGl3bopXbDbdlsW9Rnu4hKzeZTmF6Y9TfmV2ui2eKX4aK8389ziq7IWzmoOSq9fb/vbSD1QKN7
XdeUqBcP/yaUrCopfrBJ/E2BaMI8rbpRGkAXhcvQcX0REqTOh7YbW7DU9qjW70XGnV/9DFrOAuZq
QYmBkPvP1YI87dfy9UI9lDh5LwF4u1AEtYrpp95wRCDizzzDwiIGgZk1qn1OuKu++Ab+OKtZRULm
DUP3XGSz3IzPdWNwqoxz13Kph4SS75Ec6WgLfHgpmZCPg1qtOO/JStzzLqJV5ndRYot5pAbgkbAL
w6HEpA8RpU3BDzcKZFHUVcjOh4fwrVqnGDruIDjcQXHfLizDreQDHJ3fy6jtUAHW+FaYH5D9Td+m
4GnhZSGlKUswE5Y0kO33alQrfgvf5t4uuohvoAw3oPYFrNN0F27dFO40elQ13gPQtN6ho3rmLHA1
m/dNASIX6Jrh08baGuUlTHfj3jaC6sJYzf8h63cdAxq2jTfDNWwLehFx6j7e68ccfuIKBLxo1R1/
rHgW7X755tmTsLgdymbRQ48eT7pbcKzn8Soh56s9eHGZfZv7jsJoKgsMjDaYKw/kKDVPaAfJee6F
IHZvvK1KDuOcwkqknFXvfGo5d/DQY1qXDKwDapxBr4yqTtFQYKH/OC4mj1AT2KyDkP3fDrpl8VIA
Hnq0XBMdYP/rnqZXJzR6G7PLgmEoFCMYb1FnC0ayVrTd5icD6+wGlOQnRmhaskKAKjJh+lqWz1eF
LowFaep/eSdLd1accDNDNw5fQ6XMEgss7yR1RGtipKn+WT9F00lguRnDSmsmXsGyIaojvOIhkacW
fntxi0TVI7kpQc4Ljp9U2arF/cs1vBvKmO1XJWUGq3avDX1H+II+35eYSkq7saA9WEJbNRPSxYva
fbpBejzk6HvP1Zvs3DVr6ExVg+3tDbLQxbWs9+OLCzko7a56ygVjVrrRjkie3vCTQnGEeZTHLpw/
L87CLgHR5sqY0K9am/3gZLCwAwsm8FfdhGVXcxhwkYgAJr2aIZtToNqreLDBYwpUsb8yXEhz6/hE
6ItZN5y/tHt/63622n/aqEeFPIXQgfv5gZVsvLzKpDdX2W+PkUURyM1DT8BbwXqp0ixdzsLMQAzD
scd+tVVLNUe5Q8V9WFhR2MY+8C1NS0JPy7aOVW8OGCAEDraUvKin28oO5eQMNwNwjUDPnU1uNfP6
yVzZqV+K4lhMG/rv8jVUCly4iX5UaehyvYQs47E6iKn4lih+zkkFLTkP49WL66wQ2Dj4dfsJXS32
dKI+qFXXeqfHLizrEXlnZXqTJQinCwRCqy10OqnJNNLVE788MmD4tJbhM3Oi84x49a4pCBkSXc+A
ucEMqsBhAEAOZ/xpy2LKkIJguhHW4mDcjgXFSPFLW80s8iK5zBbnamiiN1ulzROjFRtSHZnfzGyc
jBHuqdfyil+PH5BiXMDMzJCTIVe/dDAHoJjpah7R2CiaVHirWu9nYimYyXlVF8f7WKzxUrSAJoFS
M2XbL88ceqW6hqNrjdLNLNsHSzLVf+q9jbAGkwLbhlCpMEu7o4Et6by7VfeCYJOmJpfZtCk3Kl7x
hPfZkupzn09/iTj7RNheBqdKj8Usj8fbnLbEldkg/2bDDSOlIUsw9ER4XhguQyITgSh7SsJxPKOv
p9aGo5oXlmnA/j3d4wkbFuuhtSGSBijiDswlMmBGWR+YRDRVJNu2Z6PAISSMAquO3wMCTYhG3IZS
u4Uf9CQPcHD/A8/RZa3qGf3KIEMRWAfrIT1ec5NWd8xDRGQmHFUf3sM6jZpVcn4StR+0Ks6hD8E3
GZyBtPln89Qphp8BhIXzZpNYHNc7nStZCHcpajgR+nzh09gDp/rz+DtU/jIH8khlDpXF68mkppLv
hxMCLgY90YJJCnXa5Dg69A2DEfbqyKzuT9H8zsoq51opm4oDYfBvC1zEvoyDQYnEXOoOjHcyoEST
1W+g3kSNWSaNs/z7drYlCbu4Wxy9kLO68nco3Fic15Ub3ASYEnGVLuSY/OySJLdIma7GDFkGlok+
zqsEYo9yhgW6KfcArK0FFLLcZGyB+JcvgFMPxD7j8HKvCKH70ibOWRrpPQhs6q5rt/rkc8uKULjf
u4LkOufT7mkQ/B9gh2Q0CPhmjUnjtKzoZRX7PdjEVxMxC07uM93n4XvCWCmiyUbrbwmkpAMxvLeB
PxzdSFtP8l/HJmqz9ibm3kL0WFzRST1P/QWe+j/qIESxvbsajVT70rAVFWqynbOBJNZ+9xKwimEW
HcyhUhimOv1+w+Bq0Cj+6Ign/pSc0IY+1VIfHmGdVgE/FT3U9Jd10IaqW8fCkR3vQAbeE7Oya7Kh
55Din99a0RQ/5f3yKAMFIy3MhSyAiMYY9aFM2W2OfmfTlpWQWiB4rt6u18j/XcEw/Zc1+u7GUktX
lQ4lggtrkn5216nin3zKspsZokxmdGtUVjvI5K18ZAfkKRZFhkhHJ2V+OAeKznsIsd05pCmt8i9J
brFM5vDi2X0ccb2nEl5xQzSj6eVe4BgVdPA5wFhYMN/9+x7PUj2Tm7rCeQT4UwhagSqLAKexIhbI
nbEz/2BeunkaK4puclQAUZJxpA+NJveqcedHbQJtuN1WRpl79QFjrd/nFIpNBuZhJe//G2w5UEhc
hNKfJDz0LC+nbCetlCU/BaYBcVQv1XZ4B26gDCb89tsiLy7KzpD0jrZ0FzAdcbq22pMyos56BBuy
y4qDddeD5a+RFgGcFmufvht/Q+XPKfcjTjZjfrFcNW8UThlrKqDQ0SoihOm0lt8MNMdeS/cFPgO6
YujsFWQCQArI7xsN6mIhLcs5LRusaSlQHD+DuiI3HAeZ3Vo+IOA6rOE0c2RnTFDCOXhjHWc50ECX
v7+Z3YS97cNlwRwBcySFI7Y2qvGnBjL/oWqIKLRUEtLDO0LJgR9Bhobu+NHTjR9kAJGHo9kqOoD+
92L7//EoJbPP/m9P43RtgVR8rWmyQVAyITd+VuFs3ny9T5NP7ItwNV8LFARZrw8CgxX9Tc5gc70I
aFEoWO5qiNWzyK9/DC0E10j9mUtW6qJ6HImmfSUMpMStKTxMxjXROTTc+IO8FbfmWnmIyLGxxGSG
OO3NVwGCVSD4lfyqGPyk1CPQIR+fUQtZFqYuT2Dc+BfgSomvpw8uEERW4KKhREKyk9OzbkWcz2kE
4iWvCVhHygb1TcSsV0SNARc1BvxXgJveGbDXL7jNKu5pfISLYsvEH9geWpF/EVg1Astqy3u9kqq8
UIOygyCHWPHw/yV0n/DSO8/QJLT34qlQdMHY+RuyVWSlC6JqAHv8KSGYeF923Um/n1WTDJ0uMbzB
/UEGVA3gzjIj0LFVyAP6Vkk2ndpeNheMaorAPfEIxrRVeK5Jx+EiH2sOkgAxcOb+gEJ2Agk+NCub
wHJebeOGg3erIEEQeDKDCTxamUiYaZHCeq27+tTGuC8QV5uImMAhjeO5Ioubama8Jchd7Ec/xuoH
6zlzTGPsgorZz4KCV6Q8oOtIFSWLjyCQMFWyzUIOie29EOYESqBRLMPqDX2MKNRbwslMVngZ5XdM
Y4hq4ByQgsUNWIM0dviBzIO0jRHqvT4yzZyyouiXg5O+cqnc3M5DiJ/53HuLGEFXn7210RTf52Rp
+WCUWgn1EA/ewm2L+/rjLgD+oTH2xbuqZVnreIFVPQbV5EF4FV6cPSuXoDbF4a20acs2NFRaDXuj
3hcchALPz4EXyqCXZIg//eqOeqTgjM5emRew68mbxeN+3b7ZZbBJJ7ovXwbQCtWRZMHjnIs0N5sG
tv7eCnCcYYqOFI8llTe6MJJX/93vpDRcylNI6u4mDYWPRClSyUY7/lH4phKh9gov0wtKnuxqOsmH
f0EkiGQfRMuta0RJ5NmX991WDf2mbjwzF1GqQ1U7wXhKkNuGPsA3sqWV+xWfj4r9LKhUBtOchwPJ
SahVSwE4g7Ru3uqvMA9bi2eo2ychBFmui1TrHijPbCe+aivx0XIw3RfId+2kA6IxWBq5qS371y10
4EI6Ye5LqLE3u7UBCRI3RtKcZygwG52e/kdEjFDHQNIHBwViT/ko3yuSdWTdSBgfOmNGXrXDzJkc
HW6wLsMRY6yApiAloiup5I9T/cTNxvm30gbV2mHVWtfnblXfrlvYqdHC5CJYpMpBnjRDXqZXwZab
InqIGNWnVa/j5cOs7l2vlpKJpSsnHsJz05bgnOljqKdEHjG5egBVLZPbAtlYM4JoNZQX3dNfFOz/
9+4L03fbagOJqc0T7lhGApSE3lmYDEnJnPEjVvvx7SJKkEHfKGsDZB5VdfpmkPuyIyIEkgDo+IuZ
/kTReKqcb4sND/9OyBZdBFXKpuIS45zanuruqy8rkHfyBD8XLv7Z6ZVawsJBnv/23IHHrZriu9Ot
2Bbam89jgzJYwFX8iRj7QJzBt5kKFzpuq7/TyJNfmuKuOZFxEK0wOltL7O9Rp/xGbbVUgFLiZEY5
TXgGIrxHNJQXPfQ/iskZB+rsqxLAeblcLHiWvPg+fgHu/80YE4b444c50UhtPe5t0udx+CBBRzhw
NgglNnAb0/zafPav9qhllVUL0sqqlY5G4f2R5u6auLWO0qMEk/uYj25v3rXxcY8mb1tjY1HR1POD
OQMm4erNJDOx6w66zVByiXk7gvBzcpyohrnj/UGx97jvo5NMay9I+jM/Wwb9P0lvDT1Sxu3Feuls
ti9BXajmp6H8BMeCnd4YtLr7nxay1KrP6mj068/41jKyBfm7TbRH9NuTzVj5cGR8UI5LenSk/sOm
dLc9JmGZ2zHZqjgrovhWCsj0QIHvVZTyripuBaUBSS0gyNYssrjgb4eG3aLlAnB0OxVKcr8kiaA2
h8X9DfdFPOCUZXbnnhPzBAshwomWLKO95bm/+Tn0BFKU7bNl6OtVRh0TqIQDqeI5VoBwMF+x4rq3
F+LvNbvHyvHTOvov9Tmz13HWLZlgWAMwhoszeJqkLs4bMewgGrwqmYSn7iAcwWg7RjyViPI5shnK
2VG1IxUTTzopneoENElAArXsj9Lb3s8ba8ony+HcM96GgwP2KwoY5ZKc4DJKkFD7fWEQgbGKjqGW
uxao3hQtROcjTNb/8k1lA/yDI7bxJTWxuXn+jpJdwZpy/uci04v+/mMmZFzpCUADU+q4usSO86BO
uRx/UQybolwRB95Ms+FuIC1rtdEfhgVwc2BchAgh3syjynzLx3jEl84E9dypYNElTwi4B/aQDkLu
7xbJDNM3ecwyqS6lu+iMkvh6I0hTXE2Fj6u30wycdleOQqHrgNlLiodZb0Os6Zq/VyiXyTClJf3J
griQKVYSmIk4k61UPsu4xVux001v0SZ/ZX5IKJpjlxxGee05GCwoUl5MT0/RAkvt4CF30KhRjjaz
emwhk3bKSsO4aebRUoV8BOgiC6IDyDu97XJRe2sSfYyHAkz8NDKHBVgpUSvmHwBnHwHk3eO9AdK/
qUN0gd2MJ3mr81xS6C1qW7METsGeJdgfdSTB7JNNhwJiQAlqD3bxerAIesueusq0r6gMiYGVTs3/
gwgAJ68+UeCij0VaWRycs9bvrLSsRGU3KdHuH5ImtyxdnsQJX4Ud3BOZWvPonkJWdgdUxz0Q84ae
yL4nqO5nz5kBd/n8ArCyjhKmAtAS49KkBGJvuLR4EB5ZTVGDWbh4UxY5oQm8Bhnlbxhoy3YGEPiE
78XrjZJwfP/RpCpJKGWOBQun0KhSDhfK+V2HlzB9tnrQsMSJQG2n56zi/RoIbgUH83KINwDTx956
bEZgzkmETN/3jzo8vROVGFa/aAaFPc/Xe+y1i0vNMwUJgQ7spNC/DIojynkAiEzcCUH/i46ei+t0
DeWTKmkNfL9b2FZaLK7yI7oMtVIrlW1nv5hhhNKzGAUN4Q24b2nzbuCMcM4Kv4O577cbdQB9FZSC
P9AwkCu4N9uzhPdv0FbwrOjgHM9CejQ6Cr60hpRvAbbamuJRLB/rUgOAtfqKYUTNiGqlFY8HlD4k
os27vKMnsBERvRM3iOf/IGyciIQGkKGV5TqhJr3buU6GlnpnY9gONgM5ItHC9dt0zZMjn2oAVH3z
qu78Zo2c3xlaBbnGrZ9TN4g0psjqnrCr+dqvs1+K7DeS2jcL8eBZgCTD4QuHmGIcBp9qKcuGPJzg
pmtejQenr6EVIVXIk/xBOBmn6eSxQQX5xGAweGBFXXYUs45aYrI6jtI2xrkUfZSLzbqjR+CKwIgB
zFUqlmF6CzPVsO4FRU3UtxUmJWpR+yK+8mkXa9YJLIE5pJYtdZ2CHnxOQ2YUed1Jvvzqq8iJ4+5w
jMeHkUjznDc8YBF9Hk14NSI9yyN2irOof6sfsSZawcPyFoMJtfGryh2sI7XbQgAPAjn2sy1q97yD
A32HTkbZVOEqi8uDHKin7TIDX7Fzn68p1uWpBfl6Ig8j8UUKsVhNkvYeO4p0LAcaZR4iIp6b4bi2
8GCczMTTpzahH10W9yPV8ne5HTwWliC3m0UuiRfJA7sTdL0/DS3NwXXCDB9ppuwnIdYvLti9on6b
IevV9VqoPmBFd47f83BNy22Vb9LkB/udQtt1Ay+7l5Pe9WrHjQD/eteY5ZLVr/YxKr/ND30kJuy1
0Ey24CGR0wr0IS6mIflfSRwxkv4brpAxgTQDyGOm6p6KNkBqvC1p0c0Ksf6j3GovfGfyyms3cult
hiwy3XZ4hPx0L42HkwNCUCEKuWjQbefVkPLxcuFRaMDWnAvLmDQ8UNAhoSy9cgzxTeFYy+I/1ZRl
xMvU6l9GFVIhh5H1c5oSp3HuvmWvuFMrTg0IZwC/z/TtgvB2iRRkKIP6eOpxHVgQq0g8jELSCPJF
Ua/Qfzl5YScKYqRMoD7wjN0N5Ou7aoi6nK6v970nYwXXHZrRbPYeXxPt+5pJP9RNFwsy4VOvQstJ
DsujFcvDF8ABRYuyVDhTD9RyPejx7WuXUiIqqXCklO/nJ4MgZnLbKBX2RtI14+rS/U2UVQGXIlO/
6xCjYfR18dvaZFI6+WHTvzqw2l88k9hRMrFcnHkCVHZuZaWmYkdc2aHrSeVEV6o34a/HhMrykd7S
rQmf0ZbZfJcAQ0p5M9pcTtCIB1fWEwcjq84l+lHxHwIqbaFncL5Z6v/cgBHReS7GV4oG+Nqsk1gk
hWvGR/BtmUJc+a1zf+AbwP2SR+z+Ihl6MDmyEUsT+BWcBXrb8yWteuVXO4WI5dbRvs4GdXYEtge7
Xw9BfWGy/WC75zJ+xYMdvaV/NH/8rrIjS96ezIF3XskbuYT6zOG08YftEt7W9gbsP8zrgrvTJYkB
92gLpSWyhMOfHC1oZxTVreI/NFuNfoJYXc5Jh3GkOG+8q6JdzHbNQk1Ik9g5T2PBRW1lohDcGsWd
KENBs0rBgMfMmmnDop8J99yRfnIU1S1rd4rksSzh55I5qpxrvU2ShQRxUHvZUck5AHEyGR7RPEPt
jGoi77wDmRBTb1JFUFV++mPRAozbMIYldxgDOm5CDRXZbAf88v2+3O64oDuo7OFDiKsF8aJqqnM9
RekLMfKgmimnOtPnV5GelwVzjn0pPWa/CsjHT8bG/uFaGYPoLsIO8LHJ6OwuAzv+019Zhg/dJ6bC
/6XyQvYht9r5KbSbbUMXCzMR4db6QKq3Jv6Qp5vNJeSdSlCwFSKoVzGaZS89Ak9AH6kjTnnl4QUl
KXdOz48qkbgTCcyCC7E5ESWcuGzx16EysVKYYzSBiwTLU6NQeDaS3kcNExPpgQuXXidwDkndQanX
8H142ZLcwDvFkXFFccBdlHaKAfMfln0crrAdLZLCaciJvnGQo0WBrrwd54OEP0f6fIRg+/tROBBM
O90tnHKU6axqowGsb5Y/lvk1sDDnps3Wll2pT1pWtwpYWhy4vih4OyX4+qZSNJnhYzmM/kT5Myxs
rBF99uUWkzDjLTplvu+cBVYU3xkBZZ8HgR7CeqyAYJmFEBOkXTik1GYX0aYZlXzm6r7MXAC80Q1p
sbQiCNuYEBeziGG1tOur7y6jFFPTECwT8PDub6nDx42s2rw+jdQ4MkJNlK0Jf+ws+yL9WwSvHQAa
v1Xwx2TkBSKq+ey1AXQYRVzLpOtNVTM3f2jXin8KpIm6fvghzuL3lGDOpkTa/i6k9KvE5ZUlsyA/
kxc70C6XtzqZGSp9ARFpIg1er5tLQBBRnoa9l/n1M2kKn/5p5O2IiVGz9XcXGdJqAkDkEC6CclrJ
fhOCNYioBk5H0mhkeRIMlmLWWiW5/6vlAbLbUOIgbnW4mCBpYtw7GUwVD9RKDaW7/yq4v9eYNvhB
vMTcd+C9FLFNlaO/+AG76/R/JrXlwUltGBtm8FMsUK0azl3XYI+X78HIrrmix8SNVLUaMcL/lMZo
0JjbpLGN0oVSalBqSIAhKAg06EjU0QTXIyAcvHi8uhd9TjMkGCeg3C6xVZjnAb52k4qwlmniSi6Q
gmByIBpKxERgw7GZW1QV5hDB0at3F5zxkiYl7UhVj29hw2tbUBY8sF1sx72dIft6aWpQ7UboRhxm
1X4Fq1ZAurh/o+/6yR8Uizxb0gQlbYDo0WMw+5j8rxpPw/UUEXTUcCaY4MYG3ExlqOS+aR84GNPe
VD+Hu8InreEJrrV4CX4HrKZ/B7Q/NR7wjF+CcKwUg5n/ZWVaNqwdY1AMKTwazzm363HdgJ5Kd+Zw
7JHzuSjPuRLqqnSyki7QLktiP9KgxWZmUu81NrfrNCD87P+0cX5vm1qdehj2KAE2P6tUHH88WoVK
Xw/1dpkbFyX+EEGZuBE4iPoFcuwYfIeelzESABzrNLXOtYs+5ELC/fJ/Zm6DgMOnh/lATDLTaU+5
kFtj7lx4vR0/ErcPsLNR6nfESBysgSzZTTnAvJGrBtH9Q24Aj/+VheD7EeUcPCo3StcH5EXOOwxt
iyNtHmsY9aCXF41eqbSKmiG0dANU9jz0yjxx/i9PaUD3j28B59/M1J2kT2YtYEEfuFa4oGfEMSuv
VWvyShXBppXoEYZaerYQRxDSOCG7E3iaPYa17qcXv0oSw+OjyAW0MsEC7uZBsFgJLnEMe/movaEp
7QfWtKJCENBSKXNU/rasjDWa4O9B8uk395KBR4H66hyVqN0aTDfyBbgZGpSQcVD2MshoazqyXOlK
ldvM2F74LejEXpcwjL9cfn9DZKNn1rN3GH4I+UOORhKI8bSqpK7QoG8dGy+29E/VqJii5cFFD0k9
cr817uDHF38Hpo+CSykP3N3W+FF/k23PAdlf5cgY/DGoBk2PQuE02+jXmCCvfBeae62Q3zySDcZN
GkhqbPmcNK2CZ3pZMAs8Qca3KUve3h2Lc1LjOgD89WhOrjre2gYfSZwJgAJWHM94T5F9loVcfENP
4NDOXwK6WjxCcO4tXGOv0j3H7O5UYik30EY8X0l1U7DBqukfjOiNRGUFAxaPsB5aNue655ZfWxNv
udKOimc5Jyf73CjLzpZxL5LCyP10YtJ+vF2YTZfLkqLz3WDgeQ/JqsF23EhNZMRRzhAAh6dyPmeT
vSdyeE2OAmMUxERUjTXFZeUeq9PQQZYSyRU4/o3iAnXcZFwfxsh9EdzUcESJ3LlE61WF0a7b+IPp
o4XkygNvETI/xTJDRE+Tjj+6HB+UJGzMQ05ZcbTSgcJaRy2nvP52AU0/GTYZm6oBP394pSCWo+sI
L3sy/VasZrZAD11ZuuxlrI3/QG9hHA84Qzg2qFDoKUTHnW0UKqwrFFs+LawnGuD3A/Q4CajnjVde
5scPmAh3ebmX21mjw4mA6Sjg7q1ynFihVGXnB6aGkK/osuVgd5d2tiP5ukcPCZ8+PHMhc77V7hZN
GJOuG16tEpgEerZru3lHUR+4ODUlDiHRuL+43gOll3RdKo4xQB1a4yM/ZsAr+jiH7isY15lgasha
3sNROTOZK6fkrxDLyifsO0xU/1XOCLWxUGR7U8AtQTxCOOmqztjnQYTjkjn+vPwIwRM1ugN6z3aq
kqSzj4tQQY7OL5n7CDRXCNgetFxQ4TRHlVJmMG459EyJy2G2kE1imtmZRlOJ6IXKEsE+P1p+ZbeS
qi6+fZqSA6Xmt232c3D5/gyY4fRK5Jo1cCTwyi4H7ttd8c188y0FlZlBsZIIYN38S+b2GU49dQgP
CaPKrhUuvtJVO3s3veC0Z9uzfYNhD93D1rwWvgib7zp858X83t2d5eIR6wNY8jM+BxzdnN35t6UI
r37sx4OzPWQb5wTtcGBrMHFZ45jOTfAiXKZHhiCBN7jaQoPQZsmrCgR4DUvuhLS37qIIKMUUH553
VUVq2AgTobgrhyGf1QqA4xFJ3M8XMDjcodJgrDw8j3T0v6dALwNh/GcDFLVLBOWKlGQgJbq1IF1U
1W3rUrEub88vnaW+yT2JjhpIA+SMYpyr9W9dV3aC+9RsqJvOh3k5sfIDY7jsvs8GLrsbHrQVZMpK
nbtyg/dtYN2FL9yh1aBr9sme2tIsG4FNG2swbeAQiUj5AW0Uu6t0k4Fbswdgk3QJHLgmnsrib6fv
6Uvym1ydogDYt5gUPFet552/n9V1TMJJxI/OIckW4OkGb82PPW1RyAy6+VNg9AIA/78C5pk+bzTs
Q06Zy6HYeNsRNDQu4Lgu090i0gStY23T9sOd/3vJlidCPX5Gx19uVrb4EayFzZ64K+vKQl66DLmn
znc9shztEp8S60ozFNRKnWf/gYUsxppfhbJpQpIaOXbeVjeD9WISB5GxIqp2CQT4H49HcFYcyU7V
fwezsrdblBRD7Go7ujTG1dxzmmet/rV46IGXtqm8F8GfQ49TNSBjysMNKPtQU4pIFuDN8kIKa+I9
6nBrkgGWfsqnUUkSG3L1Jq8q6KMvoQ7rvKPZUan/W3ULyybg89+v2jPUzxsNnTxdMEbGhHYso+q3
T7e1smTynoWAoVw0XQCVSGYVfkriEX4mWIF+9S/ByNjtya1VaG20OMvj4hxQ3wBMDSwM1c/bDNRk
TMTHEDA9rOc8pL1Zghk3qtqzULT8+kgn74lYl0z+jbZZqya3i7h35J2BXiaUBMkkfUQCXyy/YhjA
07xZumGd7dFYV2RMF0hTCChsH2c8S69LLB/2CEby11HSCSptqWniSB+JkyuA2UhX/V98FxcPCOhZ
bZspZMD6sJDbsP1RSFVAi3dTVlTvV73fY/8+egGhlg0skXXINMiOBWs/TpqqkA8nYq60GfKb1R2W
2zv+64pwcHs91XgBgq6T28c6W6aFB/2zA8C2puLzWTkY5vwtvA0GDHdwx6N2ekjQSxjzGEwFVPD7
o1dKNSknrAt5sWqDiwT+dx5KcC5y02mdOutX3J7F4eS0lZQ0vzGMmTZ799E8WmoT84Zwh28UD+Tn
vGKOwTx8uaGG+NnLouSqliq9LprXjbMxR79yDjgSjywXGK09m/G/KynYvuuKjYVLqZv5k9V4QWpC
R9mZHYPcSkT6sjKwpM+g/CUuzqBmZbKDS2P3iQPL/pSZDDO7xoQIK4OojuYJU9GZ+5unWZbUYYZg
q6yHjXKVYshXXNxqKz6dzy1g96U3EkK7A5BJWeAyAkgCtWdqIwxpu2G7/39SAZ2y09/8ckYUpeHs
g9z6964lIWXfQ8XY8W+ymHpcIla50ymm87C1HLRN2LnXJ8YvNyfYtGdB+mzceJzEAw2iVaCro0kH
vsgEljXm8AM6/48J4M8KA/Pj/hWVOpUtmCH/UJbx3cJICi64zTEQZXmSwDvUshAVOOLOZnc3gwCc
QHt68a9qntG7myes+bkR0KJqXrnQQH6DPwhB/+wnyF8bvtUUXaHP+bPT4yx7FaHITfKn7SCh36UF
ffMaBT5Gm6mbECnd0T5VtFw+MpX9vLK1eF5UlWydVuCqNigAGxY6mZi8I1vSLpksXRFyRL2ZnY6+
kKck84T8DeHjHlRlAElzcZeZd8+c42Qwsz8n9vNZK99FwK2gRcmZ0jGaOQttwcJE2sOx54XSWjAP
a45nb5iSzmlKMyeCQWksmdtlcQ9rVd1XlcsrBFq0Jkh1krFVz+rZokApS8IpLwPbvMYENnkcb/BK
Rt5DrsaAkGWcJLIjqZhHd6x3xrleMx3Z1sOzbgHk0Y72F9cwe0FdtV+CXp/5NV8RjYEA4Fy2+4Jl
zJ9Y7cQGAuIMxXzpEpYPFNXlyZ28FWS5cEl7bBz2AL+RMod4GIoLFGMx4nbnODvltf70izi5KwG5
00ShBXWMv9cFNZ2QkikexWihIlGza+gxMXEjnBd+ry9oYSIcXflF4b2W+fd6riHXS3BzycwElZut
0PIIne/yizsNnd2K+PA5w9I9NPQeecLx5Qg7nWMrIfFS9iF1GmwHt86IbKu47+V24JTvsbz7gq1M
m35184grKvKeG0oVoaKB9ueiQc3zCnccDF3+avPG2JCPcKyyjewuOf8vFpsWr5phNvKQxmS5ohO9
+1/kmEMTOrwX07/119QiK9h9PpGRgMLJ5eeYk0bjCK1EzqyLScL1bj6hlqirqpxJnMa2nwtYdqQx
uWvwxv7v2vdwE3TZ99TM6Rz0VPaVfT8wZ58VrqvXDWsvcrSqn64h2rkkR9H9G1pJcFV2OLWY6w1t
JF4xPHck/toKJaavmmcvvrXDOTZ0ERnX0u4c12zSQTmXioCSH3BnHQglcAivmr2/osfCb1V96D35
/tCJ/F94w5BVF5BzCaZ1agGCCpMYFidPSyi/rzznTb66ai+L5WnB2wouz7uvQu+Vcz2mL9eb6mpn
a73Bzfb1t1L0r7L/sng6E0TsEgfPFJnkQ5f3LJWskV1ojIniXub+SxJVmQgbGsdlqUhrLCRBUkJe
oqOWOz6/WXE26eZIx0lqxhTn4zf5nAqmPGkq7P7hNhTqVeeJFKz3jmm/u7+g+UeimlvaWI1Ti2Zz
ftl8hKfUrbrL+JjLPdSjDqdrE+7bjaeGR93c9aIFYdhBl1dWVZjONoAa/s5b/p2uXc+2Tca1wYba
1p4/otstqoKXh21nx1+k51mliGH7i0P85LFLv+idJZg50HVyFFRyulUSO9lMtL3y9fgT7VHyJazA
KY1ROd2tftgcFj3POSs+aGBKI/GtA0XDNAeYUs5cQISRU4Rk3uNO91/a8IZsxEgcxW7FL7PUdOML
jejnnx9TA2adcKvOdEnkaFWtEgGq6WEFoxwW9OUAtp73kWEwkE4YJ6gTa2G+nywIL5nbFVGqHtGO
A/wvPU7vTo6eCe7EXIjuwGg58FL9q7GPU+QZiiIQndVIBgMIrYw3Faq9iomslQQEGVkFcXOp/jZY
cRBOnCajM5F7UMH4EDnTb4TogiIuOKLdSABtMmFtSYAo8TS7UbDQunnavO2s0wyaWmjOWOIQtT1t
g2MIv+nFlg7Mx5lQ6Rga2H01njCaxYG8FuqEW+jzSuzsHaAwYswwl7vKF+Xf+5Jv9kqQRvpvyr+k
4QLkh8epxY3JmBPo3W0uG7ICZ7q7mBqYsU0YpRVpajTvcZopVeUX7WUuNTtuq9tMiyjTCxPw8y5R
b1p/AfyauGMUInYtMEy3gJefQvzpnx29w13Egr28icqxq9etzB47f7tVIQ0rjkIRLTkw9gpDq/53
JMsP+tSbzj4PAMAFUL7AihsyIrPy9fRb3ibFutcdDR7hRPTHfi5v52apWiQYhaph9LDorM8Zk87a
4jW+1Z+PZpsIbVNMTVXTtOJuDeQj3zzn8KhQarQWLbsLG9XagOeXltIXflbEccoeraDOYEDf03Ad
v0LOYBo/ZuyLp/ALErqQlXbU8nleAwv2WMHqKmabR9tdXRITrPKCCs1S02N9XDEiPkzj0kET9AYL
w103i8HRmIe4d1VydgnTvQiQh7RgZenC64j2Qk8EcuGMBX8CHVVzdUIoCbi3/aA45ZuA0FfNSd42
dpCUR0JzHKuXZcLkXywrfbg9MMMX57yanhlgHNFbRTa2Qj6J/c6Rf6seEo1BGbCmVE6QVxSUMEqr
yTyW9Nm1ScMAywd13Wb3nCFf4D2ol4joYmjE4AMHjcG28sb4RPo94+cbwobeI49f/QuO3NujdT6g
S1xWeYuIxMy/t0axI+JI3z2YwXnMk6x3tirmKzIL/mwGBySfIudldW6/8RHjf78uJuLmGAOa+4Sz
RCjkRtMPMNaw9rdnz6jROMYxCHelylLDN/6QjwRdCZR/zbHsjrsdOGURe2FFt31u4W2xNA92ALp9
PZ4JY7SC66aXkp1pAH2pV8IFPOc8+MgZVjLGheT0En0gxCW08FPzj8+vTb/nw8JMeP13Jfa95HxT
V5R5sceWFDCM0aDGOBfNXhJpEhgwRGBDnqF6DfE+s7hNJNh8kIltw9lmYTfQ3wgFj80dF18K+ggi
eNlrPXZhRBNmjErUoaiT10D5z3hjhyex7Mpd7AZKJVfd/n7FA+VobB2hJ9ekx1d1HlSciDtw+xAV
Ge4b4RdbCrijEApaSY1qbewTDw5TCbIB7ZKOSrg7uA/6mY/Kz2kbqYnHD+Wk85gO5JcC+Uukd1z0
Ch74pPPBQgPhMp/LdMW735ka17/MJfWNXIlCLbdrcikGhdRIqSCH9d46FMjEJ2AEh1Qyrp3endTW
0CKLXrtuNw4EIhD8wel6wVib0RcrxiShadYCKFGW32CJcvBJQ+VY0F7aC8gpiyTWHD0W7t0ENhTV
qdwmqVbyS+vX+cOeYCXPk+eTVKOfz+k0BS4nckYQ8p07r22GdL86DsaszXXuOHUIssObKiP9TMVm
e9WDP6taJixM2Mt7OOMcEEbbyLk0BVsDt/69bpJD6OrEZ3Se+TR1Cxm67HwH7i9oNnT+SUxpfq+I
6mYIEFSov96KPP1kM66oWobBTUgjnVhmCEFjcKQLu2PfVHh/SxAG6/zv3e9sNCCXI64fR5iV6NgO
zlBBatNuE6gnJz0EGmByyTNyh0k98vKumLv5C1NXXsdGlFsrpfxq3gzrAvm2XPdoiDWpsGoEFA4d
/QKydLi334w4BOCLt7A3QZsFalWPLl62iIZLhkCZMpyuqbBRs6jyY4659CQ6lbMHHesJ++4ctiqk
5FRuzPo9dDaDAHFzm/2xb9hvWTPJF3XsNTOqQDAOi3x/qJT/dw7af8JSaOVqC6IFo96EJ3JgVZAH
YfFGNTca8/udXmEqZAElPfzy2NSZJNAPWRHxgK8d7T29EpezEPs1IsppucSUqnzx4+gYahU6pHTT
Dg0Te9sIcmaPFldLdJY0nLL8f7lhEKYJwFbDGWTlQyw1sOAgnDnI60uo1ka8qUHAkFN1AAA/zRVx
APKR9sTC7VC60CkFTmQ2W0al8P1L6vieIim6t0lSt6eoYVUavMj3ZXTbnD0BITsQstm01H/BCQK3
YiVMi0041n10ZrKxYG918bdHpkAgk7nZJO3JbsRjGbBHoNQKIl+0NUpzpoJW09bds8pfr0ZBr+JB
2wtQDUFZ5RwRFQAe6xTEoRMRNnw0JdHcNgvclI3a1K//QSX323mZgH1VG9NVRXETSDTuW5if71Hf
N3EOZtKa8meNLwNFWUqxdwtDm3SCsonyeijsu8YBwPsoFJc7Ew6Q0RWbBPSOMrECnLe9CmU7HCHd
yhXrk6lj7HNVZLDymW6Fpvb4gYnuJ82H59FMa+GC9gxfZZ/8D5mKPypBbcDjbWLdV6iXnDzGFGMu
O+HM8v6hdmQ5Pnn++YRLJWub4/bnUDaN1zAFYxK+4izl6FQs1Ip5cGAvSZJbp6bg5ry5hgEp+j3C
zPZtVY09zGINOIYij7RYfr+SmvyWPi9IBnW44Ir9GNic714oy4G0ugg/0K+4IUdxA13dHqYpbWBX
Syp/ymYkAj1NgwpvSzvDBP+Aafxk4lYkwzZ2TJT0pInyIPvUplAVd+EMLNFOoadvYS0dIlOV8IU7
zrK0clx7+5V8RL1Zkym/4Lf7+iaWieIkr+YAae99upPrYrfYaWVySz9QUq60PkE5EzngH6NYihrE
XfUCtuo2k1agrsS9VAyckdPA8mJcJi/oO51uXI5Ez+EEwzqtq+Kgj5K0X7qAIK0i5sn1YWlhMTRG
pWGxutX1Yutet6ZT+SOkF0NtYIo4DBq8LNBl0hO8QDp0L2PV980nsRoFzssVdO+h/CUNsYX0Iwt5
XR4p306klYMElSBdNRIp8kuM/K5lMrvQSIkeJKtfDRuOTl7I9tRHzfeTo04W7PcVKi3yLeKubJBZ
bBcFKjq7bAi3uTupmlEdHKynQtXPTnz91b5ngt/ifqIFalyGe57gsb//sPiXklefoD7S+FksQ5S6
6/4wwtKm/Br8m7lNwNgrp3yQZaJMYlsegu3Mxl+tL6Ax4xVZ91OrF+6G6xZ6g3E7nt22UIODKYxQ
EYrG8Q2Am1UyTUcSdx9fHJf59b+0zeYNfho5LKDP7rq1e5Qab9i94IUrRLg/KJt6fWikOVl+XKgy
XfasMNBDF6Xj7kMh8zzdQEfhjma6awgoOiAEuDDi66V3HRcMqN8x+TuwGs/xRKXsaY+CwmpKV4hP
gVxZQz3Hdzwi9uDUhKmPOqzZlPXr/ZW9Yz23RpyMXUJzI3OAxrUgy+Rc5ZI1AU+oabijaWsgJ5zt
MQ6iasn1YIvLUmSTpc1L6Mpr/nAlFgUyFcF91PsKWWWiuqUnr1R1UmC7Dwrx4XoDi38QKGrK9rs6
H1bzGVKcpXq7bFkS8HhbCbpnmPwjMMbOL1QMK67Zk0yIBWGTJ9mqvwbeCH9dGTEs3h1EZAb9FLDT
7/KRUWd/aJaNtujjKOvkLDZaDJrVBRjefYckEQz2O3sM3dg434dhs/e5ra5qu7zcBwJUeZgJ8E9h
qLSwgvr3jUPt9wlzGcZPK+phCBPu2I8Hkwjtcki/g2RnsNpi1TDAEgTcI2aART7IQN1ZIp2ZIo6W
1AJUWzfWRHyHdrK5uuvt8dC/LfyhV5CT05+z1cnm71/5lfFUUak6SuFIGNrOWyLoc6LU2irkBIwX
kgraC6cOtbnETv22NQM9oEyU+XjLLh6RouZ56jEQIJzQ/RfqRraPc+4tMD5BWfwT8+dCZjhi6csv
lhs5PDi10sTDuU7JkFExBN0vzda61yDMQ9BKvDBRo9pCEM4GL0IU9JnpBU5/YppHSHOe37amxIKP
P7o+uYkP8p4LWWqITxilC+n28wpLVWExDiEWT/i4Y8vYfdUzDfUdKILdls6SG2p8ipf4WdXEprHY
n0/k9zoUEZQQC4dPmjMvAU6AJ4YdAyjV9pClEDB7CZX1tmktg9NV7axXk3Gyl0YEqIeJlE4ztZwZ
8dtALVsvXxEOPDz9tuFV+SEC0RI2tdXKb2l1cEloHrB9nX3Ho/ygalaZr/6fAWxJbXbylc2TXJ1F
ws+xo4ySrR2nKgKlrggDKXt1UUyv3CTD7ehnWjD8X8FFiRNV0kY2Ceq7HgNRJlAOWiIZ+I7F0MHq
Tr9Sqt1l/0xzIP9pBJidlEeboisi8R1Sq6uXwVR0EqOGimPlQdUB6C+a1h0nmSvMp0iI5X3Jd9yj
7K+FOm0tz7mm4PID5TOFzwg7ZzPBY+jc5iY/Wi7pZqM0z5Ip6UqhGaJZLiweS9G0yH8PWNPxtduO
XvLFijmpHPUJuPC32imdKBBcpATbaNjmgRp/UdbNUXGmS/TqACvT5pY68b0kmHwijKzNHRzgsPcZ
wLOSQG3CuZzXkDvgXCQ22w3tu9wAT/x/SSUS96A7zm1AgiW9kf6LJ0frOWEUwzo7fMoplUPtZgu1
ykyX7YsOxVWYvegXqOiA4z17JE9p9SPBFCI3Q5miDJYRpwaNHrZiA/zzuVWOTI+nvq5uChNPi1J9
ugt/m9UGH/Noas9/orpSgpvt42SsiPcsFOflmtkHT2cD26WhuFSahcU7YAi7rKFIq79i+MEzrf3G
js1ss6/4dlO7ELgLtJf8erk6eTPWisCuGT7l+VYM52D5as8/S/rL/lPAq2pGdgi2BZMmx3woQQjE
y4N92SAaIFf6zT0oM0J84bqFfou/W8gXFZbrD/PIHADuI0U7S4hWwp7SPlLj1wLFbyl710GQWrGG
OyWy5yi31Fllh4aF0j4DS53FlA1rSwCwAdrZpsZPbKjgjkY4ari7Kg/Y90yxjp3Zu7bs4Mj83Xqs
lz7c93CK7COZ/hk+4gT5JRcnayJjLP36fl2Yx4S6E1eQ4cMPd/p5XN0lWgH+lX7fXHke65x8maxU
PISY08wt15Ks0VFwNTwt53qKOYxmJFBEg2uHghLtUBpD8GFQ0ya145CWNbgtdv7Cc20m0IFWtPVP
RScr+srlD71qWduVplIK6hsR921YgQQFB+sCR7ARGrBbvKoEt/n2dCSr4tXvQXJyGMcf5+8y4O/g
CXQ+FRFYonUp5ntIy5o+RGRFpZEkyNFG4AYb47C06vrWTOvlXzxFcjuoipPcm2qyQPda+X7VejRy
vlzyT1pyzNwTAXH5hUzFYkCFwguqXvcsZ5z4Je0Qo3xrkV1M6ZSdsnpq/i4lVFmkHSRGt+6zHpqd
FtgEmiYbWTOd6C4ReMGWXCK2g9t+cJm3q897d8P6xpjT29iZdronvpZ8eUmax1vYRnogBuiM3Afu
2rENtMMFrxW4W21OECn1U4dppmHGrAbTPToVzcG3b2JV04+wZxmuQvMYaNOQFkbBL/W6y673V49E
gxLzCS0W0PAoC0Vh2no17xTom5KcV38V6JE7MwkZlUO7gh8LvV/Njzt0qOPRTKBXZNlCBYeeVLx/
fqxpZiEsu+/ACAaAkE8j3Lh4BlF8OoBDp6cZmtl0JOrsJ0wWNHZ9OyiUKOdVpzXwloEW/zaTaqx+
kK3w2yz4MnvsuxhEGlqIjAinZXA/FiG7k1wvm23K2pocXd0sKahRLYb+vvD6TolfXLOM+6PsyB+T
QdlBWSJ4FdFj5B5DPOFaaoVknOOi/XyBPKSHpOTDnKYx6AGaqYKEHWK/Tm3J07PT66/ofEU65U7F
bXj8EiLaej/X3849vl3Ef2Gfo/28YGCcRJb5DRqUGgsgyCRubakHrdg+dOvE3tHrShLfcNqJAhTZ
8DxtQi6hofeS1afNxYTugAfKx7qZ85DWiBI3/VS5XfeRF2jw5sb+60xVBCTVQ6gljanI4xxmi1Gw
eei/o3REO2r2SdSbkk29P83xl5jP1zbhThiuTL10vc6jhDhncpkC17ehq1eepKKJgccvWqCrhgKb
dcPT+Rs+5CmAteDAwpNnRNkSPva35wcVZVHRwE0bvAXrPWyNngFd6Zi0qRFtIrp7F/eKADiRz+ME
tN3nyRKakw0fWi2ZMduaUHoNBS430WW+Q3g60GdLi5GGH2QfCZ/HiSopoUNOL/gKMCMoyLDf/aNJ
KKtcJViuYU0H4gnyaaOugudo8TiXSWWxlT1zBQvQyrdufjrvXaYYhfKAa9eT58voHFIRHj1xe0fT
fsQrmgv78niirGtR+tul6lWHNIzz8JfyHQ4eSH8LBl0Ga8KO5M+P5KGXzlAtfaYbatBn4VK0q+6L
Eeb2LCyThdJZcap1spWnNYvPvEcLQOobXCbOocfpyDPD6h+t2pDmYNsc/PDAgoeYH1yIr0wQqOMf
a50oL2EKBAdBOx4yeoCCbmiXdLRTEiOX/zqNEdKc5PSIZbzSmINjHvVTahX0Sr8RufNpP7J0+2HD
ADVijJpmJpGFDMvj9IUktsZviqqGai5icPbvpnZwFVPv1aWbEJcint2w0urjMywlvD5Oz2EUCyAM
XfPPww//5xN92mZW8/xJVuNaRn+MeIgFW34OZEijPFwwpK7/eirsobA/bVzBGGpXXb0+rVuelSTy
ZXG+au1PoBva5WXAjQEAA9LOSD20SS9Kic1Tec9MPERnIL6bLmqpZ+1loRQkgua+710QERaLBPyn
+8caX4q4HWXYgRn4JJx3BddC3reW7l5ma/ttll3WP9Efft4IngRXDYl0fwYYwF57NerxgV0KoeZD
aEvfRKpIHimSv8v4OVbObBxKlOVTeIQofGt1yMmbY89XC+xtvWBF7LQls17jVnFF6X6LdazdBR/N
TBAa+GBGAFiLFJo6U1WtaZnYd/aqVxRvTnOLv6K6s4fTw8pcRqxRp1sufs1XeahtT/uAbfTTh1sr
v2lTl1xG/1GkZm0n5oJd/wyM3f5PheyhL0QAk6Ysji8Gy0u3CZoqjsC8az4WopcoidHmLFHXGpdy
ecPU6+seXbWSBnZPWFrCcEaQjHrwz9Mw6Tz2w8kDA842ydqKo7Li6WgsU2B0XZHJ79RflqP8XD71
wizlvWfLYmmBv7dyUlWNrCVq5Zci9nVHkX4LcHbafCxLQXbstb9f8gosQuo8vDfa9K0p31Bi67fc
6FEUVVBZh+37HhoFUMNfj2/Q358XMjTAIFTesXgZ7Sq7BfMby6ndmTRBXxbULg//Z6zTh6D7S9q1
2lw7nepR5Jf4qaDseo72Wt/1kSPHFZyl5Z5Vuqdt9CYNVsPz3MfzMyuPPVN7l6IwIG1a3EV6FKfl
E/c6JnnzosLBU7ELFfJJloaVWudbZKIIr6NeXLeeW2Fa+KocWQt0fmeO8DrRqgPSyfjF65ddhSya
QLeGoX3xa1aRAaGOI3pIpxr7YViRyGdcC7WaMe1x4H6M3vqsDm4/WePEyCmEFu3T+cz9Jl3OOhlj
YsKeb3hSLPqrH0NuOcXKwegbeCVtSMjHT1/+DIn0XQlbY85Gz4ZHJwQUtD6gzIG/WMJ/zwIuXH6K
NEQim5mEOOcasS9eEzb0KFfnh/Mqof8ap1zdAdnTl714LxLc1TKxADY9H5VtqO+/QSj0vnS59lTE
RgKVzGtnSchLevF7mFuxio8RT637xvyv/MRunKGMSrJ+O77yOeSqUYRfYLDkGM51gQHyQHJH9YT5
2CaBOCdpclfUjAX1CZ3NrRN/u8kBKQpwTFa26VYErGwWsCqAReTQEFBDWSHthtrOez0E6MnM1Iuf
wElS+blxW4a9ESoURkAAA0CXkZnj6mtYcT2CDwPYA8WcAAh41DZK9MZeGDrF7S+nFWhEty2H5B8k
y7xoJ0lRsV0KPev6KvcEeNTo+McHQiJPXveF8XRUwF/CL6lCMa09j8nYqPVmqsfrRTlUUKY3DDRy
OX2EP6hUSlHCPJSubJpQ4FxtF2d9ZSaz/0ZR+aP9Xilq7qTq5+higH4QIKgDFsEshU7iFGUP1p/g
7nS9tnWSa8eQNLLHl0tR05F9TNk9+yvppu9rkMJS/C7IfJAXrmQn+r628IkPRFeK3xEOjc+E5aOG
5EW1zpWm1EiMJemH5HtIO3xwlrAspYerKJJVXG3wfag4o7hk7+uTBWqVxffLNqpqO+wOf821quQ4
A0AZdjnaeNCwdTEvi1eHytlEawMNmhY1j+xCwX31nEl6K4sLx3uBNqqKxhAccdHmwXcHhIZ2kedF
O4UEJWLoQQflv0/lM8Q9QKLfvMh9bfISYkv++9o1i75GE3f4z2QF6EEBQOwnc1/YElspHyy09OEZ
n/0bXvC8I+tz97wBPigOaCTYpavVSv/XWylgXWekBQLxgCc/9YMl3OXZy+EHAC4smBuNPXIfGWIn
PlLrCVFtamfe9oYSpffikA0WPyCN/E8FUTTeowQp/NTQWJ1EZ7Lk+VQoUC4Qm9nMEuJ/ZwglBLvs
aY6OzvuO+rwFOJG+1xpd6MiyIJ6SLcFQgM8bLWgncbfF2SjwhmnLkvE/61FNYBw0iP9U8xGUCfpW
m817B7wn0GXL1bqxhvr7onO1KymiWhOJmk8ODsrGWEjcVPBxVVKWGwZhuJvB6nwkru5e2Tr4ER4R
YfFpxjB/y9dqkygBNpBA3XCSvfK0j/1mZN0qFH7b8Ghgl4fn7I2ycmgQN2w5kDEhcFBMOFbhXSy1
lugCo1yGA1Xv08xp0skoi95lmEdbLoYz4FLm7McAv40YmWGgvQzgToAvAMpT6jybpVvpHL6f1z/g
Up4+Bg0tDwovbHG9TD7wZKf9Yjshvxs6THgAA41c8/JQBpBBpKsOGp26mewXK4unQzJ8gje0EYRl
CaDVtOW1fkd8EPcxH+awFtcSgpzCxRpjIx130rMh9VBXYNIIHoVTpjKS8awnmhyjyZUVk2jZJAcJ
ZRpJwhAE8OcRV0qfDyPRc1O8nfrykQ7002NLm8+zMG79yd1K4nL5pgXOWyY5RR1XRZ/LzY6OJkQ2
Bjmv9AbCjkl5y8AgUC56P8bmeIPb6xL3vYS5/xt6TzgEIG5gk1WKko96R815M5q6//5QuBDymheZ
hewziErm0q7dc8g7gKWM1kRAyLzz3WQkBLrawslDmZxLtbY+86CFEAwVMbu/CqbGysVpUBOidD9B
mnM8uqLZm5NgDoCrwo3PRoKqmWEgV7Pc0DjWrP3J8s1t6n51qX7PBok/ADvrhykA2rV70pqlyIr1
ou/zEV5RK0+y6A1jpK0aqLlXJ6UC4f+YnAOEDH+YYphwAb97/JZtaYOQ221vk/k34+j6vtehfBZO
oiescA9PvItBI2L/0iPf3UicYFUp+/bFJZSB+4IoKmhy1MT6fktuYR7IV+R+orEmZMX/yKIa925u
Ftbp/i3m9oqTj6VPvZzgnKtqn/68654x1/luHWmWIudUbVaNVKnZtebEjUTNvCUGrgMi0PcKmKDX
INJ/AKqWpeItaxT79JkdJQQMlLaX7cVCSsW0rp2K5B8SiZti9eEVnm1Bh6xx613YdSHUnQpcXKY6
Ckxadzw4ELDYImkQgf1MR+GqT5lMKVOBqnmEyRCpeahx7grtQwA+Iy6h82V9R4s073lkoujF40AV
TXp3euIy5qoWNv89peU7wv91I8eLiyGDHWom4+/3g1IlU3MDnoce1ZzZK047SLKj2k8FQ1Rh3wRs
eTEKBe4yZkCH9TLYKW2HDm8HuQEm2t4l2obnGJXEoviO1bLIRfx5Xa9Ffieea+JXzUoo8DaZxWwb
5DCaRFgehqEiQfKg2lTZwFg4bn2jszLIK+KKv60APLy+LR1biuMZFPvbwyvQeRKEQmVKbtJEArR0
a8uxL9rvwwmsRNpxIXeEFPbnNLWVPLmWGJK51Hrg8aYRjUhZRlDe4E54Ydj+kwjdY6+zlTggzCYv
oy/wDmd7iNtI4PKcEPKSjV2Mlt/dK+74kfDLY7kPRphygNtgaPzs0xqSGvLxdZv1TyGQBwtm2rpe
GfdAuHa7CIHxXqAzAhTLUD6pJVhYLcNgDu7bSFib06rme3OfhN16pZoJQHcp4+3GR3OcvzA1WgKO
5QCTgCSkU3HeiPa45wvq49bOjZGZ7cmsVDoXU0l1rqeDYjFa2nMb1k1OtbjVVpinbRqk3TihTbXB
d4VP0vl+NiUDn289mAIJ4XgiAULpY8XzHZshxoCoOTCNc5zCGxDsn79t700oTuK9CsQ7aCGvB7E7
Bde26ZCimi8hFIdsQuMpgX1KqTfJlykIsxGm1J72T6ah6zBv1LcIMkKJK8CdofhZkuwE+JRF8EVq
j0Gja+rZSzgDeziBTlQr4ZCqvz2rz1EObzWE8pfQIF0p8jcEfYVU8nH0NxLTEPmcnbp7FXAyGZcF
a7SMtZt5bTgZoXUFqpD04ilMB4JVV60sTui271pWxIGzm0RYxe7IDIGtx2H3A3x9Mg1UUr7P+RoU
lyLCLwWqvGTdm/uP/jp7em3Wmz2hN8E06Xs4n0LYEU3Bgrf82higfSMW5uNZUWsRzLLLsqS+OoVL
IxFmWv3QANOn2ARJ3aiDcAr+D0W096aP+QWC3UiaMGGQps1xCap+zlptPNr6Sl8ERMJ0vfcMFewS
oQXPfoNLaVR/3wpBp0tipocJmtEVLPbovJrBx5qpje8/Ffwifi/MzLGD4XpzvDXfG65T1z6vUGCM
gPIEvaYv/e+qqsQNcWxy2ZNd4ZQuIenl03VVjIQ2SnoGdtyxH2rzo0SIB47EtMYlEZRWrOAYD2mf
NPNEpLL1VRdp0hXBWZhMnSH66QRCC8oNsgUz0t0MkQfxbqmMv84i4yeDMvSOq8zhSyJ1+KEIzDPC
tQgUbOzZ9w+YLthSOFqeR7jDxSSzJ66SSHnsL4mKjcnX/3KtzMiSMK1/54WbXbtd3SDaWcQLg+Zk
qyDbJu2/L2QpoBGheZ128ajl/aO3r/LG7Tj2vhZSPAVktXFHQity8eBWatOU2PvGdbVgOyllfEjw
fq6ACEe/TjoTjy8V9Nf/muvHPAGWhiRml9YRwwCzGYmz4lMNiyzK/w6BUfRl4tkNDJwqxWuIOOdg
XxMvp7jxytj5VQaCNNZEnhLj7QnBRt/7WrZuxRrvtKr4JjuzcvaeihK6EA9oqI3BKfadOFS99YWf
0exa3yRxwqT4bP2UeGik6ituURs19LDmjwS2jaimCL/JeiBFJD1+wyjVR2r8enMCDeL8xWvT2Q89
3EzkTXKT6mI/Pr7l8JUDUlT8IQjmeVLVPLqd44qx/2MsIzw8cAjKgllCI0sZl5osuyx/OQ3yFAHR
kSpXA/23Q1dcT9G8oPV5JLtJj+roXFswm/+ScyhvDTMzf+wiybGhsPdI6Y6W4dH5LfqcSx7MnJTI
pnYTx3uvQD2gdXyx+PMX7nC/bBKjziMaycl9GPjwGls8Mjjik3R590yvjm7GFT70dtZNOGWdwbIx
Db1C4RbGOC6B6JGdnoipdmw7zLJXoFg1NhiwQunh/CBcB94IVieZME0gtA6Npaf8pEIuCIs+qP97
mB4fUQTazoxWgsk5lDtAoog+9lQQk6jRMYBawE+5N3/1iuvDEvfx8eUh8EXITZdLP9tX+5KRMnuw
EGx8pCFiVRfVGoiCN7e4Y1kHUBZ/ocpHP/v0UZQz53IdWcbo+3Yhnkzm2elyoypUhQvBvVikdd8j
OPBT9w0Ra0GWTB2IBtHWEY0vAKTmXT0a1p6tAGz2j+irGvEXUZ9AnSh8sILhOnFVWnaou3/Effb8
wFT2h0Lo+dcBy/bYDITOJyfocNBUeMHZ//nFhGe2FXDyEZs8BcQ41B5H9JzP/4g8lq2gyMzgbtHV
qtp1pgzvw60iqvBxEFj88rzd77IyMaqecyFnofUbVVcGA51vt4g6SjZB4x8bQMQV7gZAeuo26DVR
IlwMwY5IZQfXV+efMUghwt5I8Q3V8tvMazHm3lWnf6jLdHyYAp2SAwFpSaq5K4olnYT6C3717ynW
DD+Hlk6jBXMKYS+s3LCjCmktB/81V72ku0+AI0Mgl3eZVDStSBY1pCblw00WBoa8yB3H9FzsyZ09
LvwQR/SqnIRJMH4U6k4YuSIZyiAHG2v7fRwrzVevZDvCT5p+eQfFmUxxPOxM4Y74ZDDtwh/IHNZg
rQLKhPJS7MyDEoZZItYBIcdXyG57Syaco19El+NJyu01V5X/809cUnS+lERjfV5WqB8Xilghb58h
Sp+0d8QRirt2YJgciOTWDCXw1HagNx87XXzHAarvkRJdAPQJmsRwCmACr1d5htBQnb8IYKN/UlYc
A3e2L+WFAh6dDqIqWsU8TJexUO6A1sF9sX3aaZVnUWVvUfRiMKb/IbelWOzN2Wd4jPXMDNR5b7t9
pRLoom4jvlcDgx9bm7/ntPb1VJcbe/eTcXfCSFaJHYZALXkynHyvSJZ5Xzwhcpk5JC2teLOLt1P+
OMCc/8BMNwCoxbpx8W7rgBs5qi3HDNhDJjkpsVQPZw/7vODR19NfEQIEH61GnCZ/zUV4KKMYOwno
s3GcpND7jPA6SVW89Sf1agKdE91GpF7ABcM1r6X96zLUChw50vXsTGkk3khpMHQquAgUutKNuv/m
GSzm2n022bzdE0sNCjIiYopedWlJIuC8mjSZmbn+/w0vtOlXnzeKRFm3HEA0Jpxlxo9Pps54C/VU
FQfaFpw3GfYfO861kBlbGiePQxZuaIzvhHlv1c2mpjsRRCm2RNBQCe2F41eEbEuTkY67dJ3NppGN
Bh5vt9HIlTfJdhxXKuOgVd1xe1tM7+SGmCWD+NzMnn6Vd9dnVY7h7o84ds0UNrXcH0CMN1nQoKaG
UPIOUfTJX6FYmAOi/5IvrE9D+6mJsLqSQ6nTb9IJh0Fev/B/d4uXVLpCoh8+/VB6ojckzfY8LKnA
lOrgHWEF1z+5qnMnTSTrIp2Ui9O6U2eh+p1FWmgK7iVnX4fAsgILeHNFud1cTyJERuQQT3+kUdjX
BOH9lZtPMS6wU+ETGcgHmspLn3L4y0QnTen1kRv6KfG+45aU+bCzaCAr80hwk90Z4EwDAQjVaUqM
2e/3StIbj77nAVcxZRewn74fe/MsLyj73ndK88rnuBu6pRSaLHMnVEhLyKDtXCx0+eK68lJkG0Nn
VXqQE9TrFwOWZzpIhtaaLRY1AuSlUVyfT5K6N1nQ5zopQTuBzZOUkABVGo8mGZat+6okWU3iKKJp
a4G0SNr5bdBDyGTOJ7aILJ1zbcSM7ObEyhhDduJgiPZ5wqkDo1ioNOK3WB/i4+RYuN5dC5v52zKg
4dtiJWVcO712BRTLWsDI4lmZn2oNsT5C5RdkXm/vGnc9+rWJso8xnX56AxVKgnS6/jr6rDffngl2
FCPB3hG3bwjkkzSr/lo88pb7daINX22eTu+mgMP1zvjV79Hwt3bp2kBfGv+IRksq02zGM3t7F4ll
FZFmpgKMoZoCgc8TNpywAGoJjjDo6OW7jjLeZQ0QVhXQ+kSROmgAZLVOo+Xlf3Gs7O94orYKDeHp
wlg7vm0tXPOiyWCHt7rtHpVf/dSsPKUsOVmPUBDmibN7pSQhinlA9zXElMs8CYYrdAU15vMJPmNj
RmVtktrTT13ZlIThiL921eKXu+cxnQ9zyc81i2VjZ2h2hu4YbQ+KEbkMfZHc8xQrGvI5DdksF0er
5soYnGra5cv76+dSBYlcaB/ibXrSxgBB2cIqxogSv0z/4/RHhASwuW98hwq875MlN6lhHQ7GzXAw
UOiKbXGGailPrjWR8UQOLkOg9VM6bST/0EClkOmxMTjK5lYvoARP1L1woMzLlvwj/ZX2l6ZVRVjG
eQOi+Wn5s9FEYCK2zqTWx7JS4hQTJV7PhdAJ11S8TDq9aUnk1t8rjVDoCnO1YuN3ylsr2BAXtIKg
bm/ccgI0mDZeeTJpqVoGwl9udkg7ExLiCD5jOknUxppSr9jL4SFqytBw+nCTMq2MSLPDTPVV9Y6R
kqXoFPx6LtJ+6zHaqFqWSVdtmW506+j2yqo3OF6e5bBihYNxsyrHzG29lzMeK2c6e6G/mjy7DVkV
F7uFSqMEtuRDUZXxje9Orjw+nhdtDaeP0qVQW8zT9tzgvNsLi7eGyNgHf1bDe6BwiRz1stzOJOWZ
A7rmrhcHrBU/TTx8MJItUmoPdtiApp3Y8DtbEhBx+HGYB+QCkO4jmz5peI/u/CH5MIIEZt3lg/nB
KWlRSojyb/a0EALoMivTZmEUjhDyX4A2YGeOeFeKhPZYu8rWP/KoVKBgrhmCvJVsLNVBmZnMIJju
aQ8qxkugB8j7bFpO8GriILXDLBx/2TCw3CroGYy/WUjvoGnFieBzSsF/v8UmnEOWhIC+6QbSPEUp
YOaISxpq+g2KfGr74C6K4HsrquGrcEXZjPem6aQku/ypyf5uVz4XUjfifZPKg0BKijGdqWQYQgxQ
xGwkX3YPmNPtbvGDsTsFw/SVyAkybD18tE+AHPk3vrk8CKfaj3RREyTNk8KoqoCfZY2ukbp+HKWH
gTUOeQ/INElk+VDv6tXd0WLHose3X5hgcv6pPGO2gvbIDUoaV27VTobnJ4ENINw4m4TvbaSAq2ee
IeK4tHctghQe7N+yk/F23yaAORwMpGvXSaUg7pLRvE4YhaMAN76Eawemrrvogk/4OTX85IWU2zqi
+g5GvhZn7xYLOdqBxYPvmYBCdqbFNa5QSyIS858grHFg21IFDKNrHi2s9juEcc3rMcCY08wUK9uJ
mlWlPC2Hy+1ADmthIMeuHqgW4Z8da80q0wfbjlKZiPVdf0x5h1fzmj8do2K/5cPqnEFc9UlffdvE
cpBSOqvSmPc9tiG03uasmSfb2U5OLvUSXkGxakyLi3LnxBilp0kxaaDyvd7v+jbHuMT+nDPExCq+
KuboD7NT6LCVSGPPluGU7GXgtvTNcp1+NNTS5EWxMFDifBw/kgcWTor6L5P0CFVHow0EZAw4ByUI
klV5/IBwfEd6HXB4WL2MgP+x7WDEhXRx7bwmjpr6VUsC2I80G1rqsVgpxy2CVU5zvAxkHr6Layrs
PjljkpDc2AjGMBth/XoBNftbE4BeHTa5CsaF4f6T/Hjhh5av8HpiIoR0GFUHM4WvLBg+sSOZ6KwX
UKzcS9LcL7jV9x8vfB9hdYOeoQy/ZMfB069YMfpWXOM4rltkklma214iaHhH0vYXByVVHIur1IsB
gtGpWUh0FilIMTQG9AVaV+gZWt8+KWFMkz2WLbTKCcTjrfLUEw/hhesufU1QKKzp5qqBxC934xjk
X+e2vfaydmslE7375GZpDFGwg1w93S5LyMOg8sjDlLs8Nz4EFqbxGU6PiIcwvyFEMkYy7tz132CY
4tA58nLYEO/00UluSElVsM6FSd5J9ESqH3edvtM8MbrbPX4nI0uG6XvctQ8+KM/oEGbHJ33m/G9t
TXIwyVj5tDxjtzARdPBJexwV1PWshmO34uoJWJocdoJGwaYjx8DtdrOUM8XbZICApMGQniHj5dRW
vDFM/961kGDAXty8SNdUAjSt+BjARlcHh6vi4nHrDK5HK1EPOp0RQk/Fo8myRxvGmtpFl75XqTmf
11dHMrlJ61WSdVBJ+Mx+nnkzm0NKtvjJVYg6NySNJq9I3ffVAkx0hrWOLDmG3Ew26ERLzMjyoSFH
F0n/k1d2uu5+L7DKNEpR+5mZ+hZkBHFycIPoBP/qq0uYpWIIbtGZOx/yi1dk4KBIcMwgKI8+b4VA
NfsqqO79YeiZGnpmhUjRdcBYVmySWpxnaStCs2I8uR6MJpaVxUZpD42uCxxOhe9Dzn7Wc8rNK/WL
1MZEiT8BFCPOMk6uiwAWz3sVlaaxRlexXOlBbKhQqyqcZ642wWC3+iYh2IsPvSmCTPVX/eVLdRrp
GNrrf8taew3LGq63bJk0dBFmCzgsfRFGXQzPhXZAgDNZKC2WPO4IRE7uB9GxfGZci7577OJYnDHS
6xfYXKGtq0I8rQ+81Ygin5VxNtHozygpJDG1YivTxDNST8TaVZ9kO82dMgLdRhXh4b5A7ZYq2636
bA1ks+QK2PD4jJdMBKPI0W4WNESThMrfnlWj2w+2QzXt153V1Ge+LFSb5i3FMD5rhod08M80S1yZ
DSfQnLpEuj5G1Oio+bARKxmeHmNecTRbtRqwUGQ6nhDKaS5tFLZD2cDnd0EHOBp/a1dXOHfYNXmY
n21bxyy4XzcaQfMPD57xDkiF3t0R1tq8393KHVhSjazgLhhiwnYmJ2eCm0F9NI73Gl9hBECLymSn
5mMDEBg03ce78vw4rWN81cN92F63nPNdWdfhzfEbzgoZxGyNHZNrunW2ok1RV2KJGGHYMSxkSRsm
cAXOtKCXrifqlXvTq2VtWQ/6WQDq7SXtPrF2yO6gaUQHDxLrVd+dzGFq7pK34FX0T8Eh1ZXobm/l
RDxnoGb3fsx5aqvolB778kBj8z34QkHnoAzyuTQWaB4h/qxhLC18PZG69V7dOclqbOJjrZigJMpa
r445jS62BuzoTGUv3wAMxWafaCAiwKo0rh854i0S5n44IhuKqlmwfvMajh1ZWZATfSkAbtpQ+IGp
e69UCSk3LjNvN2y+fcO42ns6SouTymmVOV3GV21iLyavV3RSjFeVuqIJvKHsZDRXLzI/3zayBi/w
lZYbL93PdCE3sCX5MfUQPGyrImAwu8wNFgNyX8+rIsC+t6sbisEsC5ZeitCGSynk4oi0HMgPhMiQ
PCLNS2S05C5wsxflCvCyxz8CSkERMd7EdfSNC60nuksQfaKedTwYTyqIQKpnP8w3ldHcxEZwI4c6
7SKwuZskqV6j4bui52NqTXF8eqF0YfJ8wQnVH44YwVOh1XNihTPT3YXJ8BE84xVI7sS+tEVKYNEx
Dp8bpiHP72HBDo9cQvvK7CQuuyoOIfLVtC6Ack1Y/MugQ9ONGtdjgzzIDjR61CvZ5S9kpdKeCde+
Ga+ImzxStRhM9VV7pt99jOrh4CisLgNbr1Ow2y3hz5K2BOw9CDOrZ8kl5JSmC01OlM2pG1aOnrCA
sHu7YPkqgUPhSbU2EWek19q+CygklRePJoqQSuttroN/AwyDLOM4+2i5J8dq0VcIcN50BoS6VcqJ
mZ2SJvyXCzgVO8flIJdlBqLWaDncLeYbQxDdI3trsAnkE6OGjB3Sx8q6B640GsVuCl1qgxmTeCzn
ix9p6Affh9wP1gYzXxruHwMQ9hOX0cNYrtWYLSqtOdt/TZYfVcSlNs8ak+ZwzhHVPUFdq2PPiY+D
HiELWetQYUZ10EU3qTS/pSkAl2x4/ic53p06CsfoA8zuKfxdqGbQgKV8x2tY6I/dqOMZVvS6fq8f
p3yqObCwdAy7KP5wQnSTs7BxP4iujBDAuHygRxGWCocQ8xbUHn/k10urOI4R4upi9ltkziwKXmv8
s9Y7Jv8MxUGLO6fnAT5nYYXWAZfcDgGAjXhD2YLkrnKE1kVZ/y/5XVg/+dvx8ts0UvC3gio3Ev8K
CnU13oEiM4VxZVsGD0gM5C+5mx2Grb6JaDjD1t2fgWJuEBwB0F3DOju6MqDIUAfHPZp9kIk2Wb8m
IWSseqQauWtSJ7M//54/tD4BITbDzRNeicS8/stbq6CCLyv7Ib+1nyKgPrXZ/lUJo1gDTTI39ILE
Cxq1kbBpgrrKAX16g1lgKmTGGgRc4fa9SlZmrDeuh2nh4XodUfDh2eHPmQuFqtRRw6HpHJnfNTGV
JGjdcAqFNP+JQkCrTqsQM8eUeiZ6dBrt7B/xhkzVDUkNNc7Qb4FnkpmaXNRyHWazuIgwgWkAQS6x
fLVJQCOkoXYglD6VfXxNTxfIMBKHGOVDvp//EgV+knVvb6XFIdVbEGzAbg7VzuHn/Co33U1aWmEK
CacnQOkcfwcGtNVrXbXv6xqkhxVdEvz+kDaMBCEcRt4pdmwhSY+UDLTuDCs3PJ3gb/d/I3i4gKLP
jfT6NsaQNszQ+4voZ7uwU/5uzjIejok/h1EO4YNa0AkYnmSxevmF+nIPzvusFvy17kw11gBfK9nF
QYn/MFbbxxQjw4OxH89568WrmF2AZAAGAdp2owev2nNyK/6YvtaeQFCGKsxSsn5WnelpYQtnWfzo
93fTBgCfPdDqRtre3zWR+PPNX1/amQo62+NSvBp1jYj30jpBGh3KIHzmfo0Air7y8Am+FPDFjhKH
LpifkJrRHa0/zLhE/s823SJx2wwOyP0+7lGzBcSVBtgRjqtHXuprBmYAXkOtd+fcfF1hmqYe+m31
CZrRTGS2QCFQ/duJWQL7IypDrsmgOUrG0MaNfy3CndUmFxRyyWCnlNiR+AS+d2CFKmbYHTQ5TiKC
YhBhUMINfbeL0M0BvUgf5oqKlHmXUdQBPh3jc1CVew76jaBhi22qn6Z7Rhs0yssP4LmlsoRmml6Y
f4x02bpeSJ8X7KGrsDRcM8Bf+EQji9HoYGzO3woEQS+I5ZHDPGdHdzxK3HZJgIj6rDxfNn4kr9wV
59WdD0ouKnXcGGRFq4olADNmKvpJ7Z5OpUS7CK6IcXlsse5H9IYJPIcdZAK1e7BlelJodAbEd0Gm
ZLkeqmuZXqSKMVIn6Li48PvcYN0pMm+3KivYX0DK/Yl9oJC9Re/ecgpQBkbaZrzhEu3G0wCk5hiG
xVMNzZpfpuntdcnxnSUSylUPp7CiQtvziEFH9A932fhQmzTU3mSGEitfSUp6cgKykvlwa8XV99Hb
G/KX1UFs9VhDYQYe7ThJw8gqgMOo1/vtpaFVxWAI9cba/e1Zw7gas49Gg29pvbivJUaa3W/X1Z57
QRv85wUVu1hdD6+YZvWb9YyvnEsuyGONYTmxDjcMkMpC/r3LM204ElbYd6rbACDYJ2pkGjWNmDfx
yWIoeftRDioC/xy0+h5l9P+CkS2J+zaIhqj7Yu2O5lVwcenq/cwEP1zNSyQliDTIM9GUQIl47xPh
+VngUUvBFQMXyy30Y1yvw4JDAQ9RRRKFdDfwLzqV/bq/ZSfBDFV+I6vDQ8/wdNJZgqmdM4LilKYa
eOpbVuizIORRrkDB4IVmXLUrp2WgmOTxkRC+uHA2rakqGhXjZtnWr/Qf2m1+J7RZ0paZ3J+EM/un
1rjlQDKqrE9lkcJ5YzVOUWASxt9JXUCfQR976oR1qkjKu3OGH4iay9d97yxG0biCSbGculxP85ma
SfzFxRVEM4cPz4VKfi2B07ohjLy/CLCB/q5mXP/irZXOw9/o+cpF2lcPdUEaX3onhkMgsHF7VV7e
GHOgHJ+RqhgXQpQhS3T0lzQUgZZ8MGVfbOplpJYPwZ0TYTFOG/JD12gVGY58piLI9KNGV5rAbA07
x4/tk5kXinEfDIDpcnETo7w1DbCU+ktJ2NVtg4WAlTUWCxNstOevVOLlFdWTi6W/ULvKIwF0iPRX
GFVudgjsgdzM0Y6BIy8FtaDaWoqz86h16vtS3FCFMg4WZkChkS7d7R88lV6PoOMTGEmpIwNsWuFO
1dnoVdBf5ygb+Tp9Ykxe2WzQIH7wQg+kIweqL0DOjs3cT0e5cdMLabxNj6+H0/GeHRuD6FbTna5T
Fnvrcg9Joga9wi0ZRX37lV8JdfPzC6En1oYUvbY/7RZKiY/yPAggWMb5SDvSR8epPI2QvmrFkngb
eK7DYiYuEqOuER0f97/xOxtZvjE7dv/RpCtGGlmvnoxBeAC/kgWef/paObXvkKGkfsj4TyNtmNAc
JET8BQCm1FdtiJ53Z9mtxbkrMbDbA+ED3LyxqUMztZX47LrPoGnZtXc9x8n9S5Ap0Q88p5+5ID6t
6CP64ElDlhKnn8b0weXVufDZU7ghqLwmyLuSrveFl6uk4nSuQ2YM/IGnvXPoQ6F8UPsddlBar1fj
SrUU8/5m0OazFlkzb/KiG1BhYrbDCZGT7A91sSUWtu+VPqcUUtRfzKaV5EKxrkL9Tqk/3o2IAOVa
2/sJCiGd98mVPqiy1thTtHhLhqikWz8OgnV9IK6yNvQnk6bRs9qdTXh/BEhTHgjOqt5rn6/PZbbg
sPPatiS0jTt+6UV9KMjrHJRpXNeQqSj59/kD0GQnhMYGWUYJy7twGW09GUTahJvn2oMUQFhVPe0M
JJE0WlMYoBMUKJ5qdkCkPYLotnds3VhPtRCDgBETAwCSHxWhQ+wkHxiIBjXCGvD6Vm5+fkPm09Y2
82fHG09GGQG0Wlmh5Va0QhqhQk0LyCdm58g6A6KpfwJITk5f2LCPF1TToHtagFb/CAkwJH69sANV
ghnRHxKjL1qweXqzFX7eV5Pw/oO4FfmoW8bBUApZ7vnE1Ix8ii0Z38Ss8XJfHI4dQxLDKBZ+hxsl
2uKr431QQAmUeWn9ywJmuENCuX+usSFnmrK7IkJBpxxerMB9hL1f1sD2EilRhsepula6YSjAxe64
9XCE89IWYjvrmsTIYdTEpKEQnr5ij2whibI6sc1XZ2m5Indb4qof1YRFZvBMB7NK4+ndfZ07qh+K
fun0p9vbrnsdsoZbCo8lo6sKjmFqCs84KhX2KD2KcEbQ7rG+rBD1kbWKTzFmY81BJqosRTjz6W+1
KyVPoBllSzDqh5XYuFJtCWEyqRjJPL3HF6ishq2jmevjUFVZ8Uo4gEgFpMBlil80k5ke/qlfhGHj
OhjTUHBtFj0yEMYMants5dbfNg9uS73WIU8aajGasJxHzJ+5wsaTPXIcywZSSEgAkblgy+WSE29R
gnPiR4F94BFKCFOdrYZ2EEF/N1r2EtJ+Slr0/WvDz2eNRWMcujoNbSy7MiZqvSU6pB2c+rdGVBQO
+c6V1BjcoyXjt/tmemWN7t2EWY0RrQxi9FKqpOfGWumPg7dZRWAF2o4dhC6buVUPzAJF7x6XJklk
ch54suTjEp7KVt1t9kPGmH0M640L/hAiFnvZ7c9pIQymCjo7CIJzD8rhsBFFok5KNwUCCWfZM/40
4P3JFrbrDdsl+Yzo15qMGf6Tr7aYFB84TDzTQAzM+TpBSGG2h/hEEXtmMVjZgLkQM8GqsRMnh+OL
Pb3Nzw5MhYhYEZI1on2VXHhQEtJBBQWORo7UT2yTUF9UnRXFXiOlOqn83URWlGSSLy3fFzz89CM5
IcERe8PpR6hqdCHIrWqGPA19/xpPEyZmxs5Q9FhjxqG3AEVRL2jxxX/yRqtU8IUTDtavEjxkETcT
ZpFQSJTAvP558deVMWDZiVM2q4U6DT4HIXw0+tCc+zJJSJguUfBdRiRdpbSUNABmFWM83+gdbjkz
il39NYtFbWvpjUsJo/Ow5uljr2nDR9p+5A0/472kAcRH5HImpwYEPqwsqOR3FrwyWFJIuakKi+GY
dbNFm/jAX0t5uSVAdAVLGXUO9QGBow1kyuh5kdCE7pyWtao8T1Wl8SA7C2/CdMTa6bRYCpZBwBfR
HKFGPmpV58xrHCUY6UdBi267xfRrmIJVkomy0HcmH9ULV/Y2V2R9t8GIZTGBgJctz8pxhwu6bl+g
bbsaSZIAVzdK03FNmMpphwlxodyTcBGN186ztSVWy/s2bYAbEE1Kfdj7nzvCr/pFNI93pGxZuGZz
pGGd8poFtO9l1pXHxXqqsRycNf2QfKOLLNITTI6SpYr/cNL/G7NCgoL4YufRfBKvaLaSyW3xc6wy
zLFjMeWcqVMjmpgnIYJoZUCWTYIUSlIpl79sJ0NdvbJDdGWdnh2Ayjx8f7IhSzbJpn5xd+Bo56w6
qlyVv32FXQdK8AOyjIib4T3uUI1l066RjEPHuQcSaR0/ZL/OtwCzNzhGeAA7TqTTo4gvd1rp/SvN
ESVfw9UBm2yYL75XEQ2oRQVf1B1259kW+gYY5BhGL7QaWljW8z3BBKgFaHMvWJJmhYjjpAPg/xL/
0cc01qRFUKYZ0dzglLHskbHU5ySuJime+yJ+N9KUXOkI8+vcR4h8ltrLD3dfmRRRVjJiUhP+8suv
/HZVhKGyE2fPx7fzBm3HcW2fmMwqxpzXFBodF07PbgfEwAcMOc1S1aS8rpavZTMQbLZJi/WjQZpU
MWrQSJxitvabzfjpIU2TpzGY6MWUmgDJTM+9S2knpk+pecVW8yRqDbpl96VAx+Btl+HUL+mTLqJb
6jIYTHkAcvkQXx+3zynSmmdQNIwoX+zg50ByigwkE123XRfQTQ78VrTng6WG2hwhVKG7/vVRc/Yi
UApgObcNyPzqADf0FZL1qNIPrSR6TD1DIad+yrsf3aFsugXk/bUgPxbTVkB6vykjCrcCPu3T5nzj
ZkDdCr7PHk+2VG2CWHxbcWsPn91xRkL43Pi/MNJ03kSPYoobynNRHtwvw7JOz1SCOuWcJPer6vj3
cUPg8erh8oRd1xmbbXYa/o+KDPbcb7E0RgaSXHbSegLgQu1qyGJ0j/Ve3NVrSJOZsYM9u/NBCJdK
u9VN0EN7lBNt3og1iCeCG3nZTklxd3CUkJ741xgYF0tjyrMwaX3DytYUxDmIFikwn5wU42q0/CB5
Je8DsuKlf/cSVvV+rf6WsDt8/qY8vX8bURzAGZiXjla1c4D+PClT19OrJFxQNOmsuT3zgWnHah6b
OGgKYLgo80hkDr90a/c/+rUnVZwJaqChyXCWE3AjjyOIVVcE7oXOy9BGOwwXdmt4VmjbeN+4Rrqj
APuDL7MIh7w2ehJoZILPrpAL2pYX7vlsQ9elsFSLaYdFNexNEn7yXZF6wKax+AqoqG0k3SfeHGPF
aWnpYBqIp5Q37UsNI6mQ+Cc3ky6LnELkUs8i8NNQFr5zJPYDjpyldArW6/3nzfLqdxfbKHqp9sKP
yAwrQShTJScL4wNybZCmO6p19/9ZG83XYzbq/duW8Fe8UykwGRfQiD/Whh+xbg2bd0Uli7DnFnQR
nztcNtHutGJljhm//s55bbzM6EL+eSOIcyyWf94mfHwIhbUN05IFKmQSHVFANy0DcaDQkmn+xAXo
tqeIxRV/XEIERCuF9rxrLx+9uf8wLz7ot/5gvWZzOo3tUxw1BYC5ekZSJdep54v8QJ9s96Xg25Sy
461UgUT8CVEQqiJboSWbsvM99u9AIWz0zwsjPxwaBPHnv36+xsr3MPK5+RF5F6gcMcdQhxeN5qMY
+e+mKdviStSa4BpNAWPRTuY2pqlkkYXIZvxp+IkOIZYifx7j4ZKx3b5uPl75gdmCJZyMis/Y4S96
T48j75fux8uBVn+9hfkuG9f0O00XbY2k4xHq1l68u7x+Uvd9qS+FEa4/zK5R/+cHLZB7RHfRQl5h
ZzL89uNAFNWsur+SfVnxj0zdRZm6QIT4NI9oAVUEKfPZkCyOJ9x5ELXv89Mo79SNNxvS696fi+/O
tTPxRz131nlu2RcH2pVyly305jIDL1QUGbyaqPlEZginF2SOW7xbIxfOF2YyzP4Lwd8OhT0K6KF4
z+t/A9UODltymsfv7IF5eZaAZHAcFbBDvaEc35ktQ1xeqpLGp0CLwJk+pSlI0lV/d26jmKVqIn9n
xSvc7I+YMjGwOIXV6jJrIvHt392cEkwh+p3pFDiG4jhKc+48dUSeRML59EOK/DM9gxxazumCA6Pe
l0k8aCUnXlp64TrboLUMft5Vc13BOaVd9jC9GHgxlsHKaazhaFXZtlslTm9sO8THE8kSV58z/jWC
gUZTTdrMZsNOdMoOWMtSRvbQqMbSAp5MNSQ45BGI+eOJ8qMx7Z0AidvtW4DNGNrWegAjZ6bNh9km
2DGhKfG38s0MIR1vQf7vKmx6Q7xSVueHhiZjPeFnbYe++cnVdQhc+zbspDSbE24oCcwC+YkqETaw
NfOu0pe2LI1qDUGjgD+AukujwzbWxiuKadzFWELY/Gq8J6W1Wjd4lYDLPCs+foxGfYs7cmcJR4dt
L/691RUB24Zpwb4uF9r5cj/5+mwzBBgFPH5Y+avy5m3XRgk3+JUB51nJqVZr3a+Va6PpDO1CPI2b
c2pnwphUmuRCehHTv0avNfsYoE3uDz7dc11mOOe4t0b7iWAiuF81t6AXYY1EZF5G/UcezOuyDwih
dkF8XzK+wfZPBb4xwiMRqJCnTEkY/mD9VPED74RvqqO5gu/Mq330Cujm9hGad3WEPTbh1IuX0fRM
XwBd9gj5moM2JidN45vGehYgqHXCONBH3M0N1XalwRIoiZ8jw1GOA3z+uEk6Xevt1tH/Kp9MsSha
nE2VC2r2fPG74OjBdigTCLEi+uECz4uXY9WIJCkvIFSPIMursXAR7IQSahpiCpSiMphJagGuDKWd
ugxm1bB3ORQTAaEZRZpYG2YEAWv/BrtE7uCLSHA0KwNOAq7MIJXWVBbBTv/Z4FET1vMkPM4TPhVB
GbH3Wsq6756FcK5WqLPCcOX6KzTyJSfeiIaC/hLLghMeptE9hOXkbnd0gnAw3JuyYb6YxQSwCRh/
J1kz27G9nZacLICXhjK1EWolCluVsCU2MQUPMaMB+jRYKI4iIHPiJhXgjQVtdLLRg9EZYLrR6ITu
NH8NcbIdmUVBuEcTegnRirF/mr1DnZJQy81KpwFqJ67EZst88V4EJ08Ys5rKAxcMpPV10IePGwzJ
rLtDmkBPfayfmsBM/cMhndZ3lWvGFFqgF1UbDAEg0kh1/pb0+owqn/4cj6OMaFvy68VrymBfPqBT
dU/fFGg/2lrxIvZn2X1WWWmLTBBSATEb23K+570uhqeHRr6lwo/wTrkTjHOQr+7JranwMaLOTXwV
R+c4vWw8lXvfE9XABs5b2dWp6HSVugPNwYgH8M/pjOdfCQr7+1SkdtfNHmW7bTrcxX+hP59hWuC1
P1Z7TdPFzFHN99ZP/0fcHumHL2p68WbnRreSSMqGG3rihPZ3qhWZYnDJSJF9mZu+DY3HzDSiuH4Z
nk14uneOUW3XLgMy44BM9fuHQM0XVm7bVXQTCm6G1yMP8+oeEHvJqKoP2cf+7BkWAreIHAUzy/IT
7WthZSketStTDPz4BInmflyTGVeDdnAMWPiwbQlo4Q2puvL1eXIQL+yUcBRZKWTGbEJnIn9AVhe0
P3B/RhDXdRh3gF8TxG2CFNcZ5xwhbHdBaPwCONrmFdPFqkvwVNTiAEpaOIUlfutVm9+niy9KQ1Ha
9eF+g1TjvPgwHehRS4S2e5D0WWa+cMTPXNazpYdFPDk0B5MwhPh2v0Q7b+7AIOVL5hQmC4JmnJlO
EFd3O+UxIWI/pzLMVLMrPkAAE755rOIdFW7rVEM6t+CZFQg+/ssXtnTWkAxlpOyQ59p3KtHF+6bE
mYNhi7ymYVHF91hXsM45TkOwkT7LF4NMbOnOLhFAos83S6T0RIyT29paLeuIPqVFZycrwNCiCP8H
3WOX9VDqzUOu5Y7jDSVJzUtGmC3eEsgRJvIzYxy2DRL7kYbucQP/Q81yxMgGHkyp/PJcALMRjI0g
19I56ylKN1+ZaWgUcej0ETixXZlkv61qZW35axtSwYw2pbhs9erE5xidCaa70kfDMsbm/+FQ46qy
lKZfnagnaWRhcLE6v/NFFMXBReK7JinUK5w4/h9HRQ6tzKfRXZOEOsEV+qpAs/8B9xje6qZ72leI
FpDiVFZ27qYcoMLm8D+ZGj5iNDoVH24MFYSrG96S8dYmLsnSWAD6vd2deqfNaqupxKj9vFQsu2RU
u2NW4bFMXLxRTzyjUcjYAlJuMGsgo8KU24IRLHX66JQ6uCR6G/mIcZ+Me5p5pK4UZaLZGcYtSdiU
buVYnz6mbMB/ZfJHi6+n+KFtSw1fUgbG8Y0uYWAQOqTZD7tR3Q0467S/4jpCJt/vgOs4FY6hocYg
M5jgO9N85MyZfM3sUlROll5nSrzfyKS4PFZ3+b7cKksB938DQLMuPNxee49hIfhQYaZ/KtjYaJRu
74BGqhWjBkYu3uEIyFc+n+2NRPW3Xj7bkQRh2T6ZJzqxvY9FlylHgkBXM3xAPW5Xbu1q4nT1ZAlF
KLMSlfOIigsVtlmhDhVP+bh/IpEK8kFn1su+sp3bYe0MxH1STUkLmIhdKdwAAl9Pzcj7t9dsThNU
I44Y6IZNZirmvahb5fZuiKSg611WIvvaaNbR6PFcoFY1uE5f+WzK2kak4CMlPIRd6cumNQSg1f1m
dAMx0VY/eg1tuaB8oGL7vnAYk2m/29SIQCMoI2WyIoo0fR/Xdlwtlrxyyx/SU0FpmEpxBqNaJ7VO
+xlWxYVHpRREBrEfN3KPO6Ijmv5NZkJ1gDnc1yEpQMuaq5RcN01MI9mCtZOs+oE4NKN+sFWauxJ5
XBLM65v0kR9s9y4T3ln6VQhK1UXmu1eJPAJNIBTM8z0MOn7J5OEc4hTYIInFjyiMfWQXYnDIjGLj
aOIVKE7HaJHqoe2ySGEqjylU+2w61gfIssoxE7CTyXKEiPBrc7vQc9oO9IlJAhZcbxuGmR2DxKxg
dCXZ7AuQjogFL55goAIqfEFwmrsFisowImz91A19HgXuGHw5jT7DI8l8cEwUTjWte28aIDfLyGcB
KvAbYqbdZHpuvNKqCB6dxXsQAh+9ZzXHcehxXvGTBad7rg4Jd1VEdsHJSyLgY/dZk6TTrwmEFYcU
XKCsiDF7GdksSYFNeY00v2/ZQj1tGQwAycEmI6a2zYQgcdBNE5/ZZ9T5I9HwkLVxSukYlz+UfPmR
hwRXmPop4WVig8DRbYrhdUIJCNbtiP+lbh8g23xrVXaNowbDIBhGeGlUcO7pG2Uj9cXustdzhTl5
oh8QaAVBdOKjgyg5gNK43Z/bZclAFyHOuBm5BwOWUR7QGcMhnlUgzimKSeYh4DAkca2y0yj4PmT/
Vhf90a1i/JI1V1Op0mKC3rd5hjIloxHxtmvH6I2BscT26C+F7Wg6OvCC3sHP948G0JYFAtd5WVHh
i9gmU2VsFtCTbMXu39aYCCZs8IQxjq2JoItQ7Ul5tw9vuvR8TksTuLMnj3/KlwuGy5Ak5CjZjiW/
Wd5H175y9PZWEodCUsWP8PG/c5u2K/OeU2Tq9ZyCVHBWkp7KqigHNhObr1DfuZf1pPjMPFmFQd+3
NQHd/yGtIDyuFhuUU4Ac8w24nxQ3XMILqtc70z7pw+bARjuyNYABdBI9taqmmDFczZllXCk8Tdsn
XSh40/jEjj4BYXLFITJCTkKgD/UhhpFo2A9UB5BdwttIFhinXZMHutBxRfD9W6vo2/bOcG2S+95Y
/P5gu21ADgOB+m4cpBB2lCfz4nbxoAgytu76RAZVrgZGX1gRpP3q+T3MDAHBIyxBN08ES38Bi4GI
QKkhK5duTkVJY7FdugEzyFjhvRtLjrDbOZsFdjlaYv43Jcz+ESiPEziy0ES8TZ+ySzscOm3EXPdz
9wNHW7RNYHI2bDNMEbmAtBaNYZWJ6cV2P/UMyCNv8bSeUtDABEStMH1vho4Tv20IeGC/SLy+eH6S
zskU8eRwvZcEZuB4qgAIXUEoXgABvWlcrB5hcCWqR2Tt+v4OF1V1mDhu57RP9qQJNX6M++jHZRU7
UvmWHaCmbVMdEKaFL+Zqgy0UiUCcR/NANekuWCvBe1Aa2Eg+xlakeC7RQn+H5rI4yjUgHtfy63am
CKZd5woffuvtQhSoOLWDHxsyFoFDHDElk5UVrNZfOMKPHiTDai50fkc2rnslFqf9IamJCyGoXN5K
pgjsP+QCPGzsnGGzXKkNFdpZ2CB+7kFJWIF7K3H/b6AeZX3uTfcnJQRSwDW1EjfgeW8h5UwK/J8X
hP0UGQSluhbIzyMTSHwWREnafLMnqDHfYRfrS5/zyDL5k6CpXGUCcu03PXIjBRL2l78fBkFXiWCX
VFkvalKFYQM6VuvacZkRCZ6YELJvuDnoannL7iL6SBmJSm+h1GbKe8MKhsLC9uW14T03WADh2+CP
dV9jAIsjRVfAqx3yJZXIcZXJqttzgt8eTeXx6zSlXyAHnoBkdG+MoXPPjp+7nqTiNd0MfqHNnnP1
cCK9O00m4ya8TOfp17T/df6QVxfX5i7WnYvxuVdjZ13u95ovj6/e4msb5viH/DFUXxlgAhFjFndo
k5etIzE6/Pr7TmOQVoc/3ra1Hbgjh73fb+EptS+ey/4sW5eyzHYVyQ7Y2LwAd12R3vDfPRYvqnmf
u+1ZPsITVRENxwDqW72ixmPMLxXbXbV/VjGXUbR6plPifIbtYqeDqFLZXAg86//gh1DmPpI1G23P
4rjJuC8q6bQF4j/A7fk3O+G7aQOqL4NfXJkMhIw/y9APc85lzGfcwoqR1hVqfAjeoUk9Ocejd+6T
vLJk+cFyRMhafD1pA0MXu/cFW6ir2w67lBc/BdQsWSjU/2JHSC8meQiL1qxMv+2jnrL7/S8OXs29
HblKDlJryiIG2YEHwqF6yLcg/OD1zKi8WXuuppzAEr0pyybZLUh0HV7MH6GNLJVlbaicJv2gi+Sg
VXFWGFrYPdE/3HsfybFxsC9pYMBCKm2Uj6nhGNwfHrlZ+fVrL9R03uqDocWx6qq2igg0UMUhiSC6
b9k8xzHtLWLFrORwrJUb0TDK87UvVPbmkS979a6c3WunLVO7AjBCe+0IoC1d2bOftIAGe8eKcHNA
gW+0T+UDKXKFoyj+wbTNxG3rxuhHnQLwUWFXUuHmT6L4BiWiHMgSagpEJTkTmGCsE1J4GnOoY2hV
fee4hdiVVMX4yHdaHme4r858L5c5ltlLUnUCRSy4lNSxqmw4Ffx/0C2/LAJX7YGBSGEKDSUzlCOY
Cz4ppB+Cx+9hrtPfooZxgvF6FEBiFIdoM42u4FNlT+ZnNXzaKIREML88UZgxuFUwUbaeS0Ujl/Ho
YQ6/Tx7VkDJk5CLDE5YtJkWhawK9b8ee/MNzgdNTygXxAMxZhXcISoe9fqaZ+pp9VrqZGZLVABbL
xC8VpYtsF6slj+gpIKjrWsqt6c9qZGNThRkhHhyooelGcJtLxAKPerNqt26SZj8Q9yXGl6GVEV+y
jETF9TTurtry5kp6jh+ZrWy8uRcFUXpXDh8kD+luLOvOb4kdB1U3xq+KTGSHBuqwMKUQoyv9eeVe
BhBNfdSLG26L+KE6z2wR6Cuw6tKqc9qNXOV976pTa0etNzY3kxEGGP/g3spr0fVnKUl8B18xRxyP
XXI5D/LQBu9j8K/FuWbZvGdZDadKy2OmbU18IzrzH0+mkYc6jdQggIHg7KT0ikp/w6N3AhFqjDen
8pcTeGjLPT4TcrPoMv5LCamcToFmHTUrYNzbfUFP9VOceEFQHy3Z2coFyhTVaLVvU5mYp8jzdQ7i
gum/5OG0aB8dkS+Dti8kG7ucOKbDrKeYH+4doL0MIbvU3cCKwNWClhD8b9X8KyV11ay5IyQkGDo8
HoUQ8w987irDBE0D17rBtWkivsAURLZqkCO5Z2vI5VtYu4XLTZKdu4MZtgWnkOzM2HF6JGnLh6pw
yl9t/HwRtE07nswPvsY4q+x7J4EY6/0h4HdybGIDzh3ZfqO0MxMLgIUc0ECwMEB4BE/IzUAH1fZK
7ZcNtiXn7WZvnvocdi9Altc7GI1vAmPVZw1n2yZrtCwZvlOmFfXTxMujG7LDMlOPcozgQqi0QbM2
bZCfi9XjlkmHIrjND5YtqHk3lK7pzNSWBLo95C6PN+927AIEDv8bW+5t1sUxDS8pceX3mVg/rI6j
Yfpuhv0viLRs7itG9se6iHv+IaSs+03M5QdjDqWX1+e06MM3tf+BqKukYpFroJ9vflaZhZlv5f8r
IXlE645HBdlRmJ1bRlXcZYqo/kXY82OXbDbEo+ayd6nn5XgbpekwCauv4xddELPS0V2e4ZWQB66F
ctwMgOqVMepyClMaM8oO8sWChhqhgt1GGPwg26zgT/MRS+UcjEDNB57nRsw3qeYvVEOiX/T33P+P
tZR0xnO4nwlHQ81x5/Xx0IREjnfvo1PfMU9ila4NZEeSmUILO17whSRtUx8ZlFIt+ouZHNogcj60
NzcGHVDQVmSKI0YMfNsoVeg8I9ZBqdiAVY6XFetWc9nCvVwt3aGPma9cnZKWWFsM0CJJCEqdHVbk
sbsg/a82toyejT/tD05xj5RFu20eGima97mYyawsJKQtmDk+yhvB3r6C0tNgzeo8G1Jq0tn0mUIK
2MZd1PFtGyk9fk6iRTVILEtSVgvBMJsCe+s5So85Wm3FbQ/+OwqU64Rv7jxBP3UPR1MW3n+YdDy5
49iOgp9xnJKMTWFtBR4WDxVdIaxxmoUGbZPKedZRN+T7qJwmYMD9V4bLvsBDN9jWrds5pDQbsOTM
IZ09hl0BDb8QHwSyBJimXAR2LISl5LM0j+Tm4n9eCAFhIxJRP8B5GG6uLfCBpRqO56M/SqLnrLY8
oe2vxmwJdRPvuBoWUH2YcBSkNmwYRgBX6Q/UoVtNKOk0InLdNAnGQmjEgwGFphCz2Frz/DmCnIFz
udub4Dx0L6wKRoA+plBL+VvXurkCKlD7s4RdKpyPgMq/X632DalW+SLcb2i17MIx50pdE9AQN6PC
zE2e0XZGn5j8uZ7g7aXEocTkqN5lTq49DIzaMyUHo7yt2nWp0mfxVj5M/OrK3SX24ZEI+l1QnkLG
F/n5xCMj4WScTQAAHkVOe+0iyl8g/Z/SfQZKffWGNSnJmCGbeY9IhOjqW3BODYDc2VbOBxu5halX
4VSU8GUDMM0x10+KezfEN2GUl1HgFINpSbTjVqWfriaWFdaw5RPT+qpEpTOw3O1kUn4vJe+4R0LI
tojUqs5XyDXO1p4CSJqnJivahXRiLXaKeCQuE67qfAlTj7n13nD0ZU7OR3QiYWwBCh/qbDO+fo8t
F8pVITjS3wJh8Tujqza+OQN5Pz5yQsrCgeUUrBaeueUkHHPSt4zdN8PE1jRXzI5UpKsIUIrjppBb
BxHkAyShIZ/scalONg+kOK9T6kO0bG704yYNFcgCo14ipydEJBLBs9EnmzsErJUjlMqSKqNmcf1M
U69s+mk9HILUgTzkhPXmSpRFEQX6Ql7+lN0QQ7xWAgnP2ulhJzdPtROHJ0miZS6CLZ9J2Mhrj3XO
tzdp307qW58HRSrL9FpdmqVVMjquyaOpwk6dO6Md3G1LUmnWTm2y1uIORVE3b88PQ7OGwZpucqQF
6eRSGzlEwjfCCBGuPYaF769vTEVOE7jBiQ3HJC035vcWNvh1/LMIW20ZQvVjW5jNZNTqyi+t7nWY
exqVxWvX2/U3WS6VEJAmr5iy9DEF7mC6bHiHANuyRrgCOVehyuELZqX6CcWa3prnBrps6lMFvt6e
cc0U3qbRc5BIQ6NMDsfl+6r9NaHGb5bp/FAMZ0tDKF5gu53sPh+I78bQiMw4GHSQSyEY+4upB6sE
T9HwxNLktGxNe/zvld95mEnu4PjGUEfXZnDdfnuhyjV7sNYoY9BTVSPQ3Fn1/7yb9ysiCYbJskcT
1QGpDzAftiMul0N4g20E9I7JvTd2T2GSeCsUg+yCwDJuV8a2iU4cCC1VeIqQCLVON/+I4hk9/FJv
hJHcQloL+fRkysUJt6VSKYArQj5i/+bRyhNm297EKfNcwULsmLWSwhJfwDobdgd4wAcYysTt+ezC
u1h4dWmkCoPzAHU+Oh2eqUIVtR8NMXTWKJD3I5slRwZIMtgK4XpBPcoq/sH5uHH77IC7Pcmrm2QK
DjhXtwonaXEuPJ1barthXd+x0fntl5+0HxbU63t52dyoxajN4tWgmgGyrpJpSZiGrWl1p3kh67y3
Ex6cgKX3qQb8Nm8WVNNQ3KyqIkJz6RjVE0gY+Mu/EPePMVx0YghHgIT4Dztn+803b+OUibzj8Q5j
0GtPXvLzSCxvgVeU8dHCOKz9+seXc3xM4tNVIOSfVxJzWYHfS1bOuvv3W493Oy7wn4KGUkGEe1/v
xTWnSvrZ5YAs2MOXqSP69Sl2KcF3G3htMYHSmyOlqjhc5pisutFWKtG49ZoMBTLk65Frh/KgQY9X
rokQzvsNUDJoUJDVFgbyhDVbedsXqNuahnZ+PvgDuC/kMvXkTaBJSyZR4S6G06vT0pY6VhgDj1xg
AehYNjFOzx8P0Ql+5griP+ZvApYOgQkwd0cxN7eiRItwbGqQ78JCVE/e/3HQAy23ynmrFt0mWXop
7mKruQp2Nc1wqgMVs4xVy18WDpGREv46GqxyB1G2FPnF8w51YMrhGi8+54t+Mc461XGZr3Uyrmh1
AFtrZBr8K3duYQ9pEj1mAvgEWT8owcbdLhgbAD6l3dQcib60GJh8KEXSBXpKfLwILTmanCVVwHXc
VIDsCveZ7l95kbwY+Xg1Hs/smfOJCY875KrHHJQdHl6aAhd42DkdlcY2ZlkNKLKx3c9J9SetrASH
8WZpTjfti+s61DiuyADPRP4MWnASrv4y4azQ2gOZvBvOLaSp0tjbk6xqHYIbCGL+P13gue4xCtJE
wePfCuZiq4Ef/0lYWDpd7IgouxwUC2IFOuSMpnCRwbnuj0hywbkM6ltXrYuXy0RoDFuYQ4kQ78Hq
agRDgf/n2zR88Q3xkab/n7lNRf39REmC3aAND+G8+aKSx6za3FEcCbiTg6IOGoYTDiznFRAjJgEB
Il8YIySipXxHxDB4fxtZLfSzHo714N65jqDsIyJuumEjkct3q/ppiaElnGP0YcQKHeiS5uWa0Tum
wbohORbgNJ4iDAwMz24Gksxw95qQ2vf+/yh2sSFuSE05QUQ4R9si3QRId1tZcVV/gH6h2TU5ycux
Q7o2IU557w8v2vYUQwKTpNkuwBeQSGYKL/J/vJTFkbd7f7zmL/k303S/hQGqayFljz1zgvmM/mL+
LJjFRp+E3RUgKuchTXNk5VfWGRNete0/txwDbzDgu2BUG3L1EboTFkrE8Ag6USX3Hg3sMAz0KXIc
e0oF3EwdrSLR5Gkiwv0ulfONE4nvPUohq2AVvz+BkTqOqeHGaKlfS1+RLftiekzkYsI/5o70XN6y
fYeQ4vjLkEOOMfJF4p7ytg84ZsOoo8YMoZOT4Bj4nRmtq0OCP4pfcW/jDKxkA35/P3CQ6gr+IBwX
KFySgKrrg6POh8teMNK78tch1tEiJvKviu1rEm6m1i25bTVzX1ZlHRrhH9WrIKVMzAXajy0YIp7B
/s6p/JoJyb/YzyaCAiNyHX41JRJUuLQKmEqQk1K7J2Fo0CDpZNfiusD6UJOj0pYhMd1+bUdr3V4Y
IS9uyR2JQO+GtFXdWQY6MTEyMbRpbAQvAC88UVT71ZyxFNZW9YkBRcAgjAfGQhoMhIJGrE72Ji3S
evrdVHxnpQfKT37nOkhPZlIVZeKyjQnx7JZ+qnG31rDr5Cf045BNIDPRKtD68q1U2HQ3rjKvlNHm
z+jyk+Eq7Rc5La8nQGWhtgvUG9HOMnyo2iyWG9rFd/+5NoHeGMXmWKDSdKupwyZSgZ2au6ZnXaDr
hBxl9aRR98pxltLKRNkJ84133AjyqfRbCXIpJYZZoZN8d8J2jJJBHnuoDToaJluL7u7m+Rg4yNy3
HjDdCLt/N8pZlGWHOLWlYOoG0CHMXYxYnP95RA5VYTrkKvqJvvg7PBHSwhXjAVBwP7w97h2gvUec
sOtzKdIGL9tLuCVarBiH3BCjpIjCKTdM5Te/4EAEj7YMFt9gip2pxRyVkU5VzIwdDa1bHaSUgOb+
NZRUAfZvA0+z4BtN8+VGUJa4oslG1CekJHQ7LSasiShxSpLwNDlKIKIOTgwkSenC3TkIVTB1RZVU
dNhY7Gf74Palm0G8b0lO7Sw8BRltSuXq6iasC8TUVBmhyDM7hHykK1lhVo8JsF0N/c+JvzAvBhUY
ClwCRUuaGVRPtZW/+SmZK5I3bG96sQQS+J+CA5oKT6Y+LX/g5C+n9uwMuLcJZ21o76yNp0ZweqnW
7R7+sYIVxUjmEAIvHfMlBrLzFRQdrLLqKYvxGIcCab0kdLwsdLq7sj4xySfvGq2JVTub4IL0magL
mui6Fh1zHjC9eIJFN/xFKL+bRZVQKlKvFId9d0S/avS0IEVr7UtCP/AB4n4OZb0rgSj3ypkhNA9k
WyhvpWGi5TyP1wr8/T3YDwksWaYOSTv09cRW2FsZ13aPYVmXmHwPh5G9N2VfafscZdNaJpU/4cMZ
hUO4T3jmW3WqGy2vSgVl3ywW3XuJ8nICj6ouUWd3ZSj8odZcaJrXYH2ZVaPrYJ+AULmRaiqKteeR
tbZD4uWAFUPR/C+wL/CrYGFzKooBKL951WEzD9bYrJGruwSU82Ex7wmaVIg4017gUMDp2Nawijzu
402mMqJBd76VqKAk3TCeQmbWU7MguTxRwjjv/RRgpesKoBOhf/w86q4NWhA9NaPr/+fFa3OjEchc
yi4Tt6oalqMy3IU1idkN8Oxw9w7UP+jumGfFolJZ4wgmpvs+KQFiFbAscbRHPk0pYP6LRl3w8Kpz
RlaSzMCFj00jvLzA5zEzsXdepklHe/bno/7Kuqggh0gItsCYqPD+LdRO0kbjfaGdF/CsJ6Eiwr8i
M01TNRk63w6FqXdGFDgT0bfIpx85Tj8aRHmRrlu8wxrkOzIxbC0fsh1upy4VlGHtq/U5qypd0TjV
y20hI5NgKtn8V0yLGaoLiBD40wsWIp4m/ZUyc89vdoQ3qCIpCMTl4RSR6iqzAjUXhodY/i3l4XWE
7bBBTldDjn/7FXX7nnBd7r/mNvhlK7F/ZwrMPww5npptpwJ+DPt5IxBujWFEHiRgp3cDhf+r7N/a
T8ZD+mEPclBKDGm0EZOkp2tR8xhm6AFfefe259iu9lGqYONbvcemcp5nXcG1OEY4J6rn8YOM2iWt
iFs5XWgT1T1a0wo2zRgErAYRgKsIcFpKYGs46FXmVt6MT0R4xiF3BYszSBQyl72jJCNKlcaY4sU4
Ih/JckKxIoucFMCDLM2BKrV1ATco4b2MSsQVLGrYWEf6qD3c+lWp5vdMKKMnbbyCELmtgugPB1m8
a1jkkSkqSISIXhIGtWW8gPw9/yNKlJvCFtQWiK6gVSVmmzyj8tsU2+GDXAxAWqbcOdwAzeTr62hT
sSZjBe8ZGBIdnsQio4CRfmudrVfTAKG5mE3Pk9lxGvEd81rVLEm7x9mgdqv4dg5DYSVIT+fn5tTS
ISDMIhTSXlmNvj7IbcZVvmuf+4YfwON4n1UoxdQBBwuJGq64MTRmmlegO1ey5LJIN4ppeFyydFjs
lYFW+cl+mwD+nhVbF72mgxhCE6mIopiL9m3Jc5kMbCAL0Wnwd05uhwKzmaUmYV1gtDF+vmQy9bse
U+kRUjjCO9JGiXTAxhNrav0JWYaE0wHELpoSUSalAEDqI8aiBC1tg/X35/zMQkwTMlLT9DtzydsP
2N3ylUHP0hBjZizi0gi8lwIvaoSVyAD0+b8V7y1EYBvwOwzDbjBXIbANDOmberxahNQ/Smo8PYZ8
JyqBFBzfvYCGexWtprKZaR8UNYPDimmenbAT3dS6FOeM1y+wRXf88fOtouK4DaAzf20Yem7ITPXD
RkAnPo4TkTfMEgGLJxsKqaIuTrK2UNgybI3XtkE+Cqd0jFVW3V5gZcOf/KJyf0MbnpWYwk6Gr92q
w2T48SVZolfwQajyCUIhlw4yHha9zoOw7SpQEhbBN5XoA0SPDZJ9g100BneIGfq6QpokST+l9+9O
5q85HvopXkB6LgfpFPq/n4NIek74hIfDIPV5/wPzQPUuU6S6rag8eq+FOx4vYnEBqodfE5FdAuKb
lvx7NILRZkD3cY3mqPQKG6171OWS46qTtMEz42tAJFmLd1GOsF47kEg5qjPllvNjgHBq+F0b6tQq
l9872b7/q1HZP5u+XCQQttYzh8VoJ8sDVYqZip8ML2LDLkxD+yFSfGkqdX13u29uygskePrzjOlM
6HAQLt5d5dhmDneTzACOXQ1W14dqXtLy2JppYiDfFRRCLQ/AJxbVki50yuexFNkOeqI3unFynz0f
fyOYjgeBWS2Z/8LTgyBAu0Uub/EvdHDgcJqHlDaWxC+8LqPg6NmCF2NfTdezhyqXfLSsXVlmjuDa
kcJX1JWlw+bomTBVAB8eK0E9hj0useEfttqoyf7R8uH09imgxpQ6gKXFtfduWIJJcjKq953dIZap
nULhAJXqd+isztpD391lEQhgURzXcqPhouS4iIduErhlSugfjArhyxZ60KwnfVu4ZoS8JAXYlRHb
nrdJfMPelnbRmqgpW8qIogkuRGcJroiggiU05D9OhroJ6jPQ7UMqzHdxn5DMII8jsz5oWvNoA+hw
j4sRBgXVU4HxMtEGH3YkD6dlqn7F83TVE/LpYUphJMzqr/6RJYGtC9byysNt5ZOk/BOptVbH2Ws0
fUT9c+zirGh+et01PBmhUVmw9CiAT6bP4K9C/DC1Lyd3kj0Q2vveFEiM6KYRAJnZ/lY/qGkjfakv
uLif9gXpjXx4C2hUTKY0JaqQyq/3qDk8C/Wxu2mKNJM3rL5HTrISXWkBw7R/2P4pQufoVA8O6dhL
GFcihhOvILNDtcRcWoHaMg2sOFrdSH5SBsE//VhsWNfxd+iyrA57Q90IhZjgN5PqFbgFheuOcE6j
5v8mEDvtUcyItmKCOa/q0HR7g1WVyTRWkXcVH8yafD+2zilKT7rouG6NS0WXMYx4jho0rWsTHo5D
DfLtzjuBCZcXDFm++Z+GHWpFgx9OSTZETjryqAbtKdUA407hTekUynHrlUgD481MeR8Rs4ACTuPa
+rwH4zeLVSRBwme7o9v4KR+PJds2j3SaHKrPwJizUqSGXYMKT5qc2/bm1T7f/5eZ+IMu9jT2yU3P
/XX8Uv3nK3d0F+V97JFbK5zsAWH9ssMXoWp2CzmdF8BqPKTbAWm7Cn7tHmCionzKspl/KS7T2h9s
0eKjkhO0akadth7czRQ8IhvjYTla5AQZfzIjoo6HMCK5E/ukFc7yZHj9nEs3JJCl7KoUzwyuX9CL
0PqUdynTW+YT40i3OFUqYU4lcxbtpa/46nhFCSTt1pfWp0pr/frES0fpcif1/IPJD50UbvbrBaP2
AyyBNY3BdhgEMPp21F8puOYT3/bB05zigvtwKPcMrQ/pe2i6KNnJYP6gqT6rhC6X/5atLUE2qdKo
CusOuq9AEr+EaXDEkWe3450yc7HATeYgXaZHGjcmSoTzn3LqX6XTYdCMpHPJXfNP4BWM91ir5n34
9GY7DfMwjaP95s10e//38n3V5RsTeIR7WKswZWC/8wJcy4lw/0Rei16qiUbwH2du5BXXTGJdJXTY
0XIbgDlUSv4YL9H5m0M7DjH/LT3aHE/GhFACRKKo3albqS7R3Yxro0IUvCalOTqVUxwN/zz5UN4f
SlK1cVH/Uaxt81yrhR6R/7Gtqy/socoq+jrAGvGnmMqysGjrJnBBNcdLZHuKW3aza3tLqJ0nMnkb
z6igBE8YkiinRpwV23HJrpXx7P5+8Z+y6O8iwfY2wRWdqVuy1VuiTTVxeRATcAKon7K6rIyc9H9o
YFXF40vbylk42Ke1f73s536mn5j5TMJtzVf5YlUJRkKIp3or5TyGJQvRg/JpxM0CVWgRIb4xebTT
MPNBEb7wcTn0rw7QyFIR9OJbChQRQ+/nRJy+oGahkiXb7vNiuTXcedhPsuLjVaImW2oYZYkB+0z/
TOqPvxKvZY9asnmYA+agtxRggBVwFOX+RIo79TOJ7g6zKC3vFpGN3IgNrPfovJZJa5RKHlGkEL7g
aPgl+7m090MF2L+N96xkfcAiDk8UewtFXAkU6auo+foksWszC7nZQ1N/bHxZJoStYWQ1g4T8Pt9E
oQcYz5/VN+Ql8HLRHL9DAta3M3XJUUDD7dDy9qZS76ieg8ypnszKcF9acq5KG6f+t3BZ3N0VW13X
mCLoXFeLrHHo70H+r932MCKtpfNuEqyOJxGlh55R/WO7EETGESKLZIqQOAV02Xfoo5FV4RXEYDRx
wywaMRhBMjuOaDp5YfTBHfTf6iIJkUF+VQv9SWuWLYEkdJ3U5Vq89tsGv1XY957zfY1GOxI+d+tx
+KZmICTcLzv6TC9bvuH2psn32o6N6RiKW0e+mbptZs7CW7qB9S+MaQ9/Ufe+58vs3xUEzDAV043m
gAD3FmBXR/1wkYj6e4oSuHTI4fkVKhGko5UqZx1lYVWfpqhqosdnBBSDxyz4189S9v/MK70Ix86Y
DKocIVWunbah5Y3IbQ4utYCRpdk8qA+XCed6JxAOfb+z7g1qBwYaHOgns5RV7bxcCoYQlgHmDNWp
InzuZIFYBbrsPK24dWj5cXnFEYJ+VryQU9kdcqzt8gRUdJaSgiD4JNpy5plqerkvYqkq872XB4RQ
JS402VRUbQllVaZXEODEL/eZszvGJiv7v/K0L5tF3sIOvSPhExoFRBX/ufbBlmEdGLxEchBxWAeC
8O913pSOepowkSIwZ482xyNR9ZdraXhqvLgTclckxdT6wZqH+LfsXwOimii648zYu9fF4HR32tRP
f+ETWTBKH4iktDygeqdMpc6l3rfPJmTqg0cmwjjEdAHuiNj4Hw6Pk5rqLfXrPxjt69JAopMhr540
hQurEgjA4zfPoQqqOS6+PVQV1WG6bWckGjvRcYnKdTh10WDOZNPzqNvHvtwRxkKns6p/YXfxjnpV
8DwDb41KC/wO/EIZ8VzgcpNnoHz5YQlKv/ob7fVknGNYUvuetI5mEMMi9aS7tnxFaaIJouz6hXzv
pJtIMPmPNMmr4imkqa3sD2A7rDXhrBNyJq7AYezhc029Xs+jz5yCPKg56BHxe7wR6mzZx7L6DTKk
Q9W5Gne3uCHo5Xj5udF7At/BMc+ZDSJz3uOJD+a3miUKbO8JzRrvqeFsSf2S0RZriHXRQL1agaA7
LVlV/TwjSgm0amn/Dj1lol7JG3gnTcHN/Ed2slcAJHfX0ghTnUOUSM8A1YF81fzgEF2GzYGuzYdb
N3wXrw41+1cK88LGxyw5tbsNANwBUDYknVtXnzoYzJh8ELDZfFQRGJUqy0f3i8ewU5tYVeqHfRzY
kUvQui+8IZwgawyPKrd1/FZP3R0zN3nfzG9uWaz7o/f52ip0P9LFRywiPPAV7qJS6lIqWDlJY/r6
6O7ggpcyMhlycV2TTzlaVdLzIvIpNTdX+VwtW0P2eSe35M2DVzfX/mo8cLjdTnfMW7a81HX0uCo+
dDg4gCS6c0k94pf+AHYMLV2Ey6ZHFq6UFpZx+gpaoznfN7ZRhlVtx+AlsgmLJb//ChdrNSuuZbGz
36irI+un+0jTbubZRVSvuZmuVhHiY4UsENzMEbyZQsOprYK4dxaCYP+PFaoSM3hnlMTQme7Liga+
invSOFh4R+wtXjwzkYfvd4hK5eqHNOD9h6tE6biqRglrV1QGuogajigTBLGgj9lIvtfws0i6i+c+
4f3uBhMcRzyoD7zRIlsJ88XxrDDZ2jBe4jzeINdAmKR8kvaZiAkpLPpKDtE5JnJbqVLyczAbfpij
6ZmSdn9TCAx9iIg6mlWbbqWMV4XIftgybfWeAcd2dtHmfgjxrj6swbBelb+iJR0MIOMsgQEQJcjQ
A7v5DzsYtURlUqfxdITbRIIAi/gm6ufMjVvuJMgbiK6qlP2eZTfTs6GZ2cYde+0C6eDVg+UQRbKt
ntau6rAckyDcqAdno2JF+OXxVTgF2amgbJR2SyqHZbRTDNPEh4pfQScPAPuYA2tuiJcU/Q/BrbU5
tGKEdGHVbC6Bh4pMbUgNdOfUWy6Mx6pbqpRGZCNz+8gxzbWo+ISTl+aYfsMpahYnLouDTwO7Tgly
wkgSO6w1b4dFNjx2leq3xEw3zbBa7mpRsPH6KSVb6hdLLwveew0eMWVAivtC8MWsWK/DSt/sgsI8
DlUqfARGtEDYi/c3/O+GnX2cWUXx3jhAyBr4WeR5b0STFJfJftz5G/YYAJ8Cosw0GhhN4QZ+p3FZ
1TapOSOpZ/EYtq9ItczFVDzn/O4abRwV9u/68ebvTwpgCkYHZnEmvzC2S8a9DynPDnhNmv3BAkUs
p091aBBgWvn7x2k7VB0uw8O426LMsT/rG5x3ty+rxdHeq86d/Doyhxp1IZmERF25ieZkCm7F76dR
4WgoY5aXfY5Dm/Gz3VGFxV1NygJEdpTBcv6ZesMkHo7VX6Om9FgetNKqiwByim3OJzfK9v2mPWTP
I75CVGoWTCzLcBBy0OxRb6OpUMX8Zk35ke/dMnsF8vXoV/OJ9eLWUF+5VnLJeiw+o21QBZn6tm4D
Bq7fx4Pais/cuERLxpnENfaXWIl8SjEYzfWQtR5KTmPImuif9wQcOZQiz/fCxRWmQQ7ICKFQ02m7
A1PXXqGldV41UfBVS3rmF4tt7Rxw9FQhz948PStKKLKrloX8jTzLqUmo2183I8lQ/RrPRIkJL+Qj
elB7OwYg1HHYwNrrh+gc0NjyuFuN8bxXao2LBx/ZH5dcerkIP2erkJGekYg/grUGN1y5MywDpz5p
U5ZQ4yiE9WqS3sr0LfCZobnl39xgPvqFeXLc0qfh3rXdQSDjsyriB8s+WErbrRrujqBS1Sr8LY8G
qmbi7Ktw1n+WSrO/yeTWInqAH2SFgMBtpYBBqhGynshI1C6+RvVE88CbpDKr+g8VMcEK754DXaWh
nL6IpkOnbEc6i4EayFvED9frhYPeWCjPwCiHsj4P4XR06NRQ3g6vkOBGBKsROHL7vaxqRPzgGvkE
mvW6hPqqPSJyMztJ3RtlwaUJHMgxd2IOkAhcFmCkaDMYNZLOEFG+mQzYsY94522TSlpdAi5GVAAj
lv8Z2O0XP/yE62/YV1RsTf1tfHofnVA5YXsxf10a+X77HdR0LxIjb9rNFTxrxg5+6sULCgGtFOzB
Gp43ae1fZSnYvlOlyppB/Lbq3lwwe66cGYaDhNOw7gCi/GoNAxBKMNb6B8brTFk1dnL3uKFZU1Wa
G9xbP0NN3v+CbyXpKSQCRLjUg74gf5vepE10O6WhH3Mu3SbqiSypSdCF5gShPgRXpJwslAB4sXRo
riLM30E8VtYgMnEoQqD4RgK1jQk1gCYp1+VsIkHEZKTGv7Jl0FwliH0jX5Egwp/VhyzZJRpqndBy
DK7t8GWrVMEDHRckmztlxfEgg/X+z6QD1zbA+bz4aeembcjpH+wvuCXE0q7b3rh5OANuClsR2QQg
HD/Kr0p5R3AKKmTQEfLUytuJagDV/wb+cq4ZTJaQqrSdm74Sys39L4twJ9cR9LfjriYVTY686VH1
YCl2akJlJQZpx8WzUpR11BaFAByizPER8wqn4N0EL7IDBsTbeanMoId9rJXw70pU3BDJJKfrmd56
fNKjmYeAG0tZjMLFRwVu1oyrKF2ym1L6JqpkNp3P6A+Zm5jWpHhbjedHihIraOL2aktjgQB8rRxA
u9LMlDOjaAeJDCzVzOmzqjLaDDsVwubkIDTb2Wwgi4SBO64HzPWYTHSf6a/XX2juBRiMZ3eiue5a
p8VYRq3ZqJ8um36HR8igAVio7V9AvEXdwxbreknU5xBEQoNJoqyKVFDaICjeZKv7aCl+GZU0lWe5
ve1w8xwsPLG0BNu6HMpfiXfE1P9s0Bi3ZPsIFFwDBH15hnjMrFQD36ciCERDrzJ7StLy4Kq60iKP
0Nnk4boUAcMkvLZo+msXBgnFyxqpXG30SdIAeMqg1pt/a4MptdKzBOvJMrykx0wMriMzsmb5tlHS
4lAsYvBJ3qIugMbQjBOiY3LhgnGpzPMEwiVdTVLyZ9ly8OSai8Y1/z5uC82akf/wiyFmkq0uk5eN
cpRvjRYVRLAggAjCoh8ZGZhq2wBtUJT0rfU/oJSjo/tB4ekhV26UUWVgU9kWAJeKH3SVdoNN2GwN
tUy9SnNBWtfpGDy4/2jtkeid+wuNKmy+fKnYqvVevhhJU6mBIwfZVrsIWrKIm2obQ7FSENAyXWrg
98Nyu55EvHPO2xe0bziKy8PXhEEoGU1zjdUsjJftbcezS3VzRi+7lULSHPAPPkEawbkM7Bo7wLkh
Kkfg2Itm8DFfIFA0eayVevEaPuCN9n/deTZDly1+7fs2FDQKBXDEmtHNLcophK2p9o6xUUlzm1YY
04XtjRj/zrZc3GnBcnDkH/L9hj3xkVH4k4rE8NmQR7r5S0/BooUctI76x3VfU+AE/kmgIldW/yhu
MgN888i8w6/MxY1rqg8KOctqfaxO4RMWAdobtD/GQ4Cg+9guVyO1u76PX1W3bAeKmZsAIJRuZRFU
mDZhppcdWf1r5xLxtEpxExsdFuqcAiTJGCdHxw2GvOZzaw5/3QYTg/v/cZqAhcPNo7mWlcYVN/jq
Q1Hv2aD5h5oOwRrQH8EftKxK1x1ctGgflgysGdAmj6vDMl8tGQXtMPNaiBO9OHGjiharoTxyQet5
yjqulSQqbtjg2DgU4wpsA/S1PXIxcIg/FIOu/0IzPXiSeFwqOA8jcJNHjg/Q6U11V1BS3Zu0QN9E
LAPKsqUHKW7k37skmOaKjHxj/tnxcG82ovrxftlT80ygYRapIBvmSyuorYhF1GP7RVNxp/jJEbTX
Y0N/eJ3edwbfLEKRHsUyNNBAURCgDiAXRQnLidyZ7x2PuAqUD9RKonM0b2htUIlu/qoHSHVdXlRy
MQqTKHFyhrfFV5dWlZ/qy61bwgRalNtL0W9hNV+HY1Nzu/GJjv4wGBdCy20g57ChLUTyDe/5DTWZ
jGmpltrEOiJujuL4xdJ0qUmemM2c27mJ3vXwnPOWSwoMPQ20oMwtmbqRCP64v2pFyrallNMOt6wJ
VI148uA2l9nZEqnJer5bbedkz21NKJyZ7IzfbqA/0QdaspaecmQVXUyk3krHS2B2E3soVVtNbH+5
3GGNyRFdrCW5TDjd9JGX3BLIyWj9ckqzVe6MmsbaRfHpNNJ/wOy2ohoqZYS/axnnEu2OTVJ3XdFj
/ps8W7wO6D5cSf9KXPADGAzHApVBIdVyr1TX9AIzF6kL38WM3J0+o7gHMYViLimqaqZ+9zVKduWa
Q7ZeYsZv2ykLpcI6HeHg6FaapMOqn8RC4fjlCsAx/FVDxhGATMax1j3tLlY3WC8oSsUYpPJ9WADg
2q04qVXtp+cKUdBVzMOHXoaP9NkgPu+0JLTuWUWFgOZP3OPZKyA4EVUBBMTtz3CnZ1MoOaFkhVdv
eIzkNraCu9yUgw34Py+EO4d7gp7qkRioXucJVy2a6RpnLMGHb2eTG4VmFHr6F8q30A37G7idDUKt
BX1jxwOYhpuXWQ3D6hDanv80WprHipUIUlOhJexMFVyN973GYQx7w6fVPQNP4mu4p/lHHMfZHs6f
AzqBnNYBn02PknLOUq4PxIqKJsDvO1i00ztbh3aGGc0KCmYj4GMwluMiJg9UQbDeg87QygNZqSC0
NhOYUSPsmCobVryNqZp2/94DgoQWokWiMDjHMb+K7kt6FFfDHQThNpY9Udu4Peo6u8NU48JlvIPj
2T0sXXvTPnsvqtsUHWDCGrMuA2DUf7ugbhydQt15ckGjT+wkGrYeOrjwkEyanKxlTwBrXZa2YNve
ntR7zr4Zy16XR8bm1aaXNjy39OtcE0vbGEgjuyfgUGtR/GIheYmYbhRlex0yt0/e39Mcl//t4iKB
Fni5oYf7b8J7npX481vB6beo3R/21xl+DkUFGYF8DtsMBlpOnY6iWDyt8w9cLiBNYFZLjFCjAQQn
GFDn04CEh3vZyA6ji+6daOjHTdk4vMrW2+gUywgI/sFy4N4Pkx4TY3ZzZw8JSa1hk0WsccEeUJ/i
fwlUQ37LMMaLnLggOHlmvpNSmKZZWKIfAsZaZuoMHYLFpTpbhqJMVU8pZSzEhXpqwEdSkuAKlvdC
95ei561K/2dAQSCXloNsgpVRrsX+id9FgwPgnqINxw2eeSksSuv/XW0TYBkW4uDAJzNG9fNx8nZD
LkRKteqslBx7WH8i0AGqE5IXn8gj0p8l3XqzfbNzyhjmDTnpgqyK0k+01WdhwplbKVafyqWyJH8Y
Kzvuwn/6yUWav6bxTYxB3xMFAI9N5kxXEvTMI4vVGk03lh3DmZyqA71BlMh8vK5+Dy6oS2H4RqPm
KGDFnzY8QFZB1Kr/j+kpJXc1Pt3J8/+cjmEmseHal6DkMfrZ3qB4d3jqDMVn07qpEKHl2cXeHzcL
cBgBD5ybJU5iUThSTW25Vv8edOA9A9Au8liRK2NlVEMdhnSIlozfKGhx/TusDBk6nX1wAdmQzCqR
S2uk5YA3a8b56IlUm3h3vr8KpYwZwvKooQon3WhGNKm9GTcoYyedbDNPe858XTpTrNBaMC8gLVXO
cOiDzgawvPCQwzkGRFeGR54OzgYzra/DgKmJW/qmhrV5ZFxuvk1XA2VnBExZES2fFkDTQDcaDzS4
mOwPQnX5PlfEgn+qa4Llizu2TNVfAg6ZIwwL4JErpNFYN/9FxFNqo2m+Mofr8iryTtEK0ylfQ9Mt
28b5S5hxdi31LIrPyLrtpJYk6Gm6pVOSZAHPPLCa5aQTJzdtQD/paMw7omq0X2DcSrhYfHHBfU6P
d8i/Ysr5niZfz3IPrSdqHBaRku7yz+xxR8ElbtKFnTkjOX6xOGDo0dikDEucUvju8Qda1olxGl4O
d01kYaLF4znl/sH78+XtK/BF3xB57/oSMo2z/mcVtHn/X0apAAaY1SJUNK0lfVgG8nIOvbk8m/0T
KSIFz7QBDH/Szesff3IGmyYeU6alpdmXvqaPUJJim9Qv7dibddg76Zf23O2IlJ7sGIXtgXnBWnCC
db7l6h0t5uY5/DtJMvka9zqAnSOA8mT4HbA3XMu3r89N8l3afujQNfL1bQyP8supkH/IWA4GJEnA
rc3ypPyG5w3apKF9SkvgzagA65PDx8sl54ItOidCJ/aoWM0QPOELDsQ5Od8uDJcMbo9TZuHPLrtK
091CsUKk7tGlcA4g9XhRaeV4vY1axDln9tH9kkGBE4EoqbZ3V5j/VTUWKJkd8Ba4JAggTv3uJXlF
/GWGBU31RTHgzCTpLOtI7yV4vjPMX1xoF3FglEXDuoVPsHfsgMvAT2DLbFKxuiqxWfmGmUBjfQt2
1UsW/mp8Y8wJoEwk2y3eclyVuu3xdgLYCDMmhFqN9VsFt6z12iWk71rzxlGkwaO4TJhpJPAzZi45
j3aLV7ZXocN0pLg4pCWXXa3Tq9JE7ufn5tzIh81Ng77u0gWSWICWit1ooeI6Zp0pQvmJ81D8u+HJ
6c5QPtnJvQtBE7MQJK5sYEeX+Jl6OzZjgck7yxQ/FnyoV+7b4IXUTw2//kvd9NgOMIlPll9282AZ
zulgU3X7LpTQv9BB4J2nGCJLs2S//hMowdesXXZiLSP1QAQlgBUjHSbgW2ZnMHu2wPwDpFd2GLfd
l0cjKXUFN/QCuVzZcX6lVChw18tJR3mOqjkwB33GtRyQZ8od9h56A8mSwh4ExO5uKubUAfLmZLYT
MKBdvvhkaWZsRHB8hOOp8SjBHyFzXcbmxpsIuHCLGYskF5PmTSLZQcnDdWwQBb6k1Rg6MqTV3nDI
BrvKjFijS4LYISC9FoQLSWKDS3e6g06Ty8mn8HMThU3+2TD4xiR9kAPJZ6H0R0VPedNV+fX9cmKR
aGsV2LjHMwjw9K+8gEMI4a+vZ9Ao5Psx96MvBM1uCHpr+WJlABBJQqFmVwmVPIp3PeiOatIsEvZL
w0Bq3DseLK8tCbOTkUOnubZ8TluzMZnidzvsfc11GaHW0sxvjcX80XOpFrIZxCYlgKBqy39YxbUs
M2W/d5/RLr6HWIflFbicdhZBl8JHa9zhXZLgc+DIEtOkUo8dPAdwzxBB4UZxElY7t+aJQ6Qq/h1J
WJhZ8ozEGYHl1RTO5QDB8Auk2fRYBqYli4dnwnXeZxsTDA027tbKoDZc+vOW0GQisqTk7EMsS87q
d1SX78UB7WE7A9tfkOx7LhU9vDc0qG1Tb/OPa1gRC6GCik649xKdyaB6Hsx6s8jFSd9ETssRKxLA
6lG/N1bTDu7u6/5yFSTnO2RtBIBAHf+v4HnQdLfCPvxTJ3R4XrqGqnJp30ctWunTv+rC2L6j9LLn
J67ZH+KvQQAceDHBVTo1yW5GwKXuiZA6yl+s7a8ZoFzddYVonrzgJ/IHj8f1lMICs1wxWlxEwoNU
CXHZyUkV5CorcXlZXOyzIGpkDiRBWRUgx4mXymnD3fy94aaMXGyTMGhLCU09HE7z17lrlFEs4wix
G9bUyWYyQ2x7tdGdmFpTRSCJhUMr6hbi9Nmm1VWRNnTblaty4QkXEraEJRmfWby1WJTgYjkRQHzb
pUUkkSiJJA31Fp1DpP7NZlZkRxlzaXk9KdQWE8/IXfmEn4rT2oiNgHp4w7e+UOoOkYn1sVs11E1c
VDCqpjHIBXvX0wXIbTI01m2mclvd07U96q3z1sw/g4fwp5HhQlvoi+BWEW40LwwaPzMMLx/1NDaH
26uGRfUr7LrXPLXGk2gyHPgPdUe9Tax97HRsH6dQY4iadHu78farI/ZALTo0GJyleDXTWmK32heL
NhILUd3/bqyW2QA5G8JOlTvmdJZ5HrUH1j/nw4HioW1R5bGvKjf6KOPdjxYsWHbuGOvU1npS7Nfk
5ijo+N7Xwfcfry5efOjBuXHjQR0LI19Mu1lLz1QMnZDZ/JPBB36Cry7r8xBg57AyqHzh9QX1NVqu
ruJKaVhQpbGo/J8vHZtO+JRf0eEN6OwBGJrMWXzBPUJwTxGJe3ICHAAAoTw/5HQ3zG4sAUSCgT9w
9OH8upg6WrV2bMVEvcMqBhBUZ1cdkaj2sDvOeuMvriraBCBI0aJ5TxJ3x+6e++Tkjt1QX3Bx4hsp
BF061Q9zurp1xbsy1+9MiVBqV79ahI5ZNZdqM9FfexhsRp1oqNBCXEaOoBEJZjUR6INY/7rwlG9C
GYdBusl/QDD1iGPbXTUCB67oU3UFaxVvQDEysTuRFXPuBYShAUGr5nAcnrzlDJREpetBFESJ2AQx
FvH6RSBSjSq13LDNQpP7wNEhlFS78F9rxCx9G7+KXyhDgnhMfwllSUgmVoOJBTfgajY0UkOjUtWH
SIgTNpKZWUz67eClFS1B2rSsJcyoWUWfZROggQP55MC/juY9KMshRt7S545eyAUJBihHKMfSnHg8
lUzqr0i5+UdmtiVgwDojguMn81GJT1GW/zTQc6MTD51X5ubRFTywE/WiSE7MD/Ao7C9QHhAY/xuJ
wdpe4UBX9e/AZPlx27OTTNfZ4HKolMr17gfJlWLLqcP1A6NjRZJwhzZLUweVfynNUEKggEsGVEHR
sGmOzxnzJBW+rdk3iNa2+ZP8vddHLaJ5XvtoZyNyGDP5vhhdq90j7SC1jupWuYMh8NEarbHrrIqN
od0Dn9yz84gCC+jKGxI8v1tx2+niBuMYXxh0DXAsXVM3Yls6RWACQPFALcqE6j5AY7MjiM6/O4o+
0507GfZOj/YNEuY2Vg3n4t1MMEo4/E6gnZZWqgZnQF6+2E+pXYt+IUBl89a7pXJjNOMj66P278ZS
R3bp9DN7pGPQi7StU2kScytFTUAaE4gnKtb4FKcHKGoKqRPmd4IXsAle8SA5Kt4tKyRjSdpkODoI
BaYvJxI9lzgNcaCobFpnk0eBkYn9yi1fNqChp6arnm6sBeAweKYdT4A04IF8fqph4h8rPS0Zuk+u
keSStoYah+SerRuGKKooCq7yk+T+wHum6p9PV2+eud97QGSrTDRNzD14gzCPjWBF3nTyXcVtJQlF
ZFS5NmfMtvnXrt7aGXyNfPXBPvWdN1klYEWXgBMgRWqdRPbWZ0MfPDweDO+TgG8ShHEJeOtRPNyY
UyWhoEw/zzWZAcaVvR/vp3BqtJzvVGGC1rxUJjsOwNfRUuav04yizxfavb1ZkWoPLyWmwqbdzSTj
Agi60l4Zxerrq8uCrdGBQrA7lx8WUUj9YjyFQEoynC2RnvCIAlnHaRpTNL21i2zsyoXUorLiYQss
Jv8SorY2TtFKr0KQp/aBIiWkdgWNIrgcgekopdB2YPy5k8LX9kGC/dauwJEr5grjimWWKSoGMBtD
lk2nevRCVdCIeX7PqDccRSrEKLo3cE6vLxA/9eWa6kMH0XwUdRAHnW7OafRKweD3rd9Z6mxmOVTj
5Vc9hoFgKwiXAayYJvDt733XRoDnp9AX7PU5ntsA6+fqG+LUoaPZKw6YyHhrQPvgM4TfFclLdBV4
FEni0nCNr4hjEQK8uMZT4DqP9Tuu9fzog7bAdne/AOTagR/J0dYMmwGNsl8VHdQPG8u0xvhJNmCm
3MlvZUKmJ4kuOIvHkMHp2OjNrBiEa+6c58EsSKPjDlLAROTb3Vpvl1vINnvxRoutBfbdnbNU2ieU
JtnWixMbdlRr+xvSikRPPJDam0bo17R+8b1ZQICVJ4Oa3005kSBtL6GEEFD9VaxBuBoACdhg8+PT
OSQGWocEC3wDfo8oLhWSd2XdhWd2iNRqAidr4HFUyC4JV+PqTHoJ2jUzUHMJgdSpaIEKijXLC78Y
0acKlzGa0E48q4m4V1n/bza+eYLP9CpLgmZgSeK4ElZVQIAR/gKX8iUDszcPSxe5mWmf/KIjj+HZ
mlnGN0fzZQ2SFhbnXrzoBivMpQDP0IC6bp8264xkC+9WyzbLO5fpyFZy3kQoCB/w3yW52qKpqb/Y
qZA8wVqtclY9hQAuoqIuZ0gFaYbd8wprLfLMhAHEKsCzteE9kVmtdiZa3hXKSar08PyFdO6OO0ew
3rXQ9XPi1EzjupgAhFpYyAdNfTN4fOSBCOKsqF5hF/9BFU/csiHNzjiffA0UiAWWJoQd3uGYXFrV
KN1OLh1muvMHQQe4rAnQOdAML+W57AXzDDnkbgU1BF5PPms3NzB4+wz0NoZL3vR/mKyUDf3BGJWo
zpJOMulvtfPrJiu+m7B7IDuhB4K4LHYp5qCrkN7QrjN/SyexgZX8Wz/gK8ZNDJeSMnqimF1fMAXG
4fyQ4xEmaCWFUAIdOGLzt+O7HdFRvKhY+oHlJmqFTutbFC4vmFrOcsY0ppGQL5DgLElV1ZxDEbkg
VINK1QXyw5lpdmgEp9s/jiarWkII0itfl3SGt6qVmv2P1qr6SD9mkCcudZF4ZRuh6aDtrXWpgPJh
+09Bz8A7kVd2vTXhUF5POHzEtfaxONLxzTsL3TpuyIyBawIGvIeKu8+xKes63f0MX9SiJTbT435H
zj48mxl4lh9Xqr99pj28pB/3zEaKdo8JujP2KdpcCx/9LLQF1ejlAdy+9azRj8sHqXbROkHI9qjK
T5TS5JCUHo7nqM5RoAwqJQPdtn6jlboEIT6Gz/JRavm6oV19U+nb7QA5M9LICjXClIw1TPW4Vx2V
D6KBp/xfTZc3SGFVCXqbDiTTX+eWbw1D6xb4IbA5sCkGOtJEHMMCyGPmITXjx/TaDxX6Zbj3/b0R
3jfk3ylVRk6cta7yKZKD9bjVEXDcrjzv2KEEmET+2dGxv36vIYHKg7f3duVn7AG+JNMFsoQqBZa2
t18MPdilYNVXR4EawV76YsvwaQFz14wfhkah2DpJTxUcCd0SA4W2l22q8CRr10mrIqnZsEfNXZ0C
eHkbWkNhVJmSMlhYibqoYFsk6KovWzKW5UQZSAYx4h+EiFJLHlJs1QiGjGltyeBsmQudg+qikfCR
TcJv6iVXbbLlLSqDGMCZQz+IxkGHQ0jn7vQ4lmgo33Bm9yp8nkPkdOJ7QDDrpvuig0tLaaUBVfyK
LLqmA0RvehK46ySL3+Xz9/fy6DCpBKTolTQ1szzRFK4FoS3s5HMtNzIkxZqONu7YnZLTs/GipCyD
ws23UsxBgHzPqfq5YQzzxJC1aa5tis9eb+twq8c492dJLbaWu7qJvnkC+Fald48b4lle2JcQYKXE
TZjfij/9f0QeKETKdpwYG1zF5+5TXNTvGM3UUnvt7rFz+Io3k9qQ9L/4GL+MD+Pw8AtiSkqOBj9O
9JdOpGGQMR/t4d3h1QxWSFC3YH5MnqcBAGliqIgfp53v6VMMZkOCgjsd9TdIkugM58sa1NoaXIrm
sxNu11R7mU14OVd6BTTZAJEh/lUKF/+zylD/aqh1IU2pWzBMIE5hmn5CsdIqE/idXy24euUsI3ah
63jywHAikEh4advE75UQyPex1V8sXDJZyizU1wwDKxmUfTPFiWd37pqkVtdNcb0b7Tq7AyZgYJ7l
LqDKAlCJ01ck6qspScWvZ0MLVHn8iVS++bK7hR9FGB71je52gEwQhslbyjdccx5nlDfyoQO/okSi
7v6PqOyWHVat7qulQdPgGMA73WqUkTeBHLesEWzOyjBmB3cch2vfFrA6YzEGSkokfC6R0daThLDp
XCPybcEaz65u2bb7Z98pylJWk8jgud9QRbR2FC0S1M9AaIwQEToETmdGieGSpWHuzd8z5Gvldlxs
aBmWnp0qajkPu8Zar5fDrbV0wWUzXTgtIKuoOP0HpruTMDsPwUBnrWSq/yWTbW2cmRvoGlsQg9wR
xRYuUXk1DPcnLWrU8kmeyxGd/RS5avh4x7on0yHjceGT6vr+JD+8WI3pVTBLAEKspY981SIyC2yN
pdhwFO5SjblaKKi2sGgMBPsJMTeBIShHm/wl0eNc7zDMd03L9w5iYzLqLWyNJexiRLUcC1/47f/R
kVhmDm0ALY7mtkuMVzfaMjs1M2vX8OweTKSqjNpRXQViIeGmuQy+URAZ5CZTa03USJBtNAjNMd42
wkikUpTeTOfMA9tRkGRDdvRzanlMFcqcRcPP1ntfGkziK1Tgx+tbxZyEVg9iy2CxBfTHjwLP/nNt
yljIACfYxcuHPZkL42ZEl8lD7aVl5j/7ZJHqGNKFA0VWK6UfizndODpBgpW1eK9SDFDOZSsrQSRX
MhNOY29Xxb6eh1FeOJ4kBEJUcilWJ8x/PwZTnNRmgiUAiG2Lz0okSiaI5Oc/V2YKyRZoYHdtIV0b
a1/BiliKI0koASwke+oaH43EA7epH6I70E8qkDMDYzRZ0qmOFYy3Q+Si2KBGlzokw3tQpaYgz541
e4KmCfRYoTC4rrI4QmoqQ9rVTr1DPA+FGCklnUkeA+1ZuUXSc6iG8G1djMAYs4AF6wSphwgMiHEe
IX43S2/EcQvr+cgAFlkLgiDw6evNxeL92dPTWYBw1PL40aqplsrtrpb03RiyI6y7sA9NlUwhaCBU
1peZ4sJ6jFYYjBuaKz6IZLuP94jfWFg2WQEl8pOe9DAhxRE+zy/3Y8HhLuAttHxVtBj+blo4RNOQ
UfEvfnJpU67kAFOVJmyMdm3AGvo9WvilML36noS6KzLLheshaLSGWweJltCqrCxLiIpo5gjIwyvx
57dM/E2dXeRrRPdeMqlCUBlyTfTjZ2kG+izgtpv4Em4j2yl4x+VgpecFQLgHoSY7ChCxFd+xU4hj
YF/kLJsDjRLUfB2tcGUsr6mQmz92801lPBSYSPkUNUO0OA+bJOHWEmhMlPEWKZUg+RdckW2dk419
flj0l1BnxQlv6lmgoariRmQf3ZLcArciDoTlqbkq1uqk/ockFaCESsm76jCkfaGz3s6hAsn7Lj5z
sDDpwxs6BSd4eOKpmKRzAZljaHYU6uvmUK58cQ7TlRwEJYKRCdRqiZ6LDq/S1VHGe2I3aJ+fv018
Y97gGZJcWVOLhO98GtcQiHcpuUqa7CqJHMOIt6XjnwclmAQFT7XJoiBplxxvJi1OLOffmtZqJHL8
BmOZ5xXPcDnvg+DK+2N8byZF+wlMr4HjXrZ4qnA8i2RD+MwYqu4HAl3yhkIeUdAwBI9Ze0vfDp+G
V8Wp/5o9SYePDxnM2I82MrykPPEYqpvfgvWkMH2YY2JhguS7KyaEDYY3wNMJG13zjrS5GW5KP+gD
JskwRxxYt5WKjjm92nykRVUGHYTe+coQlx5TPD5a0gKI5T3Ztfl95rlCG1IlLz8PelSEuYVd6Rhb
8AQWCct9CzVAW12wqF70Zq2v2yg+znMsn19bHwRna/bjAmkqV8WUB0Kq2sW/l9Au2g68k8mkYllz
w3PUsjU+bnosUDuEQVKH+V+0Gg2wAZCS2OkS4mC6lsg88ODzvCtxGv0ZpDBIcxzM3ylS8F5B55ZX
J0U1wZDcT97wvwBULSLIC8QVLEtGP07KFDTwF/D5tyUB+xt9gBDBQ+apdn9n+3jcGnUpIKX0jUVl
ls+zPDcLVf+10wneXuvPcnOj9qysIq7f/nK5psjA+u14HsIGf1Ogu0JJ2KuXEYyJq0R3wCdhH/h9
/d3hUzIvEaOUYsW8RzLiXIJFtZtuOtgagIQMD6ks7hcZv2wO8edcKjekpJgPqJWsyCxhzd8AT3il
Ul1n4tvBWldhJNw2sJuYMusSK2I+deTP1fPyLYgGXp92Cdnah6zl3MsDQKOajVUGNSJPvzaCcoeN
OwlSrbasmB8K49IPwG3Z1MVhk/bq8iJBV5yw3WUBKseRr9Q/Yz6pmaO5OCdFthFpVPuE0KG+8LR7
RsSu1ba+UtI7VYfRH21CtCIvU7A+W3RUle79wojdXFtmE7CAuY9EOC2qiWXefTRwB3HnIlngU7JV
mNziV2obf6IADZxTj8wiwaHQtYxT8B/TyhyDMRlJE8Cn7//Oyc9v8nNKZJ2Y+gyp6YKSXE1Xf6+i
FQ0Q/NtIfoBga0TdEBlihiEjEPY9ntA1ftf694tpMiJ3AZffqO0ON0S3HHfqrgWBfzqmauAOJ76Y
0ib82l73tIwKytRVSSxC5Ug1CgtY/AsPjMZ4aAphmnbCYEujk+6NJh7wr6GXYbNq7cgzL9uiu1O8
fVhtwk/DmuvLcUNO9YxWoTPaUKvnwnaq+4GVs3W9Ty/tvuGd08lvGFViL2KdPH4OSRcS+lIWjL0L
sw93aAeV2z5iWrgh2i2VM3PzXpMF9eIHir4qZRkiHtaiItVDfw9lY1z/jtJqlqE9Huqf4aV6QKcu
WvEajGsWtZDBM9k1cUKVnrYQHYPcq/cFAkFi1PCszp+K63CVxBKqNs7WZK8kUYeDDlom0EOoq74e
3nxzuG7g0L452yqtnLF3uRcAWKFLQ3iQR3Pb1XX6pN0ckyP4A4jMDBOHnUI9N7xy9cg+npAiw9LQ
YIvbx1ETaoTjhFbPdOEvRuhT+VKvlcJEoamN02Q9zZq3gum5HDRpnlHXTAimfUk4WsF/kyaMHVXz
2sndA4n+a+fp4tkFqz5HFLShfKW5wP93GjlNy+rDZm+d1UNNWDQKFT3oUqjFMPlgX7bL+GuY7meE
mJ5BUft+QOpuiS8qtQe4g/1nXEs1uyWbvHn39+vivLqtu/NrGWS1ZBEI8CBu/nFG8zCZ+g41aCcd
735dxQq3NAe2GUHoDlbS7LJtP14VCBXT+gjE73MMTHFtTxQUL63rNHAMkemrk+hL0jVJOsBt3qpW
7IVLskwxRBbv0eOwRsxYDLZeqXyZy/j2bO9yH6N/WTHf3VPTFbiBLMilsngdLMrzgeXl76jU3LcO
aiceno9NO1jF+bQO8FkNUceUb+kzbi05HtqdA+4xCu4ZMqlAbbrUYYoagVvdSGiPo57T/KcbUiQo
rZPe2fGxYjPOghAzG7MGaZuhEJ0GdtTPTZGleYsn3u8EmpaSpBEp8ycnbXDscx7AN1gyIVTls9aQ
xkdfZ6wlREwG1PRhXZlrc8m2QBuu5MeHIqCMpjIkQkLGfNlSbHLd6Rvtm+GonWNYs1klRBRET8Ja
K/2z3J43msMZWoadZMvPUB6QuRu+u1OJysBXMlW2o4IN3i+5DbR29TZQyVnBFSiY6/XY7xmgaj9e
Z+rQEbmhBdE/yovUSYrkyI9QeesSAgmoXqj3ZGFZdZgjwG1D4GWane334k39rnbHKjJrXRN6K3il
mUI19QuQrCStbaYKsjvM69u+TnATNwHbBDW/j2yH9vb0ZsVTpjtff8ZXGHWhPVjKIcUZty/6L/3H
5i9wlUTKix+DbynKJT6Py3thfb+rJFQbN3vFLPsdfifUHFnt7odT0XDi0C+ilHyYQlFS5ZLKmYOb
dYo/87pRJznv1WLUOtEl1Plnbpn3BQw5bK27KAbI28cU3fbqYAQEz7sResOeWdEu75gjUM5H7WHI
Bq52qxHgaPfk8W4W494QG3Mzz07jUtuv+k9Hzw689DR/8dSNbklt4gixk/bg6izO7Fz5oK3dKKSw
b2+h6N7/BeO1AMcS9f4mskN/nEyL7zCFstcgC/LC/DcQiGheQKTba8Xum4wEqG02y6Oul2OiM753
LZcaj2JyDnB8OzW6AjOeTZ2tu4PAcxW7PNc5gqSMO6XcFWfnO00EToynSkXL04Nu8TNkMlIgkFv5
es/1h96+ZW4wbKmLWXsp9ScWp2/01xe7NPZodC1/lI8U6lstpIA1Gsus8sbY7nXUCYPXoYY98OjX
zOlQO9sErcwxpTdewBA9xVBUWV6gNhz44oFCfgTUTV8Tcx+ce+Pb5jkrVMxBqPL1+gH9UoLjA2Lg
mM75bd1xNDqMwzNFlUuRzUR2RZdx9bKES0p4389DYIHS6d70zUWq9kj+ynVG6ZaFTv9r2pcoj9rO
CbINnqGni+eUM6CSO5sJ4tlCkQaxgLXz3kGGlSTOg03vytR0Tou7kdtWW53S3jlRjravYCMGk//j
+fYzaFZHt5oRDEurjUXkQ8UV8aUWNu0vfXQKjhUtX6bJDWN2yeHkX1HhOidrBQrTCMLdtMJa/Feq
bLZ+1kitWM4fJepbw4Y9t037yWPaZnDhfGfccNJFf+xtHpiIT4exo99P0pzrGeH/g/faaOhqVeOx
k8Kk6hYDxmDOZ+VLyje7eFmHyrXV9i645QxrLJxSl/jc7AzJRatcR9GPJV04omkhf2tkq1qGcwKC
agqYTbSB6wDxhkB+297q0RJH5yjdWehKskPPmKrFZjYa2WQfYWEn9B0HHLFrDdSxxDOEsnd3OPmv
tv+UTtxKaQGJiBT6TlecLww1ddE0nuCpsstRQzAjS94fvyIbp793gCt8ImLp3mzD0Fpua4ZijFdk
1+ipGLpTKOZM9oUIPJVXOcnzYSj16FQ7BeeAUY5VCJKed84QXQcfjeR5giPMsUqHwq9oHMMkrBAD
lKKIJ8KRxiqt+OtWaLDiVqRc4thNhIsWkjw0fN9+/W+fBKFFZVH0DeuqchlsRBcnJs1/4FMJzQku
psOVdK7zIc18kFl76hA+B8HK1vkqdhUbWoEruQG7+IrR/GR5fiB1iU8s3/l5jfzXvdr68EG9Jy9n
ZLkwlyMAocV9B2rD0OPrlcaI0sfusmhSrn/5dHQA3yPsBXG50rttoCLTsGQG1RTjbsizf6BcrSiG
1vVUM4IRqyl3NmSEENKKkkgJGv7o+aW5HOycLMBY1HLl8IAjRJ64m6nB35uhkk78VuUOHeKkq2wv
wmoniSrDX5UiA6sDqZDgxmqNw+JDmZ89GyJ8us+4leBAbvur2h1FAmtocNqM1LpJfs88NoVf3j61
ZdU1TlAOR7tP2lXjTV61R63RfOZjjSWfvEWFvejcqD9LQPKS/+FzJpulYqVY5aWGk9gWqVu9cnRZ
+1l0YDKFfcAGnpG1pd65seqRvCXdrDZffGpW0o6koX/gqzSSVODUpsuEKTpgeAjgOXOLT6NCNLD0
X2fFdUNHM0Emx/acEZoA2D4TN0JqDZ9uOMVCv8KbBkc3gFhbJxnBnMK6wJF9DbgKgQWkaV7QTVgl
E/u8duRzo0PTSy7Mus/S6N4sVckvoqfdv+Y53E/1AFDXjbX5UByAN52irwJncYH/samw2C4zf4hZ
lS0khk0Sz0xReBG/jk18P5OIUf5be9WfSgCIo13LcYpeHTg2V9fG96LwYZyuzfQbEA1zvPvsDH7s
xYe3gXrC9PSSdmXq9GbDD1Oj707rpR/c1t2PfKGVUgNQ6Oi/LsFbtbSFsUocxf2uvti/CsA/lcYC
wlGxt9OASupYI5RY/goYrwZR5FiKZmdgFG694hTlKjEffvSSA8IBb584iwBCHlzLvDu6YN1RiEfL
1VzzOHGfxlsY+5nrrgdJP3vHqXEKHOAuPR1YbLb5wj0/BzjMpq1MQ/VlTPOLlIYKR9H8b46o156b
0NK2DJFprpcNARTGnEqsy8/Wrftwc33kFhQCe+bTfPT92p9HZRsxYaboXmeUManw+sXLnyA5htvS
BMZ6X76H+eKv+v+FmXpJRoIWVbpGP3f1dO1Xp6YbYe1kbAbHFPfNPCIRmq/zbt5N/TQlYs0Bb4Yh
clA5/XLoGDIUh9+iJyZ3Gp9aDOvlcQeMerii1Jtt1oJK6SaJnFt8NV189HLyi58VyTmVH6q38jtS
oJYDhjDxU/+OO6/oVFx4cfzGBG1MkDlrWKYqwPP+HHMoEViyM7QyWHn2vRatDBvQ6olRxEmo7LLI
d6jRJIC1juPrzBepl3kuDdk0ODLUcfNXf74YNOpUYGiBQBJXeGxV8Ed+MSQ5LZ+b4oXFaAHvIm8c
ttiM3OHoeacLjKNzhCxG7kU8mkjHl52nFQBgmNxEWXwHbemDPFdjP8TUHpGqGQ7xl1Fh54uJowhO
gpJhaJUPL9alDYIrDrnBJgpbdNzskRWCmtoklbO35I+f71rfhvQIfBZupMacdf2pcAMeus8bvYWE
S1paUCMtb3AD2VeVKTVzpmlHBgDCH4rjcPuONUwUTIHuuOnUT1myurzJQQjyAaB21ymIdhFOPJK/
ghTvpWfqRPYYcVrgUPJyKRjQ160MkeY8VWY8FZtj98XicRgXhGp20bphQDlB0L9ZvWbBzlMoseED
S3xLXb6ff8GlBV3icfdvOxm9amZQmHvIpgyx7Kpf65JI2NT6/z5zvZJFcchg/qE5dLolMW2rHtYe
VyO2GDsEergOLC+PSCw6ziYJSTCGswCrFff9wdN/pwLqXu26a/NVGW2K48VOYHhvUA5g1u5Id4q2
mUev/qpA4EO3zbxO54UNqyQ664c5Ydm6MjcaqLHmgAVJaQWjAXjxe5d6jymXu2udMva5+2qikjvP
4sHj1Kw2KiKKy81rAskBnnJmvWv/Jpssi5JJVfoLjvAhv23vO0/X9YGPfrhUArgMZRiS47Y9XFoc
BbBN1UKf63h400WHa4aNTJhX/zXNNn/WdQOi+lpDGvLwuaUOSEOzq30Rac6t9Dq69kcN1KmhTK63
g7M+PFqSp6miRhyHkXYtza3JtLnuu7DEKn9ScEpTdN9DScMFpzXHUTFp/z7mGMuTLROhZgpE1b5D
Tma4hovzSJ+KhjEskS8IORdWl93WcBq2qgC51fLebx5qZVuBNl4E5HBgYFpq5TAUeY3wfEFrc/pk
+WhwhiNLGS1UPdsttbQInkRpPHulVjKoDhaLmgXirzUX2i0RsgXOhXnt+3WpwOokWJA6DS70Yiwx
tDuDIOLdkKRj5DN6lzMV9567NUngBUxxsnFZpuMwcTjHJKjyK4J/9GfSJ8KtndejYXOok4flQXo/
1NRdtUH0qdrhvgskscAPOd6mdh3DDJVdlOhwUcrf1EaWV+kLHCIeg+kN75nlhjWqE1SPlTYWmqrJ
IHYo3ygIUXagUpJtKRp0ZtIZImZS9cDmR8qUNyWqouz1Ol5Gm//CEwVoY8xIxWbAjNt1m5vHfFGU
7lA6oFcsSiEBXqwLzT11j87aBPctlw1UPXMmrpBpVqEw/iudE8kUIcNFjtu8n1s8Ul5qZsQFzYka
Vg2wlGyd7H13Dkshtrs3uwxMzkMVmWRgXnZM59LP1N5F/8elQkRKiiFiXmhkVCcQPbzw2EPnfWcj
CvWJc6RmH6I9A8C867VGQsYbDTbqEwH+9klGvSsBS6y2EN0/JCi32J3ossWReYxNauZR/PLF8rF6
togBbsvdefusnz5uv+lQ3aepiOplj3/hsCk5akxjpy8YAJF58lhp9xmVWMFse+OYymskpQxvHVeC
wEpV5G1P296MzEVF3g/FonlYI4fyAfuvkqAkVIAli9u/hO4gTqK7I18OF5KTmJFhlcMGADSyExo9
C+f2yOIALvPzWV78dIVSYsC1DCOPWrW8eKYwBLq++9zuTxTFEq1qME8LVRhiyZuEkPdktVpTuPcO
BoayJnsRUBZ1uVfkSAlyu6gxMPGPBtE3+iy36si7mj74fc0U5ocH/8oToJqiUOAsEqD7SCGkZiA1
xQcqco9A6w8zmaofnR5TSVd+FWwDGbBLa+ON3Ng3n873sE/qVQP8jMEgLwmuuEg4B9pDn+lJ/Kjw
pvhL5u9ylR0q7KG0LDaXrpc81fW68TX8j/z0SAMWw6uV3N9aNPD8C55xDwwAEY2/H8fwCjbmW9JU
fDYLIOD8pSzwBTkFC+9uEUaUiWPcjyUJHXwbChYbylrTHPMIBkvMFtqAEGUDJdr9hNFQQlNlMz5l
rH65yYr9gFyexgYUzmh8BK7w8h+PDcsHoVP1KJvKHr88yxIOdMaH/Ilj0S7X9Ecf8tXqqfLWnSAH
1SW6HLcR1lfPCJVqf0y2f46rjH6tnz1BOnRifPWik8Bl1q72u+tfwDDf5fTI8KuQy1EV6Ud+EW9M
tZrtmRkcA2I0JWOE8CQwZK+iSp7++KSpGQpNFCZjc2/zBB2cZtRqa9CTQjx9iQHnhAo8HTpvOuVw
6CwKg8SWExth8NG+qLEoqxtHe0QHTS9IajdRG2gEApuHa1Y+7CQ/fRalPMHQ2TkKAIrTxuYfVRg/
gPsUmBLV8eFrhoTF8wyNJ2OCpy1fqvHF953vuXT66CJPzoSVKg85T/AawOjN/Z9Y7sntnFfdq8tW
DH5SMy0lL38GPzE8IHvLBJxPDqkK/AORpv0XI7MXGiu2Oj/OBfqt4q0vrAWEeDRNWaf3ucTWQW5j
pEp/I47R1seouuTRrh2P2NbVZ5mVnB5Gr/FHjB4nvG61ACnP/q08xJXQnwjMeaeH0H1i38+QKNQM
DmDbsadKcCcrvx+1mnE0r3wHgR5Xt5nrsxgQzkXHrQYKbdGXHz1cFYVpOUgUGUFHX1CjOmQ3UExi
vSczItqc3IZWskTnTfiGIzPv3GI++Wgqep3iCREieDWjjkskVMgdjjB6HkvRjYukhR+EPGJ8rN8M
KmWvhK5t5TLNb92L2wIfYxVM3RaHbu+IJgR8fXcmkBsNPkUTVtE6GGpnKsVBiV5Sy8jj2XaC/JR5
BFClyBRdMqJiopSUUkrhV0v5qzVxnc3ekS7e2H/8pxM694pVsYyfBw5SNfntj2rG8foTYdEb4R63
pZ4H7E4n3AVjzPEmb0USUkjt5IWBeBRr3PxOpBNQefr6zlPz4Hkp/LIdPfan5uBSWlAL/MuT1ffl
gA2tZ6BZIYnBvut4M6Ag8P3V0Ci4PV+MSqTurqC4SWKmZqwfCSUCW8P8lG4Mnw5yNNr5Q7JEDwl8
j3UShfTB6pRkMrjfHSCGwpK2Prir9blu9sfnPz4EYwVnA/xfvHUAafamS3GG95nZ5MJNTH2XFL/h
nZwlYSBfxcQlPJdwRoYkt+1+fQp5KKLd02VPWApxiCAMIQuC/ATNgR2miffc6MvgDcfZldKX1ESc
INodZz0zmH+Nn87lP1Rnhp7CckO2pjmUizpqqQKX5ohDBI12XEp6Ddhxlhqu4Ftp8r49pyExrQrA
8mIK912D8kDSPLI5V7vYkSiLHZfGVBOWqDL0WJPVEjOv9+Xy4r9rNrcLlz9/wr6sZYKpaETnD0cQ
PAfSg5lqBH3yMML2JYChJQ2+Vy35YHsi7b2TsY9Lv87EM1Xa+R0B6oZHw5DmlZBZppxLkfbQlAZv
xNX1HGXKCU2lw+HPYwqQuuXryYB2qzKJIIQ5cc4wG1LfuMam++OzRI5BUo1jVIVoKckKcal++Ov6
xvDOvVePDRjGgNPtVDXuF1Hf1q/a4KREvApXSMbnUkC9BBez2D7Qizhv0E3EJmGMVBJk5XhhzDU8
8Z6T9hIgM/nwDtf5PH7JPEM565PfUxhwZ56VAfPDH7nacA2kRw5kGqLdYuBceXVI/Ju05ucpBUwD
8S8IqZ0sPi5tiUejIs2DQZngJ6wtbAGiuHjx/cGJP/8QbW6Kk7wUtOgqmHjh64upMjyVkI/ngNgw
q2zhf2ly0TnPv/f/Q3rEr8P2zPZg0H4V90x2bFcJDIROo+JrveX/ro67oYllEeshnoIVU7JbCQdu
ITd8WVlKiSc56wOsEXPg9hMHvMaVvdt6ExzStiNY43uMWUCZUzBJ6DqHfT9i6nxIpPhtwTr2kJyL
83KvCxwEWg2K3OAizAd3OcjsqQEILBTfXjX/XCd+FDUkxCmRvIQwxRxZL0ZTFBdbE/BlWd7j+yxB
hp12e1cfRa1gpIeE0Z/W9zoU/8+I02yP3KhxOKAQ2PykLU6vMdv1z0wTcF6O8h/uojnyEIkGNemA
gLMjKFkX+WEjMpQmcznpoPEvpyZUb5KV1BaSu3WbShmsakqmTOHJ093p03F9Uaaf6D2LSXOomY9q
3gPzHIR/5vuXjGNv1k5zRxsteeMDZh2fXDcstzIfEXe2qNvIGwNhxAOnryZKPJRp6tJwSzOUMReM
0TDjADJC1PS/IKuhRDHH2xBXn4dSAWNnERDIJ6QHpb+fKjDWnr1Z0F34g/dojR15egzcVBwiHWCK
uMEVUv/gC7iRmdTAIga6O8XOGbS2YCVJECPaY+oeBZgMovdB46lT7a5aVaYtRw2rtlCs3EKTySBx
zr7B3XfB9NoA2Dajbu2FSV29VhZPElLg+mP50fqRC5kkeU7PmWlNDD49MZevAWYZcSU1rCKA3zIQ
avQg8CLQNku8fqKUe3cccXVavWKkZ+pVF393kVN/6P+iQnx2Cmqrlm4pcCqc3E/2I36sNZ//PJgG
Nz0hI8p9rr4g/kY4FX7eBzP3D20Ft5YOk93VgU3uKPkcsNdqqbTlwZl8Nd/WSIznXVc8LN5nv7we
+Mnpd/5vr0UH+u7O+XkMcRj50ajl8OEltht7NXw5FXI8q1qW7xX70AGVsRWF+opvqC1lhi4QYiQQ
uptR0gtP8qrEukjBCEI1j5LP5cSlQcKdX+YnqG/WFqxEMiD4n2soqF4HU+uj9TtA36oH0/yQy+1D
mYUUDeG6lTXunUomAa4yFqXUh3t4mEiQpgsoXhwr1Oxdr8gi/Jo+C7mqrAliU15OXyOaAnG1ere0
omE+AtG1NqS4X9KeBGilXhPiKnHPYb7d+nevNRCBlw8qsZ1cN/1ee8pSTdnLfmNRuChnEEjEKS9C
d8EuoaIrWL9DnQrutXAP8P60NpyegK0txOpzwDuTVBgea/hUa3oCXMbMxwPeKRBHE2e0LYGoHvu3
AOrjyO8ytvULMiBhTqeLIkwSHwlWcAubGsNseBY+hVj5CT2U7azRlsPUGAKPU1tPgPxFK2RDZas3
c8R4Ma9/nPIDjmWnqfzROYCWkscrbYSzD/apjjvxbI4XQX4LcYuuDSlfLty2BkmjQ+K0IW7ma2fx
sSKGPc4fbx+mPlzwZaVs+c6G7ajcETq7LOVA76G3UYSIHYyGUzTu/YVC8Kx0OEiEWkM3O6E/jGJW
t6F34jdWpsXdCw+pOEe9vxX8E5PjjR+0OzXD6IOQ+kmwwbzbM2h751kdtMaHNPD9Hq6tDvzAakXa
pLRJcXBoFGxzFP3zhMqMAjmANZF/9u3CIYE1t6U4gItRyjcYz16DtPieDV2Pdj/E20eE9/Yn0+8M
rUk8IT9cILnNhX7+8tvwEHAoJ0jDC8gGO1VpAJOjr2E8sCg/lSRhNT+q8Woa6q2aYatPNpqBOE3v
QyZtNVBYMvX6TjwiGra4ljseocebq5X4qKPQWmOLZosv7vdHuX59ONcGQw3qfMXfljdq+YG4LKWp
u3Xkh6vhCcAYYHWBaxe6VhVViPjmJWUgeFNwfweBxcxuhMAE1SUqWwc53IlbHmoYQTl/dnSo5wCz
vZVmvKW58pP89YirmwT/NZkxo8Uak9BrtJnAXCqJdFsMACpIcBiqYVEOWIN52VBqDlmq75kfS0XK
Yiu9AGCdnJQht/4nxUf0k70p3Lk6bUicULYRZkDasvymSoyX8ms2VlkZobdOj6wiG5ZO/UeRDRal
W6vb9+WY3lnEsi3tRHayeN8lzFwRg0DNPqcvPY1ACBpQ41RxFmNBBrtEdtCJOyPZxF7Ck/rHEuPC
4fkv3I9d3wi2qz66318imyPJsaozpxo/Bf1MdXxzbhqtw8mfd1eWlnf5QaMBXnmSTJ/xDJWJJ4S1
X+jOzqINDvJxJO8MzaWP3KKmjy60h/QReKicarFjuyaXah1qSU8bCqvxJZXyKvahYvRu7sgHOnD4
i0tVzG9GA5P4uTuk/Z8q5ks5+zcMx2x+ErdWUdzeAI9cAnAUBBQ1gkTN1clVttgaC7ly3GgdM5wS
mfJfQDjSlaOzYtXAw/v2H2K6uOcZPFwBeA9iF23I/P3BdkDw1h58aTRn7VBBEolxFW6VZFdy9IcD
5Yo5OPyXaVA4AoYaoochrfPVu9q4tP2AYMkGJhR8TuDIuxbmqtACgB3l5XnEBD1NElo+eo3UQ9B0
vj5TJbF5fznSoBnkJMFDO6015nqR6I67vFIPqtfQwEYbsqXOAX3Ih8nu+vohnGiattvTJBK+OZyE
s7hb5n13gyMx6a4joDQt5SKYKdnlsH8RKQbHJdRHUGRMVS8TA3KdNd0TQdvMi3zzyWjUvj+h98EA
4OwUdGOfmg/0Gm0IslnU5EtGL5IpMY+wz9AUwJGLjmsLHwqaR+YsK6RudMzYhb8saCXLK/85OckC
OGN8M0jyMrexY8PeT0rCiv8Y6Yoe/s9OafYHOveAt80q1CM537YTyXnxb/x22AbgJcrDb5hdrBS/
aWAwAwk3l+aqTiVTGTB97WZZvLfRwuxX8u9iqMEGKe92V3H+J/An91hRURsvD35pC6WZnTn06wDi
/DW/Q95IYYWnyM/g6B3TuW38kFwE/xwY9+9kmc/DH97J+lKvl9QgWHzGhitx/Yb7ZWIBxXY69Cq7
cPBFwAMC/BzTzG0cjUKukWUoTzc0JQyZ1oKhawQ7BM2HyYoZxm7rJDK8Z4ebB84GHyrjp4eyZ5ar
yiUyeaiqd6SUl4U53291tQm0BtE1wIjWBWGM2K5daF6aZjyEnt15Z/zP3ni+PUSs+O2AfKvr/50c
LKbGiqidn5uKj47N2eO7/2nlHm+BIG+ooAbmHBEX7525rvC+KB6nuJLIEpxmcdgZ281fCJkxSDcW
jtKtRbz47dCvRBwgE2JT1R9JVwsT6gx65bKXTMqKGgzsusOuIceAyyakw8g/kwwYMvO/WGhQpqgT
tTWhX8t7J/3CQMspXESWuD/VGon2kOlRFT2dgG4vc3Ontqhcjavf5y+tz2ptB+zhA+FmYeowo5oP
x7XibUhNL8MdRVSWk9N+n9AhZNh/tZTEC+AI+tUWP/8GC2RQVBpEf51Ry/8i7isOYODIhOxXsm/t
zeRlCD5topBy/m9NdiAE0N7xtQ0vvEGWhAuxb4m3sjFH+xMRY60r/FB/iftfiSIOMb/+tQvKHElO
563/TIl0ZBMqoOtR4ZRW9R710aQLgtPHbgyf9ERGrvMUvzSEthhs7YZnVwNbzTzOJL4AycIIxldx
JIPOWA7U3T0RHL27zGaOb1jhl1m2RDfIV5UwWbmzh+Smn6W+xjgDFiSIDcRXFE/B9NAJJr91CafI
h9ck8Ldxu1e5C543EtWcdC2O7xGuyh5qv5xpch7NCXyN/RF8HOsrf6LuCi2xaA/y1KaXj1nioXuz
aw0uOG8E/LOb7ckfPHZAdzU4vYvswb8Ehtlq+nmUlnCyNX82Xewpym35AT9/Gn0LXLIijxOmb+Hc
Oi9h8E1FBFI8JPL3X3WP2umt4OHWdasX6XjTs/SHGyuYyKCrUOuMfriJ5Cs4aK9SJ2SCreYPM3C8
zdNf9oGL7xh330Mu/U8ejrgGncjYgbFznwY6rPu4B9CILD+X6VdOc6al7U81RQufKISu6WZ/x5eS
7xGZ3q9l3wfD+T2RRH1hgJsYi7UyD/Hrqq3cYybSzUqrUK/Ben3iz/GxBBKQpiGlGZCv1e9ZrMfr
fJETVD91ZbLtT4QIlPt+SHgvZBkaL1HbqxAVBiLrAaEQtIZEM3dtntQkJGIZ0B7Y983PlYpGrCf8
iFf/HKL/VtUItnPF90qmT+kjVVmeWCrebqpiW1FIaQPxa4E6OiDHF9CWnRVWvzx1iDqBxbQt6tv2
DEcvr5kqiSfCCC0VwfRsabIdyVTj8qX4fDZ4ILChOtEEf4/lW5o6ACVRl1Fk9Of+J93KJNH4FxbU
cosd0xJmhazObmXhTDugCX97Ab8Noh+uqO7F+4mfJYSN9MLmSdg4+pqd51YTOEYDcNlX6rtIIrns
JMfW1Yhd5LEAw1IYfEFQs5YfhYXrRBsBErt0hytzIjBWaWdag44BmbnN+ciOkCOsWk3ZNLvAGh8W
HNjuNjxiz0cCeHNjT2owB9/67Q6Uux8dSwfbpEzAgipSfenlLQZQdT+mVAaPo+CGktizsXgFlR13
H74ZSPXONh+p+eeD/B15XVqiZNjGWQBTbEe/BckitVWaUrVo3nRFWP1eggKzc4xbHHkNZXQKEpwU
YXMRE1HUv83ixj51hzUMggwdiniEHh6tEHpg/ICrbuHyXrIhLGOq4Y/8uHqzS/0QXqrtTrZXSiMA
vpMFDBfrTctbRg5qU0Lf9AJBA1m//f9QHf6NqRcBawUuVdbi4oqXUXVP2kfrdtpPHLCfD7aq5/V8
+TXvg74lQba4pCD39KRBB/gOmkzeZkLlYJ2zp4gbAOy4hvA+uBw+hg3dfmG+vwgwfUC3tvkmo5g5
yLW29bZdPqlGam/08rTsKz8gKNKzVNFnZUGAMCzh9S2oruLGGhwDfJDSiUSYZxF/aaLwlAJlonn9
7+k0DXDFwlQLG1FweixXPdEX9Y5od/WwKInm4d6Swe4S/dmQdLqf8E4MfM0rzarXeMLnOgEv8xgg
UdjVzsk3TOIS3v908s5iB/FDhQIPU8MOHunXQ5l3wJil6ae1TZveJ+RZ9ClDAJRomKQRclrvw3sd
xwl5R4QGjI4zEg+07GSWtsZ1znvVTxiYNWWgxU1WOuvph7wfPlKJyQfaHpEw5jpPEdg1FwH7YFMW
x9B5i8ne7Xi4/v22KDA6otBGMK9FjYkfLa7k3OGrPLY+GPFRc2dQFPJ76SblPR5LxnQAlq6BcxJh
3EGClLUtKoHMyOy69B5AzITostftp/2+RYB/nnJbXB17IQkntg0/SzUVWNEyoA8EW2xzXF8EaZHP
Xajp7iJC7v/nswjGitkVHNYAd4G8UDPhQLaZoKLPb5kd+8+V6qVImxCC2KhgSLqlSmN/wRfziSw/
AHTPz5idQ9UnFm5vJls0o00vui42y8RCTKwMWkHDW5kBz51Dg0n96lYrDki4Gwy5crt+zg/xAqyq
MtguE2j+BpxWjUZMtcAxqr4TAYn/LI8peO+K99uf0mftv+cQ0lBDBV6HlntFdsvJVdt7GKajjZyY
H4nAFQSionCwnbxzXXwjENkn4p6zCRQqpngxgNcXI34Dra2BTHtFR0lpJkjhTDlbB47+bWMfINXq
iMFU26bwJNnK0AvBqkfwiS2aH0aU9TOxVy0mftp5Hw8oRei7462pfm7gD9uV5n2+4HZoITC/MW9+
qV53pZP+1wzR/Q+H7VkCM+jwngXFY3UUf4YUL8jYuiUqjLpgOU26X34NRwQNCnYP1zEsIanNL/bn
XezwsBuyUF3lDtolG44KsXuXAP0kABymOTbHidOoHRcgm7VUvXBoeXJHzbgCYHiZi4n8L3uZSYL4
ZTtXrFdSnkKFFiMHogMOwtKRSv8aT96e17NBts7ge5Xey8VxQaolcLvlMec3KYzoPk3tHPRBTJum
5jO7CTNR3AJqvk+8OEHvIpW8VFOdCg0sS1jFfYJDueffcgqb9SInAlYD01wSx8lqGm6WLjp7pB3K
5M6CJ1yJCimfCgaDSFbAisuLH5R9zybmlTpfb7qBSAXpxlf0R3LGk3Px/quvey8r4YHLqBQiL+GF
b2RKNN6bKIDwHUq+ECTQTI4AkT/yTTai53fI74FEeROR2B/y5eGzLiD/trvaJCSf5mc1s/5h3Zhu
oI94EQIFsOW6mdUNYyKtfR5AST7bBF5YMJKDqLueUZ2iYLeO590yxxjQzdEHfk2SBuuq21GkfIyE
lu1jWkK195FvfG0PDqF6/oUvmTrVXqEJK7uzyL6e3bwdjBU4o4XD0PdelIXAazMvvtSneaJXfVGC
TzJlMbIZeEJZA0sNeAH/jRr4dfx7etE+h9O8JUt5/YAwSrivRldF9j1rCBfYlq4m8bdMUC8k+Jia
IuOZQe/tHw0xkGinIzqVZoSerfg6+fjK6qZ9EGnlmEBa50CWUzmYVw9KJhC8cJyrVOrFXLhaOZqx
sxyg2HQwa5FGYfj74eb19Z+oyScoj+JHVEAYuxTgoMx16P5FtaYZUDp6fHzjw8Jbb3z66nZ83X9o
ZBYqsU0xwHRVZZ5IVEp/8iZ3TJ4Cey5dH4zObyydhDHY61fSyK3g0i/nWgg36IwloDKiIk6B/uGl
kKUhBXnScx5+OC362nIqgT4gBQ0y0GQTGUoPQYAEvsZX83LHtVmJ/3uB7MtM59qbJrnDAWNNqpko
zY9iNJuusxcty8AjXsrKVHrlXQKeqDTyl4trANkYvtOu/z6jTs4SlC0AQDzWaBHTojeFqdOUTnwg
+HgUUf0ddzWaOgRPn5AWz/exF6n8ccK6HsktiY6UHZ1Hcyvvd+RYwSre3wwpx9NFgSQZSr2Tl4WB
gknhIykqIw2w7Sxfua1zrqqZxaO70OMOLKmwVT4JbbeEJLj+rH2JZwHE6vvY2PsKFYuiMb3i1Qjb
fQqGk752vKi/ObrNYxngP41yc5qPArt3X1LsVTLZYp6aMWwQwhIPawpW7LAfKEbc1g4IMIHvyNh0
tYTs3WTxvEmiRxkfI0+wTAXfvt1mq/Wn03pUCd//G6EUyw3SHrqBTPDZoI5P7tOX3w3RLp9ekNKV
dz3is+s6JIEM8vBKE9o9nYH5P6PbjJ8FVLbmtUeYDGNnptzDa6IVQqnvne9avTsXshUdIOW+WCCZ
tj6vnVLDr9aWMM3Oymo6BtA6OrCvc67DJEr9wp27STgg9e7hCaZ3HrTs48qfoVT9pv6QFWetQ+g3
LF4ahnjzREcKA2ixw/wDwOyk8LJUmja/Kf5OZFpaFPcH6kL9xnLAVrlA8RDQhL+YeCfoUR0jqyli
See185nr4UfxTsqvqIoVcHKUyVjHLY3GUzZQN4xm10bUbrH30HmodOHzRLStVRGGMNyIT6vGllGC
volwMgRXKfxlaU5QHG+j0zs8Fzmk8l+07c8DCJy507Ne8VjUWZyaZp1bjkZwE36PGo2QKKlD96+l
f3cvRg6t7dKA+pxbPB3/7Mlyyp4z0Y7PnrmJLIghUJ1NCr6TjmBZoG6YNxvh9FnNC2CJNWkDNjCp
PrOurIaolAaQKn1Q7frnyKcXP7/motWtCA2OiB5W9R3SxCEgiaftsiObKXwA9Nan1DYJgDfOtJEd
J+isU3dot/pajacSzOziU8SK1aK+y4uC14AiUbiNa9j2WZJZw69P4HVpB1eCxUD7cxQgPDlzCzvO
RehSlaoBEkAeUbn07ns1vgGVTXnBJHixm4Tl/0nSnawSgBuJkwCGwssdvbHRDh2rXX1wtKtsI3c6
hQVYVXiqtiNu3w8mYArsroT5DYqmplwKFE3I/TqGiDnw1WouuktQ9Ulf1kkdmyFoFVoH3GdkjoQv
xE+gDiIxvDOJRjaMOBTedBrHBYN2GzJm7Qoa9Ub8fUyj9LTRcOkD3GvWUx55FilLI8qW6pQt4LGO
rh2j2dShvW30fbstoQ8F5wlJh1g/ArnFnSJMjgFbPxkqirxadLt0+8Y1QWXkNMa2mra4C4HoO8Qx
PugkPBE9LBz/V1mH/d1eXbc8VGsta1nPqsqkqd3I6LLMxc225WRcBf0v3qjKRDmN4Tqd34y1gv9d
0bJGODkz/oPtC6Kmo/I1Gs5nSISnPNWK2WErwNWViSREElE2KIC6ePh0B5/3hg5Ci0EqQMWhUBSu
cveSjkQYksb1aiY9PiXl6u9gyHxA1IpAufSdDo2pUYnASgvY9GUu/lIkEwkV7nC1Nyp+/aJnck+T
kosKSCjWayfNophbvctvEa3ucn60qnj4eoodTrnyw8zueJc9zkaQenKdOlFMoSX7F1BjswdvwGB9
yt8KyJI/GyUFJ8QWdRNAep7SZp77S88DlmZa/jx+Et7Qlmab7onEwWoR3xFdYD6hLMDi4RqhRwYW
tOqHm2+Ch4enxAPtsg03V2+P/oXatPkPVFP0PBaxMdljjv/uZ1ZfWrlkHhCtxKFupD6xCaoU7CXH
Sa5Z7aEDt7iIwyujiYWbMF73+2xcAM9vh491JuLHEcTmcel4A96pUV7aeBHR9vwxNXlnwvgfdlyW
aPO8MRyQzA/kc7Hm8+9/ZQ/iNDdZira9QGT22OnZ5WJbfm8zO2OBv0oseALC/sowccEL8leM9IMW
lHrKOae57XVTxZkcLSvMA2Z7vaX3GZdzrkks2s3IzMFNmNZl0b1wfAe3hkYxWxWkYmz41b9TWCih
4MIx+MAn0I6D0mfVVUqlFyG7C10o7LLsyCfU8w2ln4AT2iiQdbwyvC9OXSBwmPL8HngH0sGEp3Dr
H8p45m6hwIjeBrEPA43LXuKliNOqtdIHu1iELUc1FeNJaaKGB6RUJNetMhoRxynJo/NvFyqNJpbv
NxAmfD0GOR3k5rR1cL+6Ku0axlpZ3GmIvHHaKOCRk+G2VdVJoEu6QYo0qtlbKunNrtUb8f72sgEA
3/oDVG1n5zW2u1lzzpySELMF13hcVzEeieN/nsc4gMhn2dwSMHa/hnQVsNNGUddSMbdQNQBLzk8i
/DatKCThu/Tovma0E0ghE8/bNoXLu2y7ICJv+UEjhF2xK03/8DTLYDuc5dzHCmMMk3o3mM+3s8b7
7abbDQ3lkstZrpNDsYkZxgcSgKVNJEC/rEU3IGu1Ydh7mldKhbszNlSXRx5w/7afq5Iq8PO3ohZW
1k3lbrnoIbIivSzURZRHWKzeVKGk5aahRuxmAl8bS2DyBWVcUFkM1TlLg5P8MoD5nl+4MO0fRMsP
iyIg0Ue8Azlpz3F685vYZr1irtpE5AVwu5On412mPwgILG5GbuwVy5UPn40nujq5yAoq9Fz2DE2F
b7daSsi+pEyn5Bvy8znsg1AR2RJFloTZ5FjKlSeFtImhxngokQF2W8XH+/kOLU+mVk7rjJDkEj4B
iyWTUAn3B+sYUHEobyqb5vx/4qsrOatVBq4ccfACVlOjH2CKLSVn3qbSDJ66tTUpP2zoKgq5j1iX
C/EnYT0DYp9Ygh0U2CzMEbL5IhMwKcUGKd1YkIcIbuB+PB2N2bpNU/3cNUKrvNAGq8fNrF40hP7Y
Fpq+zCU4zvZDFYQ4AP7KCP2cV8O90bC0cihcPOQ/27nFkd5GFnCBD+HnPr+238sGfRuOuceHFZ9T
Nhz5yWMPz2qa9r5xooTGZe/KXqzWBJknhdJ1YDaV5i+1NDVhI5T4mqxZh7W0B0jLII7Y+SV24e73
hbcRReAR+1bKNtGHFLSattDz2nbU+6pj6L2UOlt85OfQfH8cvDQUI69p0m3/pC0eh57vEXzFAufp
nybr1q+kDBd4CkSm17l8slIom20uRC8jPaWhNH4snf7B6O8F5Jwq1HX8R1y0kGpMv4oPqQUadwlr
gVbe9jRvaWiIwVnEv/ZSnWyaKcEiTVdmRFUIyYDyPJcNSCNBKp0xVP/7Iz+lmvdlp4+Vh7maZDwo
ueYhufLuPf7OqFBkYfJiK0n1hjxSpOzuuE/cm6V5eO7TxRsKMfCvAmI0Fr8N+QFMIm5MykqRqg0u
evHLfWe5gzHK69MwqSrd3CmUTrTZU26LonreZ5GiBMs1UmxXeN4Z5S9tI5eYoKfx1KLLaQ7N9/UT
PUUV1usjgTutnLmpn4EvN+xUIdLdV8jkAywCt9DYbNzErsms5WVedep0LVeBiwSIkdTBD0dXaqd0
evFO85zKKeIhENia6b+m9JKQHuExifB4Fpz+vIgj2olnbR0jUWL8l1DTZp5b6PabHNx/ckNChQiU
jVnsb9Gprh0S/nEsPnlxCMq4kIlGfJ5QwJiB2QJCUaCplrajqqPdsLsZgiQxTQBYaXg6QpHIe1Z5
+LtpzMtwEXoof6yJ2bWXygwNHCe0X64ZWuYlouUIQeb1w+/U5Qja51hr0A4/FVm7on5gSba8qA0K
fkSgsiVEOI7+tv0sYaBV/vRkWxpxG2Bo3/JxMkNuznhriFA8Uap/8dFxX3CfubroVhvgoXF+7xSP
JqafMLIVlb6rFh9KSvZCWg5o0TQBvEZuX9/RaLOPcYWo4hhEXuuPbfEEnaHBr1uGzSlog2ugvvf2
bJmM1Df8++iW6bQ/jw/e0magdZE/PUQMhuO4Xbm1TxeABfs2GeZ7p3UhHmASdtAegNy4fKASTUWc
jjyIwpUBDQimwX9nLTpxk+j3S+OuC7yDYMOAPXVbGrJ4wEIaxJOh9u0vwwpFyQo6wEuWAoGumno/
bdFyvukCtCCCAuTjCs6cBlg5r0CBME/c2Hw2v/DWCqSiNDm97p5E2psrgtVoz5pfsXVmWNE57k3a
72OR0UBt9sjRQ0Z4n1LebGxqIwHqy5YliByVK/BewN7HyP+P1EWAmQMh8pbKDURF4A8snpySqxNa
3wZUZui2J1KTPG4eYfAXtJbFxsozgnLgYZSia/gG1R1FE26VNXNaoAgfYR/5HN51I7ZN5NirLV2i
2oRiQ7iZPcU2evJgWCbVW+Ho9NNi7ponKs7rOeY6QRZDngwZRjiD2ltNRcfVbat2qmwJFvMjhsid
piit3ftZzzSgdWOjNtmUmdsmT2wKtqBrHsVY1938yBT69lEvxupAVi5LGeKxEhWxd80FrayIoVYZ
8TyQ958AVku0QciDAa1WKMRXGGXo7ISerPDH9L4g8lp5/GukW3hvdnQL7DD6ihlhxsRqicoJKa1d
PxQYX3L7D1XiFXzPE4p6r97yZnNS3yWcj2qzrEo2i/TgmrBea17faISZz/D2BSZAMgCvbRRyupWe
XyPps8LZ82UMy7CjEvTjDJEQYvsdWeBpvLVqWELuz47D/DfrBA3GiUv0vPeYCJ+x0Axe7BtH69sk
xsZRtnrrle3+k6GY/dR6qq1D8g4mBJU19QO8pPQC+XpwRNRQ7BX6Z5+hl/Qih9O67ukEIfkrUk+E
yQPCb8TIxRM0Z/fZw0Dh3cG9sMW4Z0raaM/IKwJVL5KxtS2ERSP8+aMlkVC8GBKTdXmxN/zWsLey
eMRmRTZBJRLp9F6F7TnMWs5zAdfO9FoqkspHhmZ/kFqXJ34EMt+BWPMOGgQQ/p8TZC9+8mJAzNJu
hLwNZIrc15Vv9mMk0jZZMP2P2dxMaZVLBTpuxH9OvBb2pvrkQSvwAg1KUyG5AXi3CTqQW1kw78WP
6Hzz9hj4nIDTcCzrqMS8r6yMeQB0CKJ5fUdp7P79h9b+zx8qdIL0Z4kuDJzOQeQas1k4S30mjOf1
j23tJE+VVCH+deLIsDzXkUh2WFrBlg4miY+MARG83Mk+m/8nBY7uHl7/hBCOC/cy9ROgBePnTR44
IGBHzbpuqoygF5DAAqNnd3cuudoiJRnH2n3zG5xuz27nN8teF9xnmE75hfkCbjmbAFMMs8srbASC
Ao5ekKQLmLu/QfcapVg7z/jVpUiZjGR910KxrAX7PmvwNNrfPgtvapdPb6iHUj3XPrAD7rt6JqFJ
VDBMQo2n8jN+M7wjE3+AJP9UOqrlG8Bt6e2mRwAfwctJzIC0itR1FaZ4mYbYXmUZB5GQFENaUe5D
gKl+Kf4uHlkDtYHEwax/IXwURrJg/OEntxHnupquYlssRY9qMm/4VCPM/BPtf2jE6DMAtg8/jy1R
LoHj+UcjZaawJSkh4G380pQAgBmR1n5OdelpfxA8Aaga+worxKOqp8xbne81yod5VozYDipZRgtb
jTwnNdwlBjSJwf4QKFOF2jZGdywk4eefmKh1qHOdSEpUu+e6Mlk0koKIGT0xUzMJIxDDqJ5sNItQ
U9aUfMeP3NxX9ePlwyp/QaOJMla/DMKxdvs65TCQPbz/vQfgaVU8rotlbiN9EtmLekOkxhFIZZfb
KCWob9ftu4tz6GaZXAe3j/YHYR7UgKwIKyENtDVzb5Gt1MNnrlj+KYN3Xb5CaNRiRUS37n9AsGL8
7nHUaswu4QiSAtephFFjgOt3cjLXIwftfWCTfAj7rJ50+UmWE9tXK9JMEgArhaHZdgeEezkO3n8n
rEUMdbThMFd9C6DkG4k+u8X2/GcZlnisq/nPgoHPXde5v9W8OFHsHxrKfvmpTfkaY1j9h2C4fQN4
aJokiwAFeBQFa3V5pqq8zggXXlDdHaj3XgapCcFT/xCw5tq7ze7CyNza2fcUXm4pek0EbYH97o33
+dfRU244XP9GERdMCxVXiZf+T9RQegEDQ+3j2jdUmD87xGV7Jv60ZXzMAB9AoVG+iHWm9yZfp/J2
79809PPOo1UDA3lppzUOP9Yin39w7pNdF5l+vuZJIkwrYeABTR+wFXL59txdv24lNohGU+boiltI
gY/1R+2LbXeSVRB7CG1B3u4B7BwsqGvlhVjWGW8xzMqEon6MDnMAtZVR2a6BZ0/7Xkkc4Lba1eyZ
CR9IQH+4FZSowf/fzYeh2C2PbDy+CUs09brQWsQueSCmhXk/M8bvq+uFDVD+Z5LiuBcV2ZSFTf91
PdwM+Sps4/wu+ohHRrGlAj81KXSAT+MCny6Q4XIy0w3gyr1v/hUHx4d0vlVcx2Kx20ChLcT0JBRI
oIuGMRdKtGe5MKHcUvq73sYXuY6lkKz/Lck6n1Tva5eUTMgN8c5hRTxupsaVrptfg5FWMZRh5/4R
T59Qy0Db/nlh6n7JA2vCX06D421Q/WspfvRXIQdhGJM9ToofnjK5o0eulHT2yA1ZwEbujFLgo4o4
WfRgdqgOeA7gjtZhwZl/v/rxJLkSdoR4qo9QWa8wfEKALFTXLQjwC4Lfq7ldAA8j8gBHO/NtclHM
1QRPJom0WG3u4tLP7tdM0dX0d1z//70LHVaTHSiRIp8lsKfFDuEJn5mqh3v2uUngA2QEbIm820eX
vT033q2r5P0+Vex1SYbSv+s9bnj6HNSldBFHE+4XOM16pmxECDDnv1BnWFLPIJXSqknaivsxeh9k
WV8di34Pz7kCXEvnrXohDc9/YP2DXhVWrfQl39ihOFzIrwr2e/LDtWm9K2AnlBUAV8N1KSZCUf/5
Vjg9sExfKaB0mIzQ25J3POG89F2MWX6SQcFG+GgEbK3yvbyZA9QWj9iBFzSrfKwg9fGKjGySYeOf
mAFQfLqUw5+3zE48xf+eN8x4HKO/Sba5Bz6xFZVjK1in8jMDY6hN03ACmvQxz9aGSe4HFhCnim1A
roZd1l0i4j46kDVibmfOXHyqZuLhrs/YEEracC8QrJzZlTnrn4h8r8xMfzfUoBm/syTPEjjC9YSn
UuKMYvDWA9i4rGw5XO3DEHDO4zaD++UmLCVPJGmEKHH6tPDZgCf1YOYMfcCM0A1erXSPPv/ds10w
nZFeKFJ/hGnq+rw/C3201KVew0tAO1gC5foQgZtOR63cbWKJW1v/OTuy2/r7kqAW5ElGs+Y6bmpu
wecbtu3/nyWpJwNq7K4ZExkR5rp3++Qo3T6iuGLIOobh4IKyeB9fchdODPhVdytOt47wpvd73guh
JLqgTabsUehzyGUgk+q22Xqn0/6dleUhdWQrTCRz3Z5Skn+rcZv2ROKxedXODCQ3lAmn6+peGdD8
kAHX3EWIGH1cvUDJJVQL6eSH0ZOdICDBWciFQ1Z4Ycrlj9DdlXLPKbb1r8uROhye5ZUx18wUvBgi
URbLxOlHLnGvm0vvuT0s2lzQRkUquH54wLIoWhy91m2ehqLkwXGgGkNlfzSORi+y7FliYhkE2a8S
yG9VR/dDNtC9UrkSbs1DlMn1auo43lxwjdU/4mm5LTr0H1NWDv5lQaUjBlz/wRO/lolCPpn6Wuxk
4jfgYQUmENmvoQPKgttaujPfRutdOLDKKwu0E20rN2A/xk8x2iuLh9WMv2aqiELO+Zt2lDCtki1B
pV/hBgWEuxZ0M8UEyTPAX7xlOkPHLGdUYaTdJREvtmv515jBQwhi+I1gCD3n70qCuNHcNQg1j7Xq
ot5cBdC+NCFOiqy1K7Seod4MbtB2B6+ICLOeMm0M9lIFumXDJ/r8nMIdhGUd4qr9vuUj132ug5r6
s64Fg0sZV5f7LDk5xbHAIyqWkvepsIvkPSsD6jAKwdgN9J6IuDQXRAaZJGazALBT0lG+kcsce36Y
9hp/fzE66XMJeUKFq7u/F6V+hXEQlHjFxijUE6MXpkF8CCUSsZkeMFKl/Nr0GNtKcP4VTgaE+0KG
mkaEadzQfXbjsnUu1JS8AaQryFwV7s69XFY0+Cwv4sPMvNlCn2FvwwVItb8ml/iW77z9amK+dI9p
yb6d+VvGCayFHvRAHPeQRDMo6ZyL8KqFR1hZbXsBz7+SZr3GDLcdkmbSDwcl7/useOJjn6QdiEV3
WuD8njXWuUzc7UfcGbhsThpP2DLsQySyLkfs3b7kQYQUJ5gtrFT+/bl9/V7r4+f+9YJIIqiV4SzZ
Epr4A0RAxzNEkEuZHHt39eOD27DgWpe6tALeROO1l9I1CKjXcYSZ9mq+PDJcH8WgweovKCGRYg1v
C0TgrJkebE5FyvadZ6ixoLiCz0IXo+c5bAL6iZeJZabV1HeMRadU2FaG7OJjpWFwNH4LV3LcwcTw
vqfuaYetwhD1tn0m6uadatapyhJxiD95ZAqYqJhQ4bd1IFlRAhM31Cdl0ROoLcGGTSevShYy8xOZ
ubQ1DjOT905AQaptbIiA0Fj4UNqzb7oMwQe7g7w7SZ8MtfBed6MubLW7OzM7JuKdP39U/f7vnPbv
/1UAAC5Vr9NgYKK8IncI3f7nviJXuvf0/bKFnLv4BKqjZoHlJzA055Kv3TlraU1CyrWdTEqCiKZl
xUvzyFr0Y6Wbz37vuHK/FVRlbi1ii65CrQd+aJeVIqciRnJI9BFiFP8oAAwFIbuoFDqp9lysSSpO
9ClCnLfekE9co5E1gTrZd6oXYCkMZeMvud363QQRLUXA5pawUmeHRwNbRT34E7p0kxDqkrFEFQRG
ZoGIVki6anZvybTAUHetNlgKXtvD3LBQiO405YyjfMguQr8OY34BiKwvOcaSTtTIjrhlaC/wwzME
A4DepiEjrj7aViMcLTfIadGVPP2tzXR2eQohmTiQkJx/ehrNfuq4ZdeMU5bxr5DmHZt/u2myrKTr
T0XeOWnxeqP6MLSiIguJA4C6Vc6ZHOEiElfkIIjLHuVu2kQYrMymASBfTtMg97XOrAi4ka2nxcyC
UY3mXDQRDrhaabd3mhpSLIo+3I7Pyje/iWM6d1zVP6WmVLlU9nO9Gy0+iXnOu8a2/gIQUZOUSygP
yd5Jw3Ek7eX2/1sionaeaDC7v8aQkPvEGnHvWGs61qwx3tO9Bl5Z0sqit7GUEVgEr5hO/8kXysFK
xYFtOcK6s5YCahSYhZQlNFgnAsK2Wb0HfSAln5L+OgONwyKAawPoVYFPnKNNnT0qkWd4YUzeEHEz
b1sZ3+HiWH248jPmO66AKN4LNR69PLbp61g4LN1WkabdVsC7qHuHyf7rIU85hOEmIFNXNrhCJjZX
2uYZ22/9Ol5qZzQbMi2tC8M4EUapQKnESEO0OhOrq2/MywZeR5BV4JPQO0cxu6PwSdhTkG4885sm
M4+of3A6btbzBYRBZmG3/fGPlLBA9MdVr0rsu6u5FVNqXMX15nZIW6fG9C7oKHwKTHk1RTZnwsie
WbjRL0eNpLa+GvetFqkYWFzlpqp5znX3ikCBmFSpjo+a1sq7nNKy4lbbOzhNVnKsBlsfkDKgTYrC
jxNMzsm07FE6e5Tnmtd86J93MJw2SS66BVaoTxkxVVQBynj5RAVfjxsLLXUd8gIWIHD5l524LIjB
K6aLGi8Lv6FARXADe82xhG3FytymgMWij87ncnibPu88J/A0jwtaX4VJUuWQucZHC/v8l8/PZi8d
nNbvfK0iSNwu3LKq7LxW8frk7bYCFCSKG7e0LEGkbxPKJkg8W1ipCoWn/lpQy3hlSpjL+9orOy2r
mr4uYu90gP65BgTHynCoE9tULWAvaT0DJOMgYyXSmL7U69arH4AkXAUuhdCl70WRuWupvHPMEb+b
fZBDe9TucWEnwhXSeB79qo1v2ausiduw9UGXyK6ddn5gNSw/Qn93K6j9XFpafuqb3Dx5EXDJFK+K
eQSvWG74mFhn3QJv3P+PMZCksnv7CDzgRfXqXOgpd62dv9LNEO26cZoz8fZbiCFJOk6dDysRahog
wvRWfT6eO7feCVV7weGNGrK832f6UgSEE7UZHHGTdMFyXER0PFVC1VwdDA/LanAQjDckiF86fQ2V
TtLHCiN+1XuluLP/6xRJVWfHuYZttTL8U1vfSWqqPT5XXHZj5X5ZPDP3S0scS3750h2d/kall/Lt
fcvHY8ruiUGOAaaMkxlOLxup9zF54a86ld8QnKkfxNX4McxQg+T1e1a3vmkNunR3CaXip1ltMRS/
26wdNM9LIHzwBbeY7jv3jwtOMFZi9t0kBtJZtN/9hLl2BsVaFyJ9TjdCEEuzdH1whIMcqwmNGk2V
Dqv2bmFHfxjeAuTs3Q1MeV97yEeSr2a03rmBJ/MmZuD/FHmryfkS5d/nuQI8J59dgztMFUCeYG5e
cd164s9+lr4dCo7f4KcIqGSe3YjAZzafW4Hf2L8lwoq6so6OC7jxSJbdfxrdIlyZkVO9U092Y/hv
7bDY6Ac3Xs7ycOYOU2rjkm+mxob+/L9U+fzygxzJ6FMcNpkZA1CEcXDkFuWOaR6ZcETW3E4eX3Lz
o/MAb+uWTQ0l07DM2npSQ6yuzDbtq2ZChsztNLZ8++fcfW7prOt3oJPp1EoNABZth4QL7xCW/blx
9nlGNKOu5R6grhTlaGr5dlhxK7lW7CZy8DoEUlJTnPvtuBFrPQKLtGrfOpmbjtPBWPkwSiPk6wBf
murjdKlKGZ9enDsmxRoSbWA7iz1B7meFvtNugST5t+Ough+BqSCwhucbvG/R0l3xRtRr9PVTtBLR
YW5plahznfTjz7bJROpzsHRJ2eYjQTtX9VOuBN72xIhOXHU0N1tRg6hNrnTIctp9FG7psTjP/ABl
VUblRkO8SYRKAcDZXVMbagsXDOZk50XfKwN7LdusB+C6Cxm0nB/sUkn99AeLYc5kZkUHM6ZXrN4O
FQQVCDfIOQWutQiKG7Ff49YSvN9rM5O0WyYUJEEh/jEzZq0qu+T1gtJsURDam7qt9QExMgg9R3Iu
iOMjhI8Yj1DbsAwsqxDKCx6DnRWhLZ7ms5bdHUQI6R9pkKJ88yfS/GaTeBxMeYk4uK2r1FIopywj
XUncDI5dqjZbZXEktW15YfGXKu93Uh7vd1t8toDBolaNtwOm1meOaqNWUvBJskrngjNQDg/Kqmz4
SlzfE9jTRdW6cZct1Ek93l9O5vdJ7OKMqAKPTF1hoezHG+8GuT7W6FX7OQLW3iHG4Q9gHYj5Z5B2
+BQZxNiC3pPguR1wI2+/33A5cOLX+iqoYbc/8W/hmI+AH58DsLgel1wsUH0uNJ1y5xnx0cqC8HI2
gBvnb4rog9pZbBS1JYnnJHpXSpmjz8ROs7ztpaB94eRPOvhlFGpn/GjKDOLYNAmsZ5ERK8FQm3ig
DUWZr1Fi1BwO5cpjJqKtaU58xLVZ8ooXMbAccAp8w4lQcOL7xZmo2NoEHU1DXpimGBaVTxEyOOpz
k5ODAqRmT7qm0Ffcip9WJL6fRSa/0xgN/2CzWbDt4e74QNcrrQprkk63emvdovBpUvhiVPu4Vifg
ij+PUkk/D9B6w6ma/0cx5NBUQgDg/KctXJodHs8sTRV2rkbspegUqzXmUwkEFLn0lq6ZRNVcPnuW
sgxvRpFto11nvNgIfhbmGJL08uaJLzYhnhX7K2PLCFYsy7PxIHkFFmyrxEYx3g1brDvxKKfbKACp
xdAZcnzONn4CngpRcnDcxjRHEJhf+Qz3zVXn3w6aPvxz15Mj2zowtqhXrsOsk2/Vo5uN6LZGpnkF
askIQpbBA/n90GIXw6JJJVE+wWVme2hBfTigcjsA0t+FOlZM1op5+md0MQr+b5DQN0lqsSBDVNU6
ha7LyTE8F00uEvIVUO4m0X1vG2BNHr+9DJ6VyB7HpVCtfrPk1ruUo6FOTIIdbAwZCZK667G71szx
yNJXWKeWGpEyhYSB3jg5fLvB2KwZTWtswBKziDC3dR/iu6HvMEqnTO0sZA6hHTbDXsJgFiDbpBWO
VmQqjoeRkKTYLRcMJapWY8PUPq1/g1tbkwEHzkaZrwYSJt4NrjSneuEgH+61gyyc5pRpIt9kRa3A
Ydx4oRH8dEzKVPHsqLlje7sm/SfsA0xbrs3+vMNYirZjP9Qnc8mAJxk5ALJD05AaW8/tX/R9Fwky
/hbIooLkLsPCawR9ojwxdcMCPJpTx2COSkTq/PDeQG+gdewGuXCS8Lheq4SvKITyci8VWtoKcSId
Ph/9iKj5W/jd3LuIAm2lw0cISCtYfZxsL7Eh6eRkK1809SnLVoUm2uydM2GFf5Ky/arVlqqHvG0z
bIUUJSud5eahOadJdFH4DEJyb2WaBV8yvISViMDG+9yVVqda7tGaZEZ2v/166EG/uxgjeh1+mXvR
8Bpm2CWKOi5cEn5TG1KrnzP4Ot3Oa7ZdVwm5hl6wJ8960Ap0t7TKxHdoK1sM+qGQTM0Md4Rlvke0
cgwiXstCTQRPaKakEHLsY4Yrx/tYaK+6aMF35aeCEQOOSLO761l4kVWrqkHzYnpgFA5gkHbSUGKp
ZfN9YXcOJDuf73orZ5u99jGy0XtS6Q46+xqFt0gBsPZP6pOwiPdlFIo+4Ro5yyrh/HWooRH7Gv1c
X2W/kr+eSnNxlPKp+B2IYjiE0ZCDSuKTgM9wmTb9wKKwHANwRqbOeUSZ1kXCrF61uK/zOvX2RudY
Sc65gt7xlFVKaHc0sR9kIcfww4m2109xSBUgb+p3nVfSwu7yAiJ6ty1u7lQEj6ecCq5iXUOHGIjq
j/1VVi6gT5klqp5bu4w5gVUHpC43kF2DB06UHKf5xFvpb3haKWCUKapzLYecXdWO469btyOO28rQ
4TlGOKXml76B6o9fqLRvQckjt1j/VsC6Ix7sVvWdv5VhadCkI9k0nYR0xoQmi57cakW+AG5lwFDK
/r9jm7D4zuoCRCJkNyfYuh8cIySIK/TE8507dGT+0uXuBOAjHY+ax4+c66mD2fyiLx+1wJpSoxaf
gtEm2j+aisIhslqNK8fRAoy6qEgL+sDD3bzICb9JlkeS9uoV8bAypACs8w7UuO9najCz53duCbw1
Iur1MW/Qxu+jmaSkkCPYdLNczaaSJIXqw32a0PWssTBxAnYXMl++uPFpvIrJVwictdqe1Hjr/U7N
V2NmyRRCSTIidH7/zspMYzTqfj2/My8CpZS934WrHaQuc4yn9MRj+v94VNw+hvOPlU/VQsGE17gy
3H4eZNne9/JaVUIEyMd2duSornWykMcKX8ZQqrwoueankqDCvU8TyBWH47bWjFd6cd99la2RW7vG
hYLSciWiQfSfcQFUD1CfinApu7r904QcQGn/JYdvVK846FdSax/2ALMVY72+kMrEyj4S+hWijjIA
Gs5JE5MoZZCJcvXF2O1HzsGpgRLe/7XD8zUJd0FkZUJbKXCXZh+TQkQi1KhfRQFkqnwVJTKcC5+A
T4F6+RdLnTH+kbn3nKhDG6pXPo4jbgIJZ9E9A38myCnm+Ll22w0l+qS8pmfOQJHH8aJMXYg+LTMX
cex934WxeYw+Msn+jBG39LSdNpq/VqOhjDCyfpN/JjLi70WdkclsKyunq0azIrmK//ocuC3T5lQ2
FWXZZdYW+K9vhc7VBKo83Hu5f9YXwDNAVHiTD2lx7v2tURXfG3xF5eHQrxzvrLBT6KDL+/ltPAoU
JwDXBndOaVYnzAswCeoQLMk/9lVt67XlKKhuJFpOH5ehNp+VqAm45XmiqYCm5ZNG/lbk7e2dJUUT
f4sqMD8Oe7UShcysrX89vijiILpQkq6DUwMzxb3bEe8zE8QiuBWvVzcY2QTVvV3AzzR4lKf6hyng
KVCWAgVwM4lSi2XVq8L2NOvq/9kmEORSv2SY28d0V9BjRzfx9Fft3Inw4q5/W/Rve+70sttQkyar
GnMmWJ0cEdORTMQpawV7XhhILsH5N4BiFUg0RCsosirafdrUWpezTNrCgwwNt1ONXB5vNsUtWIMS
Xc9YnheE6d74dCUPR/da+KwoiUSwIMHXs4ciFFfd4n7rrFGYXoGfUiavgCwe2xNOV/z40ZXyYkP8
u1jbNHLnhQT9515Fcxm8P7yYi7Ki51df6uuVw5bOEeBTiMNUVyKOLri8pYNiwgPi6UaKflpCCUIt
tWiVSG1k0fmsNnEz3vm4vZhgAGnm2KpzgeXVvTFjfWq15mJwu/i5aIg2Soru8KPzN4jSlcqmC4We
myrJmPEkm0AQXt3VrKwStZ9O5eiuia8FgC6MNAg4QH0u22qJhP/0pEi28cp9AthlAkfuCZ6gKg88
WFgEjiBNkEsWXRa3GDjlX+1mtW2ErWNdNDVml5G1tv7vxwQBWE7Tbmf8Gw1iMKV8I/4UjqKm8KrI
JdrZjii/xGoQoP5H1l3bVEO+lffnYYg7d5UZ/je5Bct2qzCeSbJO8VYCBEY2Jdz1jRgPohlaiXY3
X9ajs6oGa3xHrQY/uacj7/dRY6MRJWP1J3n8GP/5GA+1P+42darAAxdnyvziXeeAI3kuiBHqWHB7
kIJXiizuWpakuPqM9quOArd6M2w7mnzWbEXHJVQl0KPgsgyBkZNTDd8Df8VGyEDDvxeK5KWKMBzs
+NfR+aKJ5P4TAyfWh3iGC95+ExSVsbcqsf/dad6f7aoxv2GE3g4827c0CJjQ8aBx1kHq2tsNwr75
aNoqc28G/frwP9m87ZqiZFe+N9Bvx6QzAfbojHZqfjm8NxfymmLVwATRWG8DVGgETipu9CKjG43k
81J1gh7BcxWVBOuQ4XfCkT/FLgaqxIZRfsjOWV1SK1jxaTcwCrnMpsM6N6hyhnAnyCrjoPCQsrrS
rkCIuxeEcfAD7YOuKPSUoPnF28A9KMm04Md2FcZpv28cH4vbQHKJpVuJDS1+3TKZk4kyuicOIxvR
uny3ChwZpXgrvx5tkeLyzowdovbT2AQrCmeRDgSTwMOgGy/mjTfJ9ZE3ObzlJu7GbSsHiMttPngS
DA9nV4iAYr6QAjrN+Z308k+14oT6IxER+IgaRU4Wq4JRwNqWwo+FH0AilQGWHjLzbUL1+fhSkp81
HCiMLplHzfC9vQCnzm93tZYPZ4DdDLqGz1gG5CSfd9ZDyL+mXVgl0DREUclORCTY7WStKptRRZYT
dQ2IOEqoLOTwKFn2QcjOrfBIf+yPLzD7QFbqtkW8DLcqCMhWAhQ77USE/gP6Kn9S89BSlf4DYFgu
CIiiiM2xijvyn4av5eNGzNeREB9dJ7siN1tZ8h6NUhr62EO1Z0WwtKirJy+UEBsWBoDrH0+4XQeV
a4dFVf92k5UH6/kR5Qi7wz3vFZvoG5fi4UnS06xhu5wSeZOZ4aBAgbxaggOnnQGnNT6dvlhQInv3
RYvrJE+XguNcaIZRrpDYE12UVs0XjYDKyEVOFNi1GT6qXHofaiiS0e0xSsadzY/IFaNGZ8Av8hQB
tWz+7P8/H92Uwo9WpBuUpUCfAdswgKJVCqH9gykQTkdpYxoHf5vF2nATeUOjkMcQXJSWYUivSQWP
iJmyvBcFyC26U0N8WLjfQzpBgrAXmhaiJSnMimWStetBTYV/2d4z/ZqOYCL/xUGSXjqIf7erTkRY
LRyb2Fakom15H8HP+1fejkURDZeHBmC17u5QJ8QTVfOsnjko09O1A3SauW9AMa/eSfu0zRPRUgmb
hUqJot3qr4akpixR/wa+xb20XsePe6Br7dx5E0fKGYEYwvn0L7DlzsRZ0wydx4zb0r9OY8l2VbhE
O300U6pBrLKQ1pbIg5btNU9KeAeA4LeDtbB57fwGy0NHc+8wlMSZ6zKjjwDG1GaM4QIB63GGd9h/
heXwk+cs16TEHTDzoS12BTB7WL5dVcigDelXZ8JPInyqe6gZir5CtchS3xsFhCieqS2plyLKhDW+
nl01yXrf5Q84ynPq6+FmUzN3J2TvDVTBp4a4ZCIbHr/dSfza1VTInf5fr8yghaJ/mIOHeHTCOKNX
b6tol2jdQpdiMrmvo5WwLZgK3wdVqhk1JzG9wVsQuvIaKIxfRRkPJZxgFqjkA7JcqgbWamYDZc1E
XsLfvuktljFliRLlT+yTOGJ6gnwwidlsrkvFjiWhlP1TcXV9efKP93QJX8ui6/vbCycC9fz63H+z
2LFHdk2C9AfkoBHXRXkPfIrPnyJ0f3H80ySVdeSxO3MSIkpVn9z/ah4R3Aen0wePZvOSLp4WLOS5
vA2Bj5egXsTlH66fzqC9ID9dJlerFZu3B8BVcINEqe+DwnNo+tRjOgGZ072nGQSbCaldkYkHNTkb
GqPrnarvIGweyFzE4m+LJt9zRqzBIUdm9w6+U03pElozVdgNl+qDbeG9zuaRurAEhjWlOpxVdH6L
8sVa8dW127ueM3l5Uuqtu3cPy6TznI3uI0nL//IjrhwbPG8Tgu2hYATi/cTHq5/TK8f8xMuJOIU7
EVx3vfYuERivh0NIjmIFcrTaOJlreaRPDUHJjhl8RvOG832l5fj3DycIj/5u9GDTRv2PRq63hnkJ
bT5TPlVTJzfTvqKKPoCYHKRpHTUW0RD5b6M5/NPf3lQBbcDO3urb1KJLOHlHCi5JzaLnTbM+na+I
yQGlkDzg2ybu2Og5N3g89xhgprcgF++6rYbfg+vmV5NDFhtuoztsHphzUOdn8Oao1nM3UkGuGxJW
feG7jxqz/XHAVajtqqnt2coLQT36TcBBzugh/UJ6mbTomlbPnBB9o0p+67ekfJ0OaaXjRtVMBiYM
/3iPzGXjuW3gb3vBBWm0pwF6SEWOOWjkGQqD8dlcWuAXWbaj6H9vCeZIlce6pfMft6mKS34gDVnI
ct2escRiEuMR+y/zjCJNd9Sl9eCK3mPY/+Bv/5D0hE+YtDw7+CJiBZZNO9aPfjERXnlkIKcWJKus
uWy0nYSXldOPN8LyUBETJmBXo1PHcj2kVxnHLheWKvly6vre0qFw7OoyQa2OF2JpRzePlvYmDxc2
u8+903o/cQ/XKwwi2PrLgzlrkoSegBF6DIoze4b1aTQc07OFHG2RQOaq/tlQ5W1VntmgycC8ZxRW
27GnVI35diwem+rughHlKU5ujHxV5VStlIPgfZyeURXgmCCG+nowgygkt26uAfK9uqN+7SaRwFqe
gnj7rJ6Wz+nmxPCY/ma/L69D56VEvB8FkhnSuZ5xriSwL6/krMu8gjOcgMjqaC3mqFNqpmobz+i7
Ce6flfN1Nv296M5Yr/s6cpKWy9K2VnZzpVIP+3O3vxCce0cNA5sXRio+r9XVWfd1SxTb/YT5DL8l
Cb5XHFJhdK4lWjGdD+GllHahL/Y1SuZ6ZpcI5MQaz/jqt3ljXg9DejB3YVZ8JMybsq4DrGNXwtXT
d+5veSgcO3v+Ul3QWLZZuYwJpv6dDX1mjkBk9AvM4EpIqeo9fWNGEb0ESsAtr8AilEXDUsexvnmx
EKYwk0i63CAvYxAw+oNxPyX1DbGQbqg6ksnazvdVkECZ7VOTl1b9dKYZwbbke2lJE7DScIJEbL6P
a524GCuLk6T0XTUFic0NSzVOnSEnX3TfkW5vgmZwuMOHIafOnUXbRiMU5TJGNopPF4Yx5zWaUbn9
V1uxMKlCxmOcNVk7hngaRFwJL+X7sEyXxYoTzAPjznrQUzbxRdgpe7UDVvF9MqXGZOZKx8Wd/PBV
BfwdhHbCOMQH237ELKQKqP619V/YheeLqPuAnDm1b1xSBE0yMEb7tVfZPlONADJNH0U2usMB8xgE
oyxlaSlINWgA0qryyQJ0OKxPB1uLiOtC2o7AHAHHZIdtbWRvjuO1YhV2BMLG2pfyT8ryTSE8qnLb
m23SxSoYGfbDEKy/cD6ql4GcEky9IRoIhc7lL3mjKl42R8TgmRtT+gmclekk/oeyQ5vYxdJYDgDL
XjtNssYMqUY6RzaqsXIIWEjnyzZZL8UD+V+vGBKvVJmDYJ197ISajNL6ts0zqVqwrKH62o9V+Zfc
uR0BzqD2Yac2XbGZrti5j7tyzIeHhxkbItTGqTFlNNFXgPUOKH6ERoahmMTZwvbQLGyMd3vpXAg9
bO2Oay59lGTNUQ3M0Es3EzEZN1ZdD4/WZjjHogSU0vVzxOARL4lRe0Uv+/6DsR0uYjcbf89XaHpu
Y6I6p8I/8lirvh0DyYmGahwEbwX08wc3rnUIv/hQrxtRtYgbT1ayWF3CMWiPeRP+Nifwrj17KAOd
gQmk/bSS7s06er/Mjp0MUC/uaYU62aMKSCk/qH2DhF0heYav2F1SDMifmR/VeL6yclsfw6bjWBmO
XVGievy5txzVN/X1MHwwoHtIemZsnJllxZQKU/N9etlDMLLE0zGF9YCv6/+ntN20ETpjZ6MnAIuX
NbcrkN6OK89ARBL4Wa0pTjCKBWiKZo8a5KBoShMdehNc/3MbIeK570o16+ZRKsYXftpxk1e3ubdK
Zde0oFHtfRetPpjhhHJbg5SQqhNeCylD5xkcMDnjhk0tneGDT1pZ2gXVHLo43dCBVtWvUFgZyYTl
qgTjQ0ig3VRSSuBe+QZamtIbK8ESFWeKeUtEA3Vlyxi74AyqLjDK/u+f9fGTFud6Ao30F0PQ6cVM
kkRB+cSwvWV7c1/C5InuWxtVoVPmkNeV6pEQ1pTQ0K0IntQIZ5Yo3oD6LV8LE53UND3Lgy0wr6R3
b6FUBGXhMMShTSMRN87Xlv3rSSvWrzDMdU7tJF7gtehYQ95Il5F6D5KVM0WCglYWXcLQraavrcXF
mYYRthD6xbJ9qyD6wxH4OK9HfGJD/LEeK4Uiu4ogu8nU04lZFRfFzRDG3xDGadbsnrIOXkDImq8C
vMOMVj/QLvFEyrqZCW+5/VlYV5j3wt69eT99s949Pr++d6Y7cx+l++I97FKfmj6nj6NDNt7XJKTt
TebmE5lnujTc3/6G+VjwBvqVkOJ32Hg0tMrK4CTNdOxKZa7CfOnPFpMS9Qs6lik4MXyzRXEOxNY2
gRPzv5SDPyk0T9UXSudsTnsH915D5IM3sKzcCQvcjW5ns9S86uyhQKFhTKm+U1X5TKr+Hli/kWLQ
Z7y+9+YjIUJDGQ2lV2+q4iAG3MTAi6jlhFFXVUSKaV6GibcCI4L7clsp9MZSQNAllbjdVkaVu9bR
mIL+5VtaDc+a3iYSHk5btVnBAL+OOqwS8Jgccl7H+D9vrBVLeslC78u+KrfnD3oj4omXRA0QeFkX
Q0GybJiU45h6RXM1GvGrkddCFqp92c7+FrapnLesBkdEUEyJCjYD+WphgjpA7fgsMFNBV+Q7uFfl
cI2SEWRw835Akmn9DkEWdE4IAiXQMfXV4necp7tz6E19xBkEVXDNPcEVhSk7XsXoC+NBVdxioO2f
eRefJ2fW/3nIMv3yFLZF/aYWzPvRYBuQNWXFegkZwjZhQqjM0dgOHPJvpSSgNASuU8+4nw/E7OTx
j1jnUzUhqF5Y+gH7Xyvfea+Jc5kNKVzcSC4GbDc4NXE8q8GFtJ9Q/XAqBzyzTgXMEjUyE3Vnjr7W
zjCOdr81f4mI4e3umL6lbnXyGcgOBitTUixkqydful3RmDUfkovdJmdAMDwU9dobVvtx40DIV9GT
m1QQUa9AGS2PtBYOE0sj5ZiFHoS0BQ0x0xHNu4NRMx5h7mubfVIKTIteCOwhymRuDE8pFN6cfs8n
I9KpzQGe87cOep4xBYSOCmAyitNmSWIM1JYyOKCbbYBP95TcIr3s7E6db19keIIcW8z7vd9y4BxF
yBhcj15QXcgIcz9uFYQmDBZghCI/5CCAWH+n0k/I5d9tgXOC9cbU++VvaDnj75aThUuAq1OKacOg
ympDYDBoEj7qBikzjIvgGuUSS3bvE+D1LK4AnQ1LcT86puRleHUyd4p58Lyx4buJ7sCgwCLt6XRw
9WWPJ8L/KMmKmVJQCKM1a7kWO8l22iWpVZFbbHmmf/zFIy4/yWdIPMEaJ7kNbJvYuFJ1ZrD5daOZ
y+3idPmOaZf3k2LJgHeZbu5JJBYsRtB7tshfcHFew+Az6tj5FYPzlMVC6yUQpRgrgIGdhKy6RHzk
u2PhaP35W+png4fPJI84eb3dXj5FQsLpjgNRd3OLvKNGzG9pgCllQDfeuqb9dgqv2M04OHiu4jms
+tRgPh/Z5SRJVBSlhHYSiPeorr5RIoU00WJJI0efwJhuQUt0ZGQKbxVxvWFKGXN5sbdiI51Lb2Z6
N8SBGUxl5Da3zpV+wl/tFBLy+wqj2FYJaQyRTFar54q6vC16xrpQ1bnx5040yE7jlesk3G8pQU4l
u4wwMjzURVxXmEHdVnameZWoaqQC3hhImHKZ0a4mJMC/zDE8V38u8rR6Q5F9bbenfdV94V2W5MR5
P04tWRJj/in1zs04R6LEqErubK+UOiuPkT6LK6U9iBxGnFviNvV6qs8TbKtAt1hPYFRsAZd7nJAd
EiOzH0H4vA+YN2kz2jRpp5/iDN13HG9ch9pxvzmtpEm8uJifUbcw04Us+oQGJCd7JssksSt7b5tY
o/oQVirZe3EeWYnBb/P+RpNeBmhIsCmQJon28Y8TNPS3zqwSW1akCGNqFBV9LYcy5Da6rgfiUgJA
kuzOhbOHquwqy2mkaCXtt2LmO5qNE+tNuf5ZLLSN6AvNbjLDORWG8cd97ZCTbp4KFErjb3WoRbGT
7XWxj+G/jUqGO3fWg+baHmX/eF4ujHwqmvsF8+JjjpNvczxz2bDvypWFWFxBV5uf5E+zstLQT4a1
qB9BFm+3W428h4SzZlJ9YNfj/VPSj5BuFlvQu3tEeZt0od/GxdEIcmWYazH7iptdzsNLvdFfWClK
bodjSmT6f5KeqtT9W+wIqoFuIr26dFpmLATczLdyV5XxiwxLvXq3QjHXQqkbHc4rVZ7iel4ERNzt
y5MoqpoOXZpuFQ5ZXN4tyWCflw85ObnkEX8NZx4tx9srQcpGuGaKH572s2LZtmDL6pmMzefvyUzU
2prKXf9ZDc/XB2tPndkIrrbnjiBBYTn7+jL/K5NT1M+1im33HWGiNTomBDDTrhcwfIxQ6L2Q+WeX
KjFubDVNlu5gJLkqA6DYkcUJTujoD6UR4jS2vw3vTuej7G4nGupDe/aj7nkVKE1KigsD0nLbg0S2
rBAtmF0qJJKVmUMG4ZjeStveX0ocYNfffyGjf4q3+6alcPBW8HWyCSnkZrOrQcTU9LoGsoI1sGnn
F+RolX8Db/DyvEOZ0uoRyfpEH7QP55HzdEogiuG6Xdj7McP/tvHflH0UHfslj2RkMdATn3wdA206
j6we8/gZnLDnot0xbxtX1WpmMwbadFrQnGg5d2B4bvKn+z/6v3wnJnDUKSql/YnlYa2UVcA9HIGQ
AN2LBhY7ZdEbCDr1Xg/FQZ8vTkDr0E/aZjQmCoLG6gBOXqR3yfjAI9iC7tVpc8L4INMZ2H/H77ry
emZJ/qAtCmUmYFQNPu1prDVdO9BkskkRB1NcXAnrmRVMNz+XhMm78U/CMA6F14qRmltuW75Fy5aF
Okwy9jSUQhJaQjoPO9RrkIrsJIVv7XCKoDOsLNK4SB/0UMrPD4YQdOdAF5qeUL9BvMYH7bPdywH0
64lFV8dpsms1d8t+5d4Rkp9i1xHkw467FKNNxOqgQ/CC2KICtTq6wqKQTIYrNEP1q1ETNOeqqCQq
MYmG/2FvfQSjULw3siqUjRXyzkXcCMkY3ckW9iVZiFgLsv0GSa5KOYKuMDyAYjkOLfMaRZHVyYVI
ynE3lpQBtwyqGzXy06R8caZOa9xgXR/kNsem2tqnCG/MyDrlUApmtWvcMC7cSurTHfyK3FYCHQXJ
gCQAi89NsFk9qQVFj4i990APpg44dbEk4kbksyeSalFbOrT/xJribyxzuvaXYNk34Zhjz1rZhjtd
Z+W/oo/ZWpnHGjjt/gs9cs8tcF7Iy+5tLyrzQT/Zs04xDK2VFAseZQ9teCRvZfV7EVpC4ijeBaMT
JRaigghH6qPzEkUlaNAdYw8IYQAMc9FkPs/SX+q9USWSao/Xm89z75wI5qygAsxbtepE6+WBHVRM
T9mKgbzZbiopcPDbygvSRZrFXnygerjCYnCzZ3xScJf43vUIq3XPeM2Ai/G2Usc8UwwURIc0A1IQ
rtFOIYDGOQRxlBivPTU+KrjMwcUSTK+2rOcuKpoMSrrz/UGqs52uCIO9ilTcN5Mi4/Uc4JS0+zRq
1V93PBwtwoA9DUxTcZcQUMFTiukokKXMDwF5P7zxTpeW07e/yEI1Aod33BE3BgcJ4DO30I083Nsn
VV+lGWUuzXtFg4VX9+zWeqqxm8cdeZzRXRpABQxW+EhgTyf4VoXRQXKo0QaOnQHsLmu/5NEc3MyK
S6ASusrOuuKNI8FhlvT5+kAw75TSIbma1JED69FQp7KGC+/38lOaPgrBema9MDctMebsQ4IHDuQD
qCU1M2U9eo3r+96aTFUGOPCsffsvnKccBgqKIITaCA/3nVShXE6Z7zhIdXz8KZT+dH4RdEg52HhD
VWK371Z9ACh2LnvEK5SqlsGlSgwN2gzJPE5GI6WMyunwmH62hYJBiyUtDZ/d9yVncsn7TBb+h5Vb
qXGstvHcUPjsr8YZ7iK8SXNPanZqh75Mk55k3snnkkzMbFCH+LDGlpkG0hFUzrHBqP47LQq2LUAp
XIJ0fQyOVJj63UvR5ymJ3XV/WJG6OJe2hc8iPHLtxMRs1QBaLmtJE2//wpV2pIxaR6IbgDt7963p
wSsVVQ1qg9vf2sxEjU19FvPUn+3EwPi4uocDrzLHn/pOvIto6g7JGY6b+t+s4ZdvEb5xzTcU3Xum
TLi2kY2SRYb1RScH36hnldOxdPWr2QlswGcKRYrdkeLelWm05UYChguE/KSJYAsrNhIRPDjuzjHp
Bns1vube4dA/6az7g039x/JHvRhNV8hO43FAo+ejxp5byBLcoOq/hv8+quYuy9fCYPXwyZGxpZcS
4VD3Qv9XeNUbnZBzxH9PjcPPw4JMFZ6TYX50Pfg74ZEPfBtroRo5K8ZCD9Tyg0+ehsyWP9GXQY9h
KRDKIGsGaeYRAOCQbHa6wSNV/iDzufqZgl0b36RezSH+igULhYkTIIv4D74wLuNfcwnJZPgA/+M+
rgYg6XEHCOwEFkyInO8oHIw2YLSJtckRFMRJs7l0o9GESFB9pnty5MUdYTaNXGwEgWZeLqaUUqn3
B5ftUcel5k3qNBVa8VgYRIfSozSn6noJJD2qbFdQ2R5HZs5VV37IjGSFz6FDQ7V/E7DkFOjXHEoB
w3McdLcLnoFspqKg5rX72d6of0z3MlzR8y+hPYPX4jcoiTPQvS3Hyod9T/gIACSreRJOWG3YXrYM
HebXNnwa1+1xB9AkijlxbxoodNw5ZN3aVKlKuDD44F7WEJIaUuc9hzHkojicnkPzKjGC8AGckA6f
0zbG6dngprw88mYYYQw7qCbRcLuWn/YfhT06MVVGIsQKDdwORpTZrZO3yEQs/HBMrb+riVgOgK5P
VJ0A3WxSbL1z0DL3AvlBHpsQ+FDji+dnDhW8cFjWUHMuAcB+xsvLfmZUjBKV5OZNP/Ir56BqNtFC
xsuJ/19lF/1tOhT9Y3+7o6iK5MOvdmHy3KxQPqyzeev0e74YupVnqSHzLVJPViXR3657xt2y0sB+
b2AfWQtAI75s8GARGlp7oQjxtRq8lNdhvEsVoCfIg2VvJ3YS5c5Yjr1D0fwX6xaRaYkTkzhClDL9
8+wO7sd8B9+QaH/Ne5pkW9XHFkG4Cyy1yt3vp0yWKC0Vk8nHDWoBfDsVmVJ37tD0XtfMsIOTaEcg
H1Fb3EzbuyDA2WQ1uCCNM7bZ1mlYhJpgDhwEZY5RJHU+gY8IoGrbgdpNy0GBeMIk0vhcYUnkJsmc
+o62Fkg2Y/9e6UhSU9FNhKVH8YskTv1HTD1xhKgP+wcGazH98X8t1XqAmyDwEbrt4Xl7cNM++Muu
DnVW7/i97bkaJxuhALfQpqvJb2YMIbitA4HdSAgRgAf2XSLDAgi0NqruBTe7KobevJVvL4u8P8Yr
P0RScSjm9rfdzTql0XCXaS66WYsOJSedJLkzMOu+7wQP4KdJ1quyrzzrKXBdq3oQHaFPmwVLzcjw
SYqWSInRNmPOPoaYD+vnOrUzushe6PPdesLGZtCJwU7mPvAf0uXbzzYsXS2qOgHt1ug5JE0VLk2w
PzSFyDYC1Af036hMDR4LftjoI+qEe6BuMZX+QN6x8I2VIBgU5Nwd2V+FN+prhA4Fxb8Zjx6uubMc
3hX3MuTwvHfBbmp2kNP1qq7PhZmH08lDqturxXbfOXHD9hXEuy7qxBxKH3BycH/0oVdOFcAaNrWo
9XijGqJYe4lE9bw6E6OB8jCNc8PGCI+TKYT0MJSHYaXDNhg90Z+g3p7bdtAfYUk1dVE9Xayyijm1
kztRWhdqm1JhPhiPs38U6IA5o5e0F+yjkHsxfNXlQQSFBnsI6qj2kacl5S3tXGTNJMJl9p5xVPTX
oX0Q5IeirhgYads83Be3KXxUMZfVRyAG42A16e/wMJyspqgIWJ0yDpzN7OYBpWwtrwxvkV7KNYPq
DGZlYfNgelrKiTwPGolVkWRk7ZAfroftPpg5L0BRTJv7G6eIqG8CzrXDlB0OhNLbv+p59/Ax/T/5
737Uur9yeRvhRqYA2Jk6GS9wqNdLWwbj2vRAENFREi0OopDb/8YQZRAIiqLq5ugptB9xdUGhTE5d
3lm8LlAzM6rNmedSmK4wUD5GEW+Mg14/a+OVyVPfTZVCEkG1Zl781BjyCd88PgDqlV0GD4fbEM7i
gFyUaRrncNa2CC/ms1or5GAhd0t3X8tST9Hc90ChLS7pGybRmFb7XIBTCtP1idpNNBVrKn1/Nnnh
dazSoh0oVzO1JujoK+EmUOg+YV4+SolU3bLa4Bcni7feqqqCeYWvq9zctC2JQFWBk1018IBqrsz+
T1too+7mQE0GfRFIuE7aakgtu8+0ERhxjaOf4BvQ2jKzNtCXqXBLFoU4QGnE5lc2vpFXTL7jRnjz
dlTIskB63xrlKa8V3hT3p0+83iU4+639EqX7G02OYzw4SLVjkxN1j7OgMgC/WaQniFq6qSL0fSGp
TRfA9YN7nKHT5IgaFt1cc+e8Rpra43cY/UpDliEAT9Ps4lSOuMFHaE8gEAIvgg2gwYNbTVgMxIVc
YvXsp0PTlHYW60Cy88TMIQ8UKJhKB5jfA9FAUy3g3LYsR7YWKzFBgpH7iHxxYPtVk8kIdHGjb7D7
BQykjne/gy32wuy9LW0BgiX8/j6LG3xTVCTHMEVMNc9M/59dwYg4i6SuIAYWC77s6jzUZqwYlAJm
FdabmVFKFb1Zv4Hv0q+1i1SfqyfSOK/XykVZgYrptvGjivlv3YsVt7DTebPho15jYPYvc6EmpIRI
75angi4CmgpEEfSWmPkEhIFcAMeNRTuzqkQwkU0dlM7fhtuN/nBwiLFO8MpVRt6MDbPDE/HHjO+I
EFipNlcm6mJi3MYz1+pT0YS/xaf0yBwMikU300l9ArxgSLLP2vPDMqEBNPy+sgv6CzXpoHhd+6uP
9u43xVZgPoFw9FcC7vskYvxIIMYQPAQC12mpUhEw+esbD+xdzoi3m/EOWZHRmHQMvO9biUE3iU3a
42FmGNKcCbrviAHDrjlORI32kavJwtKa/t/3nc/8HKe7/mmMILxojrdY7Qax8t1WRt8g1vWmQ1Wi
0HwLUe62b0XgXMFJEhGAuuj62iPCqaMfOPgIlG0TR1JYvmieUoYJFdlzt9agu9MgTkb1kFR2gNTS
8Jh5jCxJ3rWr06laY0T++R2NZA21Q93lNnq1nenHJy8yQaSJmafBZkIXQPEQQEqMXwVaxO5DRy5H
ScdP5ae1Lb04i2UXnxYd/WgIoPSeqDTFkaUkVPl0e9zQgePK7EI6Kyio+t2ZRdN1KQOxIcYlsFYw
BSW3HFo5/4vFOVqXe4+YvYuVFUHE/oAky7tjRmbQWC/uwsmkOQnZC3LaASloMKVKP8V0aFQ2n2FH
Wk99jCfYJwuAHTTqTYFqAJbhbNjzKo3Xbx5TCfwAhmUbEgwmVgNkUmbD63Y59aCf4gF+1v6XqGCh
39OgLt1CZ/GJi0nP619IDoZ5TDqEOOwjoaQG2087UPP0oVZaGzTdLDtZkFWwY8j/8oo4wK0nS/ei
nof5F66f0Qts5KnVd2ralTB7pWk2LpWRj1FRGCXbW1c0nnbwcBOVO41JgxvqVcqgcY5CJisURfCX
bNv2Y+7xJIKOK7RlBgR0yZBU5x6ElmziPIE8cwsEUS5PqhKL8I1C/lv+JRtuQgCaRe1BAYjnzbf/
RLVQ2dZSEJG5Tof3WOGtNVrhCdx1mGSnJuqXbAWQ4IedFdhNEw4q9F733kPWb7RPg6LPuW4UVeUG
a9Skosj60/kBhaRaBbNTjAt7xZeCDg6YuBJhbkdduDziHmgujtKUSCm1WbWhyt3UhVEzt88gH+pW
66qiqoOfo0S4kJRIc+1J4ySu0KgIQyt2fCvi0vzdXmtkE1fzQahwFeyrso5Dlg4XrMODmPmjOdzw
OQdZt3KLXMm+rcZ4a8owdNQb6iumF7jFvXXJ18/ovgeYA9ntcqO74Oxk4YjFF6ztFqRM/1L6mphw
kPU5aviBe1EYTMpDtdSvO3uvymtudgPPPPVcenTFdwRiccRQchR4BYTkIUHlzArTHJdMRiGc98r+
bizVjcnAu/RVbzoKOAakbj0cFRxh0mBttOC8oKcDy5iTgEulBQ/VxPA8uL3gomnP0A7QFgLnOhYH
h5TaY/9IcXv2sKfhuDvFcJpRxHtMTIpb0h+MN4PgAX6p3ETVe8/qex9S9s80gV7F4vnhIfyH4bfq
LEqPb++Tf3REvlQOEKOdrLGdJ83iO+Davc3xKy+RBMBbE94+FOJv28IksF4s/5XAGJa7x52pgcAO
oFgn5jkf3uh50HydRL+hXSO4IKYmPTOy9cTKysLdP1cOv/mzoNWe/PHcx9hOQNljgAl71mIv7d4V
V3Jrag/QRGqwNTGu0b8ixNyD7W2ml7XgXeBT51wXBLDAPvsiVYtrDy4JX0TGIehGHEM488LNH2mJ
dAfP47o9D0uvjuOp3xxWDoNicyBVee4da5CZddjFjoEg9k2UqNxIbWH2OHW2EUxgowwPxAl6ZpyC
ewWc+iy4wYX8NaiN8hwGlfUgAiRSEPgrpHrrsVBK3WOydK9Lj72zI6p63UEUUGO4iRdhhy7vYv0M
tynKMa/CTc3SehHaiNF+qYEMWSMmGNeayVOxRAyl7CN2C356S4RImisa/WNpFPQ7I9IxY1PP26rY
C2YsHrGMQP3OrW+UkfxAg3p1NavgCM+f9p4M9ERRgPER571WqPg2hRWx4rGdoaSy5v4AAmThgl28
VPVlWBLNwir+8LQTUI8o6EKyKCoMf6Z11cNtgtC/1mNLv4rN6lsMfpP4qJd2rc1FVtvoLQ7+nAQg
xdAodIsj1Nqtu6sLFFS2AePIUxeBKPEplXQV3cL/1lBF0nKwslaKuD2hQcL/5DFWZ7ock022lci9
rY08XkNmVfax11whDDaFDhv3Ua2OJyWCKXk4ivPQSuc/s88SaWEI5W6F20NOnIHaCKvmNop9Y7TW
B4jENUsXNGZEV3Lfhsbd3RGtl2G+AubmR4ZPqGhHdqkpnEIuBtyBePSm68Swv0DSY6v82sMZaOeq
RKnP0Ld8uyDLQSMvWqKEPVAfxkRDgMVqR+1vksE0EDO0/R/es5TqZ4c7slTyRkB0V3gNKDkiVBv+
h5bCNXdOfCVb37nnLklCyp7LDaICvcvSa8rWTC1jJ1tCV1g47VSJRr5Iq4Qxx9feUo0JI2JY5p+0
t+h1aOEEUz95swoOHEWMmfWX5+CjcL19gCJ23CFjQtzoawpun91QFr+0j0YPflsamDhsCjukcUwk
l7MjufWCjfuBUSbkm6ftgVE29FuOyujR20bCMrGdxEIf0zL/XIzKUtfM2xWlIOvIisW85OeSBRm8
c51BypwlDwM05qmsh55YZF8TMm0S3fQ6tnby9t4Con2iehM05h4Z5WiZq9RlFmTGvA2uhvWk94Zj
C/s24s2NvLDafm0ZDNV7cYJ+oPN/fEJRTdMLlsmC1Hy15IZYjXjEdtLpzCiSQmQTTew5/agcNDDt
hm3MKFZT04StqzYJ581dDq6yVPyFl5G9B1v5bRZ7/z8+cYDfYilcl0Fpi4UUu6CBHlFhXniwHXKW
v4jbiRRrzHIPFJl3zHjoNnOVcPSvbnPHYMfQuR5lAgdqLJQDhkLKHUcOFn4qq+lgsU2Hs8AkF5QV
lxf6PR/aP1fEWtA7l8uFdVvnHnuAmYikxpyiHgMx75nGM3gmBTMWifI+9HJ432j2F7kCWroCZfKn
qJmMnLUBLgHvm8ZuQuiZryMUrCWmPnjtTam4VM0Nh0Scr3pI10xq8XvZS30kMCckHTlLUqBppjGF
kHpl0NaWdSppB8YdrrRSvA3MKHP1s3rfqSdopc175rNykUtJFqV1BDpXt2dn6t9xwta9EbP2bU8f
lawy2Z6bfTw2EXxLwJWxAzvfsx/iYw3Z9MoUnujNhAsYn5nVCEUWn9s2RDtRoCEGIqK1h9etKI8S
11qKwrSD0LMnmfz9mklU/qHUMc7x3tA57la/ScKtfad/xmJV7h18fLHdCMD12W3TnJanIKkC9UyU
gw9vLLyE7Uidqa6850nVie2gVpK6dOhM4lEVP2umH2kJNMgBUXN/DgzfJXLtSmGhHOIQR0d/e72H
HDzfbMI9uvE/JA1zSkmtBj/KNh4zJGeos8VuAhW4ujJ6tbhTsIDoqEP+NYnvm6/7dfJaKOTxTx+I
2mRjofQO55yscH3kErXIEv7pToqABrBhiTyKt09Xgx4wFOUboF/+VZCz3DmsgwemX/vQMTBXeZq4
QyUlb/zWDdUy0FY4612jw1E8mWNJNddzlfhIesxVWtCpK0HhhaP/qqze8MPi65jwgsRtUmUlpH7z
IMdz1QkCZLbo+c6POCh/V1I+oabOsTz55IGCzg1Xmkkyd2YGyPYXRm4H4wyrDevSwegyJovM/4Be
Lpd1O3XjypboAH71SiP1VWiO+oTd6CYKJIyenutZyN5VNi2CjvZ64ZG6M5KFIwsC+wT9oLrqwXdl
WDYf4oOIliKqh6D3TsuyIQCSz32NHx273j9/LkZlM4IFJMCs4vUgJrYuLblzJ/o5rnZwWI8hI1Si
GFhn5mRKpepC8e1fjk2DpFB7Z52iDhJk18Y8AKpVHlCWww0rSJD6cmX23ZgnoXSq5Ep24US4iQiP
tCKzMuMF4pPgnIOQ/Z8F6tdFOl34zvwu9RoPknH9ZMf1xxWpFPp9f64UaQ23Fccy0oISWgW3hkqN
YYJ1ULXUQCDtiCDCGv/UJQshIHB7h5w8BO7nKC/UEcIZJB2GG66Wlo/hsdzXWTp3tdxNpfQS/7Bf
2dUZDZWJfhyvca+tsced4ISP4azZ7a/vqsckDHMRqRcKubY0s+VK1KKYSylMQYx8iUMZ/2WsVauA
q8XWDUHD9JXfa7nnNOousoO6vDmOnc7+7LUFa6/k2DkdjjpRSRj33ifVxQL9XgS4/vMza8tzMT24
yTSs/P8cjZ10f6y3Far646AMRAQP5TRntoJf1R4R6ESr8kOKqjlglKXSVoGeuxkWLR5BjRsvw4qp
lVBuNxM58K0XdkbM4DGPNdm95ZfKqjjNJfzi8QgQHh47ypiE5VEZeWRyWHmxXLok8SD9AvURcS9Q
igWxYmg0t+ldQsZUa4YWNEqxs+I9GDbOfNWb9uR2cV/L71DwxVUhW2Gfe5tDfrwq5UEP1YUPu0gZ
hfgcosj7SiWMA7NpIs+WGCFrNgjZXidBKKK2id2C/Bh4BN8EFz+AzV+cJWorpSzOSSQC18p8Xyj3
uaOwXPNeKZhUf/1dsIK/HDF4zqEqfYej4TZadSyY+74eja/nyIcPpOIHI8TWgvDkTU0I5y/Gr3Q7
KBlL9WVPLnusAKxo84b7MzsBMfJQCYiD/6zw2rMmj3Uh/aOtFNF4ENQlf9pPNewoVyNVwnILbU07
1R8lhuLkzQlMKhTCMgEBltiZR1X761PevFt4ALkyn9kCwQtYf8Uq+gRq7QFuyExHFrFqizUzeqLa
hQbioTeF2RYP9uOx+hSbsjg+z+4s5TPncwKfIsCboRgZ1EcEJLl/4OQGMq+DGLWQCJP+3WHJUQQA
ug2VaWgyGzUuT+bnYCU/ttBwC7M7kqpnZSdXh2Ib983CC76eu5wdv7uQhkK3TqZVmEaQisrn5kz8
p3UgxysZrSfRbxjM2tTqJ+xjx96S72h4BHT8b/2ivpWh9gb+cbdS/RR1FsJl2QlpkTCu8UmLq8Z5
BWZ8Z0Zf/jW1moTl/K2nackuSu8D/25yoIvHNIerTdfehk2mM7TK6DLhYtROGSIGZPnWgqrJgnZk
3ot9A0uqZSLuyJDTvmqXxhQz5PZAkKUWWYNi4hwMCpg0pW1KZpezW/cQeMGbg9Rkjh1iBnD6TtgI
bCMTDLtqdomrjUlTCX+d1k5DDbwxuVwWzraqxwPhOq6Mib1Wz4W6dyX2fJ2//EJXbiteVotxbeAN
eohhaGE0soz7ItUqtgWm6F+Z2Hf90fg3Vmnd8OcE9hy99Ry1+ruixk2SsaqXMJQL52Xg7jKZW3E+
ViFx0ff/m+OR/ktd0Cjcp/rYdx0mtlBehCkGb44OpA//07i8XZIyKh+iPQZNiVa4Q14/TXJQjDlB
sQSUPl5sqo15SHj9wtoV+NCtm6A9fnpjIbEuQ7JsMRdKx+WPL6kO8Gv//w8/LeBp5A7BJ0Z9kqyN
gqVt9Tg3MF5cncI3tvGWlmzyno8vy2GjytzOvHgJMEXCpxakED++h57ftN0GorfhXj8mm+tC2AP/
899KviN6PwF4LgiHX4BZf2G5QagnVBSjTHqFTmUB45NvuP1aVrqs2hRiKt1YQEE5pw+9pddP9tED
Tv7eWxChLAJubk5ZNHbsJLXsnGt/8zTCticu3v2U/3s0T+wnVewOgiELsxS3sCw5wYukdnZzFH4o
QvgGOhhtDZDwuRDn6PZM/JTjaF0sYG0r6I9bxr3rIqZ3Nod6XKjq47+F5RuaUmrB+4jw5HGBr1XO
NscCqx5P6PXY2sirSrQvv9f60sjXYx6BsNdiNa4IPcvvzqVnTSf/mRw944wBAaCRLTC8Ff/i+JMs
dkX2XLQe+wradW74r52aBKG04iPz1E1eLu0pnbu8kDyVfWvxFTw1FSPzwXqLCcu+K0/ZOiAFDuxX
jOl+2oXhtrXo0L09CyjwiHCRrqX7mz3EfkD10fP1TKRNys6iwa1mrFTqvi3bculxQXIQXgl28pW1
mI43wmtWchcC5/Au2aeCoQwtWy+mI/g3aFZf6YygGhqHhO0FLlr5+DzQIOlN1w3PuDApCNj5Jf8p
rZjxNUav15Lp1lAqI3y2m/tr3qH1swZ+XXNhtDOEB9YCEfkaNVP1a4bYDSQBJ6IzkTCETOgGpGkD
3M45vmedghrlNl+RCZnH0wxHcIOVTj+k9X0lR7evZgBEnKDTEOn51PrMSlkKHsUrfGj1H9uK/SkS
2xyBH/b9y6kbHQkCxc58TmVT3sPcYStsFXJFQNu9eI/73bHg6NTBAkxze8UBYOa+WjO1WrtFr/Bk
/Bat1YIxqi8Ah2iQ+N/5vabsIFDjpuCJQf6JRiVkW7zd8E68jLpWCvNFzoclLy52dkMnp7Ct7BT0
Eq9fZ+x8sw74dNZdwKj+hfBG1GZSOU3g+eWGLou7IfK7ZmxugEnij6H4Ytt84dgfxpKCjzJAHVzg
vA/ZzX8+O2Po95BBHq58I3I0T12CF+VrgvRdEVC1NMg1URgnlY099vO7VaymSnLU3BchuVmBjjlI
RoGdF3Qr5VyQr1b4qEL6cPLIgEFnzwRwWA3LvDTsgWtwiyVkYwfpLmSIt6XksUSW+qNxIz34/A3B
+/JLxPyPnjJsoUGAlPnsli+d+eRQBxNcmrt6eRuTjJ6M/CYekPULYUB42qw6pBsjlBxFdfZCMcFz
HIXVbYYPKekRu+cQlcnBmvfkI2nGuh9fqX0v9QkAbMLUm6+pZG6eQBxaE/thaD3hE79BrGy+qTKh
YDjtnf0py0LWnQBbCCzav9o/L1T++4roozWAbzvXdJJl0GAc0/tF6kKQ8wuSMTL5bt4XTWstewVk
b97575vwCx5eb4hNnH4qkkXxPkgdHrxA3MO6eOTzsm2pfspYp38Sy87XAqVlNt2HOyHGU4LrBypM
xl119NSm+qQOKnLhzJ+dC9+r+JLnqMgDkDzouEva9z7C/BVRGrvRIXuXPW122ivfLHMFUSUZwMCr
STOSar6XLY5mK3zmY/K52h5AkPONERJZucZcrt3KS/eIkU8PIHeQVzgaDoNILubyG/v6g3uDXcJ+
ZkaiNNpoGnrTq/zlIt+Q1FpmKRzEdC7xlhCx5fzVx6KnwUkkDebUDU4T2eHQXNklJHjLIu+X5QMs
vGZ4E32ZOQpvqO6TyaHoNJLuRR19+QWdx5F3iy/Tj1I0iXp9fLAPna+1iReQXavaiQjvS7lXRnaU
zfs5/ToxlJVcUGyKRv6ewz9uL6jFhhJ7IcemEINxQXobU50+YJ+t+RUWxTeXfrexaI9i597yy3Uf
FL6iW9wEQ+mVwfX4ancxI30igYyOZ/BTBhESoBeW1Pi9xmwis98ZB417T6seyvryhwAX55H4CGu0
m3N8I2bGFldn5HHCBPYUMiKDe+TtHG1BVZdfSgQJxCiXd/6ApOvbpxcuB3624FmW9S6yEqDuCPgh
TjKPrxj+6bmhvaF+eUQD/fR81Rw6JD3HF9wAyScBUm0Muhkuv+Vydm1Xo0smxzJ1rc7SodZ5/KT9
rhcZ9JrluPYl7FGNeXv6hIYw7oDL6aJA0dQT1qXjI4zRPOF5sFi5vrOCn9zSn+++F5ofSFAhXh+p
sEK0gP60SmFiMY0cLJpIMztWsEo+FSMMPno6ZlU6HcJ+j5Vy+vlLDCq6NmixN7BZwWgq0JReyRbp
kWALCdNRQ4RWodr2w2z55QqB6jSIZmwYMdCLlNQ5R7wt144nTt/60m5S4Fbu2GAmOoqumUEtLnth
Ouu6RYm0D0vZHzNmyPOup6xvvh0exvrKvLEBG0lXoALknIPqfOBBzR5Nmd4jLoad4hcbqeomDEa2
WrrVrm0pXsjFTtoZ4f2fcoPRMwEtT4aSPeq9+/ix57gMOQSsvg7ixNabFUZwM/TuWYQUJPVE7RQL
WUhC9RYrA73oRHesu8VNlGUaYGmDTouHW+HFheXqTfu2XBSQS7KxMMZxBgchr0ZQjUr2V2/DAqUv
9E5W7VNBisxfqLREf0HIsCuYVpP0bPzdtd8sLtaLd7SVt3ahJ0oYByAPw4Mh2U2HbXdAbSaUIesO
anf8Klm6nPGTxx+AjA6jV5CDyYf6i8wvaY0rp01aP/+LiBRUYyCwLncKJxrEZkbLndhA5UH9Ar80
SUc7cXMAsScpyZTMbQp0i6fNHQPDAZa6LbBq5oQVWf5/js0H+9yOz4SgPWvWYc+ssHX9Uissextt
m/7KSJduEQI9V3+oROTMf/gZSITcVfXwRu/gKzyaaMoTZ4OcXrOEgviKcoUoQWVxrR8AeOKsdqDl
r+XC9eldmw6gjjrWynlfUC8tpHW0s3O6w2cab0T2nVk1fH3zR8O7ecoA2AYQA4pIydoZSEy5OSDz
DBExios6fur7olem8zbEuWl3fEwJnpRFauPk7mn5oJF6YWJwOdYO39ijD9A8Uhs9t9gGSoYEdOGF
n72Dv+MC86hxNIlsxtQjWMgkaYezEPWLiISwbivBsJQpseoRg+db10mzbAhIKJFxp5Yvgur/S96d
Lt2FfXLUGCIc7Qi3sdBOROxUKxmaSVxK4CSP05roG0CDZppLNpb7FxVvQzPsb8u1uMgSdNiBWhuR
kYyk+zQYppHYH1LHlcbR5TPHQscpqcJ9xGiNEvpHA+/BI55J63k39Tr43V5nYEaF9pi/kuk8s4Cc
Vovy1gjWrXnKGpM1DdeUuQ4JCyodWVcgUdzxQpjXmT+HB4gnn8B92nlMXualjgga8Mg7gGtO6hcj
hz+tfhrcvbDCHNzMhIZND703VCMKt1OjqjL1MrGPsS16zJNuXxpNr7sl4tpA5iMLXDdjinsvoXkk
ZhplBSjW2sFzfo1ScrwMpxWuKc5BQaL+k7bj3ZZz+2/aN5/feaxcbU1qBF3g90WiaF0FW/Zi+UzR
lGgou5lKqrJjJgnwnhZOVmhlDKFdLxOSGmeGczhqwvzbEV/vLsZet2k5mhOCFog7UEnqF+RgcslT
MrFMUzEpGJXL+8t7ajnNvHBAyi7OVGsbB9tU7wuzW//xdhEAikex7tqrRXPdUPfeWEw63FUXHC/Q
DQAe0L/CH86hNk6GSluNm3Nco5TYXaFJ3dt4BKla07czaCbE+gMQF+TMuLcZoncDxsrZPgyVVyAo
RrTqGUgQMiJBSCTLQH0rUytGfFJqYNqxei94OXBLnsa0j33DA8Hk7aP+i1rg9352sknJoE1L+rUH
61136RUdZr9XSI531tvbZzlobd3P5p5lAlbYhtc/CWju1PlCShEAwusswF++AgdwKFak7xFMgyeS
kAqOo3+9GAYSU0NNSot3g8PJCNMbUyri70lvdoLVP2AtRL3clshBQtzd1rzF41nGZmhLAlf4H9Ai
sUUrcwU4mayB1NCrwf465zHGWVMQs+0ff1ujFIvqvnjFMZY+Tk07vXZ1GBm1XWaLvBclUzu4bYd5
R2OxupRqzcgDle7uCSG5MX43UhzpZHzHMj0Z1p8qRCtC0SQ2tlagVG61gBp+fV+27+vCt9/jHh5W
VgSpjVcaLnIzbB1C9qeZpLBG4RqGanSi4kf9qHZQXcRFcsS3/6PE7D7pbaJBLiUQzvSow4L0PbHJ
2StBY024Lg/+aO7AQn0kSNn/uTbMLbYjjLJJVIRQxGu41YSzV/eWqCKRzvyH6t6ophpxtU+M3IuS
KTxmWRf12wu8EjXrsjPp+++8a57TN7ERq0NcQwyj25R0+vT9tYSa0SzlXjU2pfLXGwVF+nWAqKaJ
X/dvJlWnYW3QJSd85JgfHBmcD9G3wNpjWT4Kkrkl1GAUxPf8y3gM6NrBmhPZSoNQ2VP9MuFvnX55
EkONDhbRjiBLVtob6xsiZxzMmnTeFMONRF76RpcE9O/zkuFI7O1Dm8LNtA1tRxRYI0chP4P3HghU
47AcyEfZ3SfDG4O/L/04zsmgNU7MXgvkOYavtP9/SvDr0ChDqBoLP8Ff1tEXsqQOpLqwqO9GUP2B
B4XCUsSgKUAjk2JPJ/ZhbXQHFvPk0z3pEMjqHA/ykmVqYzCZDj7kNstLPfePXHQt0rdJUTZaxOh6
UtxG9hOtDWQwoS8F8jMLzE+WtcrJ7UBk6LT7jhi5uNU2FCBmUYsDwCsQeU2Bg6qhip2DJ1dgNUL4
rzRQ2sIWXLvivdGRaS8yd3/ZZFtb1XepIq3MTn7750ba/Bdncxmg8YBOVYPhRwZT5e3wwC5lv5Ag
VHmaGlciI0Co0fXlP0VwyAkhThNSXM2UyMCLphDjuTkTGkhIIrKUT/TxuzJOAZZAdphicVfSFb8v
r+PtTMDKRlctTi0MSg9zizIIl/e49XwlB67BETTTraMdNHysprUfrzjndlK9HLsq7Q/ZuLWbymtf
zbQJLpbhEZZltCEgBcL5auWMXHIZvRAaNfYeXjZagfGrnaukql3BuqSvziD08ngjuiNdDkcWVB9f
+Tt3iQ1w2NJVDONqDiPoj3HmoMDysF99mxEOqWepBOe8wOEkT/lltPcO7RFAhdvz8Dfi6W+BF4rB
za+IVgJWNx0u6G3l/7P5Txti25NTVe+WCcb0OnxeH4j5mKQT1FhlUWMa3I2d8hvoz+ELhhuMf2cq
iAFXZjreZQ2w9DhGC4iuk7DKzTXEnhkHm52JEpBKVQCY3PyvKUchI7U+xCnBGHnuShScA/7bQ1v3
2CE2FXyopgZF5d69c+O3nEADL0w7gwoVnOJA3PAeTbX5U0hPumhHYP9bmAjcMDZvuyZT3RJ3Ri9y
WNZkCdUuEGws3eujoIHSg8SR3fF4HSQ5fpsDz8VyQAbWeFdaBf93p/EBTb7PDZA5OWZYcVysyoH7
Vw5uFnqykY0WSyaVqj64GzsKkVHVyQRiCBx6/u32xtUeHG/8DFLeg9QqYhxRHzgXcEQG+DEuyQDT
2eY+Qxe2aYUwO6sut59o2bCXNdAMuRthWu8HSuO09+zeXIGxi81l5PIwQWqgYj3vvx7K2ARICFTC
dOFaTbEAcoZ2a2RyTVXAtsmFelbGuruMafz56GV7AJC5zlo8Dln08Q+Zn5ktDAXwZDkgsSu/QiCR
I9KFrp3Lr9/VQXE9vJfWVkGXnPFBz7pUbs2/a5WQn+k+OHGxosRakXzrV5CVu0QoKnzMEjxK6vNS
d/wygdLde3t8Q7iZ1k2H3VcjVDbN+dqTX2jKukVGD9VeKaxwQW4Lf4NA6poQFRYjSFkA58NOgJ2g
ZIpJ+GKgnD2FZRmcuqP1ddk0w7LB6cRlOOoQgCxXJCa5bh7CwHKWBhqw8bcMZLJ/XFTocep0P9M6
326jZ+Q9hqRuPiirwVfxnGwnO2ovbsgTGMBn9RI7Ae/z3BZWsXURva4CovodR/lkZneOI+o5frDO
vTJ7bOOkPudcK2R3cKb8XCLgU428YrtmxfAYlkmFdKQ1YSkvX4WnSYGoTmwltm35BWlkuGtFNDZp
Bcd50vAFNfQULcjMOv+mol/Yz33jmafi4nVvpuyS9mL9lmupMx0zHDQJ979E+eKXKzqoLx+JWeaE
QBZwqyMPfSojv7t90CeiXETq2BSNogGA9BY+YGj+gcOzgmNcji+vrAwriNHasxnJd3moPAaCorlU
FtKX6IKNb1iAf4/3aMsMNwWdwTmr5zroYkgkc6hIXyQMaTY70NthhtVQmvseV08PsJwAvV19VQsQ
cI3xsXByzTzsRmh7s6k/LofvKMUSUzirM0rSbrVSnYSmBDCJIHpSWabD0iuu2IPpAh1J1uIWolxi
8yztALdvTN/9kdmEvHEvLWKsEeMJsgTagr5nEFMJ130NPdPvXutYcMnhZbh8XhaMdme4SvBQvSMA
ipYhEVLEDke9mr/ElgtAlbJVmsinGnrNCo52DY2snkM9nD7iqUqQD4XNZ5dWXMIQjRMz3LA9I/Az
uvMaRmBCd+FSRkvvmfQYxHEVfY/UfCJQalUPawK73acltdt7bNY+0jjYX1nhHU47dCMZLS9U/BWt
X/daY3cu5fMItlDEFkIQav26WT+8kPIBQjj5Yt79XuTulfK25jScD2kPLqsggPOS7GkyBgvg3LGi
TNGtIfCLwg1PgtLfDWJBYR0CD4C5AyAeE6NF0gOrQPP0BVJlO8DZfW3A93k3nTStHGKi1QJm/ELv
TKAhir4OtwDAtMn+IB3cVchMpMPzSs8CINTbYPBlW6BcUp3tNM8eUxCPhOIFlEzgZpCZaVL7Ll2y
WLlcgyj2i3z9mwVhFltki0iwzdkjtwO2NGcLKG92FC8JbrN5Nm5WNsoiEy0jJjLM5owiNsQ85OnI
23tBxfwioHcWUwe4hK0vMKaAy8BXb45ntxZG9cW/dRoAvfwRkp6RWeBlKjvSwMFLpoxkxW4/RZAF
1xWkg187yKne5TWYRBJ1ORnfwbyB14m2P7yMhvGRfCFFqEYX8JAXPqo4g8cV2As5k2iOa7Jy5XgD
Saf3lLa5bHcESHwDu880rqOtU6W2qaamqoSHJ/4KEq0elDB2BzSuWEaIHad9k8BMeVYWkXkwcNSY
fQ7Jwst5ALi7qALhVE0F5g2rcKbophg98dlbUwtu6JH1YBJH+kCJN/CDBvfcDMw+0WyCfRJHPK5M
rO0KqiPrw9C5ByYQKuBM3zTzo8DIb1KpuZIcbmC+tESbW/8Uaq1RRA4FGLu3gMPn9EHXY22fFXnL
0eNkC8Bl5G8xqOxI6IMngR2AtwenlG2zC2zRfgDnmLX91cHMi+fAnmv/mAtPUDC9J482v001uPjY
AftdPyoQJsCmZFSWuv805IwcbXqJOYhErFtwfVWC5Wi9xnExo9fxidRNdLIsGzMzC820qCQysY5X
73Wue3400MfPegLfY1scAOOQG1pB1C58ZYVkT0QY1YsugTwFsS+gyiDwzoQSMCEzfRw9hmP1p7fG
KuVmfD/XKf/SSvnXjbgnD5MBgqCruJCnzZJfuY8fRxsfZJpvMX9Pk1UzIYLJuw1+0z3+DbsOvLSN
jPPTN34RArcMx2gnoLzeP/tF5pufUWy6pO4LxNjkrzPMj3QSbsHsE9VcY3GCnfRwPKL60LZp3qyX
K5NZ5f2IiATiOhSZ1QRwcboPFRlB8Atspp3dBop/nc16peLXTEDHF+2faMQMgEJ+E4+pY/a9jX9r
GXmolIs+jX1mzwY4Nj2hRhJh38l9RhnLVqufVsGLeekM592Diomjmyq32jVqCzzEJUIUNWpkms23
4+JnjqC6zCadIsugPMluYLibzXjw5UzFp49P1sRFGtPqXp+j0gGadEEjSJPlhBvp6S1Pv51DTgu3
GS4JGFON0LxGk5N1vpSy0C/uJdDVqdWtZtYQqpdwy83UT320yxqi4Gn6T/gybub4WFTCHrU6Mp9I
Xy1DNM5gyGx7+qhlmNLWdt4+YFdECOLL2rbJe7+qlBFSdforu1F/n9156+4n0Qjhb1MOyhQNxBNg
svlEBLQvVtpGHBzTs/bK1/oB7sB/kj53txxnP0elSCnt6a1/mHpBuThYO4Pdkh16xcE0PzE0nONs
XyB5HJU1HE1SvYyDgobFhSMdhW0b3QdqtNIbD90cUML+JrNh5yWikBh6aN7o/e+s6FIX2drB+6O5
ltXuPcfPOGbZXprW2h6TazkRfw/mNso95NBnsW/TsesZO/SNJpzr5zl07jhJWzpZQ+h0XAdydY4N
qpKQhpiD6z4280CQntKrG4n7/3AUpcmLMr7w+Mf+4haRyRKOfSZJvpkbRlnUnTKlY77ow4r85pSj
Tw4o4cGPd8boQqKnNEKcjTho14gOUqDsd4SO1uA+p8754bZEt+bsQ9G+IfiPbm1XIV7NglKkJ09g
OWlyG1Q3fqCSRTRx92bNiH0LliMZlcsTllIZzG40XxBfzkKbtp8aY7Q9JeJUwYLLadYiOXLGvXQ5
cFzaBrr0jfLlSKZI6IJcYStyxX4gaugQ428Nd45AVCCUBPDGckDd2RgNdT8RvrCwOg/v7vjASofk
ifnPmnFlRHKnPOhmxQjjqTGtYHPGYm88PYtKv6khnFtdYKM3Eu0emmybCeJAQYCW1+QJOEbK1fgl
SL3m1nJR0E1CgGuEKM9LXvLc5P0eOEwdkt25KHmD2hbh5G/9+5ol76lRwD06zZfNbRoAeo/lcomP
vRm/+IQdc7k5SlMpeXH2p6k9yZIJaOTUS0PAH7EwVyZS0W1ilD6XHhMOWRbdyNsWunbTAxISxpHb
lpaeGoh5NXt5scTmJaAoTm9p7R2B7n8banK1p4SdT3fWAqJJKS92kgxXrTX3wpGPptg8+uhv4xd0
FXspxu6S0D8vfQwu3CfA3f41eXNPWvYn0rH8Sf3d3I3b4cXLN+xht38DVsYe7IN4ALgUGH8Z4MAZ
UiWiqlomQlmG/5YvYW13vCjoM3RUoVmtUoDm6ewbyLwQLEyVtm3KPwvm9w1eSnh8FRsec4AsfYhr
lNKh2FSZx2o2foGL7UEJgoMQgUeJErxSfJw5Z1jniVPHlxnD/uF4Krn//ge8712AhrtisbG5Ayx4
LjaPkRPFF5/hbk6BOonRHq9Jqpu9iFu9AUpJFMuU2Y5JkNnDOW0FJ12xOqPYvyrvl49KbTAQGG8J
/Y54REss00eS129ilmUrz2GfDsjZCOyrW4BzPQRUUz0gqMBJRezuzU265VLB1aWv9IRrKWdXI1KQ
7pRarAL+hao4wlp1ykoUA6eWAI9B1FqhtZwQaecigPJiCiyXAI3pbZsl7Ts1l15uBU5v0sFdcIJQ
4P09kdFha3gZu+sVCE7H+ynzStz83DuH5dJwz368i/KswQZefwqtKHXKNVeYxz+J84qx6/apaAFQ
v9dLbiMIpUByoLMWCC1rSP5LsNLR5Ms1xnUcw35TkUdgyekeDlq7WQod95C4KZd/hV55nJqLvEdx
jk7VWccZVwhl6jo7E9ndEPM9bDHSAukjV3lCY7fWokg5UoeXn+THrqbECkFA6bTbNhvDwNFbrOnz
9B7lM9hvaC3NgFBpvyQlfi3cF3Umctw0lEGdWvEixQ2G87dFVQVCguuR/PUBYhPFy6OCdcKFTm7Q
nTQG0YPE3S8iUoYVX8CTvPVK5yKpzV8F/KfYHxLobiVNXGyxbRX+1U9UVDXOJPiPzRwuLSHz+4fv
O0UY+s8b7l2F9MNP/5VAhXpDmCEPR9wcB2j3OJ4KYiGoWEXKslBsE2faJ/6ko1oiD8xqF9/Z4fb7
xZMvUZuS3JFAFdrDp70zFWeJc8XH6KCplGXlZkCsJARiGQrqrUUHFBE3tGfL8J8oLYVrD1dEABVo
lQmFt5JG7w3L66xusjBnB8RETOxu8VDFoJFtIOr/X2gPVIf2LBfmy/9mXGykVnlZojEjna4J8KXf
LmR1denCtH083KGLk04owPqFMG89OTmtnUoYjPjz3z6CRejuE2nMoIwOzXj4SdNWnpfHb88EVKjv
lSxY59lOizDEPOIhfQY7LqD+nEeWWdcwNHslEDR3C43QojHfJR5tP1W4DfyRrwl5yK9lGthXxlj3
ptMWyvdtD3Dv23pA02WL+eQf0NE61zrGqO7o0iGVsEYWpXyH+5bCza+kxTSkl0F8x+QaWXKrsPe2
lKjDidb/AXmMjuXYgz1P1rur75LmNUyXn7uKiyowSCkS7bS6xY0MvDX1Qp3s6cMxCiJymd7INBRm
RG2DH9iwRw6IO8g5ylSj8f0FjO/61e9FZoFGTtHWq8mATU5MpxLE5t4mTlnuNHhp24eg0wAxq+6P
n6DUWHtE9QTu1tGeMUK5eYTIK5ihffJ7UDN2g64DP6mUcFbGG+DWSEu3BfqataxiGfaJdjCmZ97X
v7d7gcsD3RBWyX/rij/xcBSk+t0C0Jav46sTd56of8HriDEfNwDRKi9Ro/BGV+b2Qf82QQR/W8HR
AbIEIwQpWmGMfWii7+5XM3N49/7Bvhefw+m86frknXZbEPyzovRNkUEAhZhsvpDK18bgsLlGcPVB
zVnBv+hV66fNPWfCrx57d+ejWGWRso9gULRTt3gek8fSBNev3zj74hhNvV7odzESAnNsDOY03Cpg
4ON2efDIR2kdvHsjg+sMDjnmpkmUi9Yw+3yUL4U5kTc3ZxNdYp6bcEXyZw372JN8IGuVRBCTv40M
VuJ25DuibV9hF0w6Ctf238MVPUUpQ+6UbO8nT/Gpd4+mlHfm6CzjFABiPtAlWaRpVvVmDnQDze8x
3vGkNrErqC1g+KPsW61z2st22I/TbtkCtB0yFItOb51T5W6isy5sifcX/8yoyywEB+5iFbrNGxpQ
whOOXyWVpvd3EG2p5YyfCHw/Is42NVs4lWyMrKYW0YD7rAtWgwR9WjqH4f4Nq/eYG1FxI0sXm+p+
+U9UfOhWKCUfsR1zxT5kqBxf8qoClbGk0N577lGD3V1LDnORHLxN5cVoOJd2rtXBAaqq/XBopqn5
5BjHxwT6Mp2SPuP0t/vJLRSFlcTubPPw+PoiiylkGSK79F4J1BZY33bFENv71iBgJjelSkMEyPKe
9/m3/2voV4Dovj27J1B70rkQ/rpTBLWYku2uVY0LXnRjzvzOe8SdSkExvXSp9C6uY0gN8A2LWdva
KQA2tAmIU9oVfoKX4d6Tt8oOy1yrYcbCx01W8tZef1RNpSb5+vmzFmKEAc9wR1ELBYnka2xkZAXf
jxIvP9OXap0QD/ND7aDp3FOAUjQOOj283CXJ1nkI4LRemnasVnz+r75MVAZ/FG9EFB0eeHm8nTYp
USNJtQopCb49eg/0SvMxsD2R2lsllzd5s26YeU/FOrkXvlJstsX/XgRheREWo9utN7oURna46rjs
G/0QcF/URmw+RIovQ5btPRr3HzoZxsp0hiMOHL1FHZLCPauMG6c4taQQI4eB4XEJTq5CVDCMfVy2
ehW7d2R9ctCUlCwb49QvzfZcwXXMS+ydrvlSKsrULxFUPBoCGNYFR7VG2Ex2SGse/O4WrIXE2752
CCH724MbRPp7AhBaNBoSLyILnftowu8MuejXr1TFj2Pwa687zAOstP2QMEwPOYvXIIwqpoqBacA4
zcwGpFgG4ZO1Wsk5LLLTW60vnxvqWXTQ+xSq9k0mwOTEsnnh+PZ5gNnnZwuxpWy5HpY2DeA6avBr
uuQFuIReW6Mq4Vu4M+yI7lLD5Z4FXO2ivlMPAVdckP3OqirDSrPFywa/VooMDmxrrpqTmzAEUtmU
qNvFgP4LtKoKcXkIMHD43ImETKoM6AcmVP8yOFxDxolFwxNoum83kRTjE58P9+bJJOAyxcze6fKY
uTlwadRG4+KVCr9cZMT4rVzy7+kXyuAXIXPyyeeo+tUoi0NvcGWJHkZKlYvm5+RN5GBg1fAUGuyF
t3AYDbqwHzC6ZDwPUJasdhxIreepSU9EGpxA88+6Stm+MQ8WeuB+YOBiWYDoxJDqwJ2l7XrEa8Mr
YOgxJW5r0jz/YEQW19+4WlIVpOPj3hqPokT8cQovu0474qStthCqMX+Uej4dPcEfiCXq2MseQt6N
I53iFyL26tceVf4iBZd0f7m9GCYKVBItEf2XwU5nAFcep7u3njsfAVFtGQ6Zr/oP5nbmWl094RCE
hKyvu71uWuyV+Ncifq6p0HU+m6sEC26ryr5y6elwv8gyyk+mK6607KZvSCqrfdPqDYMoTQpjHnOl
dZdXEpYIR8EzWiQDQ9Z9IUKH4LU8Z4ks3Pbmq1htCc6GnMf9/T08CWkIiBmAieLnvPGmD88WCaKP
UEnvIMI34Sn5lGhPvXL2CxmU1djSwqRSSAbH3/AUi02VL3ZeaAmR0eYo3byo4juV3KCnHJGX6Zhd
e7JkaWXzbvc2TxjrmIzneDOcsPdDiM841PgPL6iR7IKbcd6vXhrZJzvu3X8Jo/+GVkNeX6KliCpw
AbDtboNL3OGJ33UyRGoCuH4a0GErWOfgFL4Ns02UmvFJrAiSCfidY2wcuJ/9iiYnv7VTkJmgSO27
2aDfQ3Y0CrqQDja/cR1WjzmQVucl1XeEA820DHoNft1tyQ0h6r+/ChVeesZWSHDzNfeywSSO5RfO
Az4BU/W/tGtMIG94jl8Oa6mO3paKSyf2fxB8e+q9yCbyAA6VVoMmcHVq/ZV8/jiPa/a3fUXbpRvN
Npf1FRLY8rlQxvAaI9AC003Ny+9s3HP+PCDQLNjKo+DR/AVu2yXa7XRsHY1awOEk1ZXLtEpgwojN
4rHfZiNCPGjW0xse0A6rdbc19T4QW2hpqrodfjRgsXoL71Ag6AF2XnJbOJaZ+IvbViX2Srjsori3
JKSgAQYD7W/u47XgGYUSngw8YVvfX4GRVEQWRcougoCB29OGFsRMeQLk/OwGHHIzmuJOqi4npxWX
qQS2I8c3f9c10sA3uWaKGzaDxFG72Td8ODOkRJNG+jkd6UB1ZDRvyxnadaqNKCGcO8OKNG2AMs0k
Xxvmtc2t8MYVszIZlwFnVu3wu0N/MsuUq1+Ej0tsNXJLbB8PgT7lnLvc+L9fL87kWPShcg9HMsHK
mJKLYqL3AqZdCPNcXn0QfK+DVl83XYORUBZX3YK+nHlkQ3PAHx5V5RdA7KNQuBXZM3iyQsTE7IAb
85q9XCQr1ZJLO0R4P8mDv/IVD7CT74C+nqsyhlHHdIJ9QCJuUzrz10nXpeFMH0d/O8j6PxF2IXkh
yHRyMme271eeqS1TUWc2yHwJ3JQaavmyKWqiO5VV4pBM016QnQoHMA+owdqSjB2x1SurFm2mFaus
2PS3YIavLffyIxa0y6/9SkpnLtSYhNyp6ExFi3QjMy2TxhXYpAUCm5MzmRDfr/5o39fIfQRtSivK
UG7RtJoB0v20mNyT7rLz7JHA+E/6THPWDwkh3h5XJRdc/+xO/M0DTvGHjr58hWX1W1ZOpx5f4Rvx
JEKfStRoVThVVFEgSF7XNpoAUhfP3HLj+1cBBDvIRQJG+pkHEI+9FGBkwiDjn8iniTW3DddfXKpQ
Wjr1NQO9C0VmJPRnTzChqNmIH/QXjx44pUmuCgtIFLHmu0gmr3JgY/qMG8Hfycrx1dSRfFMhlzmZ
o0HMu50PYRa3QY+Rp3CmZSw9ToIQPJ4Fk17DbFSWKWEAg38kk3Cr2qr0nYtlBf9exoVeuS1rjq28
wc+/My4m20LRjhCzGq+AV3Ep+elteuAmUtsS/eWyZb372wd31eHa6In5PeG3EHhh7HIjxbLd9JeF
EoOCyAagVDtO0gfhD2GeJidzVoxRBClOLl/kSCvQZdk9tNxjhdhwKo4u8igQJSlHtiXwaHIvcTV0
Gd4mG+arZiHzrxijU79Ri/VgzHAQGr82VFHuU4ud1Hy0HF30vCUYLyuokeik4lM/zV82/X+eWZlt
egb9pz/Os1n08d8QfZrb2KJzztyb0VPdZdTmCJkW5wuGkwtFByrKvHRiSjdTq9NUJY2yMK6rGops
7j+Ux52Yc1uEZhGvGR8jj4U7BNGTRXFyHs/3pn8x/E7Q2QdFpylylCi9BdR5mPmj8+yjefOVaIXk
Pdvf7i/mDw6AmV1CjA0echk8zSRdReVbpcq/36ZH2huYEFb0XdV53zcVWSvZvG6fD9bB9NyohVpH
YCyqhAh46RpR5EKDJp70mFln2BlgoMqTUMO+AJ2lXPVwulQ8KlTYzIm6Sa89OSac1Lo6AygNc9WQ
dH1cAiB2ONPsYbfIWTR+3FPOIo8slgBdSL6JD1AgDcfJ6V7Op5hDh2WaESrWhGiR61M4CONZd5IT
cKkSv/4QUdJQ4vqnzG9RjZX61rcfZfrbNGq/Ft3EqB7dQFxG50AC/QRl1JxcsYtuiAKVFpeM9E6u
5B1Aw/PW9AH/OQEH02q1HUsCGrzx0cfwEDIN+xJa6PJ4yNBw42N2q4zJUPjYE0d9CbAKVeKawiDt
3KyXrkJJ2HcxkfasPdB2jhNCSkZaPtlUOEuX0IapjGgdMWFkj6l7t7gXNIU056xgp7ivbbnYyUia
p0kFGJ9AmIw/N4Q2wN3umxrqT4VtMrlNqapsHmdbgrdtJiccDmAonfdkwm5qqpJFlKsCJJHmnRnq
Nv7r4JKtVHv+GeENf2wAXHG+WdXxP1CatY5U/cdOMr2JFmhMo0+HFYIVGFO/71rg7ZjBBQB+hLjp
JieMH4+Z3lh9wzZpcbFBGZ1ssaS11sPNAUla4Dn2LbRlBDx2gAYmyvSPp47UJCTrsEEqbfC0q49P
SDmxMN0zEYqJJ+iGLz5YoTVYcHgOMpd15rJ+KVjG/BeJKTO2cuLBVH0tK6xC0FGgO6z6m+OQ2pNv
1EKxEoJthP5Miwactu18bCqwKYpzuwi0TsH8CjbHqeHtQAy80Rbe27QcKcYPd8GK/ivTz+xZ1/wj
ZKtUgWgbFe2ZfSRTQyF4thH6QOCBWPx6G7une8COgZF/zRjoYsZcaMX7eW9Ge/6eUdW81eLHKn0Q
K7LzA727QyLCynY9ZuLSqlY0HJoVvkphkZ/Tc7eYpq1nPw7u6cj677ZacX97ZAD2fVCRSd+p9Jyd
jPnKK/gUs5LcSchG2WpAH816DufsSI0PpNSEhwzBPTmVrnwTUzqLchRI3BnVHY9Kgk2Q1exwHgJ6
VOy0yT8BtKw7pyaK9381jlXWPO6XqKmHicuVcagflYXL3SG0TqVensDX0CxOlvPmXUpKPKrGNOVN
2+Ox3CR+fuaMDXrqXPIgoENRT3ChfYRAXQLHDUuD9UB18l/lM8ijltQ6obpMglHsfWKnY6QJHW77
3rs41rhDspqGJcRahJZ8ljWpBTdO3G1LGG+fzM4Oda57NYhE1gOIcxeCdNp10xs/6uN15iNPjOzj
iQlarykOM48OcGWNIGMAohs3/cWIEKVLKEIUurbvmdV5PFGwfVsoZHFLAmwHwhfvP/9WG4vb+B9T
7zhFs3ZLNKm3NiuYFEXKTdjhMB5Id5AqiQ3j8YidWuBrO9tXXOzJnWMjEHmnDwjAY8t72Henqdz1
TPsiqNlUMgrdFggMoKMID3yI0JdqWMy8KpHC/QEFVSMTn0TV2gWT2LJTEDwO5mBv+BDsGdSOBwfa
E3H6iIRaYqjV33I4TTeD0lV8uGypBHd/p9eAVVjFe2dFoNhdQ9B18djpEWhUlbr0tNGPVJP6YcCd
S2Hp+AgXLVBnyiHB7Un9Y2Lt4s01vu2UBRxcRdNv3VbSOhXMIw1rvecRZV2rtAy+jebB8ERjtkwr
MuENVmC4YK/ByZro1HuPZhDoaBrV3GBGbVabd0DXOsI8eCvtpHrDMorfPcEa5rqd05OVgtSKH1BO
BX+Iw5ndk/7sI8U1j2lVQoGXlLuwsLj4VkYfjbdxk+uJv2d/1wR1kylOeEzMbdc5cTlA5HRQ+wg6
zWexzMtuoy4aciGzXXQpiGwmtHthuYux2WtcwKFLk6jUuDcJzsptE4MnUnFI9Db5wRP5wKZvtK9x
PaCx3komSuB1kT9cveIEn1a6GHKL7nRFGndfohjwn3lNYEsHosnCWPj91xjY/l3YyOC2cM2+N1xh
sCjBYURbnoOEQMcgzl7nEseNUgl09/vgwqDnDAjRCtuwGofkb0lsxXGGMBf0uOQTBZI6kcclBKPZ
PgDfLz2Uq8dZUERZp4tzJQcI58neBdEW9psdcPluMqd1QR4XWL4lq4OxEdnr8CZ+N83gF/OlPWHy
b2R5HbDedv+KzdiLmMQPzWRs8YFrQc5FGVllCqKeqsaYJ+9cv0FjtHnZq58zV/OUnvLZzqfcAq93
DL9mE6Zz6HqvSKL/BX3qLvcxGuQuH8peyJzYI+Z3AWOTnqHlFK7QpcaqCuRLjuuj5Pj8zJuF6Fiv
Jn3AioCy71EqF1s/OSNppHaIXK9QXTWYDxbgZOBnJSYT0zjBdRxWuuh3AchbsDBhFiQhruN099RU
j3Psew2zNXJbUEd2wwGlfgX8KhtbGnXLtrpn4nxQleRsDvKVkhnGcKdq/itXSj9ItQwNqrKjr3Em
uv1lrEy1rOraKuh36iNtfjrsLHH+pbVUbCHjU9yRvtCWDpvyA0G1VAPlxjCzZi+sOYupLuzYrQa5
YbWVTzi2Uk3PVZ43dA/Q13BVghZViYMbkIIPcNA0eFo9SJQtFlQyNFquSQdEoorkYGS479ZoEPBA
Z9Zw/+Mq2JzVYkoFDn5hNNlk1ODBt24rsIUh2GZTiHCLtkQUF+mF2dHx3YMBpn5jLaUI0jLL7zGF
jPBehMbKpTkCknyzgeyGlBXUs9SqWrI0Q0+dZpXIq1F5kOIP7rAHleSWZPdvSb166w3lC92WLACu
jvDdxvnQyW86BNUU8BhsGddHylYPolcC2nhQ8LAxDy3owZj++kFe9ZAnd/wNXD+QCamfVcCXugas
IK5VRPc1syGFlH2Y4xxXgRbPsc3DyA8gz4RbS6PJjwgyaaHGov+hv97yq9SfzAT/hu9He4dZz25U
ButmKoAyN+st5dB5xwwPXLckdXAQOpm54IQ28jHz+VG6tp+R/EuMgGjYrKHn9JH92uwtK3OrYeCt
SevHP6nq9AmwgdZsUeoD3pU4vYbDGMH/NOgbfl6L/63Z2xZLcyj9rtMZvnQq/z8DJOohddnJL519
PVfTB4LDgy8ZtskqMQzQP3DZ6sQQubRfyWkTBSqxBw7UdOjCjnTazwmwWLNQsG2DYvm7sf4IUegy
OkmtMVKtSZ2f9kTX/ixJ8EqKuuxs4WN+Bsv9Lm+VtJkDMNQOSbgZLqBxxKUDdbEgIv19J/H0NdSL
+8iSHBW5pW6nvSnUbhTPwmZgVGvqXNPE4zeWWU23ey/RSKL+J7hPhDa6++pm6R3xueOY+/T2J/44
CcSGpBqhec7AnzolRsVg6SBYtAOe08O30Nk92w3L3Lv7Fxa2obxAxr/annSCYPqyLIY6/E3PIPnz
gE6o9Dp8RxWFy2H8MxLNIrRlEEz/f3EXnRiT8o7XDAAltUw4OC6nL649JDZPpGNx9fWJ7min3yvw
iTIgekgJiTI5ooSgKOQyVYW1dORmgVD9plMomb8QS9ppg0pj+M75L8yce7TgUBTPWt8HM6wODvu2
/tgEzTYsPymGKUQjViSP5fZBrLajSfh3FR5iBVQ5X6uyAYIfCSRX/9wpOSs4TrfL3Je5d+YbdaaG
pVzM2eDSqThSHlnVGqJzUQcrW/DHw5XCzvFnaGjPUgem8k0Rw4RRtWySEac7BzMsB5N92VlaIOXA
5s9s3XYoG3V9TPOBP2AiNfCnIatFcPdp5lVkdJ3DppcMyAgNMwLmZzffxghNTJL+kVHwRLrP5I6+
kDxG+9s6ru/2XJ7q9CTcnhFrQWjcMlc+r1BZB+KZvjGYhq+xJigR2q4uOKdUsWkyeWBkau8tUX+z
0jBAiFAh//jbTVZNvNWkja3FASOOlpMMTiUhKaJxSnIryJsGVJzJ3YpZajNVzaZIbdXTQgLRJNGv
xR95GQIPBBqUR4cNt4a+mr8LPmfrQNfiJ6bHvMDvXvlx2Dyugl5+A12oa4aOIFfZHw1CK7mwOF7F
BcxiB7xlkKZTmhzISV6m+B1z1kApsar5FMMNNqadOvs5Xr+rTzh8eK0QklE63CGtf7ASfjZ8ewJ6
AnDyIK+7mNHePXwZWPvdgsn9m3iSyRDsNmeLBws8PDfg3f4vuNKAoOINmL47+Xh31o6SJ66tYmgS
kqI1bZOk2iLDYAXPWOTyCVYcRwN7DJZdHJfVr18rtd2Rnb6c5vaTKgTzsLiwnYP87ovSBskIechu
B6N7gQWoDbd5U193AKhcUcLrJ5CuATj4MsA0rRfIIZVHIo+TNuTu8tgEhZsB8igGhAER/WVSYwc/
lKZ/JjjMnYpcBIxxCSUljO1lQiV+o3AXoEaQmT7degwnOAAjPbUHIjSMm/0Bfy0+vsPkT4yRgM2z
JW9JL9e64U1LnTAnqQFtXC3n54WSa8pHgKaRdIarEkBNpti+Vt74yMfyDtoM3H6CGFj2CvVxkovB
X0t8ILcxWFb9VgBchuzOGGqIu9pi72KaKeArmtbNl+Mne2/ktYwCrTgHubBgF3OceEZHCBbENew1
s1ZLVrF/x7PUGzPnru23c9LbFVLC07WT9n0a1K83yplUWwLacWcOnW+XwiN+V4482hpHU1/gSU32
TGMGDBfU0PqqKAe/v1/cNXfRxtfTkp/tGTuMkZaGacFb3+gGMc7p2W9SnMD+HvcLD2dR2MW0xX1R
0BbXZROyWlnbc94J7NPMMKfVJtbkKx8E2J6dyv4BCFNAfdQC7k6UQaJAfQtY2smoIpYDO5WJUNDn
MGWJwSsosZ22Rv3wUz0ZObJ/R9/a9STsCyU8TwB4hBM9lBNpjvP45YJsZTYeLURzFXLVx3kAjrPM
tpYuIaSx0ayL3w26LUdy8UFHcNTY4UDgQm3CkWpf37eSVsCgSPJX4QMFbp6MFKDAev9DUk/mZQ3L
KkFLTVilAoKpgJX4IEXAaHSOLIMB6YuWN7xxmIdnkCem8gCLn1/SRcQv8m3GLHwFmukWXDNyP0pI
jaOnk9zAUTfBqIONDdwMJWJi4+wJmIKr0ecYPwBKcM79wYJLBg+KGf1MTEGcny7BooJSLK4hvGi6
DVh5bb535R0qLowaMy4oOUF1x0hsqHTNgNv9oN9Xf2YZETROAyUU8+Eb+Au/wFZ9zmazyKFqkKtX
G/fnT5ZzMZjhjKeegar3EZ6Bxpax5NQ2OYOfQCVkEMDG0wJINIx89wmBRc8G6TpuinhSAR6jWDOP
/FLFkX01H1qxj4dN5AItbXuFTCcmnrbkvfJftVzLrp1YqXODwguCGO87SYbZsw0CGuIhNEl6Ver0
KYPQwiDAuqgVPX66TeCB42qVjItDX37sPfiujzvVDhMP4CYuHZWaUpKlVi5S/OysIrmXsshQrjxJ
co3zKzwMr5hsxBpF/0ZBdb0Z28vEKB2blPSMB2XzN7oyUepVMhY5AbfbXPsXbExezCUhWj6SN28l
BhUlVct1PvxhQ+Hcv5t/l4Vgw2SS+G88RngxVSKAR04Tce4I3H0tGuSgAzl0K4yCpi2ILVkl0aKW
lO9HDGvCN1FJGZ0ZDRjqLGSAcUzb+yUIT1Eqc5/wGMT2kZ/EA+F490jbUp6LiEsTGqFw76QjDsOH
eMNfIc2x1RaaBe1VdU7agbzCnCEceCM19yrue7kyTAOLIZ6J+oCN92Joa9ckbcC+NkqfWAJ5fnOh
z5/zNlglE5kw0PFOBdkWmyBIbrP2VL/fELm0NRAU73u+eh6E1rLgkx9h27HvKvAyWDyDOwZYtXPf
zdUhQQqh8Ncb+I//3gZiOTG4OZnvUNdfsccQoU5VFDuwM++jE4KGITYpXcZNOLwGEyZDDGXrWLtJ
cUymWJq/xwwTTMe82WJZ1SOYiBa/vhmweVLOCXsnw2RLWjOMKAPptLVReOqAj8ZCcrzQj4OmmVfn
+J+rSM7FD3q22Lxjj98JNPY9jN1BlYqTP1Ay3dDSQS3xNq8QvgJJJtPjuUvfzGOvQr+sKi7R+oWX
C24SMiV8BgvAwRFuxbWp3HkdDH9mtOSMNF2dMdBXin5ffeIN6R+KUVOaYA8nQ5zwxLueyeenJtI7
H3hHqlPR5G+mg+AsGIFfk67U/VEwZl/OiLOyBZHsvXSzNHPi89Gge+CgKPBrMCqHigRJ+OM/kp3Q
FPEGoeLY03WW74uO+JG+Uk3wJ5aVtyP3ghK2zMYOY8oJ2q5Jk+3yxWViil1/Gmwyw5xSmVB6ZwjR
YQnVXBZB9YakDUv7NuSda6Ps5c7NgFf6Vt92Ta4nkn1LCyfbjbSk3StCyGjNI6sdxSbc2m+tmwHw
i9I0A7N5xyvoFRuulOzQnruhDwRL6yOyO7f/c3pCBJazBwUKPYZGhucYC+O0XZceyScyHAa3W69m
KED1Bp7R+1lFpeDi7IEUpzE2ZvxRGri7HYOWSaon3Ekt2fx1iJo9FpoCjrCDyoQRTEGPT90hVrz/
M1sfptEkhonvtjDpbYD0llGFTsUj0+TztUGDiR93rKRK+mckfGIo1r6CR4N9C35QJa8EFmNwO2VB
wv1lMSdLKj8pAs7lVcsYDfOaaU/rkfXLWVpEO1WRClgpjmfOjDoGGIRa5xI42tEID+r0MfgEbxAq
Yk9zTCpK9nmLmjqZ9zh/+ITV5iOHBy2iXrtj655YFxaRaA0xIUE33WvhQmyjJgFFFPleVnw+lDYg
oKEDQWvRn1A0SNMlEiinnVdBTaDpN+BXutcM2mRYocgYKGs0AjC0ATsRddrw8PaTkEkxkK12aG7h
GyYJMt24ALTS2xVv3HBWVzEGY7YpnMvMXBRS2cD+bJNkwogO8k+JbMLp+GbVVNZIfSJPSsUe+8QB
bwgzSLjHf4A9PG8Pz7blp7TahTsZIKLFAm72LYZ0yoYAt69IUqXTB3qrJHA4lMZNp/0zrSnGk4/p
TYU0pOO+0aTxU6nfo0eF2nTTnk1c1HZeePuRbuuR4TDzdNW7tzLe9aEkEqrOYcAbfpEd5KTjVREb
KVOTVtrJjqcnxIEqYvGyfsBi/XBr6avKdexokQ96VuFELLsHBCXBTRxvqtTg9JvhvYw1fkusJ7FT
PwQVmriOUBwEB3M+BJIJtSY4VEk7/KOACvBqWBMciBGGwEsyRKWsepLjuqPkAakDX5Bi/DpZi0LP
WNPn1+YgHFylumkrKy7SWHuXZo1kym26b1haI1aLK+WPiGDglPGmHMP2CLnNEeEZxnnz3HiKLuaN
f1Iq6SV2OS+8P/meeGX19Ac5pXz8ItE/BjJgFJnLKsE4U3Apk3yzLw8HzYQzZqPR1w8LmuPyT4w2
NYYz5QIVBnwSwP6ILn2s7uoru5VFKyqh3XZoPb1O2E1LmK0VCJn/bp53XAQQURPttDQdyVRcTIwC
4PFsugmcWSIfdA+Z6Z5K0mxbGhHAx4zEywECjd9kYkobforWTxVc8M1jRVC8XBGZdBETyBH8s8w6
VrKilpgn4vRpaIua6GmsI2jQlJSDi6YHkGikhuA97m2sc+iZVVlwXyhQAy8rCTBMYCHNOxPkFujN
KXaIawUAmAqFvGFPOLwxCeDp5jg6EqsDjiLo7z3Zj6TdqudsQxvIV+ZPeN2BmeN6iLlwawuS8LRh
i97nm1xvLOR85NmNqMLZI7YHCIQeIMqd9hSnmeeSQaRDeJuhpzYLumucEDpUIdSloUo+2mN6eWdZ
XSO+QLP3A2JQhioCC8pQdF0HOvR231nMb1hYMsNoESdYdCM3iX7vErRH/zJmkpbst4G1uRN2S9uY
KcY3DaNTQiaWoZFhIH8PqV0dCKCCcMTzY3kckqgprB2/UCnOL0w3tpWcHy3ydfzTkKLgS4aAoHQq
mOpGXlxtkoe5tsqDo0Kwf7Wb1FzKtVnrFU7/ApffTaphhrJbXjGXwKelhwFSxoezxFDz/i93mW1R
54HWWQCtCGLFGNZKDTE5xgtwijo0t65iAa3OucCf30mzgT64OVMv0PKxxUDbKmRhB/5gYLzXhvnz
wptxEjpoaXGbfI5El9E/9OXH/YvsKFoDeev1fwTMg6KV+qNsp7hgKCT2UPf+529hwHtMqMoZ4X6O
iWJwR1ygJsHF8xES1X0SDdM2tFrgn9/nZZ0Mp0xTTE9y2VSVeaoBWfozFHvD23HLI0j8tR4Prf0a
P7rXZGkC2NK8T0HaPgN7FBAEEew/37V8DH6QRLad2sM4vvBWjwE2W6W41LlXBccMj9qJeV67AOtJ
teng29zBBq5xpUPd4xyW2eJ9RPYeR++nHHkxm6SrjH/zHtXkEH/5NG/XaPPRRb+iTQJj3Khkpv/W
lohILEH5FPy1Vr0IS3G0x06uqxY2i/EwV9V8v1P2AtiqdgljBOSeLbLUKFak6dcPVjp12CGai3CX
ut8Al3Ptj1lnpGcEUjrPuznH9dS5HErmftTCBccokvD79SnBLy1t71y2KjrPkyTYb8OO+vvlJSbv
7cVakmk14U7OtN4HT9unDmWdDSkVE8/gamk1FGo4pNim66RRt2MMj2XJ0/lW+QofptQ+e8fvGK39
PzJY359VdNO3CjED9He2XkoSeQi/d+JmJ6Vdf0VjgzPxIHhxL+rGiwzsiWCgFaFrx7AQcPqhRxhG
vSRPPbVmKwqNA7eJa7HxuPtQrz8hLzddYNj8H0r/SNFxf/wYeS2gAOk3OiZGIr/t4IlShU7vh+tC
8S4qGXyUmgCWnJ3GtBpedLVhSBYsSJ+pvD+293qW3+NBatQTojJ0OHKokriRK25JqxOvAvEGc2lz
x/alStidcXYtC/jzZhG1+79rljkYFVpMnJzzSVH1evy8Xi6+jGnpfrUuo5NnO2m9vG2FMwhNIBll
Weyvi3bg4BaCRR3lPCTdzpMQf58Q8zsnyM7XANovsgE5YKQaN2B5AZtymQNMSzKOWyDAWhwTLrRM
s+2QVk3ilo6+1Z1pc4iI3NO8OoXFaMv3CPJDRWG+0mn1VKbb1EkiJBiqC5f61OwcP69ZAEsST8hk
+j98DA78ZLFd0zDXcK6Q7j2JC1IJnAs07W7oasSrJ+9nR7oVDhaSScAxN4hWsXRWaqa3y6TeFQBm
Y3L5oUZj8sqIxUAenT6l7iAmEe2etiWVRAJKM9YfAcmZu3dj3o44tXq5Y56m83Mdj4wbxQhD4bLi
AHHpkzxFompBUXUsmThAQlNSwKVFc2rrugdux1wxSigZIRmaCzLRZ6PBDXf35/y+vKcA1k9OLJAq
FaD0f6cAIilTT8lESPwn+MTbNMXywsxbUOL7muCqvyQ4gkfJlah5R+gziUO7CCPDS37xncuiXPSl
/y794bYdVmXEBQk0S6HIk/LGA5NQUg3QhMsrd0ZyChzep1mZfECQ+KkT3ho0xZ3O1klSz3kS+vhW
2ullka0fc/L25xcKU0tBFJwlfUIA2kOEFjEqStY249XP3exdbFkDn508LDEm0MHTZkvdn1iLkrTZ
xBuubXCUmRuey1YNtaUwzK+yHTyda9nGe9/CS39pnIexUpdpYhBGyp2eNfpibJveGxib0JgZec1V
KED/93kn9+QVGfZekyulYfWjgE5vyx7Zjp2msac1dbEMAfbxSdSA8N+s6vc7pZLSiMDJp67FteuM
vjjXyVJYzu6NJMdbnw1Yh5qwAeOMaLFK4GJVG+26QvkU4QRwbYlD+USoH7D1kjPnBRElofl8ouny
6LAu4SXFLOYxga609qZe3h8qYUM5eEGNTeUP5HjazOzmCLMakbb9twmEfSJBEOoe0LzIhLySvx3j
O0YRBdNqsyq768KnTSO1ZzZEm0qjv6FacwZe1h16bb3wzWSMHnfPIzv36euOxQYrljt6SRaDEFzA
jGND0cIjIvMlALIfLdp8okDsFUTpXnHMT8BW5xCu09yx0QczdysXZ0jHbt6Q4tKK9awNPv8Q70ZB
sz/S1Ma0ZImhqRBeBpQaks9L84dR7XMcYm353DQs3VXeOzOl5OI4kNCCVGcYDmFJeZzy/hIzAZGG
FENFUjMZd6kHfihGYOXb5Aq/F6d8kZYRngzFQA6HUgct42gwHIUVv9R3XgGFw9I9RGJU/xnwEUH9
pchb0lzqjfS9Nrux+72vJ144GOp0Ea2XG6IfmcYbOUGyh0pPljazUVxt7qL4/uvH26SXB9l8iDFo
349pNDj7dmCRT133Uy7+4PrRqS+CamptkXcgTgUYmh0+crDb1nPIhL4M7OZ2BjWgwlkAZBTwqS0Y
FwtEnEzD5fFHMVSAyqog0GqWv0Bu03ZO8Sdk9J69KAPW+SML4HkFAqNeJeLrQERi28nXiu9p9b5x
wYTR1P4bHl7Vsl6PxomQQDgyk2yHmDv+UlVFPVmueRh4M7RWu7AWRyhBfiFg8uoBPdy8UMZrXO8W
g163oe1Axvju+t0KZO+9zBzSIzuhX+Fm+oaCW2wVEsUHS3i/c2D7eWvn4HCRUif8FKQ0nmBOzQv8
WXEFhP0sqqai7l5XTzpIQ9XhHVbKH2HhN77c00ddP2elX7a08nn3A9RJdGeW+SIzWiEv+iIfUQFK
jwL+F6u0ZL6qd5jEdaz8h0aXtKceOafkjRKxRo7cnRAZUX8JmLJYfES9EUg4eZ9aimhq7TG6+4C9
t1nh0DfZvSWVahYak/9+3C6/QtVZQVxpJQV9dsVwSM8kHGPfKxyBBeehycSAzm2IULlJCkwq6gO/
GaS9DJYxXDovfQVul5kCIMJw62S5H++WK+zhqBQsc0LpaUBTMXxvl//NzrxZ8mQcIAULsrqftrRR
5A8JAC2Vc8T49qShs2TCYQ2VW5fIrpaXLlVPp9ApoOn7U6q+8eXm93cZa/WTK9DTGOzZvt3gWDhS
sR1o+AiBVIUQp29sf95pyOIwEVd5QcmHBxJ66sqzJTgHMQ/ftbyzpx47Rr4inGKTzayFkey3VG+C
PcTkESehuiihTpFxr5GcFrSKRJg2Ekwg8Cd/Y+OABfQkW5VqHp1e1xz2pOnVLM6maqk6H2ZenO42
nMqDik3XC8hdTc7IFEgDCFybRyvgVw91EKK66wIRM7Li6RjF2Hx1R0PFqFWBRY4WZd7MBJkkZHNA
ygZ5hlNviGjxLC3giL5qBMBOluMM/CFnEH/ETd9RiBTkShUTWZOxQO8fvfq8EGsa9axNUbbjDzYt
mK6CWCXtSkRHKwUkscpuuvZRg2a8CHDHQ8LO9IyOM0EuRpTLzaWGtd6tiJTWcJPhSJDnPfS7eRs9
LuZJZaPjbnF5D9Hc+M5KHxZIuzXVdTnvIyaS2qNJ77Xop/Htk6PNCDZXnm3am7Xie5ci8Nr9VyVi
11HJdg9gna1dQSX0JSec3yubz7UjN+aN9hjLVkowEw4HIhTo06MLd9jrkpOy9qsbR/8HbHWysVt1
I/HHuBul+1b28rRfJLRbpTOZMeaDvlYBNwmVzJxzQJwaBhka9oRqkModH/3oPCMMiYSZ9JHB9c5f
VJt1nHGjN1KeTWUJSOCM3RiBFrLQuy48CvMOBmLSFzSR2/Ec8EaZWHUDe8pkGK1tYAvukSm23FJQ
nOlCDxyxLfavqxyN3K5H/Tfa0s+g9ycCQNRRki+f3K6xzCeKDMxnPBRW8GISMwhJVKQdryLFymxV
QKyZ8gNEU1Bj/NJJE0pl3DXUDs/NTWGAXY7Z4APZQHAtAfR8WTCWwpb5xmOG2lgf+H5Wt2b+nuzw
eAJXGSSwjhMN81wzW/TBj1cy1DEaKcJd7EPo6pNfwPfaXav4c9gEdTf/vM32k3KAZ+EI+Gl/fbKT
nKFvG+2UTFE1XfV+uuNO7Qbq2u290Z87gr4MVwKIfG7wPnkfkIkUA+XdnG/DEb9LZzqHv0lH8QC7
NNwAxxd8EeP2r0nfUcBT0dzPlUVS63w8Yig8Hdx46gT0T9n3wUxfJ0cgBO0rKFpMLKoouS2wcVBE
gl+Um+o5blfqlvzArW3kvkQnELPE5/xiDh5ZLLgro3alcmhkirwU7goQ9BFDj9uh2lw186WwOrSh
iyQ2eLUJ/5NqGg9+zrHMby4qZiGTZN/7xd7qEyGagwdu5nxFObu33c2mBTsSHQ1VWqOwt3UGTjrU
FalrEp5z03Uq+LKWIA7TpQWOd3jcSCFNRjQ0hmUAT2Vnd9XMqKtz+2yv/ndslhk8R4U9TMg0Cdk7
3clr741VwDhT2UZPJCq433zVe9Ri265u3o8rQQuRVZymNAtI7j6Emdo3YONzoqaiUr0/Hm4gIvCf
ci6sdw5MD41icpEmGAu3I0m+gS2p49UUTrq9xXnqEGJksUuq4cZkCiACQ7a5ayNPqXKPa2kiuT13
RRD/7Bb+8oRktV2YiJQX94m+u3NXYjKmJSEEyQN9mtrwfXVJ1xq24RgxIbJFrAVIT17RyrY0ehB7
bdJiKmH68B3WRAWCIt5D8JoksNgKUR1MfpeWMmVdi7F6RODl2ouht3Q0r4h83KpH6Rw29sZW5t5o
+QtbcE2THbxcFtHSWralHwze984SfWMOiZEVdC2/WgZjuXSXs+kPSI/+/L00pxsfvll8nHGf476/
mJJiatZF03z6CzKSvjKHjlJMCoAN8cpK+kZ03u73F+MQa9ZfASpmC6e6zZ1Wm2EjpUa4Fund3RRy
GMw/N5rpqKNDbWFYjDgmQvagHPvwPB3J+X5UI+KYzSKErG5TkFda2M+Rn4omosrh7k+9jIo/Yh0c
VNrAUN4oi3MijuSHOxVcQ6Zm/SNKNIf05tqZYaNy6oAy18P/pwBQXmmh2QlZ4fJIHhIMtqGb2FxY
7Of0PITYgBHb4SuUNZnCe6X5zBl7G8Kfz4vJDPZegWsLe/yn1vlkBwgVudqLLb3UIT8LKdkytJr/
RVpsOKVkruKguNEpgG90grJFo57IsO3p3v628/4KRkNNwFBc5G9izJthygvil4f+l7zkaawDXFGk
iV2ld+9TFz8Jker6vUHl0V8wBZ/CZ9L3lNTREf6Dc5MH7JVMjR9s++EQVtI31ljkvb4rwtdMKUAD
iA9a97fc5ISFMsUUKX/q2eaxMxN34qEadjNPmjDc4aiTBOVO2+eX/+VLqFJdzc42or/1Xuu1UIXT
i9rEi4uwa88g6R4h1/J7NYRargTsczt7AwkauI6RWz0tU2sZwUg/PMQDkS+z/9uNHg8kTvcFTmhV
fq9pwQQt6zzlJCCIbATb3EBqsoPWvwZwk+rDQh7EDPg62BJwlkQu3zC4rwPFkGr53Hk77OQTdQ7y
ChSoE772YQPah1onrJ5NAsErqWDHoK4aCpHO66y4AAsecBQv7S4T3Jmc38/42GiKXz02D848c1fP
v0wxP0+IhtFboL6GcpSgMZ3uXf0Kkxo0Opx9Y33L+6Ynr6V1QPmAHGALeQW0+xXnWiqZSdjcV+yy
vs58YM7BMlXLF48au3SRLHT2ZbBHj3oQG4J3JhX5tXbNNeP5Y8je6wWX21i6oEaISRRrToN0xCl/
gVtBdeh207q6vLlOJPx36GZbRR9dFupIZcohPoPcDAxoxLUhA9YLYnA9Zl+4+oEetjdwvNhXr+gw
jRNjdcsRn9EIYGzmb2NcQAraliWfYA6RQc94p8Q34xdv2nZZf6eJfNDwKCE179LMn4mbr8L1LTVm
4Ie+/0NQDMwIh+07UFuOv+sBy6UeFL/ioGPOY6n+UXIMFdk6D5eulHOs3qOIb7I1bA19oKUGblZg
EtAPatCz1Vpjvp6lOU5ndHQwv01SeMnt8sxMuaRc/7lNo6k+ZQgzpf7ZKCqAcwHhF2hkE5rnLvWV
Zlgi1xHpNEQd/+2hL4g95VyGYFjd0251TUYzbHEO8/TaNqAu1PA4G9RaQVD7ZwTy8jhnexYs/5ym
sTEJ+pV0lB/omkluFLrWuzFrEPsFHiaYrN50FuF173lbtywkMWmjJcWREOVQLgRXmbPgbh+akJoz
yBuij/nmtJzUXibakhXH9LJzF6PAlzM1CvFOUzHyrw/6SgvxAkRywuv12tsjFZt/RrJO1G3eDRDy
3nSSbelzXMScjDPfQrDDlYgqsvgkEQVoOJBOqQkksepfWiD5rZljBePLz9l49Ef//0e+UBDlepJB
HAQhCur4NmxfxzbVM/gX7IPIiGkLTuqG0VXBvsEVcIxo0W+P90pLph+BZMDAIL70gwgChJT2W3hy
2LTDSoNxGnQm2KHm+St7UtMC6A/yz6skqbjnEVbzP0xCZYeK746fIAXosGcNZsOzas1pTcdqc6k6
F8Gr0rRfzsfCivixTHyq5SRuhx0ts7ywAXoHbcDU0ZkA+gj5QKvhOdLNY2V352j982QtF/JZO37N
H498vljxOLSvByMLViw3F1kkTzoRUr9gr5t6Vl6HJRLiYpnBhuS8RHuKN1mPt0cheBBFrtvdUYTF
yhEJoh8kncd4DN7cpmo6uUNBvbOpX+O8ocwnPytm6KzFNcDSyrZSkGyOa/E0w9Jd1INZzXFoHHx+
EyVLdxpFjRWf3xwODwZtxcdeGKDuk67bx2i2w3ZfbU2BVO4tdTfRZZwgPC/jwDy9VzZ3NJqyQXUe
k/MNan1788a82kQgvYJdj7ia/+DPEGG8Wd2tgQTB03xjlTIgVeX8Dlipj0ccKwDUzqTA5n+ZRI4t
LH+kAZ3PAESOxT8EvSgZWwwMf2v66+4RJxX9IkqRSHdBgsZP/YEZpj0laKdifYu1GoivkhkC6gZZ
R9z6J7Nhc8oLBZk4/aVFSORyv6336THjg7jiDjGhdDD9n/SAdKosUMT5LUSomYI/8WCbrB9e28qW
w/5K5wMzI/h/HaDiE469ALhTQFbcqxKLLf9umdkpl8g/loVsx4tz6kiBAuOkQhoyFNNFGj6zRVLo
ecWcT1aB5DDQBhMQD2Xf3Au0E7xYocSp7yulGNkmEuIlAohBAhIgn1/21S3Vb8M5PLDYS0LfpIEd
vvXb20LgvvIUy/42x5KLthOrl6Q/OE/BSAQbx8b5+F8igMm4torfGXkqf8emujonDUcF9judIyE0
FWxDQDvJAZrZWjLf07hEGmMUlf2exMWbJwNChaaP8IX5hNFrjtXr77exB/kR7NvHm4cFddSPfB2v
AHIzUYpVQSA+0IoKjWy2nSC4+Zwu5NCmIbK5zmE5/QRIEMUU5M5uYPMnvavBAGr0GOvytcDzFX9L
TaPA89oL6fAZMDf3LrGuG72gnBn+VYr7LP+lhaMkfxIkSwwDEAw0FAoCrHsk9vMJl5VtZXo65tcw
sLhHgiDsgl9hivl6gLkGPFMn+ii+vOjurYH+oWtmoJRny5geoj/OAuhdyjazLHPgrNmC6gyMwf8U
wRLm1foumjS5N9ggJ5xcobLZthW4Hn0YB1qhdaWeNCS9nOmJpEY8wlUDJ2un0CNLOy6H6ze7AfbQ
CcUUZ+J1NLGq9uixnSCaXRqTP6nhZMojw66kdCzqwNoPT3qF7dT01kTtKIHRR9VBLZKC2cT8Hg1u
d1HWvkmLHnCdMO1FXjZHTRkNV4hMANP5aRdVKY9YI/qoQvJ/TXoIywqF3fc/XzqE/g+0QqQeiN1X
g9FEe/+lxePXKhiw9F4q6S9WunYRe32czAnAFyO5KkNZ8/9LQhNT/QdoaiOQjGYW8RPkzRVS9hsE
vCaz4gmrnkTfKRiwkPnmI4UKoqBxxJxXgNIkQV+9AZ0Il1ju8++6DsEt/AwS7uG21ohG3LAHZ2iX
bQVds1MmK22VhvwjmvpfOCrqicv2OZwI0oUwfM2zGeIoWwPh3opgocUrJ3uDW6qvJG8BtoBqxn+x
NbI/tIaueWCvsePDxtbBO8Beh2PBzdOjMhFlRRcyjyHgsf4Gp3DNmZKEdTS6f5/nvTB3nDVgJiky
vka/4+d1ns0d/CJnjusBpkU2tL2GCY5b+o2yKoqi6zDzt0Pf2IAK94R+Me/vkB9uiGlc4ImICz/l
uFLJJ3Sch8xXdsOcICHasAsvSUc4aylslULqs5Cm0tnM7qSpaY3v0OP42WJ7Tj3nUrm2q+jtuFHC
kkCgG18Ysv7kyBmMBKD38dLXRlNElyyRplrBC9/RrMXD/pmdLH0mra34OGjZSQb8jD+9XPKG4AHZ
pG1qq1aeh3ZlFsyVPOq4gJjYbbVljiDF43ncbtuZJ03kmtPz6NCoUlMfyJ0/NK9XYTXfbMrrIFTT
gx0/NSQzMP6cStpDrY/sAeb8IZHIX7+AhcDsWIXCYdUL846glIa/nTAyGEfLdnFIHUkgrhOQZ8UP
x4aniJtxSb5C0MeMPhcv3xlEapj0pPQuNo221iMzUUx8XvAUQjpCD6EBknCxyRsJ8IXRfsEASfT8
SB5r79XKuL5mOOL+ZkZPVNwQIp4OJ35RlaTvNofRIrsT3pVg6rF083z9KAE7iv83YspzDKM61NNr
7TBQCa/w+mXUf+l/w/Kwk22ItGUg8CFGdO8ZcEzdRKFrkpXkxY4sDXWn0aFXirPYUrOtE5aYx28m
ArSw59xRp5VNbd83jOI2aPMORx/spVc3KrKWCM4eR8JkuY6P52hcsDKmLBxxzEe1Sb3UKlC0efV4
HfiuWwdOwg4ZfhE3vKSaT2QoqUN1yg+7zG0kmjcQyOvzOaBWjnSOQLxo6wBr6KgZVHWE6+/xkJGR
tbjjk+0k7M6bXSFuQIRDgn9YZhP3UBudQuIMn5ho+tO/9WWzxK0RlG6sUuifp+LxccCzBnRxbRkW
ddM/V94Z4OmS+xmeLw/cX0kp3qRt0eMBPOf2icg71bqUww80IA62lYD0FhVAEBjtrnKrFUUV7UOR
n8IE+9XK1Edc8CJbY6/lJgeOqwfjX+ach1ozgpBdFRpX4lUPw0hs4JfLMBFHZUX4Iwk2mFyjRZsR
KAD62GQxpQjLgt2QW5Mjd60oMHwwcTJM/3Y0TUqelTmCABIAHy9r45sJnl8X6CSxUvxP8yN+bqbN
y5IqhQOk14wLb/78HTN9mH8oHpLZ2b1wq+T0bTOJ7+vLfsiIcKh31WJCNgGxtLbIGVLnbbqa7TXt
dVOtcNYp7R9GTLaZV5KcQ7MtTciFNBrWERiDbjkeVlUj11jkxCOO6UTe9O8H1/I6ohOkEegpLG18
qjvGTKz7lEjg8EzCuuiVdvZ6TqE+HnsWiyp1xebyzK8cnieNIPb1zwQzPJlzXm42fL5B9xmzvlb1
tdRo+Kj3QJIyXr2mEOf/tDnBkwYsbGDHqf3ByEJ5kbiOdrMqDXuZTSB8he/lcVxpR52fh2JXR4Mg
5HMwt9f4wr7fbYW8xiC8pgvlCNRno7S/aDcDVhLWk81ySgKSTUKhizklp6D/dEhXSbG6zMezWIXi
TEiCdhLtxdcDymaxtUKFVdAtk2xPLHheLGk7C1T6/ytUoLdHUCOJdAE8LPlH7vpclMVG/+FF3LC9
GlwM9mdzxTdF9UON6na3nvH8+qQQuB3uaG6b3qLpur0KYxM0rkpvMcHREecMPYkLtRgldClddFmc
u9jIzSz+Z/97GJVqCuLI9xvRVGEqHqftoxegGfmMa9VvFEpkm4dxCG5+KMC6mqWzSFCRzXhXyOQY
eSHpRR3I+ZSXMBYQo0NNjr9DuRdJO+UJN6XPqqVLLq+TZhYr7auQFo7JX1a9GLmsb0LtwNFDXeOQ
463Z8upd1+kPrDXUEZ7gJVljrhMcarEOxXNKW7wnkXHUlXlN5TRui73HsJoS1DOgSDyJd6rFriqj
a9/XUqJFbj4vImnfGcanSJuHHcQ0wQc0UdJscCZ9GyES6zoeXHuj7mdS4tXj6j4Go89EoSdUJ7IV
kj0Ls55S7srED0koreOMT/h6PAUjJJ3O5VoNYtabZ9UB1hunv8Nm7Yuf5BGIKvEoPFG8FGXBqwWh
Bwpz85fggFpGMP4NdprKEQWOb90j0O4YyVykgSNabmrZMBYyrwaDFyzA0IN5p2ztJYVsNFVbiFRK
4Fatp8se1McHkIoAzOywka2qe2FLX8ormhlTPT0UyVkq/0qZwmTYagkdVgIlKBGKnzF/+mdAYBV6
XeuZdLPjATWQdcWOAKpgxGxQTuqGwjkDd9xEGPkCeUSWdGK7yBfHePUmvlyunRqhsl9SEAbVfVwa
C43/pczjkAE0iMGNQcJTEt9Gnzhad+d72GLNgBikFNNeeY98FiAQcni72GRJ8SEwxuBFfzghxajf
rTgzxJxFn6ucoY4vIJke+wKNztnTMTNu8Yzm+csKzjrPjknwXtZbeJN253YVWKU0zhUHwGw9E8ZP
HH11DCC6itjlD80gevxFWh+KinFvrItfLUKRU+x931/6iZYNZvDR5ifER3gK8wHJp/DUpiQtGEig
1X5BICRmZoFszXREXklWWG8AYfC2TEjapMEnoUT8zzrc+9fttaXM9vJAvroJq49uGzr8CxR6ppPm
8flF2If6fiDDdo/a/6mjl3jLvwG503Eh4QZDZ6bbIIrCEaKq9ynKnaH/2xZdk5VtR54HcAPZwd5x
Y4lH5CnJ12dxNfpr3WO2lbNV4l4JXykYXR5npzsw0RHfSopVbDyGu7TbzicT2ozlGLoWTnzNb6cK
N/oI9pnWreqKDot3h+F73F/f3z6mlPCyIOWAS9bKz0kJ+6ZHqThco7Ra31COyQJS9EMg3bHTOLn8
P47qwIyzILEoafHxKkxyt1GIboSeRtlU0rL/qiE1zuSMTrwClIjOsgNuFxw9JuLpJuWmdLtBm8HF
U65z2s30SJNwB9jHADc5Bow03gXCciMrF6q0tv4YiY+9mdH0HSnnVuDvqjb2v+AxNPZdsC0RpHjS
6s7gkTIWQiOf28Pkh1DmeKa6jtkCui0dr0myoH+avfOhFa3wxZZdHsAV7DtCHp5VwPT4mIypJJkV
JVyla4VAywZjNfvvOlo658bAUJS59ruRWMY0XMBgewLg9MWFG2l9LMUtNzGadEqBQv+Is6P4WbF2
fQ/YEjnnfDTa36qStcYWshukLsp+liw28LTEJKHtWjhiRkh17ZrqB8fEfSIVq8WC1gHk8XDNROvL
xQCGcaAhza8ZNTbLc0mkbej5aS45KxM+UBDiKCVFfttWXbx7MfH88khOb8OItCZU9gHmn4oSgXm8
hGY7VSEmGvYG1/Hz2/nT2C7/X3jXYFj7PtdAMnLeMgtz28Knq8/U+NMR4B7SIrXchC0DXwlvFfQP
2OMicS61GF8fqrdkSbAyf40YrCJeeYiDplZ2DwA64+MthXHDKFqaHNf2n9dgt7JKblby4uCgVbj+
gPQPOxgg4I+gMiQKLatZNAq9qZUJW6QTaIErOc8+CrDfdKCOb6yjLZQMeRyRZxa6Nnefqh0yAKVz
XHH9/Q79wsagyhSiBkOlQY/7bCsSfILpQvmxseenQBUY9/IdrD1Nta8E9FB4V7P9l0eGx19wo9CO
n1UrhyH2mgjBWRbTELRI3NClDCTE58U1jOy8nsNEoOnpzYOsYgLdQfJYAWulo/SqfJhe0brEl7E1
aRqy3aRDwWqgukSuqdx0twHqjWoRAhHdfhXNwfqk5msYVu+MFlW5fTd2ekJ/xhmgB/Px+eUpMq3N
IdT+Ngy+sEzKvL2FXWPJqkoGv/CdnqoK5p/pi7KM7K4/QFVnZ5UKbhzKUsEZZ7IUF8NZ6yTirPW1
5vQNmNPGWi5QJMNefb04vEFgu8noSPczFepp64m/7sQSKMVRE+n/2hxDLjnCitCS0X71LNHm0lBU
kdtty551ilOoaEjsUVwQ/DIUkNn4xUh/xjI42jbtBdG2BBRDRlfti2+oL2Pq7xbFi8YbWTMExejl
r6YsNE+I1UiweTgPjAfSKiKwvWIKFK+ldPji+yjSpu3w32jCI2rA+E5m+oK5vAcE9Q7Z1EQkiJxG
ncuQkBL5RrhipeteC0Qt9t3dyMdBVUS6mo+SD2BumvqDytmFQ5if7hSlFElSJ5R9ooRK+DWUez/z
Gaz9E5F1d8YX3XKKCCUGKwPnM81g/+7UJVz1dMNUdHBaG9s1O0UrokmR1cg4SFjdmRdhZRgck69Y
Tgt1QEnxIUvhNE4tA7o4OkIsOgMRXn4FJIPGA3FHHs/znz23l3oqBTwjmgabV2Tq2uZw0yYR7q0i
lI5IHMFyfyy+M+3xJCL+a/fijTW59/Cq6ONaUdOdUIxHUOj+m1dyLc+qqt1iPO+O1UF0H5glkbGO
OiM6YA2T9AMdRx4zjFXKuzimniGp4Do2dr5dIHpvHRE2FKT22mR1dgboPqJ35ZWKFPJFrbja/1eR
A6xP/PgwrohKHXenpUMtN8FIyv34LVoR1XwDx7QLRfQkSMzlEEu1nRZDWg4qTlCgCWI8nApc7Tha
wPqJyAr04N43FYKhRIKzGBF55rZbk5E2V0bp6WRbtme7swZYVzEG0A5fhPuMpEbsENAnprnpjziK
0IBDQ+p8gW38YG9rrbA8zKCA8vZepzxmrtvhVLgIFoVtANHDK+QKMYdbaWf3HrG41P06uVp2txZ2
Os1uqKVFikErtx/RlcFKjrvkO8Qduc1z9wWFdQn9WAs3c+2MZBbpM0O9mzL8u5RdjOP7DjIbB60g
qr1pqC/5c4zPXfVVWYubXTcrRssi+04fr7ZMLS76Z421Sak0lPAPYWhP20ejlOQBuo0WgvIc0cbO
7hQAOxI6AMce9j1le0ydkL5+dZ9wsNovTSBjpBwq03RJuFYM6osWoy5TLx6SGRyInvGUrpiLpglD
MadwmlSL5EtJc2PTPxZ+53LboruymKjP0hH7wTFgdrOTYl/2ETS5z9uBBpJz6sBxGGSj4uXpgCcx
lKdn/NaU9IsivKS6LVIwMrb69JzKlGnPIZMvItixAxhGHyON2tAoU1uwZEXGSZQfno+BwpauNhs7
tS/i610RMjeJdk0Cqld4LN+yhnYy1a30qGNMaY6qUhOFsgAdL9A5S69GTH85FXrBzcR+evKhRsRe
K/SRYYe8iXVwlQ3hyivpxp4zlNxYcKir5IQLMLdxU6mJHsoAJjbHc6xMTEp6VpP3KbDgPYR5cX5R
FX5GysRomApn65Xlzv01yY3Hk+T3uzkD0h1TPmkVEurslWrewKVDbs5Tqlmz+Vp/8p8p//u9vx4u
BBoQsWbnV7bMQLDKRDbYfpWXXO7DMiT7PfVwRjmSz/lApoRocPt9P+9kBPyaRCQEY39nQeem1LwP
i5f3L9qPGkNH4SFiZSNOvS+lDUD6S4hfHlH59ei7O3AtGoj7evA+tHbX6TpaU+4SwAGJmVyOfFoV
sABigvu08dG6cars1NDEtJ+PV8reX5AxOG5QIRUY9prsMNxk0bv9oBQYiPwsu6FR92Cvp8k6FPvw
cjxVzC9l4OWqdcwmmPuKXywcqKiRn9U37zDf5EMCh4X5gJ8cheJHiw8BMg+eKNhoyZXBYPHa52kf
lFjfTfk0J2HbzUIdIoOK3oR3Dus0mzyeE2hDigoWXDva2lCCQoPIAjtNhn23ixTVWfSBfpdb7GYT
3UiswYiPTGWVaqK2t46EheJhBZv7OcAh57pYbQO4QEzOcjFlXvN3/ajQtokx9K369LDaSkmG0ZJ0
h1QsKUPHLmiF9AthOKcHt27wtJHSSHQwXNkOaTyOiwbsQopdzAYSibI0nyDr+HWG4+XmPLF231Wl
6c43dfCMDx6zPJJOFQbDz6nN5gpblcbUYI9pgkB4WQZ4OfZ4mmkQ23h5i1NOaH78FwuJVUCbHvXE
7UfatkcohwvUA4DOjQeKUNuRKWdnLnrL6eXqYGFl+ocoYf1TScM//qicU8eZNwu3vpt+e8aPiRpo
rDOtDrZARTYK4ey9lF+X7tzyNoSxTsQVEQ4C98eMEKrGFoyLkjALV/MORKmxzZH7LXe3fQadSK7j
MqYF/ACgG/VNZ0sj12BmPBx/eHAJh/ty1WN82SFBG/FEPzdNw5Nf59r5SmeviWpW+caz/LF5jPnz
Fr/t6xdxVhYxHjYbjZAtDs6I1D0fv+I3xIIl7nDIabysnhoZUWvogBdP1thcENnibrftAUqpMIfL
/GrNQBBwAVa+zCLAn+wse9hhjhCTXpUkBqwHK2I+Sc8ygzZgEQn/YCQbAWEB85fn86RMGZA9IgFe
H94Y+Oe1b+HAtv4l32vWgDKNPU4kdRMCCDdNulIDFzCgsTpAvOYfTRHPXsa+QsdocOuvsu3u8R5D
LgAePbqn/Z2DaliuKuUcaVHdEQO9VjeZCG4sV+b8Q/Y/3d7QWutGHqs5soaj0Nh/Rsg4RQNyv6NO
3vLCmDALaV1PhlzYKVG2vpDYE0awkIqsKtNc4SSNwJYs/zkqZiyZoHlF3K9gbYuQvnMA/PUkOLJl
oOYh5gLewEvF8b1KSo4cxt3/IKJIByt2cR521wrmBL/uzeJxdU79fdCb+L+NjXedZ49bkdThHqaD
kq5vLV8LrePc9rYEHWLzish7wuoxIASGQ9LfgOsQC1dbG8/ZYoWvbpIs4SVBTGYx3s7PrjSF2Mz/
p3ofvGSVox0pB3inbKV4zCSziigIpvTZTpFaImo3hF5bEHp+qJW4Mq6VOboeKAHoDLuRRH0jJMT+
gTE3a4J04cl7rbbPM4oNp7yUx3BwvETf5RH9EUl59gDEFZc4MCmTTYdXCpdufpaHnV1FQ4buROAo
lRaCu/w8BZSJ38YJxSKXbW1XyMrqR9YWBXr9sgsC+06WoC9V6hWcEw6w0yl8yp3rH73gzKPrtxNi
YbfJ5a1hSekuBWOf1NFOhjMrzhCoqZpcHuILuqCYuhN8LjSFRIO1gy2bqj+so/xtJ03LeaiaRv1L
hHaA6gKIGPfqIIq3TqbkruJnbDaxGah6qlLo7wpvfSRWwQG11HApoYzolmjPaN0juaZesiwjh7AR
M/HrQnkTKxbdPBT2pyh1j2aSkSmgoSy05bFep2SEBaiy7WX4CLrHKW8MbjNnu2y94O9fXM+B2jWI
YM7ODyMZtHRajn2FjYPbWLRKysWiR1SXIoor9Lv5r1n5rW97xPCX9Z0ffTPXXOlNNbvbTD2rZ2oJ
0scP2XzYUBUd/H1YYBa1oV7bLyjKCj7v64ZiHvUbPEPhabgKKvxqyUTB1/4mBGV/TksjHdaYjHWZ
CG/vzy6YoWvNzOdLZ1AVIL++b7JrUZS7aR7JsAz2AyJ+kwidXgZwWqC0Xm7D2qDA5D/UeAftBXFo
zsqNamnSHBnfN487BNNMQX08N2EfoUQU22APan18eP1xDMPv+KIZfKgfWiij5EKGoOWgBCw2MRJl
3XLyIh+b0id/SapZYfIH+GpsB4Rpgw0aMkDZk4cNyb0Wa/2BL0IQT7mA9zpGtVlDoaUr360620qk
5Mao2SNH8ty0KUcFdiDYukQSKPBR643Sj2zP9gbsDfwRsQdwzoSS3Ht4XjmwdNpTB09xsnJjBcAH
4e+vxWBsEgIZ0YEhOk57U5T2TmtegG5M+wmXVlX+CZgA+Pp8ulMYyTrDXfo2mDCL/Q8XvnOrNHu2
VhmqprNLn+0SmrSHoUZm9/+z+f7bDgQvp7YStL68mt/NHPZG15ECJwVo4v0YvWS1NUsAH8iG3ymJ
KLNEh7J5GHUrVmMjVslZRLDrqyCr51X3hV4KOQebV+LGxPKanj2VYWDSRwpbYEfCrXEDAkIFKEcE
E8lprXGwENn6KUxB4wJiQ4FfvxQKvrjY8XbM23AY22Rx6n53WaGSrOoSOvQwTJuIDAg0/9OzU7hg
XsLnjH3iNNrShNrYTHmyt0epVOQZN8b2zmMuQdpeqB/nRjA1NMYI/fYZB7oQTCUQaDpJBatCqfr2
bLqBjOmO7C6ThCSTySGO27Hl3L1WSwIqioWkZ2DZsXv1LAcWvMoKCJMnctjjEuiRdWmfT+nie0DA
kvtyVd/5QuYatOLf7kyHhroeOHjuO7ZPlcJiTXJNnvHEOBH0G/OXYTRl/J4D5EOOS9fLK5ChOf0g
TzmjTZ2j8szb+ayvHOHkQ82kJre4u69pa03iqMPzIvOYi8Gs8noop2k061xGuM8fTSvoBPzC1slS
VCDEYE1sMV7qrNoRY9n7ycLJViJpGX6Wjx8GK4kj5L9iPACLqB7Spk/uJUm9eotBfBs6rLhmbWc8
bzLLU9/zBkZDThec8uJk3fx31PaQmnNY0Zpu1OPSGPWxxCTrnUfNsrH18BXy8nN4OnTVzYXT4EhX
nSQjCYmADvA2pv99j+M/py1TCtejixnR02rcm6xdMeqIapHJ/EbzP9o5U6SsaMbU8ZjJqJx6006f
FF0RjOTmQByrPdyLyPZAToY190Zcz0+1fpTxYkHRsqmtWzvDqCwXogFv8nREzpj8I30bPOn20gYx
jLq3Yf49DouGyfpU6CbC5hoL2nSqVZP0Z0G75KQy/XHDmQA5OCnS8vn3F6ggCQM9k/3WR/FcSgNH
11UrueReQTpg90yjkl61+tu8CGvDkmtaPuL2TJCl0IZyohSjfoyJTWazJxgoX6fDoU0rgkzgGIcf
caQ2zFnmCmYyUfktZLfeJAlfVTqObe2cSuT1Gyb+XfeHu4de7c/to6+0Wgm1EzA+fiUcLJdL0y7e
zh+prDm7DgbDcNDarSSJVaDYRP+TjNAdx5ZQsXjCf3H1AvPeG0LpfxLRQB/GCP3SbzKxsCsGNKw1
p3QP+gBz3YvPfMGfFsEhK2Or7NpM3VzD4a8KgbuQMRcJPoA5Bes5kUUFe4vvh8LRhkon5OZ+7038
DBvtDrTimDXpJgMRwjOKGRVKSItoUI/mXhdnqpt8soh9n+Wnn1FeCw8H1xUBtG3q1p+uhChVXzZy
DSbTvbuYpZYTsOg+TNpv3eVXlWk/NKYKRdht2M8CXnjcrPF5K4/Oea8smQRqb0liF4FeZlMcwSsa
eQM4HTFhegQpevv9ZwSKaYuJ3egBKG1Byrzmc462kIQ4FcTJGFSfR6C+oLjikxMVE3yx9kt6ByVH
XjVfmRSGkg1YrMNcP7zckqYYJhwBCGyCzss4CvDEEaaYnkDEDasfXCl6fSSpyslZtCAco7Cck47I
1VuZyzqhW5lR5C2k472J/0DDxTceE72zQG/dpP673LpKabokIvKi5N6iUbDxtbeLvhG880+03ajm
PAccsJOpyZ9DEirXsUOaf1OKSXtdb1Ns/8eYyEXVLJIbwGQt20jbMwS4ZpR1WZDNt6k5cKWAZMUu
P3yD+wO+t92DrTrVHQWQ4v+MdN70LqPY+Pdm3M+q1Hk0VhIbD82pQq0spKna1JXsYmH4A0O8LeO4
KuAaDprm1VvkkNEAXsBbP++BDqc4jcZplCsKVldLtep7HvMdUvbVM7sj0+beSSYaL3nsh0hKrQEo
3MI0ilkzA46ZPBTV3tL1/dCd4yySZbqU8OIGXXvUSHFkDT9u+VVUaXXXjM4Byh5EfOFrbcsKpSL3
GKUWjDP0bsfP44r05E06JrfKeMTw5Jdmi9vV+pDdAdI0icPbcwvH6Jr/rHaAQmE2crWJTUp1nx3F
zqPJN7tI74VHWuhKqaXhXTSrrf/YP+odF/xwMvnUJVHsEWb8YE7qXdQNUBX42X51PvxSJuee1QNz
Ifridk1Gj9wLc9zFehXzlLMcgnY7Jkg2CEL2VIs2hCNCxAmAwP7Iugg+/k0BRXMcWzQABDArgCGl
RlTr+/AVLC71tQ1ZT/LIRTrSqoVTs3fyLLVN9+PghEps78lvDUP/EfHlSeBwr0+UKSsaxDU3BdNs
5jifLf/n2m6lRFDXtpYcYqgrRqDmEuWnAGNTxfZ+d8VuWGaE+8hNK3wGgin2v2qx/Pp0F4uWa5Ll
YhAAmRcM9wG5VVC9Ah59sxMWZd+BY3rIownfhpK+Hg+3HPKaiswBZcxGTs9PhKK5QPZh8QLbYHjt
2kKUVqCcCkHNnQ1AqGGSYnW/JomIUVogcHnF87voYFIRWUCGpsUX5Fs+ol1WKs5y5YycofC2Z1gv
LinWs9uaVP+4XoKKyGwv6Dc4NGlG/AHkLHH0dx+lQkSdra87H8WzjFE6jd1/dlYXIxfnHamw+hw8
MyUziWA2++Zj/GzTNCHzwZc4vE9hJBwVZs+KPb7Lb6DRFP60+O2/CeJUOulQrK7pxsrmH+8bG3qR
iJubsUxtkmeDhCVz/D8093r94nKBt6QvsS0O5qp0apmYrL6EdehVUYLyUSL9FjYPA7Wfop87b5Ri
YRe37sdWPPwNw9qZEyiX3T9HPU/ZUOAVE9RWjMu1olKUK9KzsxsBZWX9SBx8JvBa+yRDu8DVDIar
LsRNNDytK9BfOGzqe6WgwHTeijoO769ocLsyjpy6PLSGEUHvNZeekEu4EIE5c+x8xA9ymoij+1Ww
Sr9tdM4xkCr3ycf0wc2AH/i93SpjqzaDeRNlMlPjMBsDIt29VcdF8eaMOXUz9cU5srIks4fiNe3D
2LLqV26XLpOHZmJf4PwvOZDPXceOVGsobBYWDhMbFxLiJdUKyRq6s8jfqSHGzMD622KWfRklScM5
xSk/zKfyPvc9XUSW/IpkpZCjvUOGxdWE/j2LzgVkuQoLGv3XH6UVxRXUKHAFgNDcjyv0gbj6SBFJ
UNjLJt/eyT9BC7FmRsVTc1bIIrhTmjVwEs1ArmBGkmYqtimTs5ZZLbKqPbnyIVQ1L6bab/+B7jF4
kmefINKvghIv0ecIHT6+qsZ81mnz1XOKZ0cU6aum7HC4PKi15JGflU2fYRwvOYckUxvS4qFhX0Vv
z73TqHmFKP66pQItR0/vkMOJ5QQtM/9ANPotzC01ZCzHo1+iqlQHLJnPN3NuJvvdHNY5vNPhOn10
gVjkPOK/UKJ42mOFWjplWsgBfebVVRy8E8p7X/d9A7Ity026NLBaumpchncZwAjOX0mTRSrLlkMo
RwyUZf5N+EoVZr9KK6k6tnKiDG57hEuYGmICqTauzisbRQi/Z+TWHIUSQRJ2YWuxSAZDKZ7F687V
GYOZ+l7IahTWRs34pHyBrnp0IFFPRAQ5A7YK+7M0v1XchKOUAqIYcsw8sBR/yfgeKJ/bofT2X9yY
GZRJVof4+kRuP0dINgfnejT/nhxoYczW5FxgNNPuhtyVnEVVVbJfri8w8oCEA3Sv4hAooo6fsqIF
JEafUXPNeX5odotu7u7YvRKYjU7ePHmOumT0v6xvGIprGDO4Ysq2h5PNa/gyzYCCfuBOa+Cm9vDn
bpt/9KBT8UNbcRzTessU+htoCndHO8/a2owUnKAxN0TatayqUmO9jitxN/w5yAzBw5bVbwLeWK9W
UivaMhRmeYYTRlpWbJGtnEhFyLD6wwV/9OknT4r2ijSK1Tn+/l6298piIAge4ZFxP1xZK/D5BW6R
eFWGWTU/PqqZUiSqmOOmyApTZtXHeUEsdjD725/B3gNz/FHYPbRV85LbKzNNxpgML5oFuF2UxSt9
JzZpoTcHmegW9uE+HHX6kgeaK+/eNM4kOrdnoaFx1JUKu65JNr5fZijawSodVXTcU6XynVRWX9Tq
dHFHrDAyUm2tHinkD1X+S38pEbM6j2OCL7Qt31+GS0J/MfLWfAIqTUX1hkxwd4k8j4Zw2xeaTYRa
5t6ikqXRXEEL177E7MtKNCDE/Qm4Tburryz8HCMdQqHtWoWjo2el8PCjXnhQ3uu9kxuKiy3iOouT
+9I+aofZD9cxJA/+1GlFJMQdYFhhlYy7BHZDCewf8QxQOYVYQU5KGNmCV0fw9uiPHikSylLnOuYY
u+Cg8BRA02HU0PY+wIfq7DoUAMuSzdFMKCih7LimfMdcbFDFpNpTRKp2stTSE96vXe6LiNu9C/KC
ZtJhTcLMvDCWr7Fk3uA9Bs9ahkyE3r+aJlNrci11NJ5lG6GNfc8k3EofHlId2myDg5TTLPjOzhmu
rmHcYongkVNvQ0pzgFM8ntWy8U7W6CIfXEPgdPilgsYaWvQt5VEfTrodPYCh2L/DBIQuSRC449FO
99pUkJyY2wpTtoPSqalAfWyZ2fGmBiRsn+lPMh7wodF0n3Ey9nn11XDQiKEoqmpl9NHN7Zi5Fmge
Mqr9Kl8qLyrzURaVeeSjNuF0IasVKKfNEmj+arlOhDe6a2x4uJnHdRyQWbxZGrBVHaIPE+vwqQrD
E76wPGl4T27e8kA2gPr5w3b/ms+M3/Q38CQL1QlZM+IP4j45nTbwhoD63KUJ1V1hG9IsENCzxVZ+
1LLeHcb9PFd3XHmoxeu3GxKF3okPGfaXMAq3/T2iWBUaRg13vLe0ut1AI63bnmSpnYOY1gHCjb9F
FkGZ0GxTh6CRci2/HHzvMqVPehPl545kMEf/j3kE/o5ZfQQTN8kQiw2NvA7DZlpvnkyJCmPzmmqm
71xDO1/5qdSaKJvVWTkRP3vliSNvc/paRVLXu2+3gz1RwbxFDwMaOx4IACHB97hBoy8fdXcNsq37
NR+0y/di15O1DwgbWnPdKWctuDCNHebEX1nB8Aeg6qz5Sgxakmq5QE21d9W78UfJOp84NvCT+XTP
gw/IDMozzH+WShF69z2jfXcqKKPuIA3jUMBYH9tBDo8nEnanxfdWTi70a3Z42eLmCndnr0ciMHKG
Dj/WMHL52f5YtKcA/qUDSd/fG4A2QteHQHmqmwbgzt2BFu2pAaKnvDWIApznoBEKDYP2Eqg+1Nue
cyY54X8pwy3be7Kr2Z4j7TG0cZqQJqdpFPhW+izCEj8g6hqawk7D3VqMqlbKqQQ8s5Bz8p+Izwm9
Q9Z4pbHd+5Uw0LfliAnWLonaehP5rCNy/xi7sb9WMX247mheE8sWan/r2fWfGflAsMeFREnPOowp
ddT4ENDSgPDatlcMAwRwEg1C6RH4fyMfFvae6YY51boN2Ek8dSO7AwIc3icR+fQVehFQVqoIjigv
vsc7zTYx5JLY5/Qi34B3KuoMmUvuhKqybRubYK5YBk3sy2COGGDj69xs0lguvFgfI0XjUmS3Qv+R
SJqkUyZ25b3tuZc2gpGis122NPiqQoPDscGJ46jUqYgELTxQ/zNs0Qqy4xUuh04JQqZZXIu2ZTsh
jbkyRQuXPS9K64d8y+T+otMTXkaoEw53SMGv9iy0wQblVxU6px8IinvPrAPsr5tnG3pXDciSpoVM
lYK503qQRBRID4ZrLXYx4OQtZtGzrCcYMszAYIpWUzO1aDyV2qIR99GcBOtYsabQLu0cSpHq8xTK
Ifq2uMu0z6RXS4rgRjg8eiYkwMYGGOMdikC9/qasvcK8Wkerj6TBO1ZAmp6OLJCN6AomWow9YDzC
NiFDOn7JXS/wisypDb2ElPi61YHEdlTNwJ9oIyquTMNU0D/LSPvNPsxtsYMBZZ4Q0CLvy6GxEo67
xsZ/kobnfM+B4TfVbmCystcULWPwhJ79NOCAQXCOXwJfF4BmnYQLnyM+t0lpTSqS6TqDPzDl2ki1
v2ItFY45LuBwZhOQcJsEgBBUUj+bRWhTmJaUy759Zll5Ya2wSSM3412UsfxK7qRkJ2nfQNysGzmX
8unXhAH7p7Izp3tZjjk5fi0ZmGvMS9uKWn/pQpF/gAUbBfPc6/eAj/fQ9fiZhT9+V2jdXv2jtAua
XnJ7bp+/Et9S2/wRfd5vZsMVaFfkdAv4dl4eZyZqYujQLlf49Lm27KnHNSfxXoJ01QrzIMXQSXYS
3/Sqf7W14FgysWUrGHXmep3ePfUgCXhYuJ+NBcSz3k6MYaVa5TPuww/DBKAH9Db8uAbVpmzzxcuG
9aahQa6nT/ZyVjednROejzv+F3Xv93eoIZG5Ixik2H8Vy9Btz7h4SghHKYSlxkZbzjwS5sMfFFk2
p48cgdMaT9UPtVqWsto1j5Q6LE4hEAzcSCBVA+Ejeg5LL7bTwXIoWiIp61E0t+QXF4uPcRoaFFvo
Ca9vsr5heTPXTtkgBD71ILa+7Rvvc3TlBRA8v+OnXoUMNDFdGFcE7A/39kiLny0+hj6xYke/h88v
sN1qJH9JmNKsC7TBVcTGqekaOewDPtkF6YcAOwZ0ryn/peHgrwUGn2oo79MjP9Cl7F7PBQpDg7re
eDWLYRLxvmg6wBSrzTNhjZAqGpsz2rUJ5W8KbkVz2hl1748lyt2i6NC6yH5DkowcTbriKDERB8Fa
XfbWtGg+B4Awii9qpvuIeEnBeKQtMzf1i1JREtRaEvifkpDA0GEhY1isXuW7o/qj5L30g7Nw9ta7
a7UeuqCr99YwiZHmRTtJb6sGrUuZgiApiqbhOcsvaCbxe+6faePIh/E9duKdlqgq9kWeR5Ny+uau
E5PbAiBQEyc79q0jv5w02eLD/cMbrK6io5Td+F7kkeWbzbJUAeUSpnJab4nL3ufPPdJdyZJPMlK4
X5SObUhq+FjDFMSuFODLy+XqES5iWBvBJPATIFXoe2O+Ee6lxb1nqJpSF27ij744apZNYaosp5Ij
m1Pg24AK0e9DJ/Hj0474wRaTnTkDoMn4hu6CI547C+QVXFem1THM0AYfgFAI0Kp2w26Rov1gEtyQ
b/M8nhLdZBhvvXVU3qQfoUp41tArMbakUjZA8X8a/C78+issTfcCDKH41XXog+wivk7A+BtbeZns
+9j7Wj2u4/OpVUDVKskNSAJmBQd4EIk3otJOKFbJ9qTbgrSotSrxtPIw+D7ldL7CYr5BJbPEJa6j
CRRh5ua8y6l4V0pFyQZrh8Pl1PwRYyCz+vDbyR1Lzx8Knukdp6jOUGWVDIiuqM8bNs9Xat4KFoeP
LI/FbZd4Oq/jaFnNLIfnn2VgzZHbKX5K7hJXBhPelrgdjE6UVLHNqV24BldpkMGw4X20k2uTy5Y4
2j6C9fMNMnCIGZvdEcDI/CEPSVcVh7juOIL1iECOgsPYXVDfr7po8tSw9JMkvA6NxpccqpU/cjiJ
7Csoh/Nak8lZqdLT0inzzCD/YmqXHoL41H6zP0Vcv5CT1gdu43r5UX01LPI3nw5oHpib4wEyLO4C
/XX/D+nPw1IVX0HeF0Hw/8I+uEwigDrYbis96I7h96SUzCrBoQxaCYtvmNLtbb9DYoINPRFqnv36
iJ7sfsI4ZLx4TGbFiEhl6nGgIU+5jfg2g3Yc4sjaGt0NRkNfUNdp7MsOkRkFA7ZoRGk+z/LCuEnI
DYRiHYyWjSDCjGXGuqouPKuvH1v+KKWx4BmcGpXkrfwjWcYPXD9C5OiF1wZAm5nswUiM/mpfbUAp
tqHx0DaFBuOm1hefF+kKlkQZvKKeXhvjWzWjlE/5tP4iJCamO1+Zj9lnJBwgO2goaTTkFxcL2JpZ
9HFo+MCI110yTLNxImFqlBYpQZ7zYb0M9nGCo+I8PehwxZMZQnoSo5mm61ySMBNxhPohu8qIvO9y
bxcpdxkDvW7QH+//KsZWaJMmp2a9FTG0YvqkJLWgypZshP4bcw9E8DupTNtxJIC50Seet0xzWO4c
AKLFxTLOppnqfgG9d84ge8bsWZLSz1pCaRVq6To+3EBzdxLi50Nu6GQzuJqhvrnMq8LOyhLGQsDK
FzJSDk75lJO6UkpWLa6y6E/IF7yF/cVnKLQj9sb8OrbXSK/Czc4laB9GGJDPzJ46rrAKMpRCPOCR
J1ZAzoSRMuAGB+wS4WyTJc8cs/QO/8SWwMRWptjrq+YbgXeM2OZ//pR/CTqMTucZqiBEWSfRuoGE
Hi4w1DQ8Zkh/2JS96+CjMwXYu9Ohx6xa+Z6yA2ueJ9K8KhbIz9ceVAdrq8OsOvNptjOQcZKvOjzE
RTFpUDSXhMiAO2YpamNnEFLo1ut91W+5x6eC/msBbUYz+tazoVjmor2mNSj5kVGfbt6qEg23IuE8
iSYcANvFrObux/TDdXpP/i3S24kZkVgpZArmnY9pdZQ2Kx6mMYU2QR4hWHBLFLOLofQyCiF5TRN4
asc+j30jErjJskFawGlomSO7ekdQ6ZFXbdq5YWaUyzdwAqsULQLyi+I6j4d71eY9XcdljK/a8z8v
G/92TOmVffoSAZXfYkVDsZvHEpgTWhrUpPcF8RA+dkWWDEtL6ycUxgyJGWpAclGeWqCI5DcQubvd
i8Fa15eGgyP8MRTr/FZlB2L1IpE2CxablflZXZiyC6Ir7wu7uezbWnaMN66ljZNKeQwe+0yZ9fT7
1/f7EC92N0lgk00RijYVXZO3Dyg0vAa10SvfHo3Xeb8+xl/Y/WSpMjErjLMRxZuyzKfJviWhhBHy
dAV/eXyfxhbl8UBtEjB0pXTaEGY7b0V9yV1zPw6VN/UzW/nYqcjefRrkjsY9J7LY9Rawac1BSEP5
XYrAcaTvos2bJJr/0WXmXm2JwpQJ3nLQB38TdUpXJZRbkeYj96U3Ww9CPxw7q+oHt0ELCj/wA/tc
CeClhr7SX5EvKsAvxPvDxmqt+flrz2mJFpDW23IWR/Tpxu0Weu1RWfl5JoRXqCQTuvJZl5xqUG71
Gl5OssklTCMAhOl/eq6whX3ET3fEJ5MlodEzHxL5h61NMI5jd8YGzkyhINZl2Gnguh6fRE7okr+w
NcP539v1nIiizwcqWJy2v+vGKMy+5PU/rF69s1k3A2EllTfbl/nI4Kb80615niLr6vv3RE+yHEHc
8I09gIU/+xw9mqIaTxghmiQDary735MCIPdLNaSYZwDEQXdplgV9kq6RMaxoRKj6/X5eMg2A1c87
X9r9KpSK6xlYbTXS/cXHS7/poboQsV06ifwTFkFpkTa/fU7XoF6+VQmUcJ4PHabaMZ+s0k9XL7gE
01a7k8ajIO72FCbt79ClsOuznLiQcnF8Tn/+Fuw+QYaFkcCUpX/MSi65CDTwVzONfy5zjK700Leu
Fd9eFcZbKA6x38eTsYP40m/fbbO6pkvrHuh9GNFxjU0JvARXTuvevOExlO1vlHR1ke+Lgu8AAIL9
FfViIEpAj6xcYf+n5zpu/BNluiUOos+DZKgxDXoAqL0Fn8jW215hmUpNUL5KKa0nTu96I4nxwGHk
jOLUfgm403T6ykGCoECvXdSyY6b4bb16ELkrmcV/DkGNZqWPYsJpaUJwlh++dzNgNxnqjGe2OMfY
8iH5aBAlOUYLMyJcNiJa9jKCp+v9Z7kDr236maXnTmLRD8XdatCI2m2GjrcBFweEigiS0B5V9K92
fofjXynrIBkYg/S0oDVavigcoWsliTu37KOO6QpoKc2fdyEUcK9Firjxk8KsGwT/sZhe1N7quDJq
63qaeRlnHERMvrEHJMKjZtdWQO4bmqGZyhV73qs1Km+6/uYpLfP676ebJVJLK2D7PCGOTl45bQ6a
GlS5KXMOOKWF9sgLPg48z+Mm9d2L/DYGtIvuyXgxdR4PV2tgjTf5lPrl2c3lzgLIpTGKlFRBxePb
3cdaHAPhMchesSr1MSLJb9hQ5WtMQKMjfyHMdQaWXk1ahUkVRViwq1Elbhz3ufA70ZEhVAdCC497
93cyLI9sP4/Q26iLmKSMZABs4SYpm6BKxPfUafPY0AgCyp0pol59VXH7YCzeHqPRYOduHLFKNbyD
LFA0TA6qfpOQbks4qbLXTkA0/Sn3+ZqpTTOt/E4Sc7a8d+BMV05q/Zr9Jg92OWg9kPUHBEmBqAHn
mHLIXshDauLmV9sKhwgySwdU0Fru9BVhPs1igFe1o1lVmHUbR2x8e/vjrt102WbGdHr6tIDuNL4K
acAsZATkFuFMN4849HGUn7VU6PACE/CGXCEoqmTnl46MDdK2m7OO0/+UuNi2El8scTdDo5rwIBcL
HVkt8olG58Aa49rrh33npoCJlxErUepdwEWGIhEV3wDyzkaWwqMUKkBCz6q+DOVs8hqpQ1553E+h
6p9aww7Cp/J/QCTEscz8THa64rTVPK0q0fw12fHpcmN0jokDEjY5OSlAPa2lAFi2f3uwiOZlcV3j
N/AOACbx3W33ABMk1oHI2zVndsbXY7/H2zkpPrnFi+1OvAkqmJApcDLl2OcqCNCIBrTYKPw7hktW
JTm7znwpr8X6PZzLkZHHiWoIzun0KLiLqMzNcRPkh9YXnrUBLrfDJg2C1DSzLq9si3fSO/QJn3iu
wKCSwWhhpAqA3BjS/rBHcVMc5n85yTB9/plP7/6eNOJS5kFVluHwrTJiM4b8fRV2Zuu616O+GOFS
LU9arw6jvDjjAAQn89C7xopRPUtz9cqS6dEz2ydXnYSNmgcF2gjVdSz1s7EQ+bG+ihfiPUqPZA+1
4Ua+mj5qRMukheZcCvLbu5lR3O45breu1wTh50gZDO4RHZSjE/GEwcsvr2tDJG1MrTTWDvLE16JT
IgnYNJ/fGK1lUV9yscXM7YDLHDsFcFAexzjPAsk4sdl/IQ+sgfzp3/QIbd5r/OXXRFBIEVQhvhqQ
efSZeC1O8BdqO6MFVTrd/gVkUoWZGJoTxcVibjdv6CldJ7K9jEtfcpvASCCTqVxYbB3ZKlEt9Xxd
PTZyU0Vlqhmli0ipG4iKYzWZ7PNdL5fATYKDZcK2H+kDw4e3bKJNrZFtMhWTT87uyXDnGWkVAvD0
3rni14pcyhPvuMuR9NbgZajMgIpeUPFj1zRn/Mm3mBl1iBGTsYOTgNYHymx9SQAvVEa39TkBJBZX
dUYSgJIdAsCrSj+i1DV8M0nRB352QLTsbditFgEIhEEwFCPlYygS0KMqNwTOa2UGA7Gbqwgts7XJ
s8Vo96jAXNYn9CeChoDtkv/nMZqH+2xQrXzauhc90FMgGv+r2TuwYgBur0IUgYpgO29qLMcNhqSJ
L5iqgRJHr/3+bFEHC72Eg9WSfrRVYG+V0l9+9coq5S3bfmmP1GN1D9Sr8N3o69oCohpXO3HLgm7p
qrWjF5xqEfKcsG7QjX2QGK1Cr+VJSSfBiJt8cYKKLSVRiE+jXDDy3Zr55rSx2Zr77W25vDxYaWZu
5ri16svMbxzdKusqQaWNwUUWercx8AvEBRcMxW+UlHwHAGaOdo88ZLJgClSFvbZ1axBOKqO0LGk6
iTEEfMcIRXS8REXzE5Vs2b2ROHsmJlFBl253B/0ICZ8Ml1P8t3n/zAsTvbhbkJrIsP3As8DsGlfY
j0AN9My+a07j22kmPXqpxG/PuVK57sN7+YY/Ua8hj7M8hFfLDsRvf83KHJ8CkHUT3IrlDJ63hAuN
jtzZlAMmblBUDC2PcFMJvecLMZEguYF3bDWJQ9aMcI7gVrMD0Qcs1gbXTXFOBPrXReUiNF8qpc7l
Jt3tsm9YdDMsy8yw4aYJygBvO/V0k4JGSmOkbYqOWtD6UZeafv2PM96M19lt2AN6//7UPFjeQAaC
O4BZHj0dJUICyMJ2tN+nh6XkenHpS8WM4boMO1pJbUTjQ0xRGHkIrgdoSKqSJqcspJBvfTWYR8XQ
1N3WiuPNz9Lf0GRzDS5gHK4g4Ml+A9bSKLtu9qw/Wd75WT1AWe7nWBFF26/PyDCy16amr3bQHZk9
efIKLM2aDl6v7nJlvDgEAxmFAh+Jrc4YKvGPxojQBbgahv2iAnTkzsOQMqNqRBPyEGUKMCqFLlbE
oHUGYQP+FepALdqLoabkRETucWbckStVei1Le5oQzCfdtkf13tO4sUFAV98l/xT7xcIBNASwfndg
ucAo03bUgS5JZ9/6YUJz0BgbbgsSVrAR3KhT6ewKZ/ihMZ98r6MSS1Kgb7DbvMo+FRQtF/64GwJv
Uga0x8bj8+9YlDh0nMhVUbHpKo7yLH651T3y/ucXqJ98QPNNFchgXgr8xLe9DzRku5y6gaB71HGA
zkh12t+RGWWhj0YpSb+QSd6e7RVtTLH/evBB1RHQRSriz3W4AR0J5DHxoBo+WDrqVFkM4DxS4QXE
MobtBHaiNEjR63CuNPgdP7cAT3peae/6zSX8Gc38Im18mOtl3nA38M1sNlIKhK5DEanH4evE4ooM
bdeNdX9TQvbcDM1KM1RshzesKzjs2vm+efEwPZs1QJv+jC+bvC04nbg8Td8QQ5TpXijaFEh8YnwU
50f8DyQN6nA6ooCCE4X2VjHArmIbNX7ZacQP5GVI7+WBaIGjNjWy6dSK33ty58CAy29W7DOh1mit
NDiwHZhdiSZIsNe9H58DJ/dY8gQnHLfzCBQ+jvKQg/vxe8f4F7ckCD029yBksluGKVgFGGu8dMQg
ADB0oqV9gLHVD2ic/NOYw0ps6NtQEPBNbsZbEvEdd/Rd6g9E5BFibHlc0nZphHPOtEqGSO2iFhgB
X65KLcecuMinR4ogYHvvMX3QKEN4MSilalw2X4ryh/9653XP4zNgc9FeH4dWJL7YDLaOLyKmV60b
4M9TLydtn0/HVwhm1hrZe3YmPczsY2Md7jJP5Q59CRpjfzBJRlxvb4XCvozaXuRP9Z1nWKALd33E
h5R3NlfCYapK0yuo+8R82Du3TwIYYC4WEGCkm+0NMJE6sY+DzKW27/jvYmH8bGVdMks6JlEChigN
KfgVrKaqhtKKb06YCxtL1iS29ceD00Rmvb1qlvsGR2hPlwN3in8FEkWto+NxySbp3zNXJ5Eb40Wj
FCGRudai3EkaLw2HJjI+L0js5p36GfPO60BmdkVEONirU7SkTkasOBwxkoEg1pE5ZY+byqKIgMNW
JDyXtajLjEdsP87twQ8lby3ctQx4vJS8g6UVNToYvMqmCMcB+BCnn7fFfUxzZBNIZO4UYDRbsRo+
5XuQi6XV6XLPb4b6whr1hIowXR+lHvstxMzjw5ILPBAq62S7d9K/Dk2duvC+U+CsYUdZEF2iqoW9
Ph5cAgPxPkVxU/gLchQz9rCqLDPKVH/HNS3LYSPvK0VW50kG+lh22HgqU+qbP36aC6XcWygtn3SM
jF8QSegnDE4787YVqDYXd/OSEN0eSMk1EFlfSoa7ts4n7aTLdozwnGVJLR5cX1gfzlfhKxGNegg8
TIF5fy9wRFeM+zQ2UfnjNQNO3Vj0A2LdBxMCGSvWPiFv0JZDQypmpdPYu7DY4Wg4VusVOTcYe5/a
T2UN4HHPWTkpXxH4yqwUYKOnmmddjKFZtZe2x6phOw/VrK0Lslhjx1osjpKD+LreWdjw/B/3lmOt
onlLFIJ6Oxa0/qr/bdUb8zfF46L+PFFA/emaytloaMwsIAl/Go6ZDIYbEBTB9vxcTOnmvsGvr6Zt
jcqQSHyScKyArAYkpkoXqkxosB6AYiCcL2dwaZoHIrwSQmzTfSj8gKCW171MO2hZUzxj7bgDbB1o
2UxxNFJTha4gSP//7ht5hFG/5pKgg9FfktTIuJhmdkAJ+Xo820UPNfjpzn9AI5ZXTkqZibhpnvOh
xBrGI13sOQKh10/JrspMNoW7nP91FwLjZNDWeijzBNP5uEv3PArYJBTB1krhBMXettSvhUKbaEsO
LyZucMI1Vsgq5VKxoZNbP8uPazFl12uHtLf9Hjjnp8T9e0R0LJuy7cEKTe/ktAwFuhUGDkUpEh6R
EgtF9vkDGiheUaA1bNl5IBejX+AvV9QXWoPksYqFiQDtoAoMAX3bVs7KZqZ23YrIZAEJHTauWMlT
T3W+6TV/W42yT674cxXf2r28c5j3RjLttBOuKnoj+oD4xWKnx83kaD76bzysbdZepk7H792CYNR/
uz/RVYebBzFJn8HllMHAi8CmWoHrTcW2oYxHlYivBoluybPGXTBUim29pCM57QxVYrhhc4vJCmvE
vK2fxFxBkS6MIvc62TUmmRqJR8YMuZ+Jd/QTxo3AIStBKmNq5LAzU+eS52AlNmeeNTEzFuiwV1ja
Dwni/7aO7B819ZIGyXw9d62CK2JgxKEB6C1M+HtqgCyx7IVZRU7HkKFSiCyMX7k5fo2uNHaX7o5b
2Qrc/6ZpfshfRC/x3SOn1y9Nxr5H+RbfkDBysnIJ6tCU8jEUpotaFfDeqReqMf88730nGJJe9zph
/b0sB8HDtdIHXAPG/Ca/nWBgmT0TfJZaUnGX3T4Bqhy+acSNtmcwo5ARRwORohTtwfg0UY6CvzFN
L8iUp+3oiabkzZfmusog5sK08Dnpj8aAMM3abLOpxQfKy48QhWifzIO2Fk0fBiY4M2FaKyzrHphD
WIGtqXMe7VNlCF8ozGkeECZIjXJcGHNVhZu1XR6XS6fPCpTmL+3TWBHlpfC2ggyuB0c+0lLeYO9u
ox6SIbH6CKuecPQl/XXpm1VKlWYH1kcomUQupU+yviwWGb9hMvcl4tMHzOCGEAbuvSLFTtDt4L64
J9AKQbjBfDlyRs4L7WIrEVxAfaxWv4lJgbg3FvxROzKIaNZy3CP/SS876HytQsqU62ZPE3Xlgpgt
0wnTtOFW0sXiGEcMjwJgITeUubn7EyEnSkMJmgwGFf6J4BR/YA6S/OCG20ad4MrR5sTDZq7+MJoS
X7TVhHE0vNjYeUK4RmkC6YzisNqV1c3ZS1Yq2OSxFmnEUo/aprgJYmMpIwQoNg2LEnyLuwwbTkbR
aZqW5gi+KA3+AQvKe37GsK+CGWtKKfDhYE72ivms4g1dlwGOPMyohcIC9PaMwWF8c5xRsqdm0gFK
m/UVW8Zt6/EQ9NXgNr/Q6EyM5umu+1Gtucb5QQO4WTqGHBfI+dtfbq5n8+VM/OsuyPJ/zMlJYG38
zsj632U71HwwjzEaM7PC/iNwVN7Ijq3dpFpEsJ7xnbAPKWEE39NuuLF3lhw1Cr4qH6zI9jjRtOnS
HOuoHt24cJ1NEWj35F0K2aJAEsK9NHM2QDeuTkUPplMVOiyIgYEkM0dDZplbFC+S0O4KGBvxGIn7
W0141KMkOSTJNvUdriYp4v1OlJIpwY4hj8IR1DrhWKrFCnp1UXZSU+SrppakGlXwQZdJlpC6mNY1
hZ5icOnjjl/VF7z6kvn0ACjzgUgJvYJrxpUf8qjD01swS2qiMS2ESIxcR+Z5+GoyBKK3XoiWkJy0
pSJQ/29cYK7rKNcUehezIImlMesBh6GY6dIL+V138f236M51vPmjcB9usVVFOq/czflt5YbQMIsx
N3y22Ik5g67yeO2+q+tvgj5B53ghEIYdV1Opf8LzPeDg6/QuW+I4TXNUmFBterpQFFNvAQKYk6U1
s0tR25HAIi3YV7F1eVn/WRQDoOSs7NtrhLvqLQ4AZlqTGM5b1DASUVZNU/ZLBwVWOPjMk4yD6TFN
XQV+yYrkGCKA/rHCT+2HNbhfMFmd3nYwYHCGQ4IkbC17DicQUrNlH4/Sh+rW5ukOtYcNxuqJVxk0
xbyFCmlRzuitTqd1wvD9NA8QWeOmrrmKXRS2pRcj8FSbGxOL74zRZPcjb2ObhXErEoUZDxevhSi4
wOt2jCaWWuR+g1m/ZdGaV992fa3KG+aT8Zq6JI3mH0h2XYvD3v7a1pE7SFdUEamoCsB5VDqL9tk8
xukRHMGSFYnMvU9RNX3o/o0qzp3HjwUEV3uSCpRXQBJaOvHXM0Q79q6pjmrC1T3SUFvBdHtMN+bH
tY755N96mKZSrRtqvSDEjPQL/5jnNuz5JUan/Wb0bxuPJ9zoMJHyXwiTs/JkSNPqfv6fdf06vUWn
qOnGuyIQItQRgHV1JCB2Hpb8hK5XSOB3sYtu4kVE7lRx0iS/9Tfx5pijvUHss3mfHB38evAw37IL
jEekJQ63mF+j1fuyJQdvf6DMD8gRpjeq7VvUFDPLfoJWM0ytN79Q9DPmn4Q6WUt9mRu3v/vYD3qD
5ukwyd64n1K1yifBDkfkgtxqx9pf10oGkZoM22A0wcQFScEZyNQp7hLbHMIsSVv/tRektqrvp9yT
b4HAwpyxTs6l0HNX7/u6/xDqsVDYYiYcj3EnrehzDXfAFB0DBG6Imrkqe4dfo/jONxvDZQaCc0gR
RwuSI8vlMdEA9wLdZoiv8ojqmI7KNPj4w8fWR9ZgpNa8ZdEAH50QAxgTtyKRuq5IWQ1rWR94z/fQ
UzzvNdItokBrvWD4uz9HouV92LLdBd9ltU01itm+gSR/ZeXGn0LiwtcR/XsE5oNMkoIbf1YmD2Ew
TmcxuIXSYD2AAjj/eIRF4+/qNeoTQwaToM1a9ZTHOltiYM1FyYxma9K5EQE3eqz+Cx8FnfACfkVu
HkMib8/vM7r++uPZAsVpMu/S94wxWDN4u5arARjGT5rgfqgI4wUh5dOUTsoJ+rwFjUKGpF91bexh
kS6vhrWiqN5XoHcGNFK8H5ChCaFwpAoAY15LWZn+0QSMNkyrseeki3OptT8zlNYuWVpAFcE/tETy
Yx3Wi3aGOYv+8Jzdo2raUKFnzRnYi7YIeDYORB89vvNsxp2GuLBtOY2S/B2KQFrxahtDj2H71ml8
I2krqGQnFkRMD2dzP0f1B6kfPg9Qi6GMinG3VhqDrSGBIK3OVs/bwTSJmPgBVTZFE0AtQKLlKNC8
IGwPJ6/7vq0oumHA5TEQ+GgmzkR/jHR4A2qc00V4/4rYaZJGvnzSCP3mBDxEAYS06Z7x0ZVmVp4i
dFD5fkKSEif7BSEQI+YOmdEaNbUtggP/DamDdM1tBzxMBT3iO8rtlh2Bchm7kFLIVFh0A/1Feq1I
T6vxr92zrrouBsWfiNUioyZRFvCB8cIJ7gF/3NmUxbwRsDY2KwUUKiJwSxHAbYC+HO7Z8Eq5gpo1
Epeyd0U/+9E0SQDtg2T96YS3QS0cVAfd0J/vDzC/1g4CLQzkArdtWTDkJYuSWPovMkfMmdOw1uIm
nhIiDjwqVTMfPcZkW1P7cxGDe5tmkQ0uGwMNp9UWcMIoX33gOGurrQfbRvfxN2PiRe7A0BnTRAgp
ROMLIkj1mWoSSYnWTYnTnQo8zGID35Dlqvxh6tlE+BwuocKaJB4cNyaxpTGqsi1tPF5ffphuf4tX
xE1HblhohZKD5U33BUOqvnAQNHBW65lHz0LPtW+Pr8aKcPTLW9q/Cd0xUE+AdqWMjwGdQ0n/nu3C
N07/i1emGIeMA3K3uRuEEC/hhzsf/pStMkE1Hl8VCDS8+tYTxFUTdb7LDpGBb0zDDbJANXoHqmtY
cw6EhBTg8LkgnfeCRteei3RpPmySyu+9qOc9o55QdDjKq2t7ZjsCGige+J1wCeMRY1Y4/chFJs1t
eLkV2qSw+HAvFbtSLHfV/fDZ4D9+82PHWrEH5daLrGptWFyWO0u1as7SAhMQOKmR/8hKQZYvxw3a
7HF9798GumgOYkiQ6n/lmW1sgNSuFnQrpINYauKuZxQljGE24yP1zfb4dsxSL2c1ee5pZWbXvMh4
tvwYsssZkGhwLsYhXn/Q4M+SIxj85Dgk7G4elLNNdsNUWPzEnSTiLlp2Od25i3BdBFJOMulErI94
mYKXJZhMoCBVhNoyYTk5gpS3H4+wOSkOT5rP9wFFQEC7DY1O3VtXA9wohBCzaDqymhj6+vUVPcR6
h8/hKwqzkmFaIHthCUoBaBeIT8pLCbkh2+8WjcEOO7gIiKgzpxje62F7N5YHjOuBnBzXtHeOLkeF
pEywY/KLGIbAlLtZ1d21no2oTyFitvPXdeLik3Sk7CqW24FMqSD1bZKoPXyhTqmoFJolWAWwSKxI
QiHtY/IytnC8vMg0CDWK3YqT5nVpAL6vLFaxpbd+k6/saHqYYtqKfog+c2LBWqWh6IzQ9+BjlDgC
3G5kBQf8zANpISjAVUJLFufyB6425+hQKZurD051qXuBDdxnoSV+U0+w5WPsL1F37o7Sd9Ubutzb
NDr9MXNNw/wd+UYMWdeqF8xRQleuyyulJ9TcxYfi/QUS+zuJfVNoXm1/f18QEv43n6lhTIcRPq6c
AC7c988V9zCA6Oe7jI00HkDHbQBsMvZUh8/ZOZWaJ9jIYbJ6raXdpc4gnEEI3MUH6ixeypPvAnfO
W6P48Er13U3o1fKzt6VpnLHQ90ueoQE3/NeeSiFYoRN32IGXn500oy62v1dU2QD2Yc6EZ46ugZ8J
Uwn8JBDLSLQPoUNFyWam/o3+MeeArEUh16/cYMjBwnku6qjJuVTnuG5sNAzHBF4RPpk4RX+B8qPY
mWmeNORmsGbPt62lpEpkZT7ZGP+9IN/sczALqlMyxi7mIzdNzfERljG1A5JdB0Z0/xchFYV7dUCi
DD+Qqzdk673o/we23Ql4xm3orG+QV6QO3/wSMshKjbYvzntDsdJr+mnDE7S7svDYWrQGWvhVYj4/
6/XJDwS7PiKu4lbgIrN6dZkP01auxtaNjEmBuhobdA16qFTXxg6Dn6WVMDOHJGk9Z3M0904dnlWW
E/KXXOnAotFQyc7jwvbKug0SJ5Qr9Wt7iU7+UWf95wCcG/y47QURCnj99+/oOA8VDlxKaPIL1VzF
lANJxOL7uNVZlHbYwtYnT9EpUbU4TXP8tIq4qcTswO25iJfqMSwoMRlswr//oDAMFC9VbuJp6zN/
H04dUeDp8/+JM5LeacXuWfyqhkdLiRr+PNFrLuh8A1hofQzDVhFi8zEZgntMaPIKJoJDUMIyeqKL
hHFGW5wi5nA3kGjRF/Sz0d9jROTXlfKVbBne+CTwlB6xQtw0GjDytsN5Lnuq+0rAMgSducmA2Cjs
/NgjfoZANpjVnYAUOPcEUVm7d0muWVVvYPHEfjc/psSL3+vi3+XWlS0NgiePen3ZJjQpfw1dzLxg
UOTCRXIapaNwsj3G07Pq+pY/cJ5g19iDxpOZ5QJKL6ACJBM+aE1swlnV8eRTwbmGxhKesstlX63Z
H8ifx8grMI9A427dznEdLakHeT1gCMzTGNd/4kqDgZhdeKFtTIQO7LOf7mpCwfDeuHA2gT+OhSNr
/kpcopIDfUFSs9jB1o/gvg27/H1xZjupX82yGqWY1xbmRjBhrv0dWwErbUQAMOtWCYE70EnoFd12
nOZ3A4Ql8gpulPAvfCuZaz84TK6vGSgImaKpGqpqbaovQGYwGRNSQNRXaGrjIYb3zRNPuc2561fn
cFQj8B5sOKBFshwQZavxnXJustcASty3rDgFGj5nsX0X+Bgxc9z1ojwZwqSTQ7hJRvjQBYYKrZl0
azoe1zLgWNNC2pu3iBDhOnDaWkYQxDN7TP+jASDSjciWuWE1AAG+X+2r9WeGAwvm2whqeawF9KbW
l/PATuEyLftTTzbXmoMaIBTGazpe/9/R/IiZjGXymDAalinxj9OqPKzY6Y4kZ44XOvrUbtbav9ir
hbcoaAp50YLPUzS5RF2adIOrPzaMxcxppllhj2lt2GqyeQiMDwshTyvCo1BOBiEJU3RfK8uwWDfX
VXMmjPH0szIMDW70o03Uc00O9VgPzGcfm0XOZIGd4ubIkW6yNf5r/fXG9j2LWjTWT8hbk2W9uhSo
uEblZyzY+7hHHvW5QuA7GhN4r8naN07fEoBS0xjXAaxGDPbzyqpsO9/lh/LCpOdsns1obZC5jrJt
h/sSaBjQQenNRIKTYj/j5E7rsc532M1uswQ/OtVRbqSkdYiYV5SPQy9gQAUlfoCXFBBZvhJt+QNz
qg1Fm6SAx7luxjHXmwV5Nsp1vnIWSUlsxdCel/lvkcdxRUjTfiZrMrd+0KK3YufhWo9ewcXU5Up7
d/UE4mqJXspp1KYWDWWbyffGHBvc6CC8+syWDThbJJUG3MsmR4V9N2GpNlEgviFHR2CKsD7Nb6IU
lpL94/lXC8j3CXJPwN3X4IDAKM80RpC97XZqXBb0DUVznEJKtV1J/zVwDb770he/7FLAqh/zKy17
udt266r6jlxkC99oH4gbp8r6NAmAb2eQYFzJP5r62Dkar+kNBBc2PiGEiffb/174UFwoGGuDm2/A
515/5/8FMN9rhiv8gHDbv++/w6so9p6qai7ZW/1WxuB/fa8dOrKDC5Nd3M0+khEG9hzp6UAwPlyF
OjInmgDTmi6URYpaWCC/M7mAtfhfA/OBKm1UvGxJm4O0z0UopFJ6/AcZK7r4lqrBEpyg+F/QiDkU
cKDDW1h74W44MJcNMtsiULlSnYWVDXv0BNeNomVif1LgE+MBoiGcUgHWR+2xk0zOGf6RPX2m/a28
QENAB0mMTsg+8mtISVnpWLMCyL5T5FxGcystG83vw/jYlNZqiHGVn9/feD6zMe4nKXsR5cjZMWyq
FZH6e6HBHMLGmWv7LpU1Cj7coStM3JSn4D/lYN4D/7NVPWJaCPe0L86+KoDnThOrf8UGCEMKMlRM
zhmGWoaGo/IqTshuGmb5zuJJEhe/a2INXEcFCi2qabxdd4Acbchc5/Oz2Z/qZAA1GXB1yOEjVDle
9nU7s+PD6WGaLapJar1hOIi4/JqHsFbfySFcBPvwDaHt7eheGogqzm/Vs66AZwz0wrKm2bECBDec
FccplnAyNt32I6zxiswBUuLuzC3cngybrpEJtedudWhRnVd7IQdd5Z0x0K9zIJ/WRFNefp3e8BmT
9Qjsj7Pn49s4fWyDppi21IzhFk0IPUOEGBC9HGGI04ZBGlHkgLQnjLYL8EkfTP8NEE7wvkPA+FXx
R/QLRw6ot163yvYG38XV4qLndt4WhRbK+P2nQ0T5EAghLBYvKbIhgkqRa/p0QohIKeCJ6g9bcZea
MOIgYRVVLzOCR06P7hXffRPW+N+ZE400C0FWnlhOngb2f+bG1+xph2Mx9HpAW+ZNXg6GdB29whtA
2HrST/nza1JMjJUTVzWxYC25xmrCQvdnWc00j7GdVG7wR+JpFs4ePNl7FQqa5WALWjh0DRHQPC8J
6XPTADuaEmXPLdX9x7vE/v/oIfmSTfka2blHO8o7Zmqq0LswO1CxR6sk07Eij8C+RHAv+tiDcvNx
vhBetE8FNR4P2fGZ0kLjIyRiEwy8TGIduUndT0S1A5+gjwpIl78o1j1duzfmMmOgQXMtp/aNINCh
ezMTjBuww3dqmJlIq0yFJidiT9BGlLR+6/Z18RWU1mSn64n2t6RcVn3ZZ4zmVbHjJ7rRLYM7X3oc
51ziN8u3mCDW9RUFlOippYI+Naw80vFyMryFA6goB3S2II8Nnwt4uaIR9GX/zlj3NYx/EIlou+dc
WUxDlHHi5UGS/OStrKg7DYaAVmWQaAPJtQL8A3AROVKujrfnGR6mOXNjuSJK3qVCKCXye8zM+a/E
hf8Fih2yrSoGuFd3aQkSURJ6/+PF3Hfl47VsXPv35BShc5vT3iVJS7zv5emNbr9+D7S37UVQfK9f
dxn+dAeKzNdgi6gKoQXCgTMnFoNxVl7pdCnuRc7HUI9QmJzKn8S8gGAIqclN8zV303DjKAGcG4bB
aMQ8xdxonFTGXTACZVPSVnIRpCaRtnYhyv9Fjh5WHyhTZ61EOhBcNLWmjPCu7BhC6A6FPx/5YFt3
6U0j4vN5VTdFx6TK5t+boHo+/Q5CjxSVgjVwpscMqZx/a6q1DokYYD+yu788BnoiEsf9e3F8INRp
hA+1/hUZArEYECiYaPBrELU0EkGN5phrrd+w1J5edp4l20yFTWkeMba9ILCwNWMhzKcpGe33SSCH
rUhgGtpRPNuc4EpdJtTHi1R6+IYF2atA0+QnkgYNKTgFmemtexzx1PWlDoDCl4tYGka1h0fPZISZ
AhBiS7NxAhkThPafg9AcewXoeMrf+/wpTnNfyMl3OlhEfGS85vKkB2QF6fxP5uXoOWLd8SbvvB/c
z1Wn9J6u2ng5oldXGWJUZA6HJXNEDDHOhg4wVzH0VUCAVKv3Sd+M7sNaNIuIGT+jI+luxBrjOeCx
xQpPGMbeXr4a0rsc6qwtnqLkfngnbd0RLsNcyw8qqKSTkdc7eN9pU1iVFB3ZtII6US/egZy2NZ7i
bcIKxSUdmgv0OlQ9fzIzn/rVS4gKi1U5e9ToNM+KzgIrQKYvNhmagPW9qxCV6Nc2+hwtx49xEcZF
dzqG/W+uSks3Kdy0TBlaBZWLE/kgXFIqp5EzoqnfZLLbNHkJQnYcq6lZIiCKCq4Iv3BwRWxvxkcI
FRVvf6EOO1bsBULRy3hvpJqHxwnnhTU9ClpQreVQUqauTo/WM+sOueuVSj/jddLwyDaabgRo/50M
Cr1/bWBTiuRY+q86sIBr3vLgug/q2Yl2jEb6Mb8PbwxzxxUGI23NvDOtmfhqz+q51nba6tsTDLPn
1zdO5LHXKgRuf6zXELlhaQv9mN9wkkh7lJCvytDz/0jqFmzc64z0yfW5N9MFDbzEZ8i6ug1K1Coc
I9m7aZEFuakDxtTIVlbja/bJIBlZfnUxJo9nLJpFR6Z25OOqwYdX77amTkiaIp0MfnU8soAO4d+z
VlcoDePXjTe4WEcz9xZ9/LvUPoyJlznJCRMKDy9JNKNKj4VM5vZjEW7FMyGNyZzSwN8oHtEi8VKU
iyI3bQCwRdQ02sN9W76JzQlEhMmREcuugBHHl3HY7pN50CMnvIQFWPpoTn7gGF0xJ4Vkds3FiRq2
+rAf1OoBfguE7DvknOXmVEGZ9dEYmEesvvEIc6GZclkaWkQKRRXWwcmsXvCVRimulIenCkRWXBbF
TtZ2qaatimisutPArBiHvzdVMBvlAc0Ib0/V918vrss25/DdKvyzUCxiI50z78//RwIj+EpDiKJW
ZbsSkIe/PGHlrELgWTJ2GPUTXXTt/RnCfwAC6OVsZsPQLbYK8c+XISch58bkjDOfCCwBFNY1+CQ1
kTIx30VLcVysCZLXSsCx1sr03PM1m4Z0v4ovmJ0VTeSgtNmFwqpebLtfbN3sQbFZuKYUTCOCBVNi
tWmOCqE1V+t5Wl3DYoYhTSPW2G8DXqkN1ENct1J3aRKC2qtmMfF/0QOnMfW+873HiyWB4VK46BG3
PllxF4c0bOCuJJWdZxtziIm5kKMuubIaP/2WubISnopsPN5Vod1lX8dWuOVG6V0lDYx+GMToBVuE
WuoXZsxiecdg+HR/NskrM/g5efS9wxM8b0PMuojTWFugYZ3siJzXHMDEuhhWTA9LX9MAe8QrH+n6
AoA2E+T31K+dU1KgDs4NBtxV3UPp0fy871PKH/bxKnWb2k9u3k9B3h12XvGJkE55xQ7zR2o2OMIO
3ziAO//VlvYcDuynicf+MCFvz05Gackv383G/haEngtyWnHCyR/1iEydd2J69pdEvdvQITkc9+rk
hotjjmStCIPL9X5TEgoglQlSE7c/ggnbStUVc8+pBYK09VE2cjLX0UtlTx2LD9aZk/734K84pjG6
z/8jdWvv59ku8S+9SJ/APYwqgYDESdc0Gp073oGml4xCoAALJy40YKCsb2Sx3SsWgd5ts3zrntnN
S3/bhlbO1hCV+4ATRgUI5RO1owEJ0Ydyfurtwfc2OdgA1tN9goBAs0lE7ipRrkCnWCVLIsF5LD1Z
BPb08XzlknElXgjatKWmbFV79e1LUroGsvx1kSI1BT9CQMGo/xKSIptecgG9ytid+xcArsQKLnp0
dHOlGv22oEKbsi4eyaGLeGQYn8Pt9Twi/MfX91gJLzZziIu6WjjsIS17/6nGfSH10ffzvqvA2lO9
ejTZ8vx4lBhXBAJvbcflAb7KmTwY9jFTUnFyrc46jYOHiC6HIZyeoB3FSE/3ipzaMSEFP5brOMdv
PqZawCu1vd1CPyxHg8bafj9lBnMG7GS1KQY64PYRLa3kY42jxXYA64ZTe/qUhmB2bwvAGjxTB4Z6
6FAyJbGT1+zdeqwA3Ez0ShMt4Me9p6N8HoKvGx0CnQeEscpPonltj2/zARx+gPzT8XZhiPywsf9y
+tui2mKckIfXS+5u2NaRTFbGEgNIHqjQOXV7kZcnH8BFcgq/ohFPqqEw9EnM8znzAFGbfwx0zGtL
jDWzCJEoAxTx0bC+gtcxSbSv4HhNtSsz5gkR5MmJP4AhHgP6LwhmZky2xy344O/CBZzWcZKX8Anp
ElnILGzVDhBK0yrto8rjuzjT0QKXmuHIf2mtWWD7MdCc63pSzkND7P04zEOeYcf0hAnZ5aUYqcFo
pSmlAYmZV85ZSbiavWPOnKLnG6ltb4ronh8ryG/xDI2Af0Qyf7IXOjLNBvCplqhrt96Fg6Ye3dOr
FSt05TttHinZQk8yl05b9Kt3IugLluOTh60Jpi6UuKuACcAUm+Ji5QRjKlUt00ndkIS8qra/rXwb
qnMSq65l4p157EWlnjEQvzUkA8rDr2pT0ocb+eaDnIqU8LoCv5dBhk/Yv8bVdeafk8Ob4kegsQns
wm+/P96btaJnlc0Z8DXzN+49JA1QewNYmRmS1h1O77QGq9kA5Ly5HeElxl580faOfJ5apT+pj8E9
PO8LoIVWS7aGEh/7OrTEuwen3TOlGM+JJdmrs+utoCDV0Zy8K0dUUUZgrHyeH9u7HdEt5Mx4bEf1
hyunsdMyNgfkR+orogOwcuPiJ42riPUOUaP5CCDXUNQCjGtAEi1SbhunYbjJone26xUqYAY4XKX+
4ZIOt+PkQ8XNER34iNopeGrDRz3Fb2MfnXzAFg3YodxzDxGU0IqqD3vvwvOWMmP3VNVGxNyVa3pi
FK8gHNfOQtwBm9g2UNN6xl88N1+qof13GgvpxenfRSf8La29KP3PutspgMCSQnoQ9IcKzWT5OE7J
VZ332vsuzaaG5ewZD1LfQOG7M/iivSSRjHcfKDQRyEsJAToU3yahoRHHaFCwx8t4Ur6pO2H1T+xl
S9RFtf0o2QBNR9EbyLrCvGdV1zPvUBh65OaTg8qNbjmQmke6Y+PM1vzhspYJGMY3KN3wPyLxO3bC
6eSOV8YAZuJ6Vb2KO3yMAJWr36/7JgrSvKIgiJ8JOddll3gJiKeeaQve7mQR9BdkkTpztR7Bd7up
NJ/1Z99rE5qmjbVi8Zot17cSIQ9YzHAcLPlRLB3q9oOwtwhLXc5cbwUzgQaed4T8sf4/IVcGbqJQ
SoCbvmGyovJGtx72IIi0DYOohipgTVe5QRKyOOFUccThmGxuQawKHZp6TrbBXGdiQDB5Ft49HHyS
1HDRtZHRutD5Rfjhbci2i3xgaR86RYl36tdYFiof9uKIIhf3LRLL7FZFlhotK2K0bP3jjbpGwmWZ
660P0VaJNubrq6ZbdL5ctmfaes+cqcdkSIx4xiuc7ql9oDKB4kck2kYM1ymWB5zT1v8JP2ebtpK9
Owf2wBeA7Gf8YHUc2XYxXkOzAPr/rgZRh2SXjJOI80VBYDuBrcV8+SIfVhsN+vwJtuDZCDv+U7TM
SDc9H5JK//GpiZ6bbOc/jOoJ1JVQ0o3fTPYfyd7RCObKue5aKG4MWZs/ivLkt6wGK1cDtSClVAcG
O/Va4TlyyG1DtuoUuCduwb0FCpECpe3rshruuXz90JcDIs6L9tG/yytFTYYiMP9iW0R1T0pzL3dE
yuxVyyOTiWXkLWe2A8wOKM/MkJVadGj+py7RTFAiui9ROG1kPGcYRA9H26w/L+OS9ccmFYqUgW5/
tISFqIDXMdKOq+HLEVNfXv3iKQORv3SeDA1qg2Ysa9xsBgIRqQiHKFoilUsI2m5dEla/LGRhkFy/
TNgQlc+TI7Yd4rP0jzs/v7KKR4OmT+7KF7sL+CY9q5/MRRiRC/FqNKEzkbIfAGfxOh8wRybye6mz
Y4TTKmZXQQIkxLcIjx6jqRWtoE2C6eqbet49fPRCxgr8+JlmD8qCLY94fUzykuhR/k45wPlufJkU
Dny0rK2LWTwNUoECSP1IA6n4Rx8cMB/2OwZxDs1tkcnYFIYefE4jMi7ZDDc/kXH+K89zqPHylD03
Lnod+6l3+sJwzO6IeVXBMrom53AGJFKS66obX9uOtRAxq+gihvbfKV6xeqMnQUGbvjp32ntSVUbj
z4890Fzz2AAi3KGFXMwzm8fFyShTmrTI6P62MAycY+qMIvZMz0a8gOjB/hZZ1KO5Rbpwj9qbWixV
sqeYZxY1P6nKAzXhxEpia5ipy3En0Gd+ERApbAMGzbLBO0wy+2uYUfOEPYsd1x3+P968uWFkNo/1
/XUU8vqSri6CNUf17nu+/ld3prn5pa/xtene4Jq1BDWbVrdnpWBdTDCMCgEX0zDs5L5d9LonRlaN
5Lrp/w8fi4Rw7HqmmNzLEtjoAiOx+sfLW0D7jMK1ZFP03dOPlpxagUcexbwvp7n0kUir4U79KkYi
7LibhdswcHiEw0tMGi7jajzsC5Kc5kMTwVVtgy17rmwFHFSflaMRdlmYXsQk4Lna29Seb1aHJ8AZ
cJWS/M1uyK6nnkDXvUTwpw8yMntsb4Ru+J+i4e3iYEr/uZHMPKEnr9ADhHJoIaXiT6OhAP8T8SCy
9iEkCimx43+P4EibLL2Zf2OQsbQn4iNQN0PmNiTrL6nLgXrBcQ40luYENp+oQwibTJlqeMGQ1qzI
MmFiJr/n0iU4Ehii1pFQGjF4xUQx31nR8pmL6eVcQJ072S+NDgiIXhmDypJkB23bNI94b+j4VAZm
inhZMykXBkv5athHgJDIhVK+0bW4J4uaRdBziZeoQmUTA4hMTFcGxH6rxoZglYPgjUEKZI2V5Fd+
Ivc72T+uKJH0lxCg18iFpwfx9DgOaYNqMUVf7A+n1eSnI3g3CO5gaaD8kjGBpdaLOxNj+75as085
8u+y7c4PE5mCxmh5t8p2dg3yfplOdW5uUYyJXbUokZPOe7xjLzwuKCdEwJ37V1vcPBcSdRZn/z30
pJVjaKAhoiKLx5J7CHsYih4Es6wTLVeo4B/jZE1qXwklvOgm9jHBvU9gM5rKQlTewSNCKkaWtSik
fuMQ4SWxkb1VVLcGDgAl8H+hsCDn3B1HuiS1iLltJK6jrmGuzbJsHEoDO0qIMmS9aDID+jQ6F8Xa
7lQd7TClnraZ5ewMXzeQfMGLS7/Xvu3bHa5nWmeJ+F1JMcrLtt84pjwVZJQszKXp0znqujzj591e
x2iG3zf2Jdu1slcrEIDDdJqzX1pmXOWK9j8Jcoxcvj7pVMePrv0nCgKWTFhuRac6qUSqcZSCYA4a
biCzYudeFpKpvrdlR0fY3sDIzqDBDhMbSPx8oRLcWfJb/g53Hen7m0l2VJJ7H+rTsOOms27f241v
elv0HcFIyLujcSU5xKMzxmc2yIBaEpMXj6byMa9Ear9hWNR31nOhMy4QCyN4QWpC8Du2RmaXwaHx
dzKdI+/cPjhbeFLGmogAFu73KmlxSn8X0f9uP9sIhn51IunI3oXSUYOi063vSillqIW6TXvKKdom
YEqyl5t1Rx+6co+35zf9JhV3keJeSc/zMBXLTnRi/MvrSdKcQ/XJExQQgfFWkIzTSYuF6t06bqAM
VaR2r9pKOPU2GpWk6JKN+dCiS8BFz3Lm2IZi2UpKwcpLxypw+vjf+2Opvi1LX5j0qiFyWuMdw/7O
Q3z5fhWk1GAKcjr3wtyV+XDUUCOQ6ru3cO9in0h+zOYJ2/CNq7byIUZk9yQL3Ibg6lSgcIMS6UWn
OpkircqG7R1cLBJobMHu4vYrvFNhHiawVeuqF5DHnwEI/p4jkLPltd/hkkj7orP0K0VqDPts2nvN
unGCjP5rY/LO5ezpC71Fz3OTIUPurus8/kGzj5ypnJKgreOg5dF8+kM6hQTGPNkyRby53DxwDNzn
0ABt5QtUvk8SZC7BjJ26bqkZGAda7st8FTJb57gp/EVpXzlnwTyyul4PPfSBLX4t1A9VcrQjj2RN
VAvK+/q3o47gy/BmaiuWZ3f4Vpy46/pHeVT3U2WBuOEIHDHXOk2UcgwX+rZfFuGmDa1JnndAt3gH
Co1l44yP2K9TgFBnvbmT2lnOKd7/9b3g/ZXEGIchHOzU9ZuCxf89HOLG8UMzN3ciSsGeUfIrHytJ
VcszL/+ySGrKBHFQcTrHhgcQMGqQ/VO408aS3bjr2UA7EPoljpGewbDkdSE8+jXmpAaf/6raCOiD
iLDdkddDfde0UkMDVGfLN7p0VNazIM0lD1qfDjVrRLSplaa1Gs4OuRq7kYeQtaeg/7Bq4Ow5pd6o
EmjVqo73upWLbx7IJX4EOKzbWXLJPYvbGGV9aBe6Vl/e/rx2ObPePWhUhJLTa9OC5rRrfEpcueIm
iWm53JzxE7i4otgVT8V+yutop0dGEphSdS8ZshtRtOMioSzBdLo5MIMXXTBZUidTo6dyehC7O1Fu
yRJnNDaHuNLI/uHZA3OJ56bpFgLbuUu2Bp0dbzDQ24U50+/dr3FHOIQVUAnD79JeneF8ikA0fkbW
fRPorx/2PtMJdiCwKTNkRpY0jcCf6wzhw244a37E/tUXtu1ZUP4grJwYZidiJgOVAEWDK6a1qOTh
YwtPD6dX33IF9F3XcTzW5wMhbq/bYgmZ0asNn9BDs0t+93QDV4JbILDQ3tbYuR/Bdjt+DHfqCEuH
CxO4Qp6Phkup1QDjPLMDwJ9FQZ4YGG9cYxp+q0cgTSWFa5Ba/zfG0TZgcvmUaPFDawvJKwQaJ9pN
xLLVSbgFjDOen3J/mVu8iU24SE1oXqX1B3H7V6gi9tXvOGQuLfiCUd4ynNpWHcwpEAF4/1p8FODP
DSqQxmb+UGIUPTrEypPQ2nBn2PfAFN3/1whaYAfcX4WylN+w8+3kzFPviDgl1JcL4RdMmMlTsaM/
v7tVeuWMmQi0gCUISkzeom6/VIm82WFZfQ3TLqCCQqbGqd+OGvmpi6gu4aOADfBVusE+R9x5SAeQ
hdaDWkuVWFuriEySGW4c7WuV/TgBCe+2NWj2FTASwzcBTZdPf+/uek/edEcsbkkanPmmoGsMYFgC
L3WmBIyiIsGOreEhDv6ZGD719T/+ZqMPjygrHbJSNSBIR49eeg2l8GCcqgKBGvxfHRoFXa/P7a/S
LeW8sZiQzLFjixrEwCMbRS5oJk2+omcg3inC6Oo0P/U15eUA2puhRZIkz/WC3xAjmRse3LAvj7Kl
9z8O6gPjt0DOpMjadO3zbaMtQrpoUdkgjxiJYQrQh2kJuAv8fk7Zmm8ywGyGZKqFn2TCkzzgoN4H
eaNjDd6ZChgJq9qZ3M0I6wLXoLMDGP0CunZ+jhyTB5dds5pltuRQJnehf3k6XN8Kq4+DRJu8MeD+
sBAqYVCbaY6183uJGpLUPfDNGpvTAOQGmNC9ftTP+OM1v5OD4K1qoZ1N5OiPCnzG/BwQ5VEDqTEK
ypeeBeALG9nuQYmZqtQOJGOG7k81CLzvPg6/lAcjjIgprbcY2wVLZ4r1+g7OUzQFmA0UOLXz4YIr
HwBV7wQrWEXTgLzCrkY0XuRls/NVy9UqhBKnC7w5xK+vsOWqht82cRomV0peZT22/qIfn1Jngovj
qMOd4oxHhXllWs8shnxhJpc6WcJfKcxsFwLmdYp5N2KEsi3ONVIMa3ZwtStnDiN2GeVrpX9xyLf8
GKIKfleXpb3A2oGiQKWitcnQZio105bhNyK8OUmhf8AHykvaQO85x+moA3IFRcRwhSyRvtG5OihM
EYbKhwVJvrplXSNLmvgGWzH8+H4pTAmS+KaeSd3RTi88XDwqZkG4CrDlNNlmh2sfiOlyR23KCgnc
Bfnvc1J6sENFH8wbB9sndGA0CjBkLK4KEBDXrF1+gsYLi+T6CrnHOdrDd1QNcqBBPyeS4qaceVso
IYWR16wXmboOmSN4kX1F28ma3Dx2z8VYC5tyVJs5mxKn5SfriNgd2qaMtUuRTk7i4/kvt8A4LRHG
KmN5ZM9rX8W5ZiVJohFgn6TrJ+dQlantnhWGbNWj47aEhhezAj0le54pMAkOqcPwhW3fJ4ahSm+Q
s/ncG5hX5bkBEe5Zo8oBYEsaMh0PY9qK7jBljv4WMs/uQ7V+/js+eVeDbU4gHj+3EJhUSGOIisaa
16EwQ7p906sArQxoddVgXtIJx9ikj8WZ6GrcSeIPdumKxm4CARuyI/QZJ2pTW7j79vSq01VIWDMY
+EAbrxwZe03ZT0TefsHYBWoUJfbJORnp9dV+A2b+ca9ZRAakADDmW/Et6xuVMIlSfpwsi3shg+m2
HpAtdHuvbiRhWIndM6OpN4AmtugGJxjPALFWeb002XytCXcVUsLC3jmOTWT5FFcapvRvT00WY6F4
OerVVonIYJh6EoWnFaigmDYk0cGx/nxRBAkbIg9GUgPj8wGzxQ+vEatasy2TKS5qRrBTiVwEGtiw
g5Mf2HEAF8Z/3HEBqLWorCr3DnjzosF1Kk2sJn6A3Idp3Gbam+w7shFpwsQH6hZhZV8cJRFONAWd
rqmQujAbrkfHOrzwtViaECWnvP7JW2KLqqxei9wJ/Yqtr7/Eflrhoxp7cO+CMYIbvJ1C9EYKyMUm
Q+DA8YqKNxcH/cTVyz2SIbH1btAXqk4xvDrB8rddBqaOAmTqvm1//vmDeqHgoCoa6vNUxbq1lKhN
LEdGpWwwW8byl+sogPEeCzqBiQQD4SesKY/8HWSph2+aKQwxCdapWDXcOVkRQML/YCL+9qK3339z
SK2BhJ5jvZf/3+hoz9rLKsxbkXTYGnH1QsC63I7YLUN8PRTA2pZdb8cOMnyElaj0zUMwWqtAlxO1
7GgtMa7Er1d2/4OUZl/UwuPiJ67C5s0ZQ2zl1ZIWFPKykBRyKrmKyI5DoBb+ax1xyxrNiUs1KEEN
IiE2x8Ap6PUMLFyWEO4OP+Gz1CKQzvmLVyYNV3X4DqGWNbKWhJaQ06c5Ocp3hpr8vSJV3OxDxQgB
BG9XDcdiBOJ6Z1kcBt6It3tOqxfX8ag/P6DpK7pvNs/FRY97r4gjJnnFvvT4yx5NQV3NBJ3qbO+K
G2bkhY2B8PbF6BKx8IwQrTRIFv9Qe2BThX3iwzW0i8seU/q65gWZEbRiHOpx8JZpQn4mlO4K9ff3
0Q4wcsIWXhxSpDuIdEg93Ajt8ADg7dDDG5JUm0ZxY9zKRWMSSJSB4bjVkq+BHIWOT1cFXKQJpEk/
6KXyh3q7kXudsClzjBkjOlU0ZNqC+wNA3j4/VsGq5Ln/jCyITax/eUzpSwJE71qoQ3I/IaGfDJR2
3+dg9/qDMJLLzIUNHd1aZWYNhfIa8ParzrnusHvBssg9N0RN/cilvcYVcjLKzpi6b2RPyi1WyXe0
wfLUyE0emV3GMdz0HE9K1R61gopoyWsmASMRc4ncjlFkI6eYdry2Rmtwcs6HiPMKTGhe324nBPEo
H0MhxM1v1v5nzR572plQ7/7oNYhjEXHkTYiiOAmtk9XHb8ZfNjdSlHtFZTsBg65/9wHkkUqTl8kj
BWoZgqH2OKND1YmLgNzY6/CAypzE5KWHqw+BnnA/4iZbmc6qSc493XdtuYNJQjSs+IN5R1qD3Kvj
oRNEQlI1EFQQyLmOVSRZDeCsR5uSoZwQ8uvHpMpz86BT8tcyLBHRGGQbaSqolN4K+RjYKG+UZREm
E6JPLJaaT0Uhj8SK6uASk/M6Uh3e65LuPsQ/G7z+GmjeYBBF9TXoShZLVXaA9EcsnYcjfjaaRQ1s
S/gDU+aS+PvwXkgot7yr6BPsGGCuZK01LaE8fsSKtw3Cvdn5WXR1HCPwTc+I7R61j07nWZ33Sik7
4wjUO3B/gCP9WNDZXixdQoBN3KIPw0db32IJqoYINM7hTQ+0rCmq7jQWcE9FyZS3sa2+fasTALJc
ChomlQPcMCJCRZD1kt8l0efhvylZ3pDLoLsrHbeA/SPtCpvptHXK32c1kMMfWwee2ZWtqmka1fx3
ssn08E98+wbhJzcuZlnlA3WvHLlSLAsnRcgolRTXQn91re2+th5Y9Uk7B+UGoo+Grtzw8IWvxzSs
DrYk/WPdDwOqDCdV3bVgv6DBBrcyB+bgKYehql0mXHQBDgtwjP95lFRy7BZl6lH+MGaOasAJRGaQ
jkm2Ylr/ejKcbE9a2FbqAEtV+NiSKr/qcDi2dNMeRno13JfOX47nbHYmu7A4Q7pfO8ymNyAZsTDp
uSLeXAh+fr2TfQNY/+dMftjq5VR/Z5fJzqbfDSsYHieCUDWhXHzOtflE7nLNhB1hFRJ70A3BBCvJ
Q3X2mf1AX8l2hzj3KrkfCr32ICVSmPWrkUKhj9tC7wt+1yR3RsEHhuAdhdh6BL9lLvqbcfkP03Je
bMcKOGQSq/M4fETvuZ8NwIZ8mi5zxWUsZPumrHx0oOrgrtWAyUKjcwRGv7jK+1sHMUaLR3rTj4gz
NWUOmM7MGteuQZwzzmsZRMtT/UPOdJcAC7Rc9yuNF3y44WFPpXmVerjgbAj/z+4TuiHCe2N+ZL/R
90TI2vxcGMcjOTNEKpilfhrRjJyMHq9+1i0UZvxAIQQr5o1A/vgo38ujsF3el32ajzRdZeE6s/Mc
TZiHzgB8q7YtWzZWRVKt8soZ6M9zYwf6AV2Up6pyMGkdqK5PfUgZGPGjy+RZFTSYYQzlqCbrPCP8
BwrUHIQyfllGWvuQ9W2XJHHdGJZl+FbN6ZQEUqxvsk/uK0XUlKKxiuL12XXXyn1lBnGlwqNBNrjj
7ovWt4lk0BOODeaKwx3Ske3KDGqwTNU3CH5m9SSWZub6Y/rlSkToc7N52BfvfUDdkSjHRPWcWHf0
bWaoYB7YPrnFn6GBA70f+erbK2Fqfp2sIwldnCNypkzdCfD6OpVhxFXS7VCptQdKj00UzGY8X7wd
6hNhQvuYc1CH1aDPYG4vHtP4PlO1zLoVW0w4NH0jl1RnuwTBTufPBGkkL8x7zqAGNXOm3t/5uNzW
mQZU88rm4Dpmri3WL7OTixdsa8/fRRyofVmFhHKMMqFx6p0PkS/eud4KUb3WP8afKXoyquxSk+jM
hi1Q00QXqUmjA3o9pmexRcf26DpnkSmo5Ij/+ocqctHVonTJef712R3vpCWTJowcQvZFCL/6xoYU
nCCOFFgmTTBrPWwtIxI1y+8SwnzgLtwzTceSy8Qvgs9/6h/UmciGPucBMgldKtpVPSoieU5uDpWy
7w8pN/JwBVmRawSdBHVeYUokrZin1f/yxicPhVOtsCEK9I/AwHfT2FnHC5QBk/ElT1ROQ5DMC5kw
r5UONJvYGu9gw9y6lQdpqBO4UiRGlY3YZQHaMIhlAiL46VXpXOFtGGZZGt1UdqLrb3A9RwOdmbTR
hdaToF0c6MJK9SVI27RGT1ehRAY1qkkIOwGuDNCLRAk9Le7Gtg+j6JbrPJm382QX+vVVj2tstHCP
4gRbNlXXjcORmeB6Dat9U9IN3pkIgWHfBLJMJv7XsjhHzMmZyc7nQE1sKUrBUL8U2XazqQKipn/X
UO2SaJ4smyHKcLoMncN7czc+R92HB7LPFAI9HnSFF5/dXBkMKuVTAvYNAW4G7BMc21w5Ggyl/dwH
0U3llm8egOLlbPh4t9CMTYNVsQxzXydfVBZo5bzZAJ4kP/FVP+ILSYlkVBMc/jyPxbK4W1VW8LAh
2fpKptjm2Ku23ZvG2lhSkMrBUyHJwz4oiuStnl3u4ibbDJT1NisFimzTdOIxb4hiVRezbzEyYMy5
dqrVf9A/Ux3AtvsSjPGCEwaFgIZj8vbWUp3mVT2JJPYKXE5JmbAanRrN5xtbxXCsGeuSWPTvLR5Y
VHict8LYNyMlusSp0rvmdl8svXNdOLDIr3qe7lOyRAlwVG0pKSwN5fbiNfUUUyESyq9kTCW6eo7v
ATMSYS9k+H7QqIaZ5kh6bbtpXj0iZbRAx4zpMKYc4j0NGgtDskSrmG726/qCRNoEoLn4xr8sSiPD
Xc36m3ECGUwdqq5QS79oUrrx1W7xFPLpXYMnIVdVRwKotCP4Ukez+J6v1UVngRUJ4AmpBotAPHfE
iIHiGI3XuupdrrJgRJCVBsYBsHzTiiHopAWlKogxrKD/KQux63Z0X5GnNK9Kvno6CZ5gt/tZxuqB
IFu5FA1WMq0oRAwHyw36efgpoFuSQnA+9Lp5WNmEyvsi9Ta0n1XxfUNBKEZCdHJFs7SXlhytqcMy
nio/0zcwNlZubiNquMpy+oeTUTX4Eu5WkAAdKlPsMCH1Y6XHW9qUEcDh6D1QoZ3KbrvGzocWANSl
t999BpwEwTA/K5PRV+JRRH1y6R7p7aWqvkbNn0f+bXrXUC7ixACJYHWHCcoGITWmzozN2VQig1rY
puGgvgq3IYGwGK3dUIyD/gASSwIYpxGWA4/UL1oX1gV6tUKSPaj9gHATTOjflJ/6fy+Cj+CDHqzK
mi5Y35wo5AJKkO6/ilxt+bOf0rcW7ypotwB6W8/Oft9sLNommcosR98HeQX6Jg5TFGMldAwRromp
JfBIEg4kVV+7A6ZOwpfAoogwUEovFK9uZhmFu7mjK/Wq8WLYD3GaZsXyUyO980FLX/E5uQFBMXyR
KNP+/ljuNYVp/bWhbOV6c7l2IHbVZcn4qidouitrv5PAgkLt3hFo1OV61890ec+FWpMhQigRHc8T
8YzD8WrNreRcO6/xQ7hHfupLvEU0sOuAd5WB1ZfE3FLA6wmuOcn6JsFW2mi527P0nnRKRXemgwje
M1OYlL+HY0Q9tT0RKM8jF/LThnROuwErd6OTljYJT7ti6Gd8nBx57lkneNgxLOtP8Ojp2trV7dlW
SdtjipuDxu/kYpb9DO9isz+R7QANre6HgQnmS9kPWab1cv/XpgmZXmFGMBYf+m4uV5QtUDHA8DLk
/7GLPTbRaPDzV1Kd4c5m49WNm9m/2eLt0fvt/gH3JeeTe0+8l03+mdRrBtZJGqAq0yps/j0xJLAZ
uAiGvyQ3ZDA8L/nh3JJYKwEtoooUHOjgxaOd1DUySI8iqwOjzDJw/UMZ7o+5M2NGsm+R09QxdTpp
Ew/9o+TUoPxRmOGUPiikXpNUMfEP9gC/UcOfPJlq6sr04FX4qYAL+R79oXzAfoeRzFuUS3ysL5sa
5WT9+ABwY057CR3Yri1NTzrjqTtfEMby2/ToVw47W5+/n5hb5RnISMQoU5wnfEr39LbYk+ZYrvaY
nzvgEnL08P3wo1iOBuSW8FAWMaGMfrbAy5pmD99Z0UTseNGW2SDJAtWkF6xoE9qJqxajVP8PE8VO
F7RK/FdaJATnkBJP/1aUm5KbWV0XxLi7y7MPrfUUgzWjlRaPhGb5GD4glwdlYu4LQ/hSF3COc4L5
LjT102WuXVoNT52M+teT743/cfV33RKh4dhgMXR9C/MGHh2b8TNS3lu8XJBZDoSr8m+O6d4w4+VS
viAapG5m2O4gqcxLvgk7vnmus+hm7yAWqkqPys91QWuGe8DOE/PmXnfEqlhjRj3m5oLADDldVmsh
O+CT84plwmzVPOhQnYxWQpAixAnjMauAOBw9PZBq7PUKsFPmY1PhF8fO7JpBE/lVk9eerxhvlDgr
rvxtPujhcy7zPTsx/K/ZIes61zJF7/1vcIN8rMHQ/uEQ8IkvXz9ihSRJ1N9G//tqpCEOR5FIF9Ve
2ZfEB/XB2cASbzRUKv/DlWXfQ5nG6GQsRIYdkbGLyYp/lCUreZ6pqZ08p6liVcp5UzBsauwhQ0NU
qEAXDXz1NaqP6B4IP9fCr9cAvGqWejhZ8p6yix4SIUhvFx8PMZpRO8RP4dvuF0VnxO7eds3EvxfB
R803/PjPOlRF1FXjd5fWv0pcmdPY1g3izkKxqODJAcI9MI5oMmiz6fevU3siHuCHO9zgOkikdNdz
iYpoBoiCUt8X1+K98wWq8spmDSMiqAQNnT1QtO/72HK5W1Obmw4qptYd58QWXVfENoGCYHHq7pAz
RdHtYQH/5rDrM0sMSicEovilDt67uFMJXCq7zmESsMO1mf8GUVhbWcZtY4zYQIyF4q9eiDL5s4kN
7RfI5LmVSBx8fePP7SVQOfmBnJTjZBUPuY1QpUUIA6WRFpbW0KyKSmrWkDJeyIREFdTXJBDpPJDR
xVqjNWIvVKiYZbMMqY9iLa3AASg68p5FmFabEiN8+QdaTroMB256WepPJWV8CNINaMgKBvWCSdMe
Gk6eWFU5IIzGA3sO4Qu50UBlfqs2vYOobUHvYmwnN//m7L45fb22x1gNVstViowIj0fmFkkonnJ2
2TagH7yh9qQpHCVymEQZkOBCbDcw4p4q2Zs0UFXxMG4lk4hdQ0JW5sulJ0fvH0QAAraXk3PnP+5a
LiuPPEUx9qMwSvhosop2mh5RpvdNuReQwetG0ZNUhGFrERow6k1p5THFI8Mq0I7OW/0O+5FIFmqn
19NHV9Q5xEKaPcFZvHdy6XJi4v/hEhvN5ITBof1wJmv2OEKocwNMLHgurxHE+aBEcLsL66PvJ4Dr
3711D7UTmukdLewpMjjL14ocSks6LNT35SQ68FRhNDZcc/xDqBmeT/SgnzCtr4eIGUJwdssws1Gd
OboMgLi+P9tb9LOY6aU1kOc+aMMUDeV0OEPbV6VFK3xhAesHLICt8nXwhbaMW1KKHEe9KK9ARKfo
6/0mXo9l3dFGJrLxoeQ7w3KORMySLGeJFnvjTOdr+Jtgnf7Nb+wN+Rz00p9Mnb9pf/Zkflxg9oG+
QoXW38QBsmG3tnkR8ZaU5GGbK0y4aVvINd/D3Iq2KqoDpKQOMOsacVRqiESdK8n8NE0iDjST8Df6
HPkb/+8n/31BQxo3xm147dVZM+SxzSQER39a6uB4CLCP6jrFHJ4KDIPYP1vKN74LUc0WvgmJQSdr
RaPt2k2pTdAq4vsGijIuT/Gbg4pa7Fy4HRHnCn4qbMMrD72g4tYNSXi1IsYpXGcVW2UTVkdhUwQS
07DJ0J7A7GdfzS4xIfjgZaVABsnJ8DkyxqA4qneB/5qOa4cR9vZTKb1fjtySLrFXN3BB21vbSHti
Z9sV885M4pSMu2FvRCB7tJqBVamQ+uTRL3/S1xzsxkBkF4m0oyPdhRgDW++3VYbMcEheHDpXmQ4C
dNv6nmnXv/pdpuwvXYAZtDRPLXRIQRs05irv9SvanZD+D4dfSeHGyLllYGu27SJ91dSR2HkuycJX
VpQ1f6Zr2OJhOhUlvcZEzAnEa4k+mGjRzBDJKPnCkU1kIYidQ1hbgT5+WrHi92GmEnqFoo5fFnLo
OCkvC3El7WkYtzEzv+zOl0nc+qkBLZB5fqqFzKWcNl56MM15sKpI6h39e6kxWZasHzgAN4k2yoJH
vV4nMk1EwAo8EgP/WyeVr/F7kAc00evMsvp4KSB9yLrR9Rrd5dlY5G46UT6liLhgxgbRITIqv/R9
4lVVidF0JbvcSqCad4npFOXqVGzncewDh+qzwJc2+NjiANAVlVOjbtrywE2S1Bja2q3F9j049oDv
/z2HPUiFspTNjLEHZCu2I6Y3EDd5QnEPHsJipH5GgPAmIJu8rr00BedWXzI6zvV3vODpJwOggS2o
oseG8iUANNaJ90Plk2vn5Q5OdAY/XrR5cJcB49W9OgSb7dzRxPXZ+WDfRNKjEi1JEMSrRQ24Ad6n
/zUK12qCHue0qxEQ6vEz1JKPAG0VWlsdfmeMA7+RaQldY/vFfcP14hTAJJIAGAoRREhFR2zWXaeL
T2xsj+xf7hTBnFn7m7D/87IDTwKI/eEkB/9ufA4K2pOWQAc0Fn6TubMOywxdeb1KoMRRX5Vi/3oh
ecPCkUAtgqseGYdSR9gGRgsjZGnX5OToEuhT+56WlxzmTe0EeKWaMfS060xXvdljRZU1omWqPwlx
qiCUMx64Oyh/Xz0S/rvdqmuNSL4d5krKdqRhSN7xN3j9YQzl4BhjJVaV4vd4FaFnVSaS58sSR4z5
iUmeV93eBb1nt5ziNKqsFWtcTkgFVXx3myP+ADMx8CdwvbVvUMPPC3tz5w12M2IZrAZzSh+yW2+s
wGnaY04hMr5UE4gMqXYKSzXGAZgyQuxS4BiVzOCYqThloJdfyq70QljEL/uRikMSdfSXNEQcotvj
CWPEAZmEaPXI7te7Ov/XPyJya7q6e8UKrxl8rm8k7d3RdN90086G8dRkCPQrR4+ori228yhwx+CS
XWnB/PJnqHK767OooLZG7/ucp5r7a2neiDxyGg8tfoIqlVkEzYkhba12EqiTl9CgfZHZ2t7amOOg
oAg+ptsds64nCi1ftIqssYLhctAzkanqxMyrA61cgoKEQAgeWmhyX1Mh9z84RaQ7CrvXhLkrVCdL
NqeKv7STSUcBnvjtW5Rmj3i6UtZNLj7D3l1xdm2EW1RT8rMbCps4av7ZQHhjGiOnVOosyvwLCsAc
8lz+bPeEDE9beboStohJcmQzbc8pEU/lUbNgEdSdDVf1izPeu6n6aPM6NCkX26SQicSCjeMoxZdJ
H6/mSp59yV4c9iNAfl0X06MUG41lXMShA1c1xcler4BGfCib4tUVuqzobB9Iv/k9Yw+XwYn6qrMn
ZM5sJ0haJIvnzqqd3o5zsk3cxR6L1YPeGA6udV1lIYTfDwh+ImrkXFw61Qlx7e3z5nb03DhRMckq
tLRDLbJ19kdqrAksJJ3td0PCQsM5t13uBPqmaHSyy7z7cY64KzvOjEPPy80Bkkasx3kiMkVNjKJ7
mi8c3px0K+GsLY/xBj9HPI0pWfpGdNA09Fq/mt23UKZIak3fzYA37RG0mGXdeUxF4VcVYYczGcXv
qfUbGAVGtV8BJURkRbF79oOv1G7VRC2iT9ZMea6OFcy5ljk2548ULDiASMkQdAQoG2NxQkr2c13Z
sG2K42l3E2S/myk8wVyKyLmNYY87AvInnZr+CJsl07GO/LclRpdthn/Y96djnI58ShbvKsZpquJN
zgIFyL5EGvSjC1H2WIUFX3FYUNLalpNdhcsscFKfu4AF3yDNK49oLljHFJ3u32DGjthEMBNzVGhI
Qq/XfvXRAp8N7w6AR8/6zEq7xsCPaLdJpYNy68SpaaXQFZlLJ4/v4yPs/BOqJpe3DmQwkuQ441GP
fEWD7KNBLdEOSKWbAFo/HpZ1uQvzGPqDhUmgUKgu1/9UITHJ3Z9d9WvZfa8VtSnqmBjOK2sTIeUi
z7WqP5g8C9ivOfjzgNiAY99Xsnaq3Rrv6LLLv2iRaO+RgLWOWY/rmC/59gq9MfvQjpq5kxgEhhZa
q4ElMjwFmGRvtsB+I5WbGVlFsh24XWpj9bYKpPTuhUwR19rmKAWajd6D94FQcd/yWVgMZPY+X0fs
+MBJR1lregdP7ngyzO+//oOQ7dAZKw//Y93ToWXvgHd2ItMDeCwZV/+dm/uIbqYIFNXTPPWPh19D
gV6UMJFDZG56bUxde3sZW1+JIS0MK0LWr8PR3ZfU85ZbBiGOztV/wTo9tYUJIP2kHs9DCGIPCxuX
uJSSJk34cgejWY6W29T+/rx4SBJNZ9OWH2fZ4mHKZrZLPoLf6Y2LssDKSeq7aMo05gcuPiybQWc8
UVHwmlMzkVaBevvswZm0Zh495uOimF7uFZTIxj3TqWPyoVLLSQsfEDS2uoWUJn4cPbrhig33N6eN
+5x9z09lU9TjI1a3g4cOY+EY3v9rE4ZqM9cEE2VoPrDS/4iP89oC5f5Slsd/vtSBMlPA29hw59GW
7/lVozpwHYenuHdA2acE9X4Mxsq96q5Pa2Hmecq9FuBVHbicZO6GDeKmpd5NxsR8hHRcDJ/Bcq1Z
ATeh5pmCZdt+fBImZ88M3bkBs4xmuJF+h4DkBOgNzgjXoC7Qoa3xrYiynAAI6/8cNmJrELu4FqQw
1nU1HPT/GG1dvaXL1BAkpvmlo3qkZpRLFYU1NfTxaA4oCDekpmld6ePL9pzs3TmFed7bufY7ftcT
UDw05J4L8bYmoYgyi0eivNlZhUbgq0ZaGMBHiHgpdUS6fSeXSoMLMOFmW3zDI5CTNTREaZ7Adi9V
Gw9rGY+kO/g2KSMSOu63f3KFj2MiOCh8maI3PrzHZ/YyK7tDgfyyhXMq5aFTEwrtG/EN/sIcIw30
RefOz0j6GoggETMn2ejkuVd7hLj7QUbjaEzrIHmYqslTyaAL5ovEsUTzXkIIxHLyWrnrmDuqP4Yi
HLNOx3ixZwuaFw7trbGd5mmzRZHlE2nmghrMxtbCbfhMBuvQTmtHMniHWfasfCxZ1aM/A3U2wsKM
vDtrTI19NxzCkL4x0pD4/DdbmWBcgVSsZCT+/cTzF3zAmW+Gf1xbZMgM1R0nGSIUptIzNy4dT1la
eONROhcvdXMuS+ElFjeRfhTaor95wQPQt81aB9PRlWsRHWnHIwjOXs6X13ebn4fYRhLZwUM1rrP2
5RrzjoSALrJnwAV6yEVXGTbV/BVoGsJJjFAoERxYxy7pMQ1WkDNmYDUnWdvyba35loQoZCpml0Kk
0QvQr4//0SvQL8pIN/Ah5msp5VllHTV7NePdtyC53MNfuGsxvShUlo2kVb1kRJ1upWfoY4hjMEPO
xttTUjSVFcgdS6vA2Vt40JnJcmdftkG77xb+0+ACFRp9DQCE6Mwyrr86oSnmjrxvq4uf1Z2wxMS+
YGadGaQZC+R5tb2dJIbpR/nIMGClPYLlrvd9CnGwCOSo+t0UlpVZJ9TNqosI2LNu/73BSCKSCeWf
BjaS9H+Fvv9OWCz/pL45g0sKiPA/qwnOC5RFhgpcL4ZUzeyTDzNgW9qWszrkGgRTXlYqu/1bLD6A
WRwNCJN848h2tVLxmoYn1wWklCp5/+qrRSYRA/cnji07R18e98vR4uTN/TC7JFDtn/jgUTUm7rrY
8c3HKbmpbbsN+5RXiicN+shTgyrvsPjbZJRPM6OdekVIkwFo0ysye6nW09Qf45xTuG4o2FNcu5mz
HdlTSEzFRQnFJ58d5EEqtbftECyvFq8BxFcomMT/yFH8A4hpWnQH/bemVMQk1GTyTonOxUGuhx4Y
+fntpYQjGLkQdD0vxIjVP9Cy2OsCjB1PyHJ5JW+BdFsKlYyWX/MuZSQhCWZQbl2HxcYNLmARw+WP
wA0uhmrCCT30RkKY6SYDF9Gy8v584LRLPRRUliPvtIZyWmiTW+U1V+AuiQg8/fq+mugPzfXT8pow
sMsmhFJD6udJuG4PdGpZbCoiEN9NUGOqHdvv6NF/aua0pZUdOu5WCagnmYB+fHpqxS2Q3hKk/CGh
sBVkQi/rvbQFyGPhVOvtbt17DJZy6JkZwWYF2MtTS3N85+6CQJdsdTJY2+Io6s4JGFVyUSM2N4Oc
xs7TClVXQiq45xYL7qLbQvUiK/9OK2T94lIoRMAEZZCyOKZcG8PIkN549LkxWaRpL5xhdijYer30
zmEq1wND+JguLinSiv6UMKCmHtfmgb8+Z//BZ1ySw83uqVJDZCitLzfbAnOY2lFfgqXmSg08/SnU
/BS8stHsKzLuAR+LgnJQt5fmxmjHj2v/jk1BGDKH74mzVnQK4xasv3QBtwbG9G2BkgKPeo9sRTAN
/lqox89EPW0N3Io1ebQ1oRgIsswRqiZKxnpK6Xui5SOgUiE7NKiWPuL4nQkBDyHyTNF/NH0ogbGx
0+MpEmt5TyZm34R6SBf3WL0/jV45rW495aIASRlMbzFZFtokcFOPWotO3YLaoVWLV/W2arQxAJmO
egjlj7o1VM9uwkvTZqdb3MrPGETe4Ivar+Eoh4LZJN7cK8UaxXOmrmYtHo/bXK8gEQTXafSIZfC8
RdcTXAk2QfVB659Ia1Hdpc6iW57K79m2rrMO03sY8GCR4+da4T/HHg4KZPdu79KfeyR7mVmVhGUa
By7+66eTd66QiITGqxamhO+7S/oo24U8BTQqyiCSLreFNNDGm78j+bw1Uik2HhM5Rqz48xKEo4o3
MG/JPS5X+BKIG7CVgSgzViLebdz1sJdzSIgXovu8emraQ3m3Whlp6oF6kGKcrWkcLCxYWBTmDYUU
1Ls/PKZ0ByFTfbMH8cqf1W5m/wF7p1vXEntDONUzRO7hvZUeMOHkcfhkUVG1d1wDtPP/m/rf9qu7
QMFmA7w3fDGIbv5xMlA+fTy8JJ0c3GWMcKxIhEcwln6R9KBMg0icVRAziF63UIzPjW7OsYwK/poI
Uv77WioV5PT8S0FVNQaJb9x08mGRayYEACWpnUo027r+9pQGemblcqYmRwUn/mgHd2Vuvden93V9
u8RPBlC2s/5SHFoPnK5ymqtvlg2k3Pio4jlNDH6lcKItqPktZy2weXI3n6dMXlBn402+DdVSHyiE
fmVM/LrtXzpdGfnf1PGqRqFXKtse/dQrWZaOA7OB8ovOdh0SAbTcE3Fj1B3rfNgDIE3mEcIoQm4U
HKMwiiDF/u/qUC38eHZHswSA+6SUfbFlrvCwWz1P1s1Spa1Vs0J0Sf859w2TBma4Sat+eOyUQxBU
hNhFxgcYKhsFHFcuePdFm+K56zlbvuxxY/Vfd/IWdF6FLoJwHWUIWI34mgnwBBEZ1azp3wdtI5Be
IO4V7L8J0HDn308/4Cls/WrQT10TSPLWzM0fTCAhc/BDT/HF4nPUFI2fmPkV1HTKM7BtQZcGiM1f
o/J07MwsT4seifDFHOki2cD6BffF77YptdGdBgCkks+H09qgTXfsOurHJWqLE9DLtPMugiSQNETy
19xbsaKlRfmD/V9JoOu52Mg/9WoDIHN4J9Hn7aE63fKkAn1uwGigaTvf1EZ+TRZlIKfeE7cAm+o5
f9vI5hEbs1IFtAj0jE8PhtNzXpr7K2KbtZ07pBUygJOQMPWqFFfdchcLuAToNZhaVoJ8Sgo5+PV8
nn3pjJlubPasX6c+z5B9rr5gDqvNg80b15fS99dQLRRqvtMY8V5T1A+hY/CIsgrmHyooXpQcwlpW
ZcGw46ymSWwbcCjLtpfdxp+AlrrISl0tmMeL8QnERI3DS8YNatOV/VP0V6176FJSdIjx6sU3Yn3q
XOddwvhbZXVXm8y66lhnA6/FAlDpnm0/oDKmi3VSRkidhnZgNs5K5yo0VqsN3VlgB2KQg07BSQVS
dMeo1Zya+e1tmlC4Uk3Nt0/WOWgsN37hLn4RWddoqT0ORrg6YgnzuEWoVlmBAmbhfH9ctuVaJUTV
mhv3ql3KcUjt/UwXJXN1cEAYUnYrN/XP8Jl9Gfo0ewChsA1soR13UUnl+8sNDxYfDfaU4bWTREOB
7kWxbz51D9iftdC/sj355SmWNDoDxfPq7Kl5kVjwdTz7aykZjD3PquBhQB4OrNIrB+G2QD8VPtHu
mUg04ScWyjgv1EttEiI6o+z8ff74BSAMy64Kv3UBq7FlG5fL91N7yYU65UTluEmIXGBH/nR3nU9S
LYwkbFOT7kgD6/yp85Q0ni8BuqMWC+9axoI8pIHDKE9ZrXhBVNKQ5TB7i6HOk7i4XqZcI/+gAhni
xpsMrUOoXgKmgXD2Cqou/56PQ+ATDRIieDYjj1YCH5rF7bf0HuBLpZLHUXZZqebTwFjG+vXQ6/Bl
jD3zAoFXDb9D9+2HJg7cPRwqFqiQfZB+t0kQ0gc1LhYVk5iVU71bvpzlWimBHL67RluMTd/1HCPU
71RztF46nb8+shSG244f9a3vJLm6eht7weEAnV1WI9B+O1rrFqtwubrq1+5r7z/yh1jl1G7sokc1
ihtCwFlDLsyS4mHG+qJqR/PW/suR8fS7qSC6G1Wvyg36rbPV4O3nF0dZVVd2rU+hLoX/n38OyoGV
8+VAjJ0HNcawaGUFva5hd75HXpObzJf/QkMu45UvdFrbwEP3Ic42FHrRE2r9N8/vIrkhnwPJWDjc
yGo6mwC+vdwyePjIaiJgMn3dEjlYCBU+uIkhJ5TlC181Z+cEJd/IZKr3mftFhxswEWzHFuUcyQzd
/9/QayIA6MsT86G8T3YzYuA8kQ9VAC2JLukstmuFczyvYPE9EQHdqHUtRHupci5+mzZP/E2T7iFC
HXLwxowq5iapRyxKhpnNnCv58FSqoC0EFnzccEOMKfyheJDdtUJim+dAD8TuuX0e9B5yrm5Yuyz4
Mt/+BniygE9Jq619ux0YZkcFMdAcKPl7yMhUvwNnjCNqNI5rvfLmyc/DenYuvrOmeE0toPXDfF5v
fRgMsITy1thSX9zNlmfXWEpIipUDh/Z1d77KTEwdphyFgLTMPnPdPiYuxggYvqT8w4I6JggA8EYU
ci+5ODvmvB6wT9P8QopI2gKztM5SSER08RMX56Larf8oHBEnPR2BZl/sOin/Ok3J+XqwQwMJvAQ3
n5d/4eMjeyAYEcbFf4/QlY4Cr5d8X0AINWoUz2xplK+Ff7rAsa/lSpUOfIfmvHZ0fVdQf4eKoSwN
Zuynx3izhPiPZrIPS+vgAorumLxFXdHk+Vo9vlkNI+IQcs0lghpOBqen5oIlOCJNP8phcMHwV4T3
mW2fPTRRaHPOqR33OZcpVSGQPUwwYcrHFpopN3t+SZuvLfNHa8UH97XJ8OOrSx6Xyt0jfdl97uuR
JXwIbhP61ShvH9rtVrjTFxr5km7PYaQi78B+CB3F6W18JUAhbkRu6WqeI0FeMcsrdZaTTTpPIEt4
/9VN+ol8VVhB7o0hBVaZATShP3eWqSRZGTRGOrnR6BqO27sPgFhH1FGh41uB0wP1JtROK3L+aegN
F3FJSqr8P0Xb2RgoHQeCX2bNwcihaNI/1WPwr904UgXDwn+TQXzrPy6o1LAAQgjUSYwLU1on1Lq/
VXYo1b5w1TsiDXMpUBkuZs5AJ7USFMEwL0coUR0y9opJDcAgsV8uWBRxB9c1aVQekDReU7fLU8h7
Y+H5qF5II5WjUnizLFuq8TMX16opjaBoTKAd08XvKZeiJdGO/jd8TfBWy3DrjucNTDiY+JL9sqSL
znePGkOh65eUjZwlN6pAAu9EsmmzKuvOpwh2PP3cpn7iRdO79G5HACF1JKZ93oDkPQA3gRVxCotP
6R0S2GYrgl/L0KyLapQhB1BxKc030nGskSfvd8chHKEGbtcrE0CYi6Y9d+E/nRPycwDfsc4mZKz5
DdDxhrMfldnKTriQFUzuQI0JWF9Ei8w2dJjrKVPW7nQGSa32+I7z5znQeT5PD0Il1+91Tvn0cJQs
MsDNhYHUyunm0FpQT/dDMLsathlQLWpBJV2tIgNrNl7hsiqa0F6LHPmTP5G6/uTTCgs1cl4pwJ/q
EdCc6bs7BhXiUPLlEem5AktGEbu9ugibn8p8TQd7iOdifono/yiH2Vf4//hpymkORK8bjXPMke9r
bLeJfc7ONwG+BasGKLo1yIg0wgFO2xa8kZiU1TyQuGNDaKnGXJ2xaAplih7dNEeo5sbysgTKYJPb
L4a5LL6z8R+Xsfsm4GQ+u6MhmsT53UJ2NlAvaOQPjEe9KKsGI0aZrPp3rPscTCEoScPSWnfui1Bq
hDJEXANwtZO1rCj6gZzMTsch5RVvtLD+h2fIuuxDDmOww5TkEshB8T8dxZH8+D8wgpX1Dae6/2UU
4UaEzIVpPVLQrpXadSKHHQH91ATk3YLWlQ8Cw0s0bB1cJ8mO8NSgxBmY1QbNedn56WZ7snBAaXeB
AQxAiwOo8HxPpBnGSqqDbEfgNZqpohYdt6fP1pJv4XcKiltXoihjH5xogd3L+goNskoiJAu6aYfH
lr+73ZDlvdrhxHi138mrbF9ue+zLPfJkzomBDmF5ZtKLbcvf5bmzKrNOZ7Eoon2/f5d8giqjDCqt
5rWjsYpFtD3VjxZI8FQrK+DF0NrB5AAysapslBL0OLqt9qX2n6MyWsVsYvBVL1yS2R2QsvYLPDU1
mwJxHPnCKQpmbz7ZV/YqqQ0nXe/ZkRpF6Qm8y/JXqoWt2JKxN92+mC4a/2EJ5/KK06FzNRC07U9U
4TCLr1Wbykli616bDvmKnYuoI9HhZs4v+Qft4VChHEqAI094zhJcy9mBZ99Kpff4EUIJVBbdA8yW
A/zPdLXPzdKmmwoCxgz3Mdx5hDFMZRCp9JEGG9TbqRc+upkeW77WLfBECD+E7VzEHudvJTEUpbQb
1S0qjqPuUiy/aWNL5f/BJ9txywQ5sTmvE8I3qoOdxRgIrjy6cvaH8SsIfY91gY7ylNKprRG+8tuZ
I/8BKKxUN4ivNLtzRRR+p7FKcrrOeumtCNN8/vauzlHcZKFeA0j+NtMIjRaI+tooXw8IiFJeQ7Xp
m+67WG3vD6TN3N1jA0rtMKow7enWH7ynWD0zdOPzjYHkKV5da/ee65hM4ItvqZNqNjPPRJQrUk1E
DEvDNwgWTyhOgkhIPb6mVjRYxAXFDMc5t5OypeCazoD/TXwapdny7GMfUprAARcbXl3xpK2qGykR
EniK97iFiWqrfCDUjQVv5XeeJN45o4kY0NkgJ0PN51dxUPF/uGZVod596XGKLqZnaedBs3frdpjt
QR9+I0AkUmXdeFwT2mUz3GHLIisi/QTIQHLbpDekDpB9WAjEBxZP5MMhfk4ofvZ6zLwlZHYsYDG4
bXaojK8IV8Ciy0jkVYzvWM6nCblXjj7mKbod0ua3aCyHmqDHsyKy/0MvldnPCTyBvnmxkB7N5Yty
Gd6KrCyuo0ya0nhjmLhcgKEg5H3CmrzyGpcxo8U1jBYwguIegnNlmUrXxHSWWLptiwC6eAcWakBZ
EIPv58h7EU2TLpOMpLpiyGNSalOcbuXnlDsTAOgEBDbkL8jr/VhCPUpa/gswydo1NZlxZJ72lNhK
HFsq53rXHqphX87Y96LMEoYm33fBOUzcdkN1RQ8diA3FKzfk3IU37aHyA0EimO3tEmOdIFv8Fdu0
g5eoox1YCcaI/bNvAmSzeWMBex0f25oxQaol/z7oFKNDZhpbGQsVOHJEYmQM4FvbWrYIwVSex1Ja
dbPPVHgjLvw1KkLra4r2/cfiofuajvjfonx86T3VpDTWb1UoSpEbfqaofD0vWy/MWYVlll/TY8ZX
JR3YvUTpnE7maHXMQetVHWct793UJNM3DCrjNZ3TtEYf2Gt3ALkjcLDF0xLahzWJDMhPWm7SSWqn
qbLEy783MX34Vxb7f9xpz8ssD9Ycy+KDyFNwbfiF7/GcY8ehn7YZB2/+uZEVXbemjMnzu8NoHsak
hEItfzjZUmolnWnv+4GrfwgWTZuDUSmk00qmdNajJkgDzhIbTl58ctvyAzUee0eidVT8SJyoPY24
xFQu3M/mlKj9pWH5HnSQeQNL4o9NMS24qZ1UwkP8RTh2FIbIPtKrie7jzhPt/vH2ZszJCSOMdzT5
3wrYYX/KgX0LC9l9LK4ArWgJ2tA6GO9Egj8SDo8KpGTNnSkykqBR3RyXs8V9M5jkPR+8TE1GTF5J
qYWXmT4mHQXY2z+Y7JxMx35MdOyTZ907nALOZKVQe3qCDi8JLHP/LIx4+bisc1+5uK0QpjcEwjLg
W9ShB9dy1vwCHmZItkzbta1nowa7VRMTChuQ/QM1XOoV5MnnJ4w2NzU96X/yLeYmKVExtmNphGgN
ftDm+ag5rG6z2vwZLCFfvBWIHuEQnHyDxYR+ds7H7wjHt8/X8i6qYynVuY9WbaPZO1WR2BR0qvi9
IDLeSrGZLaWHYaJST9bZU59cJPMaxxIOEnoyg/hjbr7D2J49Rq2dUPfagG4ML3/TU1GpZM+or8JF
t9vPx0SuUpPmLtDumdAVA46dNnRBaEYqs7GucvIy/oXYx7MwkCUUJ6GaZ4h3BbmwfEZ0+ll0rTsj
xPCj18IXE45H/S14HQiKmfN3H9Ec6BHL7UvmrB2uGSq02WaVwUeNCiSnYI5D0ORBWDugjqWsjhXg
0hTxBo1z33k/l1mHUNWyN1YVb9sYz9eubGC/aIcYIwvZS8YD9Yhvn5lA5KHSkWADJMmQz7XK2TuV
kjS1ILzhxQ6D2mygkR6ad4mYrMhwYJfp1jxjZ3Z/wa1iTS4sFrQqeRxvn8jh98rsedofNqAXpFeK
hWg9GdbzY/LqsUoc7gVSbiHoY8e0OM7I1iwIQw8LhAwzGwJ/j1H9pD9DoD4U4yjz1lJE/9OYVs62
Y/iwlUj4MtfTfYosa4INCl8TPtNdSrLecGPZHQOtLXGVPgIOwLob4ZwsKbOt0arojAxpY7xZwtec
aW+nb2pp6gSlWtnpR5jYTUEmWDphC7lGSMNO6EzOFWerRDNpwarqtothCQHqUj6yckpx/xqQEbiX
n924w3/98Y1fveZhY0NSDKW7sZ+wLqu/+3iv/1Nk5xYuHxMayEfW62esLoreEtIWKs93oeHr1FXd
PA8jwE2/0rRZPySW0IM4Sx0ZD0xr/W7UguucR+wB79uLXT1T8TKOym8mT9F1T0PyonucJ1JHXpmW
mC7GbQrXIT3IWj2nj5H7NCL1xwLIy3S8C1ig3iJdeFOQ8hdkGNRt9D3r8YejtiXwzXOdM+jbJHAP
jNxVgBz8janQRiErF90qQk7PAK35YkWo/ukbhoocrg/WRtUFuzfJaMGOoXS13CAkBURqYX05Dem8
9inz/hJqE7yP+PyIyvT+g7MciCxEx0X5HCeptQ63Lybm3RTXO148hY7/Gbiq3B93uwEAmPI92Qnz
yblfaBgTuU+/F53wpbcYNuftmIY7ppO6efygOKGO52JtT59B8jGXKB/Ghza/uMezGoWu2vNSjtcw
refs27fHUF7hDAFG1AcczMtGakUVLUrTEtvG43YDb6nvzF+X/Dq9UGQ7WK/F61kBar8/JSsRYoeS
Gy+rPAdR5FQ4tljb5c6fhSCLF+RhPRFCZSPZNcLM9r3efR8v0zIQO5pQFEQA2f72nH7eX8r1qmeR
bCQCE6SVNFEvfaeURAVJUALBiKnu9woKZNUx5yHoTvJId2gX3VIECPF4x3vCFXF2fUp3va4k5oQQ
QjbGJSqRsnh8vi5Zg3IAdYSuhLdKV/lQIjA4hNuOWUbXUAfcRuDvWQMNwBwIT2tNKul1oJu4vpUY
RnEYQz9IUYGUSITWhYsI+B6Qz4Hy2txre7n7uMq3ylV8k6A078xKeNMg6VhwA/m7hWZQE9u9pkmw
B9hmtnh2FqpNFOMfwPKYCATezAUubd1WrQO8U4I/93IV6CUimcVpnmVwJbKhhBsVnwsF0ZZ5LzHV
bNd0+q1UBzqPpbZCTmHspOwQeors3DE/93amRciE8cdj6XM5TyKZMUjHFIcxXoRaKC5JS1hQGn2N
PoxlQ4MHDxPKTyTuPNAKsbIZJPepA8lQSfYb+wEtNnHVF1edrdl7+/cf7FP7+OZzPPnJXrlO57d/
24jbwxwbVrwEgdBYWuKMkW5OffhRPTj70N4/YXLz7GsoJGYfgwGPDOOqdPqOA8oVQPeHbGlKwZHr
mzO4nbqLlqTPRnf/NrvGuno9aPBUkdvZrLpPKRzLyhuJ/dg4v1ESA6c6uF2UcNzcCwx2CwDEXoOf
N+zZBTWPQ56zQ/Mo0aNpHB3bbVONRN4znU+IB0KsTLhcuS+YRjIf7jihBDuGlP4TQQQvHGs/iwxR
9A4IKAxM69wfBHxpjR158btelhrJZRSwEtEogACP39Tz7xQ5tKm/69E7OzUs0UvXjPvYyUFIzJ1Z
a+qDuj/cWhZcPbEVOzOYpO+nsSmprwm2hRhos8kqSgCxq7yxfmHG0sWnADy+55T/VgFhRjPdXoTF
c82PAodQuKpGasXTc/CFm3NvwY7G3YEGFUKRA+IsLiRtLIraghrkK8f1FG76mQuxhYOPTwZXWVqd
n7iE2nPDXrS0oM5EiTYgFdnRzeyAx2B3VfTvckxqe0A3L+Fu4MlnBwmck4USLPt/AL0CPAmjeBqA
uMq6BRZqMubUKOfwAot4nXDDEMDjV6zGmceE35Emw1Qw3JJP1v37BH0lq5dtQQTckX2kLdKAbuME
bF4Zf1OE4uUTxMgTpEMGohOm29qiRhmZpAUacJ3QCySG2Xyt0A9Zuibt32/rUv3bZcMa71kK6VoE
ecIkrOm/ee8PT1+sTklyjTfPZVeiPduUPjQglmEXHQvkFXjnL8jdJOiQo+ZGRFKjNutNctnjKmeQ
7J+A4VYDoyAgQy39FJuwA7atRFzsyAgldksGn88HuNBkV2/UTqGl7SQil/GKEDj6nixZsqnAm717
reHJLd1Jdv9VaEQD+53gkY6Hm0ZU/ZVhFEgqja5V/6EZc54iF3Xs8K/OijoTvIsQ7Nhlhh6m+ZVq
Vw8b9F0qX68Ltt2zncGX6ajbGuurgceBiAXOLEuTzgcpJYbYnCcsNAIsNccWN3JK/QZ0zIG54HN2
UUtibIKYTiGTC7HnBqJ3viNpMg9ynPXmKQv7mCEUQhLBx8XZU3yGu9p199bNzydDVpdATnH8d/uA
ylMkutki963cXJdiw7Rer6j57kOblsJjihBk8C7cbN42YsOuBCiJSdmZ4A63FqU7b6g2vxzt97ge
YgJtACe3vNELuky4OZT2H3Lua+ijOovb8MEnEQoXsaqh3o4E2v099s1gMODHAjZZbel84c/QjGoN
EyAvZvbjnXgVYk1xQHw9OUiG5IEhPPGcmO+5g+4ekSM9nIgWapg54ZM/GQ3DB4YJZvXsVSZmeeuk
UdEhGORQ4LgjMmBNufPObTddJef92rGlU+5CU3AGgb97ObGalVkv3O64dj7y3ypP6Vbj7AbLrKL6
D2jKbAG4f1yvZdXxvfavl+Tf5DiLsrgrs1UxQael/+rygJK+dfn7pOxIG07S/X7A/x34/JOTvUP+
fPpjtjBHHl4tZmAPSbVKbb2pBOc7/inFrWGIRQXYYCc12jcDdIK8xZ9qCTUXNtvVLKezuJ4IsTrZ
uIbDEy0SBPjl4yfye3x9PGzxItbg6dEVWjqgfNtiAsuW1EqvJ8ALdWaxgo1sAvFnn7q7KVQDVov3
+fcfCyWIzKp4acxWz60zq0O6M9tk+5NgJFjNxUbmTpmyN0Z3W1bxqGlR+qN6HuYQg4eno+aG8wKy
c/P4GYoXUQYq1hwERTLGMF/ywV9tl3Dg7uu7PgF8VPVTNasxD4L23DFdeqlWxPLZ1GaeEMe9qyNc
x7xxrcpq6Yvq0nGsMqQRcONSGx7wthgLVIm8X6lDji0Nkt/3ShROVCCtMi0XXF3uQut9Wj8AZ/kU
dg+N8z+DTxFefuE2BDSznryqZEUfLy1xWr5Ox8GEiMfpCtTef5f5+YUIE08+jraHDzutDjD7qP1R
7N7PAGGB543x2WwdB5uQ3BNBf2f6BVKsuDZqgvk6Yd4hn7JCkLvo0XCXnzfqYf/+xxmDsIHHAKhb
smDXWeFsVeCJ/bKLivXH5WBBvJopuMtLs2XxotGH1MzOrXtXMiKU8rFl7kRAJedeOR0PQG0FWfp+
AnkFeDWo6X/K/lCChGTGQMRB3oiUvopCJd5S/8uyYeU1m1Fk5x3qGLaT2BAsFUzzsbTNYBM1szj9
ZdLBEGyzkdmiQ2cV6dCs8lhOkWzujOzxcKB4yvtP54EUrAbUOS+DvqetXfkuN7DKIHPAz9TWkGMe
szu8O5KhZZG96Gc1TJ6p/CZjzUM3LNz1ClFiWituYSYdeX9iZ4RrFYbxWq35+DbCZmf86mAj3tpF
x/jCr4bKa2GeDNFPXwvjynPdaqFBVJ/fO83SEKbeuLCIDfYD6YZk4RHdDVUWEQLaWqlXylGx86u7
fuctlI9w8lhdMbM3yfVxQuLrKcPlamJaQ/bh2oC80TgiMdh2MXLTijzSZCf4iIx5ruFoGeIqN2X1
njorI1Zt5u1opOEP07+bsSOlmAFfnaE16QAWzBBXU06IafB8c4DE8kxreG94HOwh0ppkxK+BNgRF
virA8ZTychrdQsvhAkYfajno+aRSIyzLU/9wa7BF/PsyJoo8QxQPJ8qQ723fyxFFSiHnv78Ag8O0
BGYNNFauDr5fDRYt4bIPRZ6mDO6Bg2b6goMmUTSttjfDF+7XBD3i0uinm2XoMfGcSlXAZ6SKjNon
h2LzSBD2vJDNQpAwh5ISD+WoxbUlV+KnossPPNVFRuGB+wDBHk934yJB0p5xAPWcDBT8NZD3XTqj
JiwE6CN8GkcCxhMZlHIu+px25RloPBgUv7P6iADXq/8DDXpuPWJydRFerrL3nToRDyA4aJmX9XAH
wmV3VkrA6Pn6wIQdSbhnGFJqhB7Lm0wn+hZ1FhKJK3/WNeovNfJvXyu+3j/3Ip3ZdqI/+tBt70tG
qin/Str6mDZ1zue9oC7tHWXyZT4vnuoGtaA4bKUF6LvHqZfxGwYxkqZAol6015kCSc5s/UV74dXV
az6iWYfyE/GW/mCFlZbscQX5dYQfVeJbbzgDQHb9twiazV6sLcs8j2qR1XAvc9ePMZqR89wwjXgn
O7/SXwn09Ih4hcHQsHVnIm8MkzQwqsdx/5GdVoc34Wm2mdoCVNhZXVukybD6fMVnJk9cDxgRdG46
Nf0Z64LS7U05xj92LuxDSgO78kS9O1uSXa+rYOOF7jbklq+tiXj72+hCEnxqlbZR3tNxPNIg6ZDg
Nv55gVKds3mAfbccancKyPo8YW9Oh5YvokAkRmSByJcwFQv6apsi5o4GqSfUZ+q+oyeMUC2OUbfe
D9Oskbhc0uXgmdpmirOkYFyJGh9Ba2bq56dfjlpG8c5Qu2PM4JP8XlYe9oir3n5PI//Bjg/vLGZt
zBdAK1dfKnarJgp5PElZTQow62rloWfyPjU6TBETrmTdunap4cjCBBMmTGn4xul5TtgcFsOXCfoI
LXXMfLXD7Uha/SiGFvTBuc0vITNfvzFjsXHA01nnu67rNIthW4bGkIJ8hHT6wAhpbJDzZhUeHx+a
TyXGjSmPiw2ZMHcDNLDKwYGM0ouUBRti1FzCOYnpgpTKBnZ/180ek5FAohBvnmZfQgRnYsY6ZHFG
u35P9ATfwVyDK+MxwCafvcEk/Z9c0db+NiCa1eeZAdYWh6NDa5b4/AwVjlkCQb4rIqZzvfYpiBTE
15SW/HRR6SghDGO13AlBp4D2aHl54FZ2+lcVH73r7s3jJVaNapNJWE+wB2wPtQ5J6wVjGoyRBcjq
mAQbxRgURk+pmB4oNWDnX/JWhUq4GbhMTf8HrnlBVuGzjk7Om2pRe1aQ2IxHbN7xADlzwR+Gac0j
D28fIvwE3pXV3zbNFCAFrJ0YHIBlDu9QaPA/yCaVvc1KTDMi9Yce4D062AepKme2hZAybZpl9jUU
TivGBcaHrm0W9HYb/Rlp1tNMpwv4dYu6E5RR4NXAXkhymsjgfaqfpx+V8mFSYD4JVyncIvHqmssC
028HH+cpt0Ar69YM6TNO8FV4U4wl4KWpMDho/WPAQShFX7QsNIiSjKO/2YOvKwA4WfBCuKFhYniQ
FKDEDe31Q0lLV36fwO/f5YgFW2PWX1T7Ek22PGdIur+7DERka9I4tEHXVgS24I4gxJ+NdhNL9qOp
ndtBwnpCgJ1uoxNHeorNcr6Yv7G6VCJjnBzpRQumQ7nDS+3WC4xbDE06tBchY/XJw0mqEYPwzYoz
bfHPDKECAnDBBfqq6LPdwn2kJoJ3KVbB9WmqHAFJkQb8zNat7f4xuVM5rXKojCFpo7cxKbfGmeK0
riuSosY7NUnh3ZgppDFFRzCVER7UKTDNLzTvG/o0fQ7fuzQFP4nW49KfPG5JUWvo57KDaoRjPltv
1nUpZGM+KPQrGFm89GZh/CONck4P7iDYxxTGgu+zhHvgAjhSMc3xmLDusvmjNbbxNlwhrwVO/g3E
hiT0s1JY1d61psJBjPqEnEczEMTjufjK0m1rV9IQiLOWk9WmlZNo2e6rLDOBJGP6kRHGlgJ2Qou6
EKnw5MIYooxHCYkkyfT58aIesZfkEeknGnXtgz3JF/0MjapgWMUhyzWuIRiPd9g2TdZkaoHk2Rjr
Hmm6Cc9i+uXxO6KLaO/4+kqJ69WREDvDxwR4TtINCTd+mp06PYvbGqAWGe4sJAFXpdgF+2sf/tiW
2/D9iA5uKlivNXZ6p50AfvyrJPEfDu8fWFcSR8Gai+5JK4vtOLBNl+rfieqWU5Igmr4lM52cXS5d
cJEEjkCzAZVjpSPd8u/SN5Z9dF3KkYHAq1ECrT6gaBp24Ea/SVNJ+rUf18e/Uzgx/oR415ojiWFT
uUOTWEQT1SVjb5+Waqn96F2bovlD0CVjyUVY29v+/k1ASag3Rphvde6dzs+k2Dof8Do5nRzoePd+
C119Nmxq7xSLJzTWDsksaaPdbvFsxcoVcpJXanqT61Elk1TQkb2L1UvY7LBsNRV3oWWhUfDCYAf6
CxMATjQaMgGAWjWdMuYvoELsG5QE+DyEgT7Vi4RsH3gIkIXsllAnOXll2oLySdesQ2HBWVJTURuo
H34ShWiOGD0iykiG0Eun6WwiJiZYpNzctZUp2OssmEdEyD5LYUXzO3oYrmxNVrVdS4uMTBBiELYu
vRY2wXC/ygfgQRLkVITeuKszzj9cXfO+X/FEScLaC2Z/SeIwJtu65qoyWPoRyfhzRyNA3qig/oD7
95RpiGHHorORANrxmyYGtsjjQLMTpSzgywRlBA/K1COE1RyotW05qnbKEZVXeLfVgTUh2vfapmbL
NHMgj8tllB8V9gWHAalbkrTok4Spp+DcMR8UbS8O2yRg5Im+Pvf/55HaReTzmEMKKVkd0zV3BoGD
N2OwwytV11PX9e4M+/fohWNZT2Hv5AmTE5XgqbIsAzJ4TJOsN34sY10/h/paZoOAZgeo42SSGy6n
DCrXaOyX9ZrqG9OuZySHAlCVQUBoujHwSONU44SpcZ2WsstER83LQJC4hiB+sVklSZBn32U6l05W
vDjvGT2KmFfsTvTbOk+0/OpHRJCM3HROYDMVnS0U5Lq8HW0WnJs/qqPTLRaIC3zJPy3kXfUDzP4E
Ps8X5DeA7tk65rNOVw2TX1d8RQQh14MCfhv1oWHXWJFu5U7rvtr9TGd5is+zdPODwdceQLoyDSHY
iVTe988R7TPX2L/cpH3m/OLJ7m9uXF/PgHTPWlqWgKZ+Rgm0K7YDZ67Y34C6ATenFiTO5YzMVOlu
A7FjvwNZJXSgoK5o6KQKzUeqUNA0A+v2YpVXTp5vDWhghcXQ1zRnDVIJpPMAj2q0YO1sXEjeHNg2
TqmX+ajSve4VrSbDATleb0i7a85fPm+2kcRPFPpR+wBZDj46Eb3mpgkzuMZstyhhz6oDxT88lwp0
csg6rNMhKsVLSRehadqZYO2bgqfYibpEDXHnudE+x0ZcKMoAjtyAF0dqdGJfBJANcxyzCZCH5272
AMsJij3i+9C+Wn3K6B/ZvYzyQszEHPbO3BmAp7ldM7Izj96NbCBaBa8Bibryz3L9la/+8xYwLnmK
aeAe2ajqhq8xYEPB8jT2Aw2Hm6218vAWqoVTLc+UHfpoKfS2iHcEapkCoaySbctEhwwVMuWE/eUh
Xu7aVC+Pcz3Vrv3OXh7fumkXH4HXZeFnCAV9szLUpQLKNjipvmZ06wQBvK1x7G52HUdicynZRqsO
OLzsoOJgSPvcXWYFCIKjXZgXdpgw7LSKeH74ZMZIdV16IA4fPARSuJWGDUVnxYWKvAGCYlL62B8v
+Znu3gZ94eAWZF1X5TTXQ6ZWgSVE9YfON/FGvXJVJI37WF6M7o5w2AZFKDRq0mPUr5ZtgDNELQCY
EyPS3+XRZcycBnXien+mZwGYya19ousnEmkAypLWdcwSGUbVzrrExJeewEOJEY4vUYt6v5C0nJFu
vQX5DH4n+n+4p4cy8tqOAKWpU+jpVnJEvwJRr0itIUTvTqqi3wozAwdlXziB3DwjODVM9BC4IXrv
MazNtmwUF2eLjE0eHeB2bZ6epW9bNg8m0x7/VQVL8PxCCJHf6x2mtQKKzb4MqrxW5wRInfyhB9Id
1c+3hWVnJM/21xgwm0UHEkdySC98vcNk2bv6hmdkM5qnA9Eys7NtVXqoRBYLJKrHvUMY57oRWBCE
r0hOV2CURXNm66vma9iNJAU1tIVb5WxFoftHXbZC98zgTnskt996HXo48igbEQxNvtuYCtpfrUPb
Ee8A0Aul8re0fd/8TQuQQVR5/D2nZ7KLtGcqmlIRFDytnhCgFqFtM3wmxTUcyNnT4aPFA08xcHrE
KSZIAGg8Qml613Im6qjXNfE70k6HoOygb+MCPUvG4V1hzKPU1W8mhcqnre6f0pyFADxZpxShbGzT
pqOpi8Xjvn3A3W8HKJsXWrQLy85u5+eLMyJsrJ2Jc/7l3+bEf2h/myrRDcMRFMCzbjETqvbNVZLK
lUg8LBcjcPn+tydroUd6eSuBUplLbD5q0NlRG2H+4GWLk+cdrzrjRS0xFLBd3dvq7686MAImmgMr
Hzr+sLCYt5Pp2zKW+xy+EfstFA8cCutm6Obi7UCFBP99hvhMsxGva559noN1o82q+PdQXIXj79Kp
hS5292NrEmmgoKn/XFy8EtYPRAPOJ/H30BFcvWvxRlUEDIq6U13yKyP+8y8vAk/M+8IF1sQkEJ3w
9E0tSx7pILEKDyACMst4FST5woCF2qLp49YxA0MeywSGpTT2m9X9tkwE99XVUCI6Bvro46GhcG6h
b99qJmz+v8eg+ImeRfUKf5Y/qoPr+Ph8m1q+qKeNkADYaNtdkaU7KnItY6mZLxZ1tMCoNqEKqZFG
4SpsGfVHWuKzuGTSdxC/JFybqz7+sxpI6yDb+K4WVbXZXHF5SmewAsDP5cN8vW82XBt/NZAKHzPG
l5pWl9oMDPCg0oz7C8cxj3AcG3iQ/Mc3cyHJMHk6UiLq1Wm/t1iozKYBk/eqnkNvynyhBmIKrqMN
mVQaMiOHGn28DrA4F1lXgJqaqVAKYRzUs1VyArZdZXjwH/WXCFHjbm3Y4oGj5IPTtXhgAPOE/umC
nN+OE5u73XWYj83Kw8uBxIE885Hubadt3k/ffw6OTn2S4hM7abGE7SQN44QA3fJ9UwqqRYdjiZwE
oUvXdSMEh79G8CAsaYtu/1x6CVhEwza8nBcucqzVpyvGVZitvYH2rAtM0tahUqpcmDhjk50nyNz8
uWbWfM9dX71MdQVIJKWKs8AwoR5bsnARrdUiYW6KUjs/RNcLSVYb8j95gQlW+W15q3dbluwou3Xw
HDMwRi2mi/3+h4IiTIxadcdWgyGcvsvuVnfREhVtjsyAvjqQ/kJ4BfqjfK/KFqLnN1/L+RZ9ZxHp
Lu1+8EeX0ShDbieS5hPx36l1ZWNovmGpqoqulT19G6zhjBhowRrb0JQZfbBSmQX2dKA24GrSX7mM
1WVA8DfPPsK+nhfLGkHbg30Xo+GX847rvgTEVQdLHMyfR/H+B9AgvcmO0NVgPfxgUyyqu2mFRJA+
gyoF9SxPpEuniNrUdPDc0hAH91t44a1+LC45VtdxBUS8uYVw7AG9lLyZ6dkh0SBAt0C59V2895Br
BDsAUQwtuBJ1+YuxWxiHt5XCcVXUWnqJ2w3PxZuDd1MSEKtY+n+l3Z68islN7+P+aRsvxDhEPZeQ
7JHbzlmuux02YmNWA2QQ4ccGzt5Pgm6EmxDZU1Qgx3sNUM67lmeDvT7ljPL3KC3iNaqD0Ixw+zfw
UHbUn3MkurGJ4awOp/vMDlN6e7U5LR6ryYI9BcRHHnpMgSzxZDoGXXs8WHmur6h5QxK8T54WzEr3
LTFywB/G06CJ1bRNIFCUFS9M6E8ymSeSrPTjHcX93yrF/Tgh4X3GQs+OXDqoi1PJZPSDEic2Hxh4
cLVkHRvmCcICfDFE9Gye05wuNomr9BnqCsK6VwcZQrbmZ/1UoXc+a6s7Y5/GwfuvVQrxUKEmHfa/
4me4sU1W1GVAHoFuRPV193u4H1cRaZ6IumycuNdGK0rtwN/k3xJ8aRTlX/S+PYNxcfYcwlAMv8Aa
hw+hFvELwKE8Z38/RrKpP35NQhlp2bEcjbH/mH9eNbdHZsW7kFJMdD/bjSCmui3Jnp+EvzSlVSK7
sGriJFnM7pSxoy0voplUK92P9oEDzgqPys3Q2hN7ftAT+m4BQ/8TJRbybNPbvdfjj/aX+UwkHahv
o4Erz7gYmjDph72/S4BTAjQlH2jjPGDMjY7aVsTVCGepTOtWLkZnaxDa2GEvYa7jmd2xiucHLjDz
fJOtwpylrcW3RWXqdcfyJaEyUwCAYVUSHlOrN2SgL/+dFHHOPh5c5iZuajSrFLG+FMenj5hxu8Qy
i3lZL09rBzuIiIUDCX0x9ze2KhAhWL8hHB5BLF6yoMq2kzGLq71XeB3rRrRsDQfJSF/Yms4kebPK
Eb/i/8yPEhkzGH9a+V1lqkl8ULzjiBSrDDXXpu7Dxk2LNCGuAXQ64VgVYBdfRj37TFsPYjeJVpYX
sHsUtFxJyZUQoKSlMoY9bb2hjxtB6iWd9rRJYdzK+mpfpj2R53m5sH3g8vJszCbbX8odvxVtDWDu
k+EcT5g3fCV/P1qapsZVKkdSZ5mv3XFpEmQDMSS2QmxjpNnYKYXhBbbnCfZMNDfhJITnGvBsV8z8
tSL/g+wOA8hmbl/gK3I7ROS5tI2WjheCd5iv4NjS72jPzfOKu1fHuF5nVwQbGyo+TfKIoV3YJP4d
GEs2XTxUeEDnvxJ9nG8fZMhuu0ZawEH/vq2dMUKw8y1g9xYIcZ2yiaCRGBlT4H53geBTr4yJXSrf
SVApnrF8OR/8famaosHLCmqaOHUSIUgBXfCHAxL1aPuC6oIxBmFZ9zjhUldc/HfdU7PO9MflvE76
pF0NVdvkh8hkAlCJXIVudxr/SA2/F1K5cAqhzuaYoJIzetXO3ozyG7OJAjbZMzkMvXqOl58DGPcQ
KROHEcG64qj1MilxnpJyhFNK7+qPV4lxdmVVP9FHreW1YW+N/3okcwk5xha+m9dPI6pZl9QScn6D
AuTegWpOb1xChxiQ5N07WqgIKQj8OcsIUzjrE2piRIHdYLRYRu9p6qCkjdvA8bMU//u7p0A9GZje
zPQ2Ua6AY1Tw2niWhE2s8XSQY2lfZgr2GNoMNnaYUwYnU2Iaj7MpEuRuRalKBkqC0rscNmkCeSLK
FAO4/taNDTXU1Eoer4Qe0zNG7qetPfbB15C/tO6TwBzK75tTEglTltISYQsZ0/WRInb/cynXdmYz
WWfJ9wya4/JBatygZdZ+uKkwBAKi+ep7mu9S12s1HEJVyxo82hWkng3XaFTsPA6WkpeQGE2g6olv
38SNQzVfIkfWnGWlnSrtXSf9Y7y4d4sUgirASqLV/SpkR9xNE+2X0XQjtpETqUSKYdVzjHGS0Yts
pIqYZuXl3JC3/C0yM47AbHRsT0HsKsZ8vQ5nby/oe2PWskxqSDhKvHcKlotUTwAvz5KThBKYQ4Jm
TmeM6Lk5jSo1T2UiuW5RsWmt3KO3SiJKeYlSptkSNspbsnaOdBR2+mYlj6b7m7DSAuvtlt62NhMX
czrdsFRKt9+zBJIpWNwQku9tZtD8YUkT459LJxYAwJiulVP5CYxpxTu98h+eFYo31kTsi1Kg2nv9
dlqTbWuv9+0GNWqtZTqOUcl8MzdMVbutU+9x5exmcoW1T9zETvHH/ogSrXkFI6hIpLkPjm/JuKYq
FzQbB5UQyF8jjPdS3nz1GQZUvc8Z8h7UewI1BQRFEgtA8F1xbxPkCjQstk1MsZw41HTmkYb9f180
GBorxbFeuMcvEXOo5p6qLwJBhVWotQVdzFIHZL/SWc/cl/NTdd1jZtzTJo7oNbU2WW+gW40UeQAW
HIeirYgPQxavx6Flb6Bvf4d14Kd8Ou0fLb7ec0Y5mpT3BEVNK5QCmMKOpMY4DCNGjDay+d55N7F5
rD6xAqDBJnabPmZhKmi2L4Wjeeztb3zURKzsZBHUDv9KCgzazbCKIbSeT9yfEst6tjfDKh5bDmpu
x0orsE7L4/zJbMfyBPHfUQEltObRHrJG4qIHSY/pCvpWSGxFvLfBWDXDIyLEji31YZEz+vOLBrqO
pyiR3oJ7tAhtdbJLQwFceRUrFNkD/KkUOyHtaMB+oIUF0dAZQwHjRZqKP4ALXO4r3NILZH9s15hc
vYAwAf0sxzz03RUx2lzrjO+qaq9NPS8msEZW3F2WXIywlSKFgJZVXeMcwlD54wFszRhniBATbJpa
Zc2TKGwRT8kfmA1dhcbgAejLbXxPRlwYWPpZ9/s/DTazdc12P08633WcbsvjMO1EsHS7hCh9AhBo
AOs/aQ/t0vAhWfmLMeicuOddWU3XLEwVQZsnAkr2lVIKPMpBQvvkTr/wt7NDNMHU1IjT9tHf6F2H
vNTGM+NrtCUHgejzCqnIyRbS6u3TPRWd1EqP3blyMDgOi4QDmdg2xdUuhZQGkAtmwas0lKku/+qE
UgtufjGMLbZkSzY6Eu1QoHZM7QOYzdivA4lJfliZOpr2zAUbNZMpj9K/ceAwyhaqaEUMAvnS4FSJ
fQdQ9T7mIZvs7nlqpCu2xCTejmm+j7EbXZnnSd5dvcdqsB3ixXC89Z9E3PRviepyjilLeNF0W2Cy
HakwXnxfUK4N+psugGNvJX5VQcLZT5CYnUo0ozVdgdrY7pSp5pKaP7tyK/hmApOmmZD3gskT9GA/
N630gUPzEUGDKYEP1rZEGN4ue6qRCAec1C3aY+yktDaSDITVBn9pTpCJHOVPzOsZjMLO/sDOF+VG
qYe90S94ioSz5yOMVjvbqhRgF5H/M0tR0PUGYWedpcvxgMyz7IWR4GlEcWYcYJS5dgY3ugjtLUau
ij5I1QGsL3E8ECeOF4yJvfgNAwTgDpNPT/KnzFfppvfI1tH+ngmCNohKREpi+6cNLNO0HDp02igJ
Td4ypvFCihacbaygej43R+LierrDee2FOVt6Cmx87zntvMwp2me1crhRkzMseKwHtN8fZXYJa4Mh
6nY0zAuuvqvOxew1tkjbShHJU5b/4qR9SW91JjSpXqkA1aEjnq0ebsLis1ok3ez3sSFMhRhErN4o
63lctB3yvgfMi2LUueuoSSPuXLIMJVu1qhlNjnyZliAt+EvXURk8pOhb5FQW1yItbP0hgYiLl8A1
kUDmp/7btymQkfj5LlwZuDsqxGn210RRZx9I9to/iF43MMF6KUNtKiUes8R73kXRqRvUNj5LY5I2
knyNciXI2mDiHkxyx3MFUiegRJPQCud2aYDilLecbSev+D4A6wTDjvbLlH5lvk6DbMcsTwqVj2jN
ZLPYUtj0UTfvP1H/556OaKK6pFRAoAvNfnu0jAzrJ7rgyXywD/rgE3nBmqS+lKJn5Tfa/FAUSphf
TRdWyifAraIRFQkhlKtDmgNiebOz/3Ev9s8WZm4yDljdwBgmhRd26NxfPMscCgTOirsQTRSy1G4T
3V4hW+FLfxYZQEM6N0/rPz1WL52cfU+nDK8lQ+f/Y+wEvuwNsycTAxKzsDQ9z4mvtRbi1GgWgRZI
2b2tP+xV54fCzmXjJ1yEClBF15ThJaPQ6j38/l97kwXx7JRu0DEDzZHEgjeP3JfhcvTPTVRDhAFM
s+vrXC9gjXBoMcWp5sOXxy5nX0aRHNdEre4TYK7ptcze0v/AhV1J4f/f83/d0Segzjhw4ZUvfjre
D+zatvDrIM4ogr3GsEN+xwOAhPQSHHP52+804ExMHegSu+Gl2pyvAVQNEehfDzqfNigMWeGgUk1U
Ze/dlmbkayxbmvajOmWqdi61IGFca0UAgJdJKBFUhdJBDcobKl2vS+l9PPSndttcc0MKQ2Jy0WLe
LKVn5cWVOJuE+K3ttAwB3nKImFtgb/5bFDObSpTJcJxNDIx4XJD0CimHxUzb1L5w79y8nSg1dQZW
SspwRDrOjqFff9Hz5wNXkgu1grsCe57XbotoTzdA0FR9Ngwvz2gobNtiJ0tBo2mfuzXPLxl/EdHU
kOkT6RNUJFjeH82OE0Y4yOxGcZg6KP98VgDV7hDTwff7VD0nX6fN7BCnhPt76HdPvjgp0CF5VB6h
zuF93mDhBh29h0J0L0ycxmn2r8qIRhpmHQHBKIxI3qbXysT9NkkjVJjbMjVjvGPDdTyuMmQLRI2J
FSkYJaS/4K21D/omtKG1nHyxckJVrwbC+EoW3DCI0SkOMD1YbsGQTaWrv16aEjDxjoYRXFIj/MoH
Bv4l+c5ZtI/7N9RKZI9OOyVNNpdMZcMYhPBv0GSZj88w8dDNLxqFKarCdwa5GKuyFNBkzyGAp10l
pIilQ7js2UY6MZcxzYmK3p3kUCLUyZc0fvnSUGSmmHYXs3FsUWb/Ctw0OLapTDRYOd6CJZUZGbrD
xiACuQGwa+HljjxsJMOmPexBwpoqJrvsr9suNafvLco85TXXCKC3MoWU1y7HtDlHTEA0dxjOGshY
T7fjow7ZNTqih/2WADwHm6FAecnLIV+KKxiaoGDXlvzDYbVfQ7wrqw6qHSQQbFLsIq7dIgLhUmK8
5UAtGHns9ntdgfzpkM/qh2BO8oJCFrEyh1e107YzyeEpVqRPaLodMD2fn9d7F+2fQFTHGNk5zgKn
Hs0VeMpruaoKk0LqG244TDj1/MyXMIgQUN6uAyG3Z4axyq2bG92mV1RJ5nOBFekF92n+Qi5VCTNF
HcLMXpY4D0Hc61UPrU4ayjCUCDQ3Huj2AzWsKW1sAs6A9faNS12/Cc0YVTGTXrfE/LsqPdTeAiCA
zC55drxNeiU8Zj6QoIXYS1p2Obe1sEtXy6QPvfVtIwxtYitfJA3o3VTmL3zj1CBEupnGGtATorn5
AFnZoRO4zs0Ht851iezIKnaYRrNvzJ2fUiw5e+n8oqTvJ/l83Tx7fs/izAs918H2qWb+JQYMqcx9
kI4y2zoLPVql9fT5OvjOQBjM8bZPgxYnZJhx6mZpzKyWwUVVsqE3m8v3EoAoQqHHfUHoeIl/YBzX
Yr1BNFwLwxqX/7V2DHerRWUM6YdMQ2Xw4d0bvpDVEaTWpgcpzbqeppNaWuF8H9Lyw+jGc1e+V8ld
IExj1n8A6zfuhlnxdw+JEddO9rMlfqrh9aXOZV/Z4v2SzOOPchBpzDyhLcUEeO6xI1HR6Pb8zbPG
iEQIKTA7msdFNbTsNdwaCFVZcmOFUcZU3WbCsaiUWj4+x4ysz80e6JB2G9nzxzdD6pMVn+X6CXiU
RsJGQXE8WXbfTrT7K6JnZUq7r0osTHgpi6qtVL+LHBK4+kc5AouSAhjmHAOxpeuituFqVFByBZ06
LXzF7pS/DAlWBCOlpK493T0ZwS68qVIWltVjibvTdrd2jJDJARsITn2IGxiCUUV9X9AZpFJUm9MV
oNmmJ1dyefO1LOG0rCTnCjOMDC+hOnF6cV9aMxvYV5CTMYPPPZ+AEJ3+XGu+2fYIJhvdmoP5uS5j
nebSXDamRQXN28lfBk6rMiurZxMpP0n46uAgpMZ/ghV9NDDOlFR1P4Ycw3W4IybJ24+dKBRI6ckT
YPvSsnN0QllcUyQ+1VjANk3BB8r47krSWKlK1CN2it9b+WBa6SwqgMdvenLWNNgdo28RPSdSEpaj
UsKm7WxF5p5GHRTUYuxLNag5tScZ51LJABZ0Qt/VuYxWeSgaJW8bnXam4uHPkkvQioa8BmuKe08z
53+uPO3iIq5vrx0zB7BnLJPvJSPRd0HfQKur+C3hCzrEicbK9bSMZCMUUnA/BzE+7mRmEWdFpHKM
ZDZs7yv4GfzCiw5bDIedVXFaW2PcQ7wqQALfPPXWn/Xr996z4nt/sQ9ueKmH/iHLE9SUfCEbC/YI
6OMdeg70O7D4XbgY5kRwmGP8vxoaUMbi9YFJk4clMQaQEsBEkF5KtD7WalLzLhRBHZi5me6aR+tg
3n158CicvXteMOxdGndL7Yj4z0nUujn4X8loRKfgpQbIwToPJ8gdtCpkQuvIpselY7PCEcVywJVa
RgydUuca/SEAQJv8bGXIzArMuIWELrxRrxAl354Dyh+xkx5nA/SEVmtQZuu+CwLMloynRtEwVX4U
Pc4KkwLEyP1y4KWrx6hdAtg7JPMkWdN+hZErq6VdrxzU0yKU0duMAcQMRcv6KICEChMtVXGlzAiU
zROqu/t8RDbAYxehtdKL+rHETzredZ0henz4oNXQvBOn1G9e5QIXDF1sWFpmgCMZSQN1IeEQWOc0
dJjryAgVHlOUMtNML3u9aqjlsxGtgyYHFYkOwO/rWuGhExGmquVqWtoru5I/tUh/gYv/U3xRwebj
M+InKxmM4eZbPsI/qdWnPkuYmUwqQ27JfDueyWZ+2bV7KDIa3RXvSYyFibyiuLJJiE6hfT5+hVj1
/VKaRuZx4s4s5RhZtGAwsNuKAJkO3P8fCswz5whVReHcC6fQ+kivvZjrvS88JPFL6BG5AsgJmCgV
T+z39ESzSPu6YL/ATV7hK5Jf6La63gQeq9Cr3XDxKQGjuvRFqnaWeNqnn6yCSL0grk0vCpr6DXw0
p3pn7F93qTwX2RVisEQoLN0BjKIkNXZ7D4RMNIJhyPNNoYc8ZqDImPnBX50Dzym6vOMSQ8tIZenk
Ny0m18WC9t27QP3l6C+1KiwXknH0zDuWJJZT8fiyq5DUHudDUuSOU588nc0gqIuZ1rIYLVPzC8nm
+wF4m5NJ2ZgQN1Mt+rSR4MlUaHUxRrb02c7M2pconOrbXiYie+QRoljR1P224CVLY6NJkR7Gn/vp
zxv3/rjBYAN2y/flZBFto9cJbcZJuxv4FXwjYvpjK/lnpARKChSDIuuMMARXxvy2k1YP99fVzhtU
wK6OF/VH9VewX6K07bsM8rh8MPWljTI3BKkEnnqkd/RE7b/EypgRwD/tG7nk5RW56nLUfdUCN1/N
V/Js198ER8X9MhYuT4lqRSsMLEji8Uso25Yn/YoOX8xB2dwvdW8X7Zi+a+1DPApfAubSTziKukYk
P1ePatjNocoOMWVId6Iny3bD/ta1pfRjbQCDmJ/enA4ABlYiMQui8bZv28E67xHDmm+prOU8+nsH
T6escQALt+WPV4VVpOETfjCarmAlHIYJutOj7vUly5kbQMJTQs6z5J+yUpWGnYEpuMj1EMZPtXSd
QCACQTu3u143jzMxCkcaRYIYiPshB+z+CXs0drb9lohpChEhcQmkoW+z/uSybX48NwgXT8YLXYbu
OcYiqhh5e2l4AgpCG8BD8gpjRIIRCtUWf1t+vwHE4YUNGaOZNI3y9PgIC8hxPj5o4tzIraZ0V7hC
bwmAQsrJfpGX+batmKMClUlTBDyLYc3xQ8rUK86UuyMu4XlJslz7S3tHlsUKzBDjNEfsnBGLTlom
NEQedeoEl37LwkdQiYU0pFnKs2RL12ARH7khaY6Xc3LG+uSmf+pxFDUxIC2zKdXNDbl9Ly9DVRUt
ZgbIlU76NogiWqcLgGxiZJyUUj0Ys1KJhyAFYwdvAKqx6fFXUSKqSK+PE8nm9hmUIdKS20x2lqEo
nZnRD6H0X+fmNDXe6Q++wtaMbjCRAE516CjNZQGKVcPCsRR/DxoWbiltliZnTNCHPd5B4g9qAO76
UHvKN80AxuWLT9o53NLvju7OZBmn/C7s9AeAItwxyktOavMLSKSbbDNrR8FraFCE4WKxhAQD6AlS
83/YlObraFfdpKLhkmQ4YfmV/mdVSA0g6nvMOvkrYW1W37g5kiflv9A3GwKJuHJvo7fMGaY5ijre
PVaJZtoBWpZUG5rtT+LHOE/9mEfs0kJUjs6g1XdNJ8kdjAPoSXxzpfae+5pkC0A4MJ/tM/e60snb
jZrZtluNnKIC1IST7Hy+utGCzjc6BjmguN9TFo4hUbodcdsDWmsWkaW41NTORicsJnMhMjubPWXA
m0T/c+oxDlOAoXDQEryhIPqsGFxsyP1Zs3peXSBB24smSFrhcj8Bw2ZLD8PrL01bFQf7Le+B15xt
2dJGOOCSMaqnxnJhdV8vhuDQoucTA4s1aFDDrQFCsvosfE6oikmJFbEoCL2whtoVLEIlMHys5rKD
6Ddvg7lwfQGdlnWzXNFcRZyKqMio+PS8bVtd6bOw34k2TH3D6h1i0tyJjUw00947fU6baMHG/F2Z
xyHbIAjVattP4uVZbRVp2YbJXGkDIvvCgor0B0+ROnAXVO15kYZCsJcOWKuHGsZmedmiVBV/x65A
HbPMA0r1sjnF148q0vphlVg4PjxRnB8D9vrtP0JKV3UlxwYNCUo7bYQ1s3J4nxfQnUpyg+mntX7y
SeI0YCuMtNkGq3FqXcesATUhmbS8JQ/gzxen7WQrfIOcwX2iyyDzOh4OR/DR8aAqS7TiS+tXi9u1
y7PQ8PmJyHIgMI9FP5/p2yOHYlk+APuiJbrlSphkIWMrN6abg4KtNnPbx11yD4rzoyWZBehRAKmm
YgAO+CZVeqOd+wPmxggwXqAqHJ3b2J91fnY1CEcWeAnmQryph8wudI8k2pdKT5UysP4oo6wZGbqo
D7X/loCj0E/d29My3SqTrJdaUcC/ORDDFhahx88PO33nL1PpMAeBkfnytRxoXrOJlQooy9uTAqiR
8VniW/r4QJJVMKtL7ps+ddRUxV9toMM/yZWn7ZfHQ2s/B3gIvXmygG0vcQOkGy+XGuSYQp7Brbk8
F2cCX/EL11ZpS9hXw4YkQscslJOk1tHWpF+v8y/waoX/Hdxg5TAAaCM7bVTP7zOTBbXLKZ4hnqFI
wrPJ1PVMm4GX4n/pxbKzg+d+XHE+4LdyAOeWMDsuvp+5638cSA5wAABD5amGs3vItwz6qGibSUDa
MSBqkGOfFmNx5AKQkHitxn/4VlIsJAdcs3oshK2UgWSWg1TVbTdMpDtkqhYsOp+rSPDb1d06GcC6
LG3aATokYWMJ/H71eZtQqfiJ4bC31jaVQOwVoJSv2ibyW0AtsvQGEbV/xIHbkLm6YyINW9CEyKNA
cpbI6rHlKd+LaqfL1u6FcqYZsrPrs79ODaCANESt/vd7/bm68MAi6YJNVX6Ffpe4NofbFJ/qlGML
Tsr7cMRV7maRDQEog0BbxPtMr5ZTXnlHPp1rgWFZ5N7z6/fbtSOOG8orgVLxfHeNV0rnj92YMDgv
rKuTDVWBZYVL2Sxs+0uQi7L//NIeNpvNoTbvkB3zZGpuAwOBaUelAT9nTnOBDp7qRDXyohJfER0i
Y367t4+gDOHVZPT/5JR2JZ9hlxmT/dGJM005dpLFjkpIoJ2iiXvmsggtwlG3YL9vPYyYNR0+X4Z0
T6qTfKT7Ox7lKA61DIpXYpEr9tkYajJmwdbST8lsxn7nEClkn+GpaFootSfXDgrAS8p/4GON4zgj
C97f08RQD+AzR/9Rn4v8NwpjYkMHSflv156H/sxIdA4+sDQaQ7QuciqoXpxTQEkLJcAU36zjuNmI
dZBx3aiagbjG9B3Le3T98EIlji6maKF6ANGXqeVqN4Rw7vkiRevHhItfT+KLAQjR2yZBPc0RrxUC
AgxgpDVHpQBgEtQ3tO/cbfaF5GoU7XqUNwe3xInhL5JWmRZQ0b1+ZmTZGR4gtXJJRO2TqUrjezP3
PjWcB1FldGcauOMty6P4IZYJ6nMCJ2uP2AiwvVF+8wxK57hv96c4yf6aee4DLNoyoFCoERfmdcK6
ULL4ZLJr/q3L8AoTWyFmkBjsG1Y+B++n5HB5NhzPRsHddA0bVLx+axJ8YMfOvHl4CEkiXHOcc43N
nTyepIj8SvKX4gtve1kVbYGEBD8TfxcYuUJquGpePsxhDlVbteHeaw+OkVJp4fE74oFrw9xLz/bQ
CoNSRfaC7XgXUxKpc1shLAbgT6q/R1e/Yw0LBkxXtRWZ8uN5wXZxSNbQyDTCKFbGTxp3WYboGWAF
XxeFDZ/KsYsvF/cyLYOyOOen/HuEKxeD8pY71DG9WClkLhV5t9LxWRaYIocVgSS9xgvQfKdap+pP
UfhB1GVWA5EgBvexJY0lHR/R8pvwb6cwmEl2Ra+/bwXoF8Xnq3IwVmATV3N4uOqv79KMDJS3OqZ0
04sQZg3DTW1AqMCCeN+nCkDyZQ4DJfynbRlJ5SVT8+x8+z0eSw6O0/VUdPl5ykLgT4U/SGZdRLNl
CKkwpbmi8OmEBS9Be35BQRxoqT+vpl86sWmaSWGnoTDDww4mEXOKCMWJ+CdTBryxTFfRXI9mRp2g
txNjNNoqQYZG5Mm/nOO48bOT7/N0XNG3WnF9dNaId63bsH6sM8HnpVwGjH43RP6xEZ1XBwSo/3WR
bIQZJx9DnI+oKaejRhp7AIMEIBnT1HL4lGxCpHB3aF49fcRTk9EgyW6s2zPGq+ULvcVBv5akjY7G
QYnL/CMBFSZt1Kc32UxVNp4TwhxvYMR1hEgZsYWVQZsSt6OiM8VhG6w/g6Z2pynxzi9GQlY5qB8w
w8EnIQu1saMK6qF+s6ICFgcGFcT5pDFYaFhUhqdre+iMam1+POYEJ2QY1ptA8tCKf+x+DtAwuTzf
xisT0Wn6KCQKtSIP71ckfXuRmjD/WmShbH9wcgWcDAUa9OFTKBX4ibNILazuR0xKfqYKG0dLs7fT
Wbi24ievdxQ4VzSX3VlR/WnKkJrTeInQS8Dq6RJzurc4veNyrPTP2zk+vySd6R3WHiO0M+RgpJ6u
i+T44UpSZieWEQ8RjST6245jk9AH2lGvG0v3ejcEcsKxi3OjkfwCsBDYT5Pu8b+HkVxyVor30DtS
QGN/raybEzfMcaotjXADweyWWv6RzSSm2cmA8JoXbyXGKth9Qrf682C08W1bFW2PuUNyjJDaLYM5
XMnxMcH0Ae5mE6AWDFS8Wy3qX7TqqnpuIO/rRtYHfrOGuL4ftXBDuMVP81L6b++WhbTD3ZGrb12F
rcyfZscApzScHpDrJIU1+L+zFG70gWlnc90IijRjbG3iQQXZ7Rg4BU1bLIy0UopX8HBytOk4SoeJ
kWFSVsmHHUPo0GqwnwOoQllvlAZuJ0vX6gG/HpgfXzKC1ksPFuJPObQh115sQ6BNZVGdDUNIBmi+
rOXv+4gHJ3MgSHQu3UaDsCau/jO55slAx/Ucwt+sN+I8+NbIE+7ViI4pAuq7gsQbT1+W1lk+B/WG
WuMraksaOot2UEaVqf2MwQ2AsEW11wk08yGh33hq9KrRxXgeWca5iMULvGQqGvCIy400EWEfkl42
H/NOqEohtlmcp/4gsmD/iZKa3ypUq3L/ug5NlS86oVn/5PMlhononsxhIc5AaG23hjjH576kMNcq
exe6UCy6zvK9kH+Qlj71btQgr3Pq3W2lfgnqQiUZKiitvnnTip6usubz4Wi4Gq/J+M42LJuayD6i
ugOYF+g8BsJ5l7xBLfXUjUvWvK+03XrLQVVcOxbjl0aVucu7mphx1f/FGndFA9dqNR6AEscqb3St
enH2Z9GrFOBKpJrtJQPLz/bAB4zUJcWEBTgnxzuKsUq4Ep5kFQmZOnCobAf9gYC0d9lkquAp4iQ7
fVrWvkxgnXfbyPYC02PCW0LwW2qdI/t18WYMESbsJcPwNXsRQAFx7tZYZl5Nj5dsaBsr48l6Rvgk
r1J7s/Kju8BG1ImMzaRYklNRj0wplQn95/FI4VA3x71fyqJpywvPPMl8CuQV8KQPwNXYV8+URl00
64JXhrbnlb/s4KIFfp/ZGCnzOmV7G9Rr23ReXg7VJ2MWA9sTKGqi2Il0XYf9/5Plq/2zG2HpjvIZ
37PNo9lfUpEV7Mo8n65VNVraOcP0X8qIZIGBCw4c2lMSnY1MSwNMAwRMGqNJfWEwSVcDp4hkJnD8
eaBLZDQOcCeA2lPr7pSTFOS0KqqNkBPaWM9JYzp0qVxKtKLZdi4DVIDolaYy7VM6Dg/tNN4c4ipo
U4+4ASHivko/Vl+Hd9H6S8aycH+iEQSbEQwFX8/rxxyyTscUKvQujKmKzo2ExVu1SWMmDH1GWz57
ns/NYKiua1WRD+rVqhTg+OZfCXZ3VJbbxSN7f8DvfYsgXMWe6ymy4q1YcJhUOkqmJ3m4Ff5SReqy
SmeIn6aYvjbdHjfCNCm3w7wvO/6SCH8mghWG8UNTMgkWPwnMDfY9B+rI62vbAf3udJ2xbSvgwpEB
VfN7T5afOkbqwtb8jjc8NqM8y5SS3y+BkVk/zYwFnJKQKr13Ny2b12jNo8a9RB7n1zOApN6Fkgg5
cQbJ6pbOjyvh+JN8JtwAfO6pkNBpmi4sPPBvGc4U10CtmPMT355bcd4mbVGcGA4JkahFg4ysZv8f
LcDzdckYgfBenkKH1/nzoN/MrCtYEe0KKOYmboNFRaWiVE8ur1gfIhCwNdOLvqBxf+NG3eIjAsP4
daOpVEzKCtPWW1jKKP5Lcvdbeq9AJV3dg2EOUD4n+PcdCPjUbTC9znz/47DXq2yBq4JuPYN/Wf7r
B6J0dGhs13ZuY4Rtr/cAcpZFYah/qVF58fzNKX0QGK4ZBOybn75Y9QE3vZqzGzNL35xkNYQSV6Yv
JlJi7RQaN9rcYof+untW+P/pMkR+r8iSB5ODyFqhAu7+w8vWZsuoCkxkbmuUNyHNt6vSRRMiKay5
w8Xxi/hfkl101xdtu3tTjpH4j4b6foH5vaDkaOeEuuuYIPqTs20DIfJy2mcAhR1ZpBZCTvkob5bF
UbJT5D28D3ia60cvzT8sVOk9Of/0o4QyLir41GlmR4kWnqqCtlLJ4nRZNB9ZxTMR2g07+XU+7KFG
jghYDluoJJ26z1IKfHo+T+3ovNcrQXqhSbxap3f+rsFyFaYLgCl58vxDdcg7BylW4/fec4YWJ6eu
gL+oc8iFOBx+VYc3T6ZCaf8gRJ5tptf/F7+6EVksHl4d83uBY4Mg+egcnhm0mEv52q72bmeJkZAT
1Od+2kiTIlraWqC9lFenXYC5PkMwju5LgMBvEhkE5O2d5B0lJ0FXWw4fYsPMH0lt6zcAuTrNGlCV
FopVuQQASX6YxscRHWUwCzH6+xHQI49B320WbJFBtN+Xqv3312HPTvnfaUY87M/Gsrk0mWa8rOc+
WGUNX/yCvxr/jTdrb2HHwiI7HgWRRNPQBslXcHk11IqSen4ZAjfaDl18i93jxC3E7ADwgRDxjV72
hFC0AJGvUzHbkGUxdhEZaPvm8kylKhhqWexEEJXrk4dyfYRvZfljxnL8EPJ25v5ITAEpwg7rBxxu
uD9f7Y9gVKxkF6w7eUzzS+wPduSbX+7q59ZddZNmsm7g97TN1IXPDAAX49mpwO4enJCNgGV5ilIv
GevbtQ8f40dRHF1h1QfTHKbIaMw8t/V2au9NROnKcvwC0NOteqjB/QL2OYQhXUwm+MDoXwdolrKE
OPYXYdcR31EPKJdbQzz8LWO18fjHrlDFLFC2ZqKla0A7154G3TOcIHIXXs8ECcygkfQPialUPZyz
fjqNlLRcOjJM1+YN4yozdz+THMS3IMvQ+2yk4ZNGN2vEsRaES9kupvm9lCN3NfC+1mDm9fwG4pvl
Gsr6punqdAHx4peXfv0yovO0FryqXgNiA+oSyFYAUZDZzboFFbVTYb88410o1LVOnYMPWKGrd+Ps
AvzBnrZ1FQSnj0ksrPBrUPxwaTLbzYHc4fXZ4XFSOkG17FFAAGihcnAfIHj9LbAfui7fNZqAnW77
EE3jwUTlW5exLFFPmfYalsT+X1wE/Q/3pU18BNU0DPPX5Ikb2+Hx5lK3CnDL2oj49XqzKIXemCVh
w2TtMCCuqrGZlyvizha6+nCc8gze83zpB7068tNpf83xtuCg6H0TsQ8iAoFeDoM1M48AFR61RLxh
waQARhdLK6GiOuYhNT+BKyz5WqW4s/XlmRRDwFjT0q2fEtZZUQjPHZwmgMrC0FvPpqLpLiEV7Ozn
qUUvaQrV6sWJq1AJfzaXIkDs78ujj25RJRf8jC/P07Gwia7Gz4EPovqHbUVFAw+xPoVyZNA7wM92
1r/o9bbzX5e7K+6tKPUXMuJ1YVi7AbmUw0qklC00iX+dQ3MINUCPDuxUNW9l33u6zSdT2B76Mumz
OgSrvcG+VFnAhjar3YU6wzOtw04Xbwn1iwY1aPy+NhDDprG6TwTuIsxC4jNpgpmHWUNz+FjDMfd8
9BB8+n42y2mdZUoU+rMR1zzG49fFdC6fE7pZHpuEEd9x+j7yuFuxmUJXUE1JUIquCuHbT7lE2bQy
5gtw2FIZsvLAyCuyjGwIeENDM/TxQxj+UPs5VkYzDzw/1KbCkOYAcG1KqM0FMwYYzLKFW+0alsi4
uh9MoBGXlOWJNzSjqpy8M+V44TcNBmBzMRQ1v9wok9Is7uTtl5F3vX2EOFKewgm0JVpPE2Qw/tGh
JLEFZnw4SPIsKiJ99Annu4XO5HqmQam8tzDzH4/zgBUIXUndciFcfUKOXoFU6RDGwGyjtJkdlQpZ
HUCt5s9LCR+1UAUQPZJ3woMXMiaMdGTJuuhdsYhQ3fUkp/Uy5dXT5lUouKECYI6m4HvMLMOJzi/4
TC3o+BdojxzMd6VcbkgsMZhiEK+K1N0m7tzRg5FcEJI7AG/qQ2bHEx/0Bn+J0yb4I3f7w+omsg5u
feIqwbKJ7ipdDqhztuSJmkMN6rnoCqjx2uC24sEwr5ratku1hkuxYxYj4wGuKwpxj7VBTQui4Qtx
DrHrh+K7ntnIMYfUlTX4X52v43viG145pzyhqWDc+rqOkpZQyL+U4tyNH6Rx7cAyL4JCrmDRnmjE
NrWQ6wF8HafmX/bkMR0WPq55XyyHW2NMrkCnEoVA6k7ORWWtLODqMFNQcwg1MOjcW+07VqaC5PPe
Uz3YSIahSODQVwTm3+jlCnfm4x0/Di6BNoC1ugj7OSxZhUkgjxVl28/dzCaAkK/N1DjjK+mPYqFH
rfqLGK7srN+xnUQtAI7LXgdjJcN9hfIabe2neMAuNWyGSAfI3kyuZIMhHHtq2Kf/nDxXQpMVPyGx
vN711SDaZG6+9d+6l+9x4XQDeoxTppQMn6D0a+yXFxVopYiouDBQPEOUq7d9llTDhmA+t+lJEv7L
NaUKWjmcZskcV254DXdwLbOTTLvXyzKDv4AwZieirAqlztg0wYOuvYHmQeclAa1L+xnViyfIowbv
l3GMu54q/+9DZuOWiSfiq21+6l91FBHMwyIsEs//sxvYSDwCR9bP8jkI8AK9KgpA1uEhq+0oTVXD
uUAYcWTJFukYW47JQdVLw3hPOAJkg1yIaY8uI7SDp31CEh0nA92JDEpExs4ekmAmUGwFeGmHLFyA
/Z+XvzNQNWEgtKsIM2SwjKqtZjb9Sgjf793IrWs5JQ8+fQQZEKiy1MKtLD5NkUh3pIB22H69YA2F
LfUKI4Kmih5KWl3/Fvr+FlnajyjvRcx8Q/1yLSszSwgqdQ8amM+EQWlpg7V/mnyex6gUdV+BcwPA
6mFdMdOl14QDyUhI4sHTAa74WbK1TvHL1xUmzUVmA983+BjKaf222sx1zcSUMKZRSpeCn2L57ROq
uM3vXtoJzQXJQCH99KxaIe+JDhTVdV74/6BYG1BjewZLVR1Ela/B6KuP55RzeU0vZZCiUFEeweWD
Kl8sW9oYWbm0NAN7JvLHXsqN1vgEyhXWOuRBAuI+TnBbnpdLjtCFpyiJhvN9KufHPJGPXp8qbpLX
IOYrrYdaTFedgf1J2jbwVI7tludV34iawhcvX8GwNopcLfWaMoSp0n/xkiLK3fSrQnacjaMXCj0u
98ttBM1ZLcYNKMYXn3aMyNGVaHT/ClFrXuRCGsJXbrZWgypfSgvo8WD/uObqE0nAHVIkPrIOGFvS
q6wy9CN1ObY7B8a2wZgo+ao3/fYURem1fFZAv5Twiql4LcgJJ5DZjcj9VdEKPU1I0fT+N4s58yoK
6QIizQlUhtp1D2Tb6GbvK9McErkLmewQGOB1EUE9rDuH1lTg3aWePFY9Jw/4mTYPpIBtcgKfmU/y
32xFO9yKzCWCWd22UEmCVQHfd/y7xmu7EoQgZnGorTQpT7YIkboQ5KvMR5iKrXW4zpLC1R2lD3L2
A+4oDHyRRqmfTzWkA8D+HyFLT1n87eo047dW64bySlFznxnwUs2+7t9gpDinbJGKy4MbAEnTvFLY
8gia80Fp/D7ZTXd69riewE9ewnBU27xeKPKzWyNJ22A/xxyHf4nyUv5WHdxT1ZTWwyhnhcbrvdLs
PaO0Q2ahg9RDEQUA5IcKhfA9+TH30aYoagBSQQUkx7rDeCxYLxG5dk9TKyxuafehz4M3OgdJFKrD
fFLs626heq5JQya7jG4E7M5eVuTTM7FgCVa3q62m2aDfjlTW4lYvCYJvZUVmAYNJt/TnDQ4fLpV4
78aBMKiTAY+5LMDM/erUcV8x0DRlea6Qu/CfzYUmC7cq/2Yp2fq1SI9K814uC1YNW7vh50euc70Z
CSkJKPXIu+q+ciP/1j/SNphv6+qp34z36Iibnx5wW6MtNj5eE1RkVcqVbDbVssRlO6k6qN8OLPd4
TTtM95kqJQRyUvBU9vqVo33kWw0DV+y2DQMsG6Qfc5uz59licBJOr7KBbiVawUV45F5BrzjNwZPF
qqz+dume4le4fc0/sUsbq6CFgcAmusxCd+LcO3myGpd0z/NjpwV8yJG6Ou58d0CzXe5o0zDHtpVZ
EUCU+7GX+HVjoQUTG6OAAcHGXf+SSmcWUZ4cAmbX2cqnSLUHR5cQnfFsr2/GkdU2cuCWXFC1JBo5
x+PAqNgCwcrbcZb6jt8EukuxlVRx9xGrCSQgYeJc5ds9M7QgDcXfvARwFXfSF0oPZo0Y/8wC4tXQ
XJsjDZQVBSWvn+GDEvS3EVXNlORDjFqMAS3z95XsiyNsRa6y40jkf9v+GFry6qrOnACMe16DgL7w
ffetQ0f/wWARSPoEAS9Ludt5x/PjFjpZZSj2KQfGFvhMso5fNCPTFXDDcjMK/JGoeKlPSjcmunXl
FmYf1DKieptbFgjmY/N4uN72Fe0zJ3NCb0GjBqlROu3liY0jCLaQqaQUSK3f9omlFDykXgdxifMk
Xyoy+VioWAmFVjA3cv+Pbm8m2OnzogCQO1y1MSqpWU6HD3i02oVcrlf/RduAbcd7sldiBK9/cufr
JoY2UO8u1lBFpuQ+1fJLpTsXdH5JxvLIVXglLCvaa3P5NOqHNy+1P9nnOXPRK0vuSQHutdJlZvGA
MS0sz7jpef9KhGddXzvfgwY3XwlaUl47gci5MCwcYUuqw5r4A/cHvYp3kpGBO5g2dWAu3C4sEmW2
vIHUafs7vVqIr3Mzs/CzJAchCSHoxwgHWpmVIV6CUpzdHFSAlbvTo1rlNynYY0tWCD4lOOjlAHE+
WGzPRjIMh/L167UarVzcCxpVy5LgEMPo9rwvlys/JK9wwc9Fv/uH95PkRWHxL73wZE87shsWfwpp
qF+Gpkyglq6bGbeLINifMAzu8LRFhs7CHtOHvL3Eqlsh2jUQnD7MHFTj6PPy/3CZzZu7ibM2sB8M
ljilB1PE0Nb8GX4HvoB7jyDm3JzlTgR0N5qyeApAZLg8rmlFgRQZu++39L1EPMJ29ydJD/lL2sGS
+ZtzhCMP9Ws2ZAJRCnWeEyJTfBW7LEDih5e2tEQXIRtEdh0WO6UsnUFcftYb/Iakz9VPkqejpUf0
cY1wGGCv6jD1Be+eUsLlrQ2kNh1WZprINH0xZ7O62w2CDg+tNwnJ07s9s4dZY162TZMHizZV61LU
JLOU64+BWj5eC9cODYpotXsyk+J5PHetlfU6xdsTIIb4050VACChSaGMHgnvHUiGpmnG2HFyTow6
f57ipNCL2uIi6gwbXAfD0awEoD72n//vOLODJo1qjF9HeZo09/o6d6Udq+g1GlpJlaODeQCD3Xc5
asGIk2Y7wxvQZQ5z6NACD+cGuOiEomWnxHIv7OTBzdbE8Sr92NFHQsjWL7Rl3Y7oe9Ba0lqEywXY
8mjzb5XwT10GRAykvgM2SO+UByaFtmWxcaw8mPwYqP5Ju5Mo0c3HfPTXXL9FCHQDVZRcOpOGi9ow
IK3HOvMSDBQKjaeo7yHGySezlFEBvSyW66Bcj2lV2JufP+on54v7oMfo88wI56eIba/zVg3gAo4f
o379skaedBdnkzh/rKa5MKT7SogEu2T05/5YE/4usvhT5n4tyiPELeu8U6vPX7mMsJH7my/b1l1+
rS359xe/dwDUPPdoo+VL2WMHjg7A6CxC57e3dUBYRY0J2D/XrULhT1Ie7N6M9OfJWgMcPBqco50k
CtjOFtfeTBo3htC3eOW5bpX9KtIuKpnorxsNUg38Uw+xTyadEp1NAfl0lg/7RtFJdGLSuyMEME03
paGtRFhqvFiWxIM04oDg4deFJHfJ6AcxruvtkAJcGcMUmh07A8bFo2uFNA7IaRvDluBOMHwnP4z6
No0NSwxmbhHcJi05tZlXGHoX7udb6T1xLYegcgawf6Z1U2oHTrHXkZJRhf/LS+73BjeVKmMLsPa1
bwbu7uguThIkmxedERE6d4skzPLAaATj9mxvifz7ke43Vd7XSFwM4FLtEcRbdNYKdEHBTBb/jPYS
QACcdbFv4X8YOyr7ta6Eb1cjEBfLVgNOI4HSKup8SyhqIj6sPHV8jrRnFsJdObMTyTO6hdeA2Yzt
ksGAuzjBJdi0tA4dYfpiLKoN8N0iqva5lQ1h/Ytl9zLSD1iox8hydOD4sGZZtmySHouH/eMm/DQX
lDMMmB+PXHUDKmzav5vqQT/oOsdwsr2vWcf8tSv08zflCU89OZX2OMx+jqeqv856N+Umi6ov1hO7
LZjrqkReon1yVWSTzbSZrlpgpmWnm35w/WmQ9fr9njQcSx0xyPmLZ/A1PGecUQ5/SUMmESfDvVdY
rejm43WuEs6VvELDrCpJ0qEATos3Dxq67I24QTmwH7u+JnbzCOk8SPxHJOeZar/+LiwLZGW6+/Wa
o7Y3fy4glat7qDQsS/ZotzHrtZeZd7t1W89BfU+LEcraJFnIAq0G2pqb7QWWiWYKJqsbsb4xQSYA
hK7LqcLgKSJB/hOVoO3nyeDZEj7qh+W2H2zsZDtgdpwfCtWIZYhnbHtdwevOlyOijcHiMvpsmzSU
t2XOLDBZ/JuO6jk1dS3OjFEHVI4siKmZTK68ilu80n+uX31MAe7+O8cQ368YNsWwFzvzZWm5OI2z
KLW3FcoRQtBg+X0gqbG3P62PkeKx1W0bDOOL6MzYEuDlDghcncD5fBNV6i8S51XsoIn1qfAmxBvO
ml+ePFb9zrG7DRvQO/rVz7fG+HDE3tDV/EdXKDSNFRKT2msffWzluGvQMs3ujdc4ue7oYzQvmk7Z
ujviFws9klt6e7/16ebUFvfyZhgcLfsMkCouAhWm7a9qqazq+MubZ1zeQJUM5rfx/mCyub7UwhrI
HYGZXIaz6usruQnv/TEdG+VyE67qsX98y0BYfIGCtEryxmiahy56XKtlfNajmIKgRuDoRi9tL4D9
cia34bCJjIGiAVtHvegmQriFkpnhI0tdV8za1oF85La2QE4Ngd2kUAJjno/CzWlQ5TwwrmZ20hOh
EXp+GA4RyxsdzsWBOvRXzIYhPQ/KM3sHn0Y1CCc+dDIZGTJr+t8QakAadCk0K2dbXVCTmOXmrmnj
ulvPtSZkEUYGHz4/99LLWG8ezxXWM1Vl0PONPLgUYAC1gCvMFlssmn3GCnMtojxPGxukycc+Hfjv
YTcMu4gbthbUo++OfHSwszzpuXdr4fvTn+jFbP/qkkoE8oKXpJUSiWXA4T5R7uPC1bLRPsaZXzIE
0dAyIF4JfWGqPkh9ADDOCXkVB46E43ssDQOU5fwq8dFJ+7WZ8kZo9M/laez463c8RV+qOk7InpRl
g6oBx8HIHeJPHCzqoMlsaIHLJS6IL4McnoU3q6vrNZCqmM4hbg43swzRFZQVf9zsYGZ6Z+8/pxVT
mKDWQ4txRz+ooyYk0MGH1OIHiRh1wMHKGltMpPc9tr2BdLTJbFUiu6Ue4dSFGDpECdjFc3ANkVdd
13/LMUVJWOtNwa9C3Czd/IfHtLUf3Op54X6ZdwIN+QNCGE2M919KzdJC0rq29SkzOoD/xWDHjw7P
JKGM8ln3iPTEiemZxX/iwRuWbqYB5jr0pWSZ/lC+5pMX0H7mwIdGpMYmw4Fft9+NX5js0BZuHqhs
JjzG+9Rh8KuBAj1iywDhQY+4/eHbYrPjI0xnhUgDVNwOzBfl2IilBC5PLcUa7yyMv/IQs8XSSRXc
+koTe2h0IQ65EejPceLljsaAMzOuUACKNZZrz2EcDveZZwDgRKMUNoESNI59B2gtlCdOEXYkrUVD
obgX6K1Gengu5FTM9npoAVOI/BNY6j5rOEP0lE+ktJuR/adFXYtwhG3QKKAiKbBEt5oLZAXh6T3n
CHVhGXkX1MfnnoL0NPlzhjBKxJ5QWfeQPqJLanlFb8QbVs1G3wEd/Fit7VCyUoKBcAU56VaXSx4X
4PyWhQsC091k688O/9FjpX+22VFBFNqCzSk5CvC1SlLaAb1QslUNJrg/45dxSp6UFYeqTZ/NG42/
65EpjZa6LTSf+m+tjzPHDUNa/aJAJZBBCWO5NiSf85nkJ8ifKyhT2NYwrhvyiNO4JtmcVN0Axcjt
0angJOzvKtxNgotjA9mNhC2h5KKLU39YT0H+JI7tCQszkvFaNUMpEA6tXGUiXb9Aamoe6U85enzk
yvsCJ2fwTVEAaiphyKUmQEgF1d10pIOxdEnzLB7dgUWTDkCFEFWa0P/+N+xM8kbYVHIdwWEdZplm
lufBgzUPPlrh8Ke1BBPMNX45ky8m3Sz7qXrWx1Y8m2UU5srXY1Rf+qnlN7Qg6K7salYRmvtTGjGg
bhDtC9ItoKjhVib/vI9pTSYAhPOdlqd6JDa5w11jgnqFaLMn3fLuHeAC8pWtpdf3kKFazPsYsrw+
qM8RSAVDkDjiXxeMSlBQb2i7GIrJTYA9JKtE6GKwODJdIBgmZGMuhKVP5tcie8vdQSGtjT+mfQCa
hj/BZTCOWzUWZcYgdR/bFnuhzK8CokD/FETBGhFrYbjgMopPigxjW2llm+K7l0TVQxCGG+Gnm7Ch
/gvvD3o79x762rGufsO8qv7yEbPDBvaTR0VnErS/oFHE3SUkg02NJyp216p8qnS6g10GRfMbbnTb
wtXQQpz/OMGstuWIYaGgVY2vY3v6ruH6PkRFg34kkTCQz0ixwa3hmHh6TIUfPXBLaHvKscGcVvfj
Un+eArvh0NOL1+O+TMF5NHLeZxTyYsbO9hqYgvx6sj/WIo70XDBPwkhIh9vB70YehGX0zZOxfuoj
B5KWrJ/JfelVUMHLQ58qboeIYOpYvNq97saV9X1FUllaV4N1d+mPTA5Cb6L+URp6wOFZbFtVec4a
3PHNyep5MpAbXGWGkorVzVO1d63mjfejQVOXUyde+qXGrXDaG1LbWSRFbS3b/jJcuuh4I+C3rW7l
9sVZVUQ8vuKxvaTFLcyldio0T8FN4fn6Od2Zqx2VN7ICVCdHOQ0o1oKc+/R7ltKnOBU0viSf3wIK
LNtTTY3zzS5jMykYChnCHHy2grZ22tHyjoFTp8YPm34H64Iq4yh237z4fZyt4xDL6htLkc5JNZa/
vToh+PGwiS3HZUlQEzZ9MdqjR8sPEz/tHjuoMYIJ5CJtf+AX8gsujN5ha2fB64QNPsHezHu4dEd0
8p/e17n8bz06q+yFMU3wHDJs+tgKr1MyIEafloycVd0zr9uqoxgKhcQJaPWc/KNuOsjv5k7KkYru
gFxcDshYejSs5IoBFjshf4IsyCMB9qucIPrxGOE41ivHN4GYSEMrujIuLXwvTYJ6l5ivjGc9xADg
7yI2KH0wcj+7HroP2H8SPdZl333tVZ6NbSUscaMGdZreaDLUOH2fX+BLTZwv1+2z4v2qpyCKpUF6
bnPusd8TsFNPpFxO1OcTssGYSNNf93rKLby/diyu+JQWV2UCC5T/1Bfq/XXXkzT01PhIeRXWEjbk
usS6Y7PuxFpK2zz+EYdoV9ww4CGIwgXuo7Qd22NmsyIu7JujaxJUfez5Ke/3VEzfF/hgFWvbfpbG
VbMPqIkvU9vjrIcrAiVjDnanrkbME/eblS67TNK4OQg6zLS7OekLZ10QU9Xqsuv7W5Je+LiGqnTP
OILDeMFkxDNHzZWw+5RQf3ND42GdeVUXXF+U0IjUEtNFHW/DAACIFfd+6BNreImr5BmW8Zv0LJoG
Fy/utjQ186COsBMQfdMajn0CsElo3+jUxqUCjzbi282vaGTvZKx5hls6kfImOirPXbDd91dJxeeq
BGB3/CX74lTPKgF6oMmZXWXKoS6W4toPYhj1tVYRiFTE5jSpoD6mOt+RMv2lLG09142IXy3j59lz
wWh+RFunAUtAo8H7d4if3ogJ2mQCAXcgZHFnPFbm4qzrkp2hn1vNAGgw3z//pZEkGGE7aacpUhoB
sTxvkTKMC7Z/nkU5wniRuP2/OXplCweKCdWR2vcq4GZuIkXDDLLviIYzluHqbMyZve4ll+2wBPo7
9FEY+fHoa53R9iW2oMfW9oVLWQWutTBpOOIsdYW9QSz20GlNhO/gqsT0sgRMva1/aOAeJVfbEjMQ
3kS2/QbEHETPczplkPWb93EDNVCluRXxU0vpsnhRCr4JT0QgL+2dRIbDDah43OpH5IpxgbgXIuCl
uwTDs8lL3u1Csu8XOY3eEvwZe+DSVuTns8Nr31jj0xZlgfEcwHWsT/fCGDUzBK4wxBIgtjm6n98f
LHYJR3N8rdfAsh02mZ+kbd1PWRerwhDzX5mUF6xF2LsqkQXIBm4miFQvhzHLNCCA8/gSmmXB8fKA
aNmSJN2acdmd/ZnIp/kffXNbhozqI5HIu3CVbNTkrOFKhR5leXdyFT+KZz3noKHCp5fySe3ByjOL
XK3JjlhOBXgcOTHmUFIaGWD3iX0pwjeD2qYNK2k8r4gS/tr3V8UfYjj36EdN52mU9jFtGPWCbGDV
83LjdtgaGb9uKSgsr3TWVxQZTqYuvnqkxagvMHaIXiMXycSiraOQgri/xMRAMQGc6WLW92AhbMMF
QlAUFT7J7yKIt2Q0UVswfXxytwbIvIlhcSuUkHjIh55PNgGXLP9u+UmmKW4sGZgyn1jGc/cWh7N5
+l+JLif4wfYEWlJyhLQiKWj/RKdZrXP00tzk/g1S1rQZJBr9QgWj3HXfuA2+nDf/G52PhnehT4rt
I8gwhwNqV2cGB6+hzsDTx/26QwTxKhEMztLMI4vvSzp7QSGMfKta5ugCP7uVLmbigE4pyyeHz2rl
y9hQULthm9WSzpikPyxgs6UyEpQrkj1n3jwU6rUAohEhMZNJ3LxnmzFu2xrocb5NE5PdPabolDbS
rw0sX36LX0OG/xIWnZzL8q5ZSzwOVDlA6dOBpLpdirWeYS6cNN9Qjeqkd3NbgX78ojkmpV9iWchA
fUpIP2Nkc5enYnW1IieYou0tcibGzy8jdMBaYEFrqrIDsDQsoZWKmrwDmJK4PFpvETTP4lqttVe9
z+ZidmNMJIuusiu7m1YisKx4AbEJXz9MhL9WKpoIyPdDGyBm837bBMas7OCCtEiAOaDUWn2dARQG
ddQJromSDnUmLd7PXkCMJKh+JRXjb0qSzW2DVbHYm2B9SP8u/5PF85iHh/UjlQsPpB3lkOH/OI6g
DBPZc8jR7nrnM5aigIfjaRBSGzDuWZFR48TDfyV/KCbUaebFwUQ+13BgDWGWsfiidPdlA8gOk4Gm
Q3XVEN8BkCg7xUq9REoaLbdaLtCyo6EifFL87xQ7jo3pZS5RntcveH/ENw4HPCNUQ2tjBYFvDhiE
HHfnpb8u5ku9Ay+drpMpR07aMWG8fU2BWgKexDTHbgO83NzmXuVjC9CCfDAXCm+bvpnceem0s+Fc
KzGLjZsFG83sbhbvRVLGIangkLbFd0TFEAHeO/IR311fdfGZXj4FiO2fRTUBQ0jbr3iGLOHi+MNu
sIRI5iJAEsq0EGlb1WF4n0JxUd3LwmsMtRnz6/NrEbDfM+hlgMS7pHb0/9j14f809yE4fkEu7//x
ezlLG6bIOHvmaDICV810FLJQkMVkCv2dlaCjX97nTwICRvIt8wxVWWBoHZxmfopDnuVhQLlQhMrA
mqJTzeFS+6r3pWPHJADM6lm8t3Pv7o5tYLjuYXeZkHXJvEWbbSSdpwLq318wKjCHpaFnH7PWcPRG
b/1moyv5e6GlOlHF2bVZjxJgbR/EOo31Nnr5xx9wBQB8NZZTc//tW9pvLsgoPI9AmifRzp/Rv88q
xx1nnKToiDn/QbQoMNmXLlDSSS+3u+hntYEnNloN30/c3QlEsAJHyXqbOK2vAESQhAF/SEqG7MQ7
2UksYOAI+iu4PQ8eWQR+S4RgEpPr/KnB6u6wuV+J7jwlVe/8EVaB4g32X02gap7p6NbyHSfA3kwU
00bkGxwXNI4yO9vv1lxW/AblsgfnUxY2Pe+Sx9/3ov8S/QLm/geUSkQbiWFxwQUa0BZI2B0F6Yk4
KahfAVsdQYsn5iw2Da+awqNHXf7V8YPs/6cFM+5iZrTsjb2g51XvBcppDqSJzNmnh0t0UtppIVrn
+63tAkgt4JYB7vdEZ3Nz3g9u/hOHKAsTu/QMT8ZLc5cAQa71TKD6rOfcohxK4lLbj3xnXrVdRV4y
QpQ78jz2sv82Y4JtgcLf/RXjX1xKOUXyAdVR1Tq+3TXeg8dG0XRvpoywEUzSVbVdRBrggmEDczxH
SjGMk2zUXpCVB+DLRKBhXeUkpVleqcuH+dobZkRBQe0iGi9pV03l9Lk/qBOkxP99xdkNPQGqLmOd
RgqWue7MAuJZhfw1IETQxfrA2hC4xd5KZu1uNvSgNbv1d2wMNZQ/Nfh2DsUGxSf9Fc+OmvAnvfmx
7kgIoz6Y9PFabCeliLJYyX9IX+4YBhNUzrjPP+pdfwsway25m7ln/bA1xEerpI7tLutJyvAEA9vT
xW1Iafh+T9km7ZLCcQ/i25fcYYeznqAlqvWAXFGvkMQmKO8cCr1NYnScOK+m4sXKcID4Zh5igqNU
/LWyGzU0+n6s9CDJL1ued3Czz/R6qoHT+UjDQEuPaC3D+LYNFnS3vWz+1YQCiY7e+fQpGZYIFDim
a7+P9JW6xIpCiqbquFcxtx0fj64woSSlcB1T/k/zDD+koWS7hyYHi8tQNh09yhICOdkFrLghAXje
CL3jYEhte5kWg2u++F4cft3svgcpqruJoRt4GYu35b9Xjo+tSL2gcN5MCgCTcITHaC2/mRkH5hhd
uBxGdlgYkIZA+KCTof1oXL9pgAdSpkzTalPUZrwdlwnQfbAhy0iYFkH5WQHn4e2IMcNbwCotYkjM
pSO1LttwIhda89nN3V5Nd+m9LPQ8R8xpv67t9qst1B08k1lsPkLfhfsLtgTcbCBSYU/YxjSUlbvE
m3EoIBuTLoB2DOOozHuTgw7pau1I5D4uiJbQWv8zE3APbVG9m3FJZUIzhGswW4ECFBDgGmHu43Zm
honEBS4T97TDnxpbYNyKNvyR1l/yWGgekYISPI55uihtM9/eAZhDPQjB+dqPFwpSnhUPckbOnME7
Cnf8/KpH5l9MFCBaF8qbjsEnXonSn8DWV7ATGDFQolRh5Vzy3OxovPngVcv95wZmUPdcXL757GCn
LVrD5l/XUrxlDFrtUFl4nF2v0+AzH7t7liyrJGGN+ekTBLcg+XuOUBNA2IDmqWVDTVmuMD1LBlpT
7hsjmDotzkAheGUF3ZvG9+x+sek1AsU7n4gDaXMV2++EPpK9OJHOT1qttN6gTdTLs0uw33g/86Qu
mKA3dUt6jx9HAdsGF1KGJiD1poYY9iUumLXHwDIQxswed56vvabIMFtAYrvRsR7uA8AV80mtZnv7
QmJkp9uLqdbCOQHFp0p/pZ0y1rk5EocKaSNIk/ZZ8JIb+Fv9fowPO0C7opZk866RUP8Y2dFkbpKE
PQ8MYjA98QYlhOL6KsZez6xMepr2BHwtZitPik6f0WmeflAiEBNi/QlBRVADMN+8AI2sAbT0vaqP
m5VEzW9NfaLCJpBEHjqoJ/apVdAUSMOiHd/AtiQpCSnuKtguQpfNWGQq3+Tg2uWmuhdq0gjfKmHy
r2vHMkEiS3briSIxX3yPmKfi9mp8XzANUgr4DLgDE6Hfjl/yB1JpCO6cr1DsTcjdP/bTcnFHnVqx
LnMpUOfLPKYy/BBeH7uRw3HQ4t8u41F9XyElEcZriuBvuWLXQxEq6ivGqsUvlr0MpHufXkqQTX0L
WFtxXqt2pS7G3+CI2hJocryfqRWhSrqLCEOfmcvR+q823b+s7AUD+lCIUJ6l5IVaWwHPs9X0KPp1
ZAy4BkwSVuNLzTRbzGeuyQ5H/juBurt6XhFRdutETs3Wk4A/YAvNhq78V+tYeTTsUnIXPzGQU+YY
qqHES3SbKieW+HJBAbcW+NQlX4w3Ozyg3pI5MtFBEK0EOwEsrkgSstWawG5H7kw3mIYcTJoFmvxu
1cgM9ezsu86D26W4gtTx0ToTTGJQ+fxslCeH76tJyAYTEDs7AvVG57TBNNMfEf5K8HlZoYX1Zv+C
wiJBY9DQI9pL5OeViUi03cUrFaJ18qhpErBFZ7VnKPr3wQ/l1AzMQpTOF5tw5Xvhdio9pF7l4+vh
JjHUih7k9i244XbbF+IdqK2Lw23k7bvWXk6Z+UesQBinMLulBLS0gsj2YxbILG5nqsK0MWgMRpjc
UHVgerI6bbsYQEMNlBdnxYC1JZpOEuJdt06ynhA5VZO/kYY4h86EZMABieqV77xAZ1Wt+GquGt/z
bf6NbY7qKrc5Pqubqpra+hcDx/tl67+7DwxpbA0yFKeAN8W2EQm1nl22+pRVWJFXH/UDuy1y7egw
aWF012nmbP9SZgKrvmwmAx5O4ZYAaEKkfwL5BTfhSMAGIygYxjnk++jSe6qOzIOR4OP2DBwBW4X6
tRoGvoJbIgSw8IwfwfMUBD19dC0VGFfx0aTqO+f74goURHb5l0RE5krfxKpWtbv+1k91rSp+c1+a
YP0MCmeBEfYAG030GHai8+GUttjyXjPJeYf2KLFYsmQNhKgcwF+ssPi0S5yKm9lzATXs/9oJ4Yu+
9p94RF5541GHT5zce3OJri5lveJ36H4cdA3yQxjRj+DcwqgIOPSSkqD1mQwZkunCrh6sTtRFdlxt
63R1yAOjBp78KliEd4QaVIbQha5fp4DsfpUgMmTVwI7Z+kaUEkG9dS7OZNlDqAhkCGzLeqoltc3o
7ZoOlVmwseco4BmwC5V8w58mqUcaD6iYUOLbwglR7clpQZbKjySatp9KgQu9MW2vdGHe8rglYyWx
oZSRjuXo5EtY4xuEP/4nauBn+nHH9+n4JYZiixZLj2giBnhfFvF1QTv+z4Haz/pQMLv7hU2WGAM9
Q+7z9YudCoqTi3DyoyrDG41wOLZ7JOAEkovk4whsFOpdL1PPfB1kDW9CXWcJ11F7kpj+jCmt7yZN
8RNz2DUW0xmYRkopUt1TQ3DtQ6Vw2noPf84PsHxcG2NYE7+jcYWy1N8jzNx1OcvWLWRA5lrOX6Vs
Sfhqt/PgzanMD7nMm8hKjfMxdfPN1HWzj9a9jwQbAZbQ/SwbdKvMqDOhEvs083nfoQawh7N3G9Yy
5+6lO5e1KhPD2R18xMEu5TewaTu4i7KgUZydii+ezbwVkjGBxdSLFLTtghrdBO+tBkvTBImbHQEi
bRkxcBDUZGwrLd0oSH6pkhznsKZeS55JgB10fXBf4CUPkvqtLsMoPpFwc90y1+6gWU6Vx1bzKmdG
qOhC+qpX4UIGpUmxpnNGjTcwdq6vQQ09Tn4Qie1YE2zaTbyIbEOIiNREXOxYng0pc02ULOHam9Vw
8nK0EpqFZ+AidEMw5P9DxeURi9qpoBTjSQ16jMIOcXQ6RzIneggAzvn9UfC0TBPyhYIMoe38C81M
iMRqruA+8P9FLpRvWJqnQoIhPuDRME+myyd1DKBcMqOJujQWohaj+Fk3YTQIi9TF49iOfTmp6fTW
/q+XHBmIfdYx54ft1qQoVs9/dShDL37ONmAXZ7sx03hldwv3eCo0zFGeNlpWTjdbEx6oLppIZKyx
O1kVTTKFpQO38V7RgTFfZNhbuYXxh1cZ7e4lxnrFoYQRPdbh1GL7R0ZfWxXT41c1xaWH0PkbKlJp
WD1j/BOSBQg6M0+mMu/t6z7OxElQJGUNGP8eyv5Szgrgzovnp3hgVAi3sseGdg7TwC2X3pva2mfL
oQJZbbqyLn9BaQNpQi0/1BBlOvVT0PQ3dIUoj7y7vl13thEyG5qBGV2t8rb5lfDkoYx3GrzmgjP9
aMyQZluDwx9MrgvTXWTWzot7HhCwdnPVoJddEF2qljm9WAVDByyCR7ZiWc+JsWj0nbhB9uKaDE7Q
aT6IwHic33ZruBfcO8YjfZ/qZVcZ9kw3YiqXjDfrSZRuIKc1IHtzdbQRsAM6aXK7ES7T2yEmlWre
k0CCttMqEAvv4DVsUhbpJh68koldbbDYMge9MLEGs73w3zELkluNaxKha0pnhsw5zWGW0r45h/eD
q4o53FHW6h2yQ7qQoM29Ue8yLdPOVYQmpCPuANMt3px2aB87HT/eymiSeWK/yiCB6WZv0UBgEV7n
lqjbLHBto7NOyNtBSp6dU4pBYflbv97+UPAZaIAHu7NNewEUlF727MQ3wDPQX4ffV6bSVVCPClBw
1T4f72jJ0KOTZlVSWMRCHncD/LTr3HbjwuIjUsfnayfxw78x/hfdVCl+aBWNJ2HdShRZtrL5KRbE
WaDWvef2/o74zHYveGWa8/qKq5nOKPXRvjysPIfT9buNTguZ6kXqXfH7NyyzyoW/3f24fABc3BCp
gupXUV7Uqmd7f9XNnWDnB3bojZFzHuxS63YlFrSTZEnHB5XH3TyqTAENuHBRKFRlCyo03ojC2GXh
5J/k8/CxMfqk8DRLgvSwVV7TgshDSY5kRPpqqsopPYJ0lDSg8NLwKOPtI+MqAbQJoCqfGepfb4tZ
fYZQKyYdTuL620NK9dmchMOEM1z4fR3lQao44JOr5lnvKfLqg6Awq9CqNdINKlIdbvYBVPHsOsbS
dqKiIn5LCQLYswSD53V6YE4j5LeH73zehXrJ76L/t/PzfmDnLPv+O6Mkh2pdUDJELfvYkGvW0MXr
9/mHqxM+vDrUIMIF11W4xRgnVW9hezIFxqj35H1kS7FP5fVGGQysY2mwMFuf5uPCRjnY1ZMrWIP0
gFqu40er0W5JMB/JqQG9SZgPYqd2i/HOIC3vzS7d8OmOVNk4PIM01v1ZgYvnrejPTXUdI7xmH9N/
1cGCbC43dN8QpuS9Das0buhXGrdD8WUQgBtxlZ6CbyZ2Y++1V+8RV07AAcjWiPozDqEcNlZDDJNK
I15+84qUkTQXSlsdZFN9dVEwlIOMuqJ2H0OrrKyN0jDNLTlP8aniuQXk1SKCciXLkphusIf2bqME
KRxYt0gj5975V2X5xztZX3yFzb+2GaTxTD/7h/UUW8DB5E+yvWKdYWb5Fw+wt1Qcu6/d8qH/EC/d
Zl92D7wPWcz6s8IJEZ5ObGIg5u4qiw5R2q/VLKo+kV8fTbDtdu0UvtWNr1twBomTYD+jQ3inO/10
0GchOxIShDgkRn2UdXE09J5T79rFaPawAAeTp6y34LTfHab1B88rTt7izq+rbN5ep/wxL+aUVMcH
VJdhxXeE40aTNEvt6ioM0dflIUHyPM5Jefy+1ZdWZ8oDwyHDQT3sLBdYEMPSyWzDg9Gb/iHObaDi
ld+9syRAg0enDom9k1mEu4Bq7TtS82ihebkE77pqqy5781Nxjt8PzvN1Q4z0XvUbzjseZ6uhkJJT
Om+8wffpQEHByPI31FkZ3Akf8kuqqSEdHorvBNbwj253MdHwpuTFZzQfNpPSIsgJnVVdoU0qIhcw
Y6xMB+v1oppCw8qC1GvNZgQr3BLtzBgPfx1PftgjXa1CQPITnUdeYMz41tX8x57i/qdfTluRRgEj
ukBKYIrMYv71LNN/KdbHdFqoeRzxUD02bQ+EsLpF6gzcw8p8SYExG874gigJK+9Ezmlx3HnQF3CL
/+hwF6NVgkmCk6M7OhcoLxHTQCU1eDcIzFKs8Leu0GSu8UUvm/1fJWwu0PZEK+1F6mOsAqwRgVBF
9OLekUnW2NxgOrQj+U/T6J39Zcoo7Wowuo4k+SzQtWONOkeNYFihBXd9W8Al6A55OCAuyX75TGxb
GbCMc/bq0OAHlGJ3ILFIg5mpd1AznUEJkB7GUxI5hIW8dO4R+brsOyhQgbMdSuaAGzHna0a+A7wW
1nfxqrxfm0xMw8U5eghLbD3CoEBoiQnOufDJLC8Kk8GOgitA/chkbwRVNIU5aUlC+aDxeQ1iPz4O
2hbZW/Hmcbky/h4cmsAVqnGJwDrI+RGyKD+mubHdIYyH8v2AgflZBs+mKD0L6hjaekeKYkn1hv7B
CeJX16ROSr7ht/51KL5T8qzgz2Ce4sVkpfI6Y1nZS/oF8OJIgTZWP4gifyj1hhsGiTxPDduhat3K
m2PVNBBecM0EKfrAuNVi3sJfitodYrON3LKYPWFe7rWBWVAHUaZGysZxpU5b+L1W7n4tMP5HRFNZ
OVzDNUv+rdLEJMTT7wYK017rYGjqwZaBQcIz53Is6pUNqY90NxgTZ0qa25SQ1HuAeKqyuSfegdM4
A3tVkyKkX6esWW6w4soNzrz1EQ8uv13REMXgCiKOPVVG59tgkcmmafbqw4gH/OB7LoTrXTKnopBi
p5Yti8Jc6v8guh6I5jLmJiw+YLYSvbHZ7Nz5c/+BO2bajrn72ySwxgGQUGb/bmYvDC2AsCvdvUHq
9REKyy0EJGF1vUl0UbVrqUVyKWb1BXbP0lWaVdR2FkqdDkAeMV+MP1HkpshruFJ1DKWMD0JDVVHi
kAE38bDEl2ZcdouqVFbKHDqHNV1RBZ5MpIq7XccAM821ryQpZbtLpK6mR1g4wKxZWX6bKQiweY7G
2C752jOdXQ9KSxN7R04h9lodFQyFDiAykrSqP2tB4+pK7DjKkdqHND9SBsRy8OtFM/gpK545hHFA
MNXjxbQx1C4MmfaOS5TvMKMr4a/Tl7mzbUb+VMunMKJgGgxemrzbe2CbxrvqaEnIkyKdaYcHXZwr
kz9A+pRwadoveSoQDuSP/MpcQLviGqay5Vp1bc767G0SffXuOj+RRWkjDINKvE6iw2uKNENLyKmQ
KpzhgIKnRVqh+DR2xIKawlDgtDsDRAhA0aInLC+jKeHmgA7ZWCMTa0ZvGOVyuAlJZfA6ojPIRr7I
nkEPQuOEglFwL6tQOQKliaRVpFnN+bVS0fNMq4KFskayIeCkGl3OTZe0EiQJrXpcqRNU/0qVcc4+
ztoxMjeQ+7YzXTYsc5VdUl9FGCMn2wduEir1goE4Ecaj2Ym7q4hpX07C+5t9W82gC04KVB0Bm1V0
b4d+j9foEyO/PdmJrOORrj3Xh8DusDeLvhl8swjSaWkFXh/gjOF1joZxnHhnvlrm9WDMyU75AJBZ
euSrpOB4LD2VgKYpuIRgiRBAkW82JitPqv0+NbPAGM8j8C/y/iLh1dg2w+Ev3CfxiuCx5O+uh7yf
6cMpqpMvKy4WRYUbum4pN1y6e/Xuuj91w9hTGUzU1a3XBBq8Srna+my+VAa7tiDXNjrAbAi5WwvK
ZyHFvaCFmInUIpRPSR8ikQlqqE8co18lBbshK7eEZrM9oj7d8BOY6YLdglYG6de8PhN9zWok47XN
HkDZmCfMzTAZ7fcVhr093ODA5vlSBMBSB1LdBq1i6KAvuld6AIzDVPW7Zhv67QF8+i9asaduhTeG
Sb/5KO7t+fhnK5F6UD497ZW+JXdVwZIr6a8UBn4LxOYbBQ2m2J0n221IXjYmsuQRR5s3TvGG7lf8
FSTqrqc4g+RS1+9uoG3/J00gfgMKncmFEd7XjlkTtq57cwOo2kqCFsxCuCnT9TTkSXkep+MD+gvL
eemzyNKWX+LL+T3TIkKkl0PKEBptx3lxF3th4ZyTBHtuD1sb67NoFpcPis3mJ4niXndLX0Ns3w0Z
xNZj1sJ6e9De9XWkemLqyc1Ex1CJb0vpx5WFpbLg12IS7z36qJVk1XvXFy4GHbUpAlJOpCU9O21O
uQa9/FwGX0Dlet4gIAItMYUzFS0tbKqvxsvaVxvpo5J9pWmzJXg5UnryK/VWVeTUA1YWK5PFf63D
uMGEMJ6ynIkkg9p1+wz0flRbzrUdKHPak/vJXAIZKvsl5mLDh2NkOpYkLDihS/ipxjlZ1/ZI5SnI
ZMRXNthGSapbKRvc+jdWti0Dbo8tnaD0DXcEtsZBQRrbEwuKv0fT4U14i6XLdVSLfUxF4GY4kbSu
eEFjgaG7Kz6wzN4YIRGxmGVfzlFeiRrt1SPnBltLzCi7wXGbw0LkHWNpbSS9iKkRr4plFFAgXU1F
SbUVTtkifS+Zuc49LKqr9jcVjY8eMPXQ2DCTfUDRzOetpu0X5+qptTn/aMyYAgaO6wANTWOGbYnj
p6Ep3OflsjlyCAjVoKg/Bq6jNlROw3se0YiaS4Ir2uBK+2212qtPEWOkCPN5ppNhho46fanHGBw+
Lnm+5eEVl2himtDoa6FlAEmYvyh5CoPjWNibjPphwZ6ukvEIz6mpeLlsvLs+HFZtuAqO6lrzh1HW
i4EY4cJ00iYOSEFr4LXct0ztlZgjHK9dQfuA9xHU4RuC7epNN5nf4IvJIhGfi4xzj3estzJy02ub
hL4n5ti6srG/QjclCZyZSG5LZQkD4+eee7Vr4+CYvkO2TMkb9tDuk2s6ayvTJhI4Uiwg5INQylan
TtReKoAInYYxoBkX4sg1HtYJuCum01I3znUzq8kEGGzwdpCinQShqJrh+UPM+2qKHkgaZud/g2pG
KiiBjl+xpSi59yDge5mnAKq8PZOQAr8WL9X0AT1R5mK0mbMkSk8KQ70IG/6t1bxNSFYlTRP2nW2e
OZ7ubLhygamVnccwQarp53acmGSsWa0ursmQOUsYHIlpvewceTcWWUvM1iDC+F/GS1wtHY07uVP9
MteDUKwKyo/1LIVfqI4hWji2cQrG1AmQcXEcNp8oUDfFgjjbDVgVyg2uYn/W/7c9Yw+81DPcc+nj
uUliTCNAFOw2KRuSwv9rZACvBUwa5/xCpxuYboyZ0yI0vgvO+Y9wG3Qy+k78+9J6BmFQ1ZpOHJgb
AK2qCrIbe7YF74yww27GcDbQYYVzH6cYXpkmYBmi67u1m8qFCMrbKp1UgWR/Y1CjICiss62xcXo9
s/dSH9p0ij1ekXNesJUwsI0hZ7TfYcKoRbK43GG1W2yeFmlEMNx65BobmRAlcEM6p/V5INsFnwb/
toEq1/eFsJ99Sl3KMoysjLwQ98Jg+syvzL2jytUTg0u6lATuHne0fXbRomLWq+iwwFiwIMCLu4Ws
tPaiJOEOKNRcHDvnnHra9/Y0FCcAprQ4TM0FPVYVj5aFHhBzwqLM/8CxQjhpQo/MEjk5T2TAHQU8
kpXqrIi1pxixSkVGkEjY6OwdKGXXdQs6KTZMFVhdi1lsDbSmfyz2gu9uCbTbg8pme+W1ZHu2Usgo
+pFo91WSNwjMsK03l4m3lI2rIS5Ge7K9FiI5HtAlbGnO/FAT9gqLHJ6N2ogaB+ulq4r0IGwkhfcl
9zpHQgha5Kg0IDUAm19M6NcmrnTiHNTw57d18NaE445KSt6oICubN992BWHxiSX2WTlDq6yuNpZf
yG0+hH8TWtPs8lr4MQB4hbFUk/wzTHZD40sXMvX+d3TCkF0j5n2u+sQKvpwSVwD9ihb8EZI4897H
ZIjmXsHwEEnoy3NINTJtw+qvu3Vb6/wItCs2vm99PcbKLu8G/CvNjs9zteoGPjKLwNkvyqEoYDJ5
wBTLxNvyhx2LSmdYUzEEu1nhnxRG/DFa4BYh/t22QXBN+w84GX3UrFH6b9n+18GlC1ZWklEk1N1b
ayWpaBp6dBHEYHbYNpMX08pA02aS7lpzQvOBeelMnGaxyGTgNNbd0kJJL1oxQ8uquWxmLLGDHscW
MsdAP5OBzu5QUL60zUbNJlTGzibyuvyqRkdGGVdQ+WpLgOe2aJj5DmkWzB09PrgoA8RDL91x6Fig
hU0Z8CGBBl8aacKRu/7I/wFuqhel9mm0Yh/27Il4WPWMlshLadfleq6xd6lwt/iiaYMsOrAsZHaU
i5KtYgwne7SZdwCbDQ0fO15/IUx+kzYow4tklSb3wZw9CvpRPpqJHWfScnwGSCVYqm5fQrNZna3z
O7dl8a98iyfnSEGr2sdg1chSN45hwUwxf2Jxh0vDj5pXzIgGV7A1eDg5IwYaehOXIxiUUptIakjE
09Ofb669w69GaNp5Y6eH8ivr8nvc+A/64kxFFrK0TZsi0PFvGhi8qI2wUEH4t4bi8rxIgD1IqCpx
UnWp/GF76JGGvfOqs+jQ1cy9QJhztCgTYB1x0tu/z7+6gmLrP4EKeGYwLrdAi0wufKco56IPt+UR
ZBO8dyoH4x7e5FgCydYdhx4GFLf1r1R4jbnwNU8gra2spD/CvsOYx42MCICc1QOZ1x0v199ERBFc
5O5pSBH5zc+YwDInQmIfO5xxxbo/iLnhAk1Zw8kmdhG2isnjY/wHOx7U3kWNPj8NXVaLX0hbjmE+
fxkCdkNTJg1NDmE0sQkfG2nD1KbY1Z8EGTeb5HJzu7NyVSl5Prbzuf1TCf9vHiL8InOVbKhQUc6A
2r6AWWU2bCKuvue7sk0Z7w46PpmICRFozhstNmvOGujp7o46llj0UYq9fBqgCTAh7RWsS8alfN+C
bIRbjkAjQCahn1pe0tbUNCJFiQowFMjTX826nBe2QZQF8SMawCCaSaQMvs40aLm+kk3OgtlCp6At
uK29M79cPYpgutwiFdb0whasd8PpbsXDny9G8QTfXIRxhaPHyrPxcAzyU1j+lLTF1liPRS1oYGnk
ED76VasC1STY97TUaVKQhEfaOcuir4JZFrPB/zKpCG+R+ifuWWjXFRhF43zeFCtuWNw3yiwcWXcT
xOhwXYp2FKBRKagHpgiOn2GtnY9iD/h7urPiPq284StDMSi1AvP1OTLKeXNnNr57b7A9RAZcGHMG
gQOU+Yv46zY4YzfVVazaDTHsHZUmG+LdUn0T96r0tLF5UFUqW4AsohB4z0UCcz+imfU2DwxAgY+L
VCr7so6R/zbMxBnQrpPkAjW+I9wU6FUNMQLQ6G0rThaIowEqkO9wkYhDiQ0s7SPvtQCdbf6u+Nhf
fXN048CjjrpwotlQ7NMejIRfmLVkzAat9k3JTO0HXag7KXzKCRgNuj434QxO434934u4kMJtE3jX
ayELASHtRLeOHUVTdbD/ldzEpk8YlTKo5PQb/He9TsqxlRcA3w8Em0Vy5E1EVIhtt/CrXBDZ5EOB
CNX1M9OmvqS6fuqzYslOuVPefzjKZRJqUGjMNodSRSu9TcP5jH803E5yjxM4w9uWSW8/07nmW0a7
pa5P5E6VUY0IdDwqBLbgLqFTCGMO7+SQvX4MbwCESrvrTn2nXFf+1gMkG2G5GRYFnjVFv5bV9rec
tsTzpV55TPzeo5WWLZexVWSiKf4n+5jZ3sUI/IAFH50MyaedfYrf6Fuf66HrfudPfV9yTpYPXtbE
/XfXzWSwWCvO7dX7YkNyH0Xb19vNWK5XC3IcxX0S2tRTkXB6RcB4UOYYcFMUqDhNdz5VdPGXwenJ
TXyPvpGxLM3wpWrkMnJzBZ9G4/dj+jQeBYwM5V+5YjNZYB1ccie6GmA0pCn3wH9Aie4FsMjh3tGe
uDmR3Oi1NrWIcqMsFizbqyu94NAsnq91y0qVLZR8QJ3P5HTvmWJ3ZrfBqKcQaiMRLhDV4xAYw8IN
zSUPFP7ZL58RxXt43xL4k5ATqBfFKTuh2HXT/5PF9WdxFZsT9c7GlY1+fK+zD6kgUshXSqSXsDv0
zpFDcq4X/eP6GNNuvRFniQNWWdtiJOHo9oY5EIOyUmyGNLJfWyrVwDGyOg2Dpw/yPW0L/8q28BBx
0JWAXdpUEehObVx8xiS3aRQtKLM820w6z9FIq4x+W+D/O51iL6au52UPCyc5OOEwVs3/fBQ2yUnQ
s2xqufxBbDSe7AfDKR6pmY2odRbtqYVRp4PDvDgnwG/yNZCoHsuIJYqz6pFeUyjUG6Lwvo0ygsF9
CrnNUkYUkxHeFNpvhdoumH+5ZGDdBt3+cPAVMdY/CIHHPof2+Q4udd4jMov8os7S2TVx3WqFFxSA
PCPE2imGN1aaTEGDB+VZvKmAM1R0aBwzKQeBH/OUIcu0kCJKA8ORNlda6AnUKrjn0EYRyusEi5MO
kyoPM0rdc9hBoyosQKyC480w8eLj9SAdhsK50pRdftlOIRQh6LbH8Xsa5ZRAmCXZM0gPo0jy/Yfk
Lm5dN6KGlq+4rS7OkM+MeCBOIue0HffVz3p5rCNxu2+0mqerGDqJap2XwlIHCSh7hrPR/JFV3kLs
vqwA2tLzh3PX5PTBl3c4ZR9InaUyS0aW/PMq6uY29175PDj9r4lsOH851sBa9ytnsFTtmeUoGuJ/
gfvuTD9Gf2s7xzME9OYswAuuzSU2bvkndUSxfVWUs9pQkGR+EEmiUprYBbseDTum0mzoKD6KmQvv
JlgxlpYzVI+WkHitQsMAwISv4jo0DlVn84ijSE3Mce2glJblIiwKT1W5PsmqIXAW+4erNzXAbiVL
/xCPs7xHl9IXhqiYLc/guVir+y+XJP9n8n2x9eV2kxhTpin0rmoXvN5mNLw9sEp1MFsulJkBuEj7
BHKUUrvEYm0pRCrniu/xtyLS2JERJeGmj8n3o6HoI5M+ppZt2hPqm2ifLKfw13zOuzmBay/+5he9
gZqYvFKbfT4sGTYXPAYU+or+DBjZzs2e10trhJkQnB9hguCEUSZkaz6r9LgOiB7UuyJrZElX17w8
buekzJ+1n39aRZdTUdFWi+k2tpxnD9eVJvEGJBRwhdMg7wZuW/fsuXZSsYsNuKUKqiqTQjuI1a6k
jFY8aZEE5MR4vU+pHFFBt9A15hXEZyGdliN1jHVW6+TpPwEMaVfXSjn70z1YaDEXTbScvi51qVrs
LbfuZt6QV3V8g70dM5Lbd/7Ba3hBV5unV5EsUlFCgO2wCkQydeiVVGn8XBb8fJvNuUPE+t1M8tU6
MZrccmF+mvAyL0abS1gklXpBjxbf5bbIDVaFESZPg2L/86GqafSKBoB1z+EjPVq26HctcoMpRobC
cpjZalK6gqW7kpWyfl3sP57NvV9jkhTDj3o4jeKobcW9I4aDc4JKKi9lpz18ZMfRK0kJQsF9O9kV
UEt1puqYJoBZojg3amb9GwNBjPo98/4HLDibxEN6baqFB5VFXsaNIXk1JNTOpD65zLEBn+c7w3cj
SNbt8gGUSpq/FwnxQicoRge3K76zH1/1FjNup73iAyTjS8c4WushRXbv+dWtB0g601zQNKj+G8DX
y978qrWM5vIBXqRE6tTMzaftM805oOFddyeJGke1CDBqjvrkbPpBGDLvNgN3NufpIzs9DXjlZLwC
pO47e/5xgZs1j/gW8zWBBMv+RE5xw/aPscOUn068D6Ix25OnU1nBWVIlseu6OC7Erh2LOZrP0rJ+
IlGGWlqhEBx6PwQIRYGp/6ERU1dr9ZHiRR7Jc8HajomQ+ds9HVsfwjB/ce1u6s3jiTudf3LEwG2c
LO47wc6h5bWXi6x1mRm1WPzk771Pqntd24wfB/06RR7iPF5ontDjE+r2HCHz8DiBskTG5ijGxi4G
FHsXTWGkF+AZ/bzbySNuDQHOlZFp/5/jiNkV/+hMGymaVwlJsJa0c5aYR8pSl65KpHWS/DqVPIal
F9TUt3T47Rsj9WJLlxLPXS8O+cJcQYqj/jFpnZ4x/fchvDresMh3MG4XaWh5tUcvmgSm+lu3yvaB
fbfIm1nhh/Y9tltuFmJv6tx+8H96G/9BYKYa/lel3064+/bfRPtT/cbJgtEyoqVx8oskvtnGZm9F
e5Wx7sNhNi4mh80kWIs67xGU1EdmZIN0e+ev9wnJ9Pc5RbRJ1QVYOeAVQLWZEHKiDDbe4dml6jEq
6W2Avjub38gf9EZIrw4hkP0H8lQvJjXmvMGbC4H8UTEgLqWPlv0awFJcXzUPteZ5XfnViTFQIrLU
DLipK7xxFz4PkBqfrlLjcdEtBlEaFd6wM3Vt+F4ysp5+ZFip/K8ixngmd8eOsb9mDKFXRJi16Lvi
21aPK0Sg9BTRe4kIY9esNpfvgOM16rLiTAGqnPcxmibUa0pjEwatp1si57/I6eIN8g2NBJ9ESq7k
UaUym6HWqq7h2RRkDxtX+sk9PA4MeHtIrKC7a6bdSWntDP+KhGIlce7Zbt+CS7FVpOi4a8druExV
wlROkPaE4W0KVnjhEX8tUuPl0bU6GtUMUR4uwJh6d1ayVeS7rY/PVreT8wC9zTNTWvUevrQznAWj
aIS/o80jeKoKsDoh1omgaOoIIMM9VZ8GzpLZfM+Uk+sdxURS7m5iiumYUxqJYSU3xCj0iChaP8sT
9+9CKzSJ+gVnQtzotF11GKGL31lPNeaEg4CsQBuWv2aa4gGqQQ85yWz+Ufaz2g2Uq2cqzJ3Q/xdb
kF5jn9k69KwsEkefz9JK3VeZ3asbNCuHaQBoE00Hme9WmoCo1quK3UbvDy1kfsgkPirqvad8724O
FULe9hIjpSxSloBVzKK/GsrqSzD8omPUlEEkr4maSv+oNCWpNe6uVNloeS4w3ObMvzMw9BtF5bjF
2+B/RPXB7fsztYDDdy4a3ifllVhoXoA/QGsuU5sg8I3S4Y36NjT5hmhspaG/wxmmw/be8NfSVxmZ
Xq749O93hjBMgAkWb3leavmVdbTf0qOwbdondXSt4XhFoxI/VHXaE9LxroP2P2ADtzOuy+n85Gaz
cG1tb1Bm5/eq8H0eAi6N+UJQjicxkzzDirhR7WEx7CbzLVsG+S0wmCBcC/tWy4Z/jSmMUKJ/ZVmU
nHT+RbT5PnTO09OlMVIfB5tUtYRyAYNCzKxZKGmt89CEnCWnDNAUBoNS+B1hSOn5W3N8GpfElc9a
8RK0hd1ciIjwMCWAInWCLDvMA4j1Hd59ynhwpXlAowZsEy3xgAsL/UBZ/ZmqNvUWSgzb3Irc85Tn
zXySy+z0x4aw3ab9TIEYPXIdHYaXer0ncLYvXF/Y5qftJ7FuF8qWRtOvZD5a2GljOQrsckxO8kYP
o1yV7YOhMLMvjpifTtvxAXWns+obEHXbxp1tYWBxdo/NFBTs8j6RJxoDiJAFLDsn+9VwgfuWXPte
SKet/pnsgoiBHh0RN0zGj4RCTNPI2gYE0O5rsyf2eDlQB4flQFXKza6jYvV1D1vtT0kydSWE0/Dv
Dk39MBcl75hvBmDSAEdGw0Nk++nmBw9V6SQvJI7EaFgYRMUs4ZDRkuYhGMRODPfDQAHARBPCdAKK
YNt7LVfcFwt7Na89jXK431+qkiPTNQgABYG9o1wt4al/RweBQP2I8dTzwtn3/T6V8dLraG/qLf2E
PSSq7gBXNHyaRnxaAoPaJwkeuTTN8WgyR4tB8fsUaFEWmqXx2wUwIITXvS0EWWf1v9q6OyQSbKlY
kvJZjiWg+TkuCvoEbazcpmQCrCSuOJf1sksI8DLrBIssYGBMWO3y46dvtaaYMR3n/v8I+7mthNlG
c5IptPkKS0P80u7PV99gEPe/4WQT3cnedTCB22BnQR95qlsZNplyrhUe6soUK9Ca9x96xkS7GY3I
4NwjgvExXJWZDg5yxGsMFLoCzWO8Q9YY+6xzY3/Ymfc51USaIqwpkS8HO+9X79/Nn7KlmjbNie1z
2yhMrlN5DCjuFIzogwg3YDbyQFcnj7rH+ee/Nq0S2POBHWTbxM1cqQtWlIoQOp9L66Y3LnlLq0T8
dyEFdU/qmX1qEjKwpnuRzNZqehHqBLrvuWmuS08LzuiQoPCEYfLgGlKM+HUQb/nwYONyHpJ1bBWH
uYcRTrCSMB/uOPduJ9LUB5NYb7/hGDynqrnjHtQb6OEKFZD5HmNR+dlvTthSB6vMj36d41OXHRW3
R3wCqzDn0Yj2F2vBGmCAPNDnEh7sH+8YGKMYYUT5Z8qeun5/VqhlffAXG0ctr2oxOcuuSA73tffQ
zKKnWiKahXr6hy6GU1h9+g7bCLagNIIWuiPnHy/einuD+hM3CV2vajDVieW8mJ32U+PS4wuqHQP+
LNjhA0M2lFaBKDwcfDjSy/iIQx11hrv/n07Lqt6kmmkOTYzAHgdLpwDpnowqTknIwl4TGCoxkpmE
emD6CDcKvi+Ze2XyhT9dS36igvOFLJnTHvjAPhgTqCrUTW5FuoniDYdSFiN6mSea8O7GbcyJsJZo
Xrneujb8UQU19pweG7L1t4frgCOPJLHc9z5eDJo8z0IQffhgGgi4uNQqyV51mOojW/Aeu/Njr8PG
KhMAslsr5fW5MMixmkRaJfqG8vqlQbNduoTk/iMkarydEwqwRvXImyTjn3FKBEJ79YLOf3gwREGB
W+bzA6gkwnKkfcx/gGG8Zag6/RA+Zu4p3Fx3i1y+DygY7JGhSF5KHPhxnyEweAwN/BJEJXvtpPb7
yeRpQbVz8jVRxKDh/PVZOJKSas9aKxurEWm9OzVv6/uvqZiP3nhkggXTd0WySzGcdKkl7AWBSplg
c2IQrMPRGEjGmM2oPJ1lljKbNPzXEEJeRU4arPurAMdwBHBhu3jFYCOfdfBG4S+Nq7QVzoilgbFZ
xFcckb9JiI1tD+k+EV/FBY+ZrB6cu+AWQfZsTCQU1urkH+ElN+uLcgXWLlEP7ZN1+lyWVajOFQ0F
WX4B+KuWD9G+w2BbowMkH8EtvW8NroMT135cAbbHL0CZzCijEKekxbJ3S/t6L3DCW5yKacM6gfxA
aUBPfP1Uv6+r5pTrzbqs5hub/i6Yba0EQMp42NAmesPDIVSfaaLIf84sNqz5y0zEILFoJ/xawnQH
JkHguaO2sPZv2UDQn+Eui8/zAid11pSLyixpJgOPPR7iPZDv/OQH8r8K4Jn0xmxcfsHpOsiii2mM
GilRGb0RURei0bDbOPKo9USfWK1Mmg+sDU+Tvma0rRs5FjGMHcH2E5YonK1NKW8kDsCDPqm8jDRe
OQPc9j/exufPLxR2EXcHXV0pBgKAYiTP/qRhBEmcpf6/+JsxIQYVJQXEiPR7tpeaLbjD3GXYSHJF
9Hbb0ASJhgI1RrOFoZzO8a2aTfTEEDC79+0SgtW4EqrWAP3z969C9zxzErPeEKGH3i1Nm7mnnju5
A8KTerBts5PDlVcOgND1kWumlLemw1AZ3wJoVpCqCqWtkPsTBVfNCrjN2F+cEk4p5WmqlXST6b0m
sm7MHrITanfs1j7JMEHFKVakCjtAXj+fmmMcu/4fVU7StuIDsZAulE3iXXTbdJPgQVNIdRHdo5+f
1smMuwbe6/lZDgfQh78l1Efi4nBjk+lkKMFTf106gHN4nFY/I3pf8lbnZTp2a0VhXlUGXbQ/HHGR
EF3BbhZtYvrXnBVo02ofoJqFsxvBxZeXtp0S6K5VS5GxEbEM4Ky2gG0pskuumT0ny0HHVccAiF5T
PRibV4FdMvH/lg0ZH5wnwmJVa7/M3huDBZ0GePe5d5qAQHe06R2Xjq2y1YMURxI43z/g8Q3rnrwP
PEEXbeSjVXSfpjSv/o8yx6J761eg0avxP8BZxW/WthKxmA2RPYmRASCaczsGKCDEiWR+vIeTc/z2
MwuwDlt3To7P/eqnb28036zSs219fmWu3I/qfs9kc/6uEyWvVCI3VvebfsTvLCSoCCg7fFCHrXBQ
GJayhbYnMGgpg6sPSGMF3AnhYiuvS1dFDQx1zw4NbfyRbNzl4J01Kdf6ri92qx9p1d0Eh8hWf2Py
4poLjRkEMo8PZBDBWMqZ4DZKtOZ82AOPxXpYSgASMQpzmEWIzA1mWozFDotyeQA0fhKh9/x2v2k8
DEjfx5CvnQRffH83G6q4wBCJxVwLysUCSqhcLSa4ppWwjGTR7VJBD0CDEKsA+y336uRnw+ly38jF
qu8vLQrbtax+ZqCPhLqV5LqhOYXXEXnEyOjIWP414vusNuxvH2iDSeyd0k/tRlNJN7VndElUFDvL
2wOBB2MbUPDLRzY/AWmw2ZEaspUxgKrqvqekz7VayG1hrwM2eKU8cKKw9nzTWL2q5OxaVP0XY7HL
YVtfdsmI8/QIBEBmXQ14gwx3bsyCxzgk45eNFSR6pM9zzwEsxfZhd1j/OLtt1pcJEiqLOVTi5ifl
lHZ4aIZf2ZsKpzLFpXa+Dt97kh2cM688dhYSlgQ7elWuOE74JGPMPf7wf68IeJPBeGVXtYoicn6w
Lk/V/ogXwZC14C0PmvBWMqo0sW2T4962DdPDtZu78MXrLPFPkUpfWvW17flv6Y6dCsfAN47CoykW
CfYF6kin80G9CE6UaNCB17hIKuFkx7iB+9oOabPWNgO0s/NXpRMPIRh4Z/xlqcMu9IOfR59JRZri
8jqKnGXxlm/9ORbUw6QyNqkPFFcq9zG0+6R06NRBml+e1tgWlwNatBQ4KlEso7EOA8TAE+rBVEoC
Zf3fcTFkcQNLmW4wE30BwA8JDtjSexc5Oa7tHHOoedpu3fpQ46iOPCv7eO8SpJVMuBbYmcaIH/U6
KMs+MEkh+bVwZryIO8dq7w4W4EN/XoAhMT6XtxIoAlV23Jdl/Dmi4gXOGe/FtcOmnrH8D2SKksvq
2CrGZ0JPWwTRQBw9wm/5XvF3aGhvq0clNzh0aatOnJERunGMJnSBFj9Fhp05F/T+EC2ZTnUvQuoh
JFDlAEXGcWRDeqcHCTc84/SiZxNwHFLkHZwQaCT8o0hnj54VomBSSlJqymhN8KJmfnYe8L34Qn7N
GWIs1lHbR3vxIDBES9aCd630cgkKXNpHw6Rdm+6e2pBNr6W4WqrP3k8+Yf4Ba9lmx428aeJx15BM
BlZgNrqfYfPQFnxmgnAFhzlslwqmpXfYR/qWUGw0imv0vnDZdxIR8CjJuxNVw1JJw7CglFz8mon8
OUX6Dyd+2iM8phDigKu0EWYHq67Y5ldpqz3P7N3MXHevq4w86lAgHg8D9Wu4fKmjiOha2ICQ2wvm
bSE7ZBPpQdXOvwcosne3Dj+HQJgEpQIVj0c/2iWLAP9/x3XTLyHm9gQvkNVLnyVRSaD95LOLIb9h
hV6BELKLjmaGYK64I+ZL/dk6oKgS2SKLwIy/Rvfi/Wf3FTQC0GbNDb2qFCpK2dLbIWX2+SX/OroZ
9vo+huW7zkFySjX02yOWCMHckPkbWaj588OqP4lHDQB804D+qhEctWLcMqqBwPdHHIuCXk6oeer4
/td4PKsTuggyLqhwt9AbV9ip3vVVBglZ6vNo3H6zrea2fDSI/2UJIFVagBptSkJ5DPyfoOcmbddT
5XYkG9odrVQb2fImgfwS9Si0PDqvHNARl2C2EHs/HFjdCQHL+ImCQNJUBMXJMplRJOCwYdpLIbGM
YSPy/NU9AlIhN3CKlviohUmycyWkP3sHSJLQniKVFNkakPQbEbVYMfCRZHvqwUg8klGUPVfB7IZ7
miUYtkFR2nyaRmKAKTQsToLVZZdCVngfXb/A0darqsTyT3deb4VepDv1rGyP6wcn5Sm80Id1odE5
2Rq1lull1n5iRdmDdpfyQ/4jxC6modmq4G6f78gAvUaEEBh7c/kUwX8bUyyW6fB6cRU5TboownXv
fTZtmPAqNZu7rFmfsT62/h7mICkD/WFASXU8fY+X+WXMESwgZynYGPEy4enBFjfwlCTpSi+ETBi0
hUtJFLFfS2fAhYLmroRYAGEuRP0CZHCRYouo8G5mqMUQjQ5t6bBdzixS2vATxggZtHLExG/P845W
cDM8ZAViHigLCk5XPwL8XUgq7b1BkpwBh+V8s2571bbMRvxYHV5utMN+4vfbP+lr7aQDF5no70Yc
Fs+fZLkL5qEIK6giypv8kjCjeSpnR3nDJ0If0O5o4W/wAscSnSmO7+0n0BNc7dU35QP4Tlx+Qi5X
cyAP2BZv2Rt663hoSZ5nCqxxJ9SUEI9jUsFBqtT4dPLWY67HrCPmVw5AFtiuiT3vk5WhP3FUPy4c
fN6yJes3YIWm7EoHTG2xTVzRVN5JR9ljmPzoci0mZZtvPRmXaoj3fcu9jR1I37jN5tfBvUFxXP6Q
ammygdJSTzgmgv7V0aX6Qfc5ZwDtJc/YW87DcRrG/n3Z58lQUI5RhNz/lBgeB4AsGvRbr/k5t02U
D0xQWi24VkMK7pOeNSYF0O70vpeKs4w0dDOYZKHItTdYGa85CKj+z/cmuylt1BU/yIU5Hp5osKVY
EATMq7fJgYuPzd9GakCR4aLoQmY+dxDd0WCi6EkpdvHaIyKa052MZfm9ySVOnktXC393FsFgjAxa
v8AnpbSLMs9Q3BHCLOU02HhJpm8TA3nuFKgodPRnbfPVfZ6wwEuK7Vv9B+vaMArfn1X5hWSkF0n/
kVjO9Gt6GP7vGBbjAOrSiw5x1xx+UhGhci/3HSb8azKMloQOh7BqxzkjeiEL2wraRungTPX9M5t/
157eMrCCgonNoPh1b2lee9hdTMVS6zGniI/466GbO+gOLynWTyp703E9XHM24O64sJvKmbF4Ubz9
Hcpg0bjDwgJW8aQX10LVAtSllZKMuqquaN+BTjKvF1wJXI03itOAWLQzGPbjnyjmkZdND6wS50zD
y8YIN52FWxXx/wGRKek+DtByGreFFiSkjMc6fZb+kuVwqyw57rPN2zV0VLU0n1mkVU1hzRfz+EqQ
y8vEe2XjojLE4v2RwOb+WqJPHQCwLPJhRHh0IY9jJZpTvmAmAYJlCzipiopf3OuXDWTXg0IVxjzl
+bNlrKLYtU6LWsHNt+PMeDQCHU1JbP0dk5q06Xc8wTxAuseeyrjo9pUcgA/D2i8tBbb4mfCIITka
wDxrv3houymkzZTBL/nfBV/xl0idLQg5Fn44QgDxL0CrX9JFK9hmUg+RFL6JY7tiRCw5618fNskt
0C7+TLeIzQOwC6311g7JIDgkotvtjnoivQ2FsiFsSX1qmYZ5q92UK7hSp5GxU5sJgdJXGVwNzQ3o
Aj5qAQk6a58D+ZIkfLqWGvnY+guG75BeHSRUf7jtYhHd2oXihTaJlpc/vqU3gmw/lQTp6NPdxXFl
Y4bZlQzsVdRKHLEJg9ZP0URpyXDFiJot5+hGrFEmJv7Su0vFdyuadKB0vyIm+llzANf/y3YbHMyL
xsBae/5PgVCJIuD2Nh28o2Uc0gLza14p+jQLVxw7AQOYYvzvBSfLWXKuIzt+/6pVV1c29WtCb27E
7kpnawJBYtfiwtMA+mDubn8YnnD/92Wi5p4mE6UA6FEZYkj8pj52VRXXxIYHkiTxh4DbXpNFFNqK
ZyT9CMJsAHw9l8SzVXYuaRkWwG24fkPwazkGhm/ndI37pJgXImb+xtVok61u6n8HLVofs4barmFV
WF+EQwoCLDgEVhskC0+FuIonfYyeh8FC5pVHUuiZp8TviO5IGGnQkvborE8dUshDOlDKFDAXMVRL
l7NaTmcjR3jp9Cd7BTVvV+ZH/iPZ7uJhf0pP2lqRVR0/oTUhbQLFl2b+sYp2MrYnT0RzTdZTFf74
VGfeE+ljfPEoQjUcIMMqBysbi9p8K9fVBRSM6zZr3WtVGmCNdmIANRW/shAhQbxILGWWMEq3YiIP
kKExa9CwhKTvwdTEvi3MX2KOcnuPyMoAuINiTjlYeVuuykiyt3H10nL5YeHeSSkpwbuUTK3YomA3
XveLHnuFGoou2RDgUE6SjlbjxvS06C7/pxF1zgMlRaYe642w+MqgqqP8oaohwm28rJ6uHuAs1WqW
qOuaFbOBoJxMIRbojjgrjPCkG9AQv33LNYY5/vB4mI1SHnkz9owT7zFiHIcD4RLNB7SfGOfaWdKk
Ffu/ztZEmb4T2UXNpG3YA12lkRIQ+2cDNKcIDeeV+g4Ojde1yzpKnwNprQGfu8ByVXibB3HiQ9TB
DqKMBcBs9c3Njw5brsWPM418yVsDV07kD/4qru/6jxzZD6/+4oBxOD+/FsKG7op5pRCcte09Vs9p
/fnFN/8lnEWqUQOpuip8R8jHGVK75PijPuaCWom7HhJ/maBJDyvPc1aNB2Z/4OPBs/s20vcw2RKd
ZG+hBf5ZheQFBhBx2V8eblyNx/VZGyzNEv+X+/PgJPYqgs5RHWua78s1K/D3D0mj4XsSArm05etI
xkUzvRWsqutgjHl21mgDdk0mksClelgsArYXzfu2XPcnY06+rWK8s6c4tzdsT4ClS88FO4RhDn6M
dT+aBtWZo33IkHMaPw0/Uw/ax9hp0A05Pk/6+TBlgiIB/WqQ4zRX33fkFvs5eZPfEhUq/O8n8DuA
eS95uaUk/sh631gi9bxG84P/7PWihoJxY5INg2yoxW1RqIr9Es5HVYBzeL/qjK7PuFGLuGX8Cl2J
51gZJPd11AmYr0doK7sUl4VhMu41Ay4MU2AIGtPw8X9Rz6ReqCU5RiZPNDfKb+XwQLLZSoG7JUMr
yWFLLRulc1rTASZq7ogjGs8RUOVO/qxHyHOCEKlEqeDVZ70/BQinBVYW1R/1cSN4VLkIeRC25QgF
bLewUS2Jpa8Ogn4NMFpLIUgx1kVevI9bFOaRbNYSiQezGwMlfGeFKeq4dJKOPrZcTzU0TPNgQ/yi
dwVsoMLss0BChJVxrjgkdx0wRNeb/41muOtI/3V9hJOv3h89cPTd3Ur9DUGW1dcNZydx/p5tgVIh
hDoNcF8qn8TJqyKzLB3TdXB7NL6qeaE9gKj1h4U4QnXU82kN8vM94slWd3foBajCcOg3huX4btNP
uwPQ6+zCGB/XdAxUblxwwL6v08npeDe2Cz15CNjFENYmiBArP9Mos1XwBBdnuBdcTBRaNRf4keXZ
ZSNJlcJutfuunl0nPr/cO3MdWQPY/QUrr9iVGsu78tmEq3PqSmy0AAwKG1owcUQXeoe+r0UkpOPG
K5WGe/D33bTl3Rh7DG9NFYz3sRjGhYJoRGo+lpJh6uIYVzmyiSQm3x1pEjOZkAknk/YTFYb02eT7
3N9xPXwn4j4PQKFp1tpKS34dp2PdWPG6P5p0ypvwzNYm74VhOM7P1dn1TuO4xfymvzM9KmXTrV9P
b0n2LGHfh5zEQRxw2YNy/EepUOUBTLPUTtwW0ZRWcCA4/GbVV1NjG2wmX27c42YASOGOqH4cX11e
TNcXMmktJx1lu4PKR1CA+YGZZYMKEzQzFAP5TkDlERDPF72rQynMVpkQx9Yboo+s6f1uazaeUueu
9yYj6BDlyuAP+55eLSH61Zz9W/B+zwmjPXRkDvCiedUxmyX2cUUPKXUEOlZBGPln0SPAUILtPDsk
jFnMRXQQ9ChP4O80DsD6Za0HDvfgqTwLf6VArzCEaGjw59Fjz9g2k/JluuGt6GPkMY2wNeHYR29M
j+LcLZ1VycE4oQtI2D9l6qV1edoqSWa2qqJ9VQ0A+9xWW96wTyDTxctZibMmSyOZU7tV1X91zdZh
8RKXNXjgdBEt8po9LTP9g4oSL1OV1mC9wcia0vjFQ7/8rod2Qa6upwAde2OGSeEYSpQjKB1v7qbD
IMzircxuRmJj/B7wyxfLgH37kWR++Uf8S8qWWa9HeNnhMkXqDQ/HMqtTqP/g2r1uUw7tHJ5Bqa3E
pziRnJdBjm0XJ3JWG3ZxKwsQVlpcLC7pyVWWfWfHFc7n1+T9ZSex7NiU9lxvn6eR6p4s0Wl5YWny
XQUwB+lGPzOFTfUvkhG133WyM4kA7El6iT6yAy2C/GkDe+fJ3djloMQQnYrh1ir5QZzSovdJbxOl
yE6oFJd4cu7KUCJUXMDLkK2LS1E2QVFTtTBHeLeDrxqXK0YAx3wz+RethsPLt0rrCkqyUi6zWpL2
ohU02xjdz6C8Q8KI3aqMkzgvPvnZW2sFIqMon35QkGYeUAtWxlJnTkJvNpjdgB3gK3ZRuZO/YjXX
RkiAl5rlXA6+evXKXcuh5la+OGgNYVpOa7ufmyBlvb408cPPEvBsk0oVsmU496DbH1055/ZBXqJx
ui2zHahUkRBAJmlkBamEE8uEwmagU1V+p7jvFkgIIvjcKboS/t7KRh2XxI/oYpAunqTU0h0d53Yb
PsXVOtG+7hjojjwB/o+v62AURUv4xt82+V3J9UKnsZq9nhBip/p7hOYDmpE+oSlmcvu53DSZzage
q9CTG0KdpIuZz4YVxbsNxIdjsQs3LW4nonk2pQlazNqeB4TRChr11fP/oAtp8dXBxsatsB9ywcDC
5Nwu1/HdswOYsdkdkpsefCbZnzjBlOV2/a49swe5o+nU9C91hJ6vG8EChDOiVEkS1QL0tskSTqmZ
jnqt31dxZN4jd68FbiVecdgZ1gxkeUIuBk5zrrBmVFQ4YugRjUyivg1eyoaAqy2apk80j2RdeCE0
+RjDaK9eK5dWUHVjgyu8kj2jiP8QvD/TScPYVW5j/ZtS1XhGGiGKiLLoIBk55f9JeCdKptTD4rLc
8m5N/BDxCiXHObr1a8s/6WWjCArDmR6vZj1oxhI7INvcVHpVbd7fooTVZemKVwLl5XGWYv5XCHLB
mAhr6ON6M7rKYjX3bq08pJuyFB81rMw2o6AGb2pHi642cwPw65ISUxjip9Q2rrtNTRZ0sFRQrKae
H8+ZEPOKxgUGai171RbIkS+jzw5qnHWgDu0FLZZEPTM60GW8NM83TGtM9ZIDGWEI7A9t52d6kadV
ZhMIOAgMzMCkAiKDYji0Wk94qtDm2mH4c9dFLWZohGX1/TdVx2TnLGv+GOIcpvsqR1uGV58Qp2nS
B2ptrPRB9wkcFEP3uAVcWby0lnk7kR83yGWyHUdXwNun9tnmHvXr7WiJ8DKwnrOfcj4gZiagFV6A
wijiTvU+ihkFgFtL8Pa8ahYDUVwVJvCDGVBVaQ9OP1GURqVy2QfmA1m7h8wJXh0WYBDwCVEm1kmO
mgkRvsMnJEjsXYvjnfZGuD73RzcvwmaTBInmnAdgRDIkx8TqRaNbqHYrGBtZEglnoWpigICok+bs
96+WPwWCYOlEunJY16zvX27cIqNNqe5/WUTPxC6LsJ/9k1ii5fZ4OO7MlA38pkpGnYm+Dwqswf6z
hFi/hyub+mx+w307ZB0BIBaZjR4NOPIdnneKqrxmqydjBcT+3S/rqPUzdXej1KU5DtfJvYBTlVbA
FmlnoRzfWb29yOEGe/Te2zLSP1Aba6sj1LpSZd8e0jNhhnxND+yn+mrIthpCxoovXq4Y+SzP+cV/
xGyzGCV2L+ZeZWKOJ44XAwJgsZ7wsrJilyW8EvmbiXog1pAOcRf4dEHTv5kPT77yk3ev1rmWB90V
pSq50MrrytVSwvSHGOA4s4YIRb0lQJv/WTKwozHtstCtzxpoDntNVATKFOahqgdsYTjbl+qUGVNR
/KknOoRfmBTXsRp5yJD9fgQeQeGxw2jmRrRxSMDZN/R7q+6amv76NUIaLFh3867Qe/Oq1hGPIVZi
jcbhSU3Lfxmq1qNZW1uKBB9+1Ti5A/87sJchdLEOq6xDknHvl4ZnA3sIqsiJ+77BRn/4N5NMIMVg
ufdl2bH2Kr+0QFiU/w1CuJbmO5UAf51lOn7IpY3w3KdFp6bZB+CNzrYWcJze7mbMirB4z8DSc2MS
cd4VQ3XxtppoW24RQ5WjNcoP1zK+AWQ0ZrQybZ375hMNJcESLlWfITRYTyglF1v1L7lfOKCoZ/vv
vHeHbS0EpKjf7XH+mohaxLBrQ2PTdjg+TRA15+kzp+AWjJkZrTdivSpnAxLpOG9u40C9okU28WGs
pc9CobxXyyMa8DnxnGJCuRE2v0tqUSAcch21+DuMlgBNdC6PWoIiiCUq+sH6MmTEHhnFcjE1eIeV
yxpAz1v1bafB32+a6kEvpujngZFhJ8fQGldL5xRsQYqaNSTeRMTbBfC68ZrFcOCm4i9D5aMSaM7T
dGNktgDVv7OYDo9f7ORNe3OeqCKb218WVhE8U3hfnVORQZXzT0u2oNnIl7VSw19QiHNu5ZModKtZ
Ft9JY2+SOOQwOzgwlUtoyTYmrRv6s4tRAtX/s2tlXVbx/IlHYeV9swkOHMeY69MCM3VHpQT0nsDi
TUIobGCm6Gt56BAcPLgVMPu2qlbfXse1w/D0Xs66hjNagsyqWl/iObQiTebeS8ZDOO8F38fQkACc
E92I2H6nYnYUIUeUHC3/piXatEjk8yd620Avxrei2pOMbuksD5wT61nqWMw4kUF4Cis08bgkZ4FB
7hSeyxdnNfJjKI/TeGD6cBQ20VXPIvncB+aNtXaIzbvASBk5GBDxvFTcEOJ5nxh4IS8pkGxcXT8O
G9az4zDfVavRoziLJS0dWStuVj7gQLXtde/TlHhWwUmaJTJHAM79yogwhq7Nigxite+Xl7WRZbUw
DKTkiNjNbEn5JGr/byYYmSTS08hVVKiEO9Q6li+7+hMUPCacjxWZ9/aMMpzouoFs9tA7MaMsnbZP
DqiejF80UNt4ANTHxsaj0jGI1Kc3zh8GPKabA5LCENhLVAMuidK0iaugGsli90wqe/0OyFtBzg2A
xQo+0En85s2+LSXgbarAduC5eK0jUF7c3CE1E+rcIfJc/NyypaHQ/Bn4t1atW5WvyqXEdMOCTErf
MyKIaZNeLAGD8QqfMT4st5YqWx86hLJz2soZOeD4FVj7KKBRCK7q1OjZlxjk+l6c0OZfoEFv9ORB
bshOrlZT/4kHLnhijDy0n/6Flyqw3hnDtyDGDOxspdZ07DWOJUwUlLblvqyQk4JU9uroDIiishfa
tA1vqRcSDA43/G9joGEB3Dy+TLWOKqshmw06dYr8F/0eQHqguTu69wz53B5vxSW6/T5JM00mnTKn
9PzrcookHarCv8tD9ZhaWWsGziiP+Dakw5HplWM0+GVnk4V9vwgnevXuanqiSvDKlcAAc2h1Ik3D
4KBFcd7vmSQDKYAh02D4fu4eEIbQUzQKrOeQyojFjdDvo0pobxc701Rz3hAz70r903KEIO6t2ugl
st+dBA3+xYq2jynTDxbjjdEvMJqSNxj0yGXD3y2LY2rgZ4p4q1zmNS6dA8MywbKDHxXf2BBef8s/
xfC9LapYKba6AEIFUbD6luu99KGAL+86C5Hm33AFpV8tbaBTuI1315XdPBxTEgpTKykAdWedzh9U
UAybgn/olwhBt7e58pWtIOOif2NsI9J1KP0Gr0B2fz8QvmmSsr49dTVxoK2b4/bt+zeqASnVsc0q
XcEpTpOSB7hUyscgpomVooGLc5c/evvQJgCLZrix+KpmOnuRtnoDrPvmylH6m3E5P4jfP/8EyPmR
BGLj96eSnpiPwxjamniRCpmJ1GFkGy12uWOIrrBuCK/AQVlWLJ0CbVSP7+X/9SfNrdMDmTdQicCv
R+9vK4jTZr0IfjKY7sfDWPub3LdHJpg99I7sf5+U23sds7/RA5mkDy1tHV4AKCxISXMlv7/iu8Pu
DIRGrHiS6D34ncdj7rkdtC/HQKzw5px0SGvoG70H2YhE446uUIdjrIj18LMCou1f9W86nZ3Qc04P
73jzOEqRg/P4uy8famGGpgoBJlapJGQ+JZC6pPsIVB0CkJUikcrpQ2h/GVeFH5FLI5Bd9JibHUhh
gxu9P3otsOzBjwxRX2nDUpPq5+nd8hqG1f00dQtmfhJnjgaruNmjbghMPpGW2D1JaAVF3oTxcMj/
G/eCXSnkP+8A6JGSkdvSNJxO+RDHyEBHH3ND80Gcx8nO9Wcmm1F+Zl3qonOH14TOrf+KG1oFYEjV
vcvdM/V9Dr08e4/UvqiGSsjnIfphbszn6lVCW6TjT49FsaOxnn+y1GSKDwTyj8QZnzkOnO3nTgGY
sNb1ARRB9v2qrRVTIHmTOgfiwwCFkVXWb/nPETAzPnZGf1xIma3vXTxFk+zrF75QXu4sorwxWDN3
qCM0pfvPT0n/YCVYMjSVb3IqwajEXrgdnxfPZBLeKcwyan7aFapMHLVG9hHidxrurHjnQUQ5mRHz
FbezlxeGlr6125WLuD/1qzjXqxGgonqW42bPd192/QEgWUpGL0bMqchuNj8Jk1LedC485sO+PicZ
DZHn8G1jDHuj6yEaivzzJHX8PvCxoAs9de/U/wtpxhR1N1Wy7DvoA2qvzt7uK6PTADVSjoklhzmF
yT1IEXeS2c+JNXsro1D15LfN2YW49Gh4QGjXZWBJ8IPmsbMh6K2Zuw+IzRapS7wdw7OVsmOmn9+d
ac73iKKZfmKYlbdjOJj9Ky+LN7iqxGRjXdJtrFK6W0o1yAJJVep92OQgPfiphnkLeXEdImvx/KHe
ibp+TWClBnJsq00uaq2Pvf61h3gmP214AT07k/qnqTZm8xCW4gNKDY6l1uE0kfz6UqQbLX6XVhAw
vr29tR3gQnoo9t5LAKW7u4TRQtmiRRnwTHbRmd9vHYU0b8lkLAtJRXwwAiho8q/RpvHTiPsP2Hmq
Q159tJXtEjEsb2LMDSWir2FcfjTupsL2Og4yCYgroHUgZOTo1dv0wy3wNEE5+GLzNBcCxIlt4boW
EzOw6CfUANB5W1tbfcQyUQTHA0k9YJko7rSq6/kacQf7oO/uGfyPg1j0Xg03v4l2NpPekgHL1Sc6
aylxXCjM4FQPOrjiFcYqcPkuwKRLQ5OOahbI5GKuKzgbPJC1K+jZOxLAg/SLitqvwRGTQ8SPW/OI
ihRjuaSm6RvgkbG32l++YKGSwjDwvDvDdS2yi3NItnrJfsfNwLKeChWSeQrm6gtphptPCiFvqZ4V
sW05vRPTpcNUBnA90twhbIX3ODjI3mIoF7ROiFrKCU8QMzIqv6W7ZkedxIT7Iw7xT1gJ80mW/Cl3
NGAB+InpMcfzYNAjk3821WE8DpW32lkifbFXRbNgxrHDXtVAzLugYGRB9othL6v/4ciajT6ziqPb
Wfg5A4S9yHEiEk3hvpOS9fTBFME7/4IvbwJe7toD9fTqyW8WwbRVY/EMvFG0HDokKqPYyHibXprT
S7W2hp6LNjJiFxT8rCVTypJazguAck74t8KliN61AWG7asdUKmIckm1YBf58x4ZpMQA1cvVaDYWJ
AxvTl0YgXAXrcdGwJPsjUWrPtXagjHqUSlQKuCFvkq3VM56o1oe3aR+ZeHD9LklTWMZXHrpKW2/P
FedVVBT95W2qWwscBXl4++eHx9lEFaGiHKZsktsiN+732z9Ce9XxyJqNSSPAGpnFWxmeIVzvCdTJ
R6t4sLeht0iL653s0fyprca5nOTMDDJpkfCf5J/aMpLEEPtRqtp8hUK4D3FMBKEFifiVYGBEmHfA
IqSiOJDDPb9bC53Lh+F75zRfQ0aU8zvRdgZCFIcLeLnJdpx2VLGe7TjSH1se1JQnGiFPrVqyzXVD
jhI8853TvUa6IABRMNXOL0T6IB0V2h6KrSiv85U/4Z1p2XuKfTGW0l1Jfd3BKkwgLgTneovqKLbk
Ell0R+1x/TjjKGMKTd8JUdw2kFuhQHvFECohDmnrTzbRoUDTMebAKRXfyW0fc+PkoDrsN38jfw8g
ortaIS/UNzUHKs140bXgPBCeAz+OSibqgnqGl1k3C3Hi9WsG9ZwWNA09/qpaTyIL04g84isXXOjU
r6nj5VN06uw4T2+6EGlPNzg0tdXAxMUYqzKNsprZVfTRp9xgf8SaR7/eypsg726hptf2dNmHSrbZ
RRlJDC06wvfhY8z2Ol+HhR+ivCAxfImInNzPqf7tQICXCTpqcsLWSBTqPpw70WZGhFQqaT5phuRI
YZKLA45G/q7KZS8VMtk8s02r+vrCQa6vGflGk8F6yeMk2P03X4jR9PWeNrSbIyZTUVLuy+5jJ8CL
dI6oFFVSrrgOzcHhbzL/2/vqjdpL82RgMn6ZiPU9peh0CfhJjqbepJ5/yDXwHNDXIWFVTJGmXBQC
BfO6Rks60/gXbs7uVMk1HRMnmzsRtjA1HoVp3T7N/171/eOh1MvWES+krd719/cZtRPBkBBer0jd
Q7fNE1QWRJgV2zrGU+YvvttHxh6tReGCMJjhAroaOTaEPAjeXLMOL1dtUMYmJduWCWCqDXHwFII8
BpBfcnauYvRujzFpnx2nkkwhC2RSk8/t/GX+l5Zp7WbKB4xchloqYxXUg63QiLPKLgPcvZyNbvF7
b6pEA+sZXLahUH1fJpGN5mexM3fDr+PnolC4M2bCiMgcqRkajDNuZBmNRyGsZAKVVJj9gYxa5nH/
0hfzzLzlsg6QBL0UAKwJwl7ma3sOv6r3TzJwHAoyyQTGTFmcwpXuTxzyuxYw64r35bCi5fW/ccxP
riQU7OHSh3hkVoDF2cEJlHY0E04HTDZ/RYi14oO36yoaG2sdY3oHu6pjxZIEseN/a3joC+lndqns
/z0zB1QASByWpZMi2KHDXJpY3MayMci6GzZQPV77ySsFfWxCdvr0fw6WVJCks2g7tCDUa9HU3YVE
pHc9V15EMYMUKKZFNcOF7xzfUvQ2xv0Ac3SAizU81Xcl/ZvoIPkEQ2RxK9FfoV74E1rvXOqS/Hdd
c4wF6EsW7tr2QxEutMdXeEp8B3PEe0/rra2RTtldjYLXdf5LL6fGdTltLn38+NE7M6/LOMWAmQ60
X3bPvF5AaFfz0En3s8h8D7axR/jUjp/J4CeX8nCclUv/oopCfdQ/vJjMaNYb3Cw8Zd9M5gbt9/pO
Zs/8LWuzw+IwcJpYjI/cPBnhdRaxXMxGNWQ0aOd/XtlJk3142xkKpyGgFVc4CpGblbLLZD+cTTIE
oXr+1diU0YN/y06lALZsU/L3b5qqiKBTVZjzKtD99uhLiVFHWklDVpjbUmprn5HxKhV4O2sXjVw6
RH+4XKEl3RkW6hi6CMD7rWshnOtbh/ATsqjAVoTJanvkuglswsXz5od/1gqPWp3vJs9gBzTrz1Qj
lr/iGxfk05GjifgfL3q02PYErBGRBUwWr1zHC8BCRUsKoSiqVZbezSvRYUqcB1ickfJqHysHqF9U
EhWcnbQBbIYEfdmwspb0gX4d/kDPyszyHdzUtfsb2pahCJMpvTFdBeP4Bgvh+F3A6A8dMvSkk2sI
/Mh4Cpqmu/UfBJ8E1hVTqr8fP9kTVPu//s8IooPgB08QYC9+Q9E+bUa4XeL6X9qJmpCNIQKNkxJU
xQwwD1DBpkUnLwiESVxwPkWNJXUDs21lKkitMwbnrLSMUngzyxsJeqJS20JkVZXK4yc+C6sBMl3H
NzEo+TS7w7vXQyNONm32rBOTW+wckUCly6xDd3x2QOIE2f9pRe+THTLQSkCsPpH8mMJ3jg8pByPB
aAsEuXsXyb4/3RZvvgyIhReoxxrK8ypN+796L34J77MQm/MijkL7vmGexbTT4PBrnu7TETwz7+kL
kkN2/3saTjfsOqqNREybyZSdLfRJ65qCyYmOrbr6hY8L8IFlwc+2jfgeFHgK7/5vtKT3jhHnb9Im
cKCu2WyiLmn6rfkdiHISyMvDc2NWFhaXW9LdLbDjVL38J8MKDvu/vkpMopjqBVX7CYXtlHfk0O60
Zsd+tEQpLr4RO+C4IslWxlamJfyy9/5OjbIOIbBwugvAhZgQ1qQ9hv5PQQ5d6XLsc1Jcl02BPSWx
JVi+s6CO0m1xcGHhE0NiIJc0GhZ75xatp9HGZMn8OV6Kw8IoAzq3EZVtbMGCv1CRl3GxIX33RdtK
sdLN2EvPKXvL1CWhd9N3JOTmqLVwvg7anNMoF75K5Iv3ztXzJZOtFLmof9a/3br8aTC5+m3JwGyp
3Rydqv1YKmyflQGr23ksoWLk1flWJumlT8J25whCg8WtOzfnhObfuPhAidsTzVcm9qPofpHUkL+W
myft+Vu4flUz0OAVaeAx+T3eQc6M+/NO3GtFxwIX8wsMyv51CgaBI8d6/lnpCaOW//9OeOK5X1VR
/1obzcglKgiy/uHiG7Ez8K2BRcqLTH+7Q2QT3/JDSyHzXROGuVoP80sYcgf7Qbi1J9KPB5mXBb/R
5S23XAzMqhbekG648BObyOrUlZcpxLpvh7lMW+O5YPfimDpS2bmfwsatJ0dhnromcZS+kt0u0Lqi
4lBiaC34h1X31IbduiMeNDB9XN90HVCjRrTZsFCpyOVEo3H0IkOOBWh8MSPm7Wckpor3jwTXP/5J
cqHro5z0mpD5GDFniEJU+zo6+VjOxtB9Uco542gg1hh6XxC53rQTRDyL0xJkGOvlmB2tTsiwhax8
jgJOsRPKknAVbnvNBmMrPz+iNNc2BIPYbiU7TGueKa4LZsBJzRL7s4YCmFiiokeANdUh6NftHuES
LROtvuSZk7FYjiqULBZ+bSWexjnht4vrF9VatjaSglRZB7WWiYcT39rrHI+9KrdA84X3aAcr0S+l
2XtUq6bkjcv0tT9pYCVA1D5NyHIDRasHHSK2iPr4uT2U6uNwX6bXgXyWszraG0gRKiR1Pw7b5ZSP
6TmLr/foqHkfpywXe3/BpYfkwYcwWJuAkXcLyq5PD76FhBUifFvd2IJyEd6sYlsAc6qeQj9Sml+o
IfhylvcMZ401xaeu3aHb5rtqTe+Aqku3bF2Z2UwjwgfPu3ZynQfMFV5G5AlEcyfTpURGZCPsIkJy
MNXdoT+qcSj8z/0dr7QLrwJSwQPr6Em1YLxc1rKMSYaewPogxLXFoCAAViWtBNl/1+vgzOCuoCpJ
SYO4FxEvnjZ6dktOmtkAPYUyhEEohxoEESK3j4c81MtGMxFmnDnOvqucPh7LjfsVq8t3HfD4zsIb
wBLM10i13KU/5xHwRVdiaacbDGko1O7RLpJTgwUdAuS+Nq4p8yMqsDupuSCmDtVOavpehezYoahP
Xh5JhHqHokvYkZtROvY4M6zHZslraK2fAwoGgKCD2eSoLvoN8N4QOZ+/jg2u7a1L9tE0FMRO22wC
nRHX2MyQGz3aDYn/pA9Pjydh7UFDiF7wNQIH8A9KsEQJWH35zAqY+8dQerWwAA98Chn/kpVss9zo
9PW5gcvOH9CW43EOLoMNrU6jxs999ts5xJiI9Nu5LUio/vZsLrpy6qVNyF/Cw/+Zxiug3yWckGli
XkUUaxWvbRojyUZGYh+zzebgLl94pJXBkMcWRaikYdIgKWXs1ayv7SL/eWtGuCW8UgoovjdFWWlT
nppVZkT1ZN1HO3l7PyWnNd+TjLzy7Afh8iYYdchmjuF2dFT5M3/CBMQ9/XNoAOeetWHqxVr0SEEA
LGRJzufUeela1TWl16xQG/ExFES5bFCZla4dJSh91nfvptu1KS1UJIE94pLl9TgOTyEnxCuiHCX2
1w0LHco6Jf0g2nx2GMV3VXxa9PrIA0PbcI/IytTabfzba55ci2ReAUjYDeyqUoGWxYX14Sul1kfG
ZO4NhPJp9yULekaU4ZNHOWn8A7HnsDQA0EVGgRdFRR8oK2XLHSdpEZgNZ68hwRZSjoXinMKBwYjK
WyHf8rsHfeN5RwR7wcYeiBlCpU4JLsRFJVYFppuQqocUcoau5z29Dv+eusV4q6OfATwehwsCnMFw
9FDyc7N3w5TLk8+1v2q9T4Vo7AeYQB24JR8YA3jGkYrPyGKvfRtngBeyOeokz9L1zHj9eUMkXy+v
oAnfS+213pG1CgSJCi0FggfzI4RYQNEQhQi6snwQhiWg7AiiNbPSLP0KnGEC4eToXjlkiXEhq8EQ
du9gpsPdlFan+mo/aGHaS6KxZaPU7FZv9sgIDQzxoKAOtdx0JS0cErTZUenD13z1AmV8EA43gP/O
81HyvjjJ4+9QdTfMZTzFDyprU1FcJp6brbR+0ZHcbmMBFbDmaQxyWLReWRTLp3IlL9kewJwWxPqX
sK6caLBc4nlDhcD9yrJq2q8REKtY8DDW94cg88m4lSQeOqPggrC7xaR2QcttuL1CYBt+l6hLr3MZ
8dwaedHgBW3E+XIu+5koykxy2JuD62nv1Xqy5uKxVKrY9JYSa1GkpC6v3WS7cQqdSHHXQbGKSrnw
w5q9nhqmmvLoQxr+LXsxYVv4HlgbQqLBClXKcJg6d7PhXWWY6MlbeQqUPtc3P72iQ4kv35ZU8T8O
vMTrdJ2sxK67lfzwlm+Ly9mpa4UZ10/ubp7mYe/X7p/zANO2EPJb29babkK4y5WQqpYxiEW07S9r
4OzPQE+eWwlFRvgpmGiRD3IQOUHBqn1pWQHiMHALWjIt+rRS2tPvo0ugg/PeoxLKCYSnsmgUf9Cc
gP4+PzEdimpH1ujZD9qv0vMQU5n8iSc1kF/CA4vaFsoLPnkRsdjNDj8z0YHN/OBW84JrIIjlQUR/
sWVmjdDeg4ZVIb33ooAc5X+OyGW553l2QQMqaRs7ogDeT3xOFyeiE8Xmmq1TyijuQTa4IgikACbd
TEoRMlKtU6dyqoWa5Iq/R6tVuVlb7BtI8qn+FcYAaURhzWPIQr9Dajxz9Nyq6UMBAEKKyHzPRFKF
zSrAHYIbbQfi/Ni3dScp9/JPEKvwHssxpaqH8msl/buRgeqYOKDw3hg9mDboXrZ/GkujpjQaNEB+
mHM4dyFvHKnbfVQBcf6wiFz+4pMnxnITsRzdC9CoatjsDlboNnMVnDilp7ig8QkP01rYmL4H+6fO
jc1FyQe4d7ZVG7/IcoNsQ3HIjOWIFAANtb7R9/pRSNL8niqedKBUQ2HWHcsB1K9mVGsPBFIIk/n0
pRlh4xCx+cmJlrFaWYft6XaP+kkY7ApmDKTs3ReU51EqYfbFlzBDezavzOgxlSYJtJaN/LcYAZOb
S+V+y0zhVf8DtGBcuriWChEgWInNBYAxQU0D4/i1e4JI2NzAXQka7fqtkWGXNF324F+XsAck9xYK
zY7480Tw3tHx3QzxS0C27IOYwhsAnHzG46eSLtZLaz/8/ro3xuU4haQjkLxQKyYeiHgvsj4mwjwV
jYg6k34+KYHjJXtrnA3dTxrQlrvyfgRIPpH9wy3KAdbeIe6NAfXSFqMOCuiMAFQstn/JnTZMQb/T
ieVPJ3uVJbc0Jc6n8lpb7ztLNmfjS3Ta/Tc5S7S23CIK67Iu16FHhiKy1kNA+k9g3Lz7gELD2DQ0
6c7reh6Xzx3N0cK3l/2y4mJJht7VVHmRIREjH1egz8H450gWS0KTR0cPnpc2FDLlRi83AP+9af7E
kMVGiHBTAmN6d/SRw4j6t+0H48hh+uKUnpBcXsl9Qdqz1GDerYCcum7/n/lLJaMY9WcxNn8J06Wn
/oMKSQqt4VtskCXxfD6TJ7lnVZ6uAnB2vbyRM3dw3YhShtBpt7AqiBucDsW5sfUlVCML7U6qKNKt
UNFaagY1SHfPGVvJ5ExE52/1hwX/a/6xmD19mEaQJldt+VGkbpFO+dn2fHITxyxEwN+1wN9AP6FB
UOV7l9OFzvdx/MEX/E166SB4hAJgdlnKA9RL7DaWYiM6ITs4SLe8gAS8yz/BAyf1eZtXJMdR/FgM
o3IhKKxSLRN3uer1hdm0y87FQr6qviI+vnz8sWfIsPkuLt+NLbi6o4XdvjDJ4IOQZqLQqfS/VmrX
2eJJ2Oywqn5LdOkYGVb3SUOMShDaKXxE/8RB266NNvLsTQknb9XLA7PzD02o6+W8kDS0yyDqgMxA
Pq41vuFOOwnrhrglgWAR+hK+qq1C4SP9co2GRfjTtcbtUTwYq5BXW6TTzyFdX8MVg4TAGQ+7vo2T
KpZG6kwZOGIGx6HA5lpccDxoN2XRDqjFSU3BrFNPur254BeSdXZ7rzhU8mqmIQxcP9862inqd1LF
I6UoVyQtbuJO0P2Hn4EO6cZfKlJihFNg9hkzqH6bDdBRO4pO2jSglzg1Pah6cDGnVI8hilq7z1ix
JyvHNDBk/KVDqT2fAt7Fbr7lQyhClkYqrB65jmyXTB46+OlhboJNBVgCtuwmobvRVU6AHJD/xzbz
L8T7lUs96Jf2uEXh73iz9fbfFLxUk8NgIHglH57BsRXGpDNZrG6pFpR3jCUKh5mfHW1ZddPWk9c9
3CB6681+Who1//JyQkMIe/oHEjmZ2qu91mGWDlWR1wI/B4Cq8oy41X7atXHJBggqAAmDyvVF3hzH
H/PxZUeNH4UgAlk4o8ZKHUXAMI7nCMrQpyJ84Z6xid3JsGuiJ5Z1BQR5kGmR8o1yhtmuXwVy9YMR
vi0Hsv7ea3fvM+BDmWW9aKt6QSnxGthnNAY01iPbifG0FVuj2oy06AWYSBYk80JpIb4NQINPcQJN
JmiQSE5EF9YEW46NlGPgmbfv5bHkAzoi5KGkR+vLwU/7Cw56ntQuBPnY6fR/8KCr1PKBXlV81mdn
B6dgFvgrYwtWrodeTQgCnVKTv3F6IMwzWLDZW7VzrkhW2ERchytJrzjWHR7LiZh7KirvrZpZ7BBM
6va/ef2f3evqtC0gscyMHbn354cRyi/emFfVnNXVx6AZoybpnB4HR3hqM3HvwMvmMJ0wBGjsfR9Z
iOM+NtV15YuXP//a0NX/DryWVlqOtR+seGN0Fat+p1Ts7hKo+6NYtbqchIBhB4hGTfhO3ASnVamK
saFWNCJfB/TaIitpSVEmqm9qo7Yb2FqH7h595f8BBVHloh5wCN4OSuRY1Jaf0VF5GQigxP2YvRuA
msOPUNCvh2vC6hx2UoMWVP09j5oy/qnJenftW8c4IRWs9RKUmzEhZVUZXT+PSrnSUe+9EjWOktkc
SB92y4adlzgl23dTmAD874g/NjN1YyIiYWngx3qzSqC+gFe1nvo/OtrjL5IAnSBjKtTfNESKF9OA
IZFZKanghcIg+8EcNRLWLssd8sSvMeAaLEzOiq6RWlSsBOWp97DINV/LzqDZLOKnnQUnHQaVnhio
QnvhhOAGxaMBDEf8VjdHESBYsdq6Niz0+sb4Q38F2wqf6jmojlomzTmmjMTg0K1BzbaGGYLHb4Du
zbDmff8v/samG7xd/dd33SIzUETPrkxiquPtyz8olrCV68kcnPqNuGrLxnxukFmpl6wZ0uh1Q2NA
VzOb+VeOpXUqZ6cddk36eCuEtEDTSX2N8wyS9z2NZuAVz/PEfnPMbCkrO/kAw9VUXuu/YSeGFEWk
Hp9YQannEuag2tKKQVuDxCP6rsJc6LctoK3ztZ3S6qz1fHkEDnNjmslBa1MdywOtF+60Ift6eNDT
Xm9LYECXl2IFlbt3TSR1WMqR4g7xNqHjQQMOn2TAIuakCyrJZr7k3Ipawpj24l9XvOAlb6Zbrre6
GS9zDO2GjFagW+9sgrD0uYz9BvlEb1BNNGGHJli14MD37roHqsFyVGGLbyW1WrXoQmw/cw2Mv6gc
XYdFzmYP8oWi16nwV/HwiTqC3Rb3TTF3J8jAadnQQxdoGJaxIpFH7NhxdioYKHhBhMEtmsTxei0c
pHHcK7XUVIuW9L3lWodZAhvpuXUyaHL7XwQC7jr9frSsnipx7iTTJQ/dVnOytWX6EmO/cwzwekwA
96sDA9sfdWAS7S/idOwJ6ZoiMEmXX4Yi2p7ySr+A9gguplNSod+jT1gzW/RLr1v2zc2Mn+sVEyLP
98ApxVUE3DZ9T4FIJZB+0bh67WqXhfDWLVDWCsvr4KWknj9MEMerawo5WRP7p9y7onNdepz5VS2N
/bRYgGAKsIP0PXt3HAn7M+u/0ZYN76QzNUhVaapU7VeHkqIGldNpnLrqudkP3dq1dvDaCrqXI9xd
PTgzx/hkz4vyKQtWqwDQ+t+0YRrpBEq69nnQMFPkB6MVhyvYWXe+lK464hQUU/Cs8Hy1cKHA6j2j
0dmFjvupdMiE6Yl6XfzDcUhZm7gC6farjXBstFKZYNFVewOhllhGFmN4Pml+qMvBdiETd48U0YnO
LLlPo0WAIxQHgI0D96BK/t/36KL6R+2caPMyMtc2UVKKDf0lZNaQ7Mj2I5rQyAOWJjxrl9/aDD2n
Nf9x6nBcn5wpM8HDbDZeZEHbe5jSsFvmXX3AbD+TSZkxu43v9QK2va1JwXSd4l2z7Gc1/7vx+OqU
MPV8hhW7r+KkbpUXG9KxnkSHFiWsZ4I7eGttOpIWvr6PvcGsv2t9yLAjkcOZZQlEgHXhYp3yfMtL
v5yx+Sggga04hKPqNHRU9EAaSdcvQsCINWrN3vv3lv6LIDLi3Iokcj22AoXXCRrqMFRFeerPHBoV
brAUuFvQ48wHrxrSlE6+l8+YflDmy1eXQ6wBt/saIzx4zYJjG7tLqQBPV8jFbkHH0KcPqfqLcIk7
EL85HT7nGuqzNNMZuiKxZvONmQQU6fslx2og6a3eQ510T4JG21E5giSSRbnety8Y1vdVkseESKi6
FZCnk4qgFx/n5Dr5s3Yp6CaL/a+6/ySG3HuYAgSsghp6VKGp/ILFT07llyod3kLK1hBfWAzKqrVp
oI5kLUUPKk/Mp87qnRmicVtLyhO5BRJdaDZWv2hAM+ALqiWgUZN5UOmnwogaZF3pl7MsaYJ0a57z
65Y3cAgRbp4cB8TppS6gLwkdgY5Yv9ys0nCkyWvkYSzXDo5XCR4dzG0OwA9AZMW+LwuCfQ3Fz5rt
pehTlR/PvHtye3l5AciV2hPKSoGUpuKtdVqKDnye5peyzWNIyzPXmhLLqL19+gqvDfFk0+fMLa2i
dd6kqt5UaIy9PI6lx99QBZBgiukEXxdR04HT3vcMqXb+e2yyqm7aRKpyQhZk0FwVtPmOIxTEcfSz
187NgbicjD3YCYiswtm7Ox/fJoPNPuheJ9oo75MicmI157uyg2KG3xZ4VErq4YQc5+3l7wto7j05
PXha3DLYNi1eS8ri8i8IeRk+qbQ87krJCWJw2MQHUzq5I2W0/xw68LsLOxVv+wslmA39a1SyRuVe
37r57/+Wwb+w7GIoyP0qeCLBu0AWEDb6kCJqL8bueTzraG/oRMsBY9O2vhV/TCiJ3qsyYaiV5yI5
rOA1pJFqO8iDNnu5hs0E5n1AwoBCEtu3vQa/xMHZ+aoyb7omHsosLMASie2mEMjWazg4+GxFL7Z8
Euccf3MqZ3PdKKodYcmSzoyhwNSXT56SdJ+h8gPLScnG6WVvxPw/MiYqvT+3pbcHH5e1WneumgJA
z26YnBb0UE2mYFXQrd9sFdchU7OcniIZU+OdP74FiiD/jv8h2J4GdqDtO3yticBw3rv6ET4c6qHP
n3N/bcuyShhtKcSYjc1VJchUuDP/NTfS3VTnFnqlUjFJrnUPwI34Rx0ih4B18IobUBie9RRz0/mQ
kEWFE/RpGRCw+i2j4VdAixbgyJP/7fCa72e1nGO2eRPAi+a5sSQ/OTvRTSyp+YmVPQEqy6lLZY35
tv/loyrjxarbSE4h19mPG/CpfH8dSkWNk9lLejK7bzRXHwKc9/tnRoBQMzCJv1mNy8bxRzq7QnNG
blp2yIUBg21CPMJYDJOvvnAiixLykyaux9T7thydNRSPoyhGmqoMvyOMKJfEGSNwt5FQ/uUw3tDO
Sc1R6FhYtv4CxLVrsFZC+h8S6NRCanX/fVzViK88hNTat4yB1Jsb4DeHdIAOe7ynbWQr2JpcHhq3
x2L6KJLR8vt/cp1UVUNtUnGnJuprpEEYWHh+SPACIG76XJDRMYqIKmzqS2vzJeenR+cnckV5cJmk
pp25lB1Dzn2ZXrpknDKlfEz+ndAySA1ro3RVrgElmXagVSYbIxt7b2vgUEUQR8VHbmu9dk9734NU
xNC8D6DuW2LTEi1X6nlnDdXU8kiGzF8iiQ+o9kMc+M9cv9n17ZmkPEV99isKBg0Fie96zVs+t00k
HTqBVMcO0mneTnVroyQ/inYRC36RPOUw164avJB08wHh3laAKeRtnKiX9jGcPDzi0zKrRMdDJ+zd
WtebCKLbOkeRjWpTlEjSTRMbOeYQxChnBoyrdBVRfcDuCGe9r+KxTt/wF8aoVVfv6bTTW1xeUMlV
lltxQKwDJTbL5Iqf4tM2uk+j0qQ17ZLZsiJxkpnG12iHYIHeYfADYzid4A3RTpNrIYChlb+AoWrE
9VtCuRmu1mMWKXrOYJFHCrsYrdBWb5bi53ZRBjzqbFyifAh2grLLWryYtRgM0OlPOz+Bl2lpKrUu
/VaTjpiwJkch4WpDijthGrSHkid90SXDb1t1Lp1st2OzvCJpH3lo30HvGcMU9XnKfUPz59hB8lnm
XkywB6Cjg0XZShBDYEdQzDAHEJmHTIeMyQbBUkkuBCUc34l8J/cIwzFo8ICtdYvWplTOxmvUV2k0
JIaScXhhbbUVMIltJNw2pnRW5lUM9WqCFci6y+186GEfVHFWVbBLWm45njrwx3I/8RQXm4Gwcofi
Y8vp3xJJw4b8Nw9ADb2gNvs2lkI4EVttJ7ZOFRdMWzRxH7AxyINfZWn6G2RELu/xUr1WDarBtVEr
SYhOTLa4LlfPsFVANPSxUIwbyJgDb0kIyCM6MVmzeiNfxdgGexwjB59E3ifv5RtLSGvU4SH+3vjC
EDue6K1PqdHfhTv+3H9yxRoCyOVBtSLR/pu2gS2QDW1ahECyhX2safXw3K52VIMzwmPNzNmhIouA
xh9BX9bQt36IUFxhIPUMRSCC7tueaOVM4xKFC29TABtd00FW/C3YHCNXMFgw5nfqmC0pFUgBHVpJ
1hra2agwXkYQigh45eEL1tfJazG02LvhCsEQrkotmiPQX7IUBH5N7Tob21va/XDRscdEYpxa8XgE
vP4//3ZGcwEX1pZNc1uwZ/oEXEEQLgP7VbSphC1PmLcH4TnLq7cq05CMM+ihHzJ5Ufliw5dj2ij8
/y60+QB8AmfFuVV2TSc/zSRpivRsKsyRsWrK9CdPJhVx/4oiZpXf1yl39PryxCTk4BWHOLJPyenu
MM8ojS3Dy/lL5Gbg0QyyzKM/5UpEsWhoE5lkBawSuU2Vk9KidNUMniZztSffZuFbm93uxdu72FmI
0Cdx9loWzKEpnBDOmEzPayr0D42LcFeoduxA9eQeS6+3BSk067Wm67JEHtjAUYQmmhdOy8e3zUJF
3bsFnwkREewZC+ikNbL171g9uc0VkKWovt1RMnc7gAbYvmLZmeZh8Fn7UaKPt4IruKNljIWuGPk2
0r66JCvGYsolSEohzD9C9Kat7Oy2jgDNVJEQeq3rF0g9Q/osw1UpZjCuOEvntjA7ubpIMrAQs2JH
tAYZxx8+LIWxFQ76dZ5r2z/ORl37U7Bf59pY+1NAOvbc4hbJh+vFDWJQ0003nsLZjgLopv04z5NR
XbbhaCLgLxMBy5wiPa/8+y5TZjdxZptNdiipuovs8p+NlZUdJtp+iSz4eehK2dQOf5wO2zsS2LK6
ThI+wVutsIDhZP+OT+5Zw2gwUyv+YnO7jpPqX5ZziaSec8FVbdiKrziSW+8+s6muCec2WaStgb7K
mhpicVXesG6Omp1HRWReFAT9q3re8vtPfBIjbM35unZZiw34Nw2F5a8eFj5Nq8kWJ3CbsrKnJtXu
iFJPlP49mVMW9hvXkE/r0gpxQuhmU8gfAlDll3WJcJW71WcLq4DoXAoSJD54UWw4M5lCSv/YQMsP
PU7MsENSxDQ0/Nnr3JI48ZH5cK7fzPZhKSKubmFdlq2GOwM3ApdohIB963/zeaCU5lV4MPYWiKcZ
uqq7T0EdTifRPXHRgULJ430wlYsbY+cF0wC03BpaRHmP1sfkBzFA+XyE9HgI1iRBi4vyHv2V+b8U
1QBUfxynyN5jL1QiPxoYLitv2e7iE80R/qATYd+Ld9u/wLbqwOhcfXCr/YaoTuLeTHviTljpxmB5
qiHTkBBT9UT68nj3GeuZz8Zsb4cjlolcSlXcPqnBOqWL71V5I+cfhftBBUZTJtjggR9SlSkFQQK5
UJnBzA7dzsiG4FOtR4DSJa5sSb62OL0CjiyYMfR17bSEPjM+rouWCAymuaMboppcY4xu6TxiaJ0p
s3Y1Rwi/SdH/K/OB3OtXA3CcVbdbXUzlvw1HsA2+E9ZSN3C7eji/8q46LccNmed9LyVeTPZopN1J
a0ypDNmcp7+jBPXPvOyg8K7z8hsP67SE5B9xJNX7jV3CNcWjJNiX1uRDwht48FnVz+ziwlzk3jop
D5cV0TSdJnQ4hvNlZ8VNsxt4NN83gRUus74ZvCa6SMJQiod1+ft6saFjXkIR7wVmpClcHjut/Khy
kBDF203siEtA2ga5U3n+YrpzC/tg/8U7Q8KRLPYtHuhmcyqSD9R3wVJEHoLdkZtW+TpfA8rema4z
NJ6nh6w2zlLqrdBAVyYxtk6cWMojebHhQU5mUFd+N9CRCiuz/BokHrtWe52ue2/R70PNcyzMy586
vIrJXhBG2DFcXc7CtNUobhVejUOgxVpHTtKWvAMeDmS34zCxXFq++1vraA5Kip42DAZw2h4RiC5b
7XpPInEEYD7NrNkT89Piz6j2aSejhT58hySmBBKCOK1lXlRSbT/pGdWAsCP4cngReRCBneez3Mop
MBQR4IsA5YxKSD23sXjefELc/A1xoW6DT76B9x4Mt/rvaxwzpwCSVYj5nJDB3BXpaGwgZje1Jt3l
qsid1iFQFRBvB+bugTkt/sCiNr3X3XXmPQ5T1usjd551hHK/5uJMAt52aFjeJEoZkE3CLSDBVKYu
IjiINb0r/FPmekY72CtEAMV1BSmtaE3abYzVA+sIshC1MKGtdsOJ7NLZSsgK3flAtqlFuMy7eDdS
l6OeoBGEMeR3ACJSTDMURyPwXS/GJHF+LZEukUHAOA2pGk9b91HMNlmHzDmrx/xcnN/7h8dBHSZF
uVs+jYK2PxxMPJ26Xgd0b8Zuvj5ITHj74zmajgEAznBFTN5FUsejYTqwb1Q7eKWYcZ0GeXq612gO
pHs5i4aEaBiuqSDIYjRRWbZ/heQjfQZfOqOU/rEirG0x4tY2v9ea7n7r86cMSGyloZY0GT4mWHeT
TLkbCe6XZPqWIzZcbRbBchqVTT95piDev5Y2tJUUTctx2juC1hwxj7dk5s8DOcm/T7G/FX6NynXO
QjCXnd6xszrOOWouvo8/QBwetfqLpvCUrwzucbu+KcN7wF/EiUmhF2v3YqLzgvUEDiARUq7lVgoH
t3PqgZe5GYCrG9+xPZ5UYTpOyyeaNlKdwI9H5DhDDrtkMZkeTwPPMAnO1NsXpqG6XxA2xqKyt0K7
Y5oEODpelpuLuU83JO6j+jO4t+lNWmsq1cPnY0WWse99rQXv5ZqUZ8FKreNOxwFacxmC77WSmaFZ
7tzY9Fzfbj3zacn7jYEOcaA33ISasBbCwnWoALl8M83onoQYHyIR4Db7H8lX3ubbpmUppSbYKs55
6P++UbrAsGh6O27abT8c4RGk1NFkI3ikm7u0eK2SoWyQQSJZhICHrUSaOumAsxBcHSAVSHT5A10f
QIZdDWa6YG6TxdqfQJlnXRQmBB1cYAoz9mxKNZFP+gx6VgiXYfdkZj6ZmWrxO8Ait3xUi4mBnvhB
ZuTzjpYcSGhhIzJ2DtbEO5E8fjvGlQcroj3DbwV0Yqbm6pokERpXxlZlOaDx4cMaDWWYoKAzLbxv
snUlmtZYZE9ER5ntsI4D8HOjwH3D27awpK5mTrZrPNIJeRkiP68nV2Ehcn/tgxj/JDyit+o5dk1X
pgEbRX00JvLj1LaafVunkkM71gbob2Fy7jAaWLkKRk7HL4ASwfegEHACNEzq1rQBobKxC/PsykeS
h+EEJpJY4d46Jh2whRnPtifTJbxP/7NKzVtzA1kQwQww6z7ii9dkb9GGEyplgMpqdhNVIjkTR3U6
ee0qNJEQ5+eG5nKO6nWltEEtHuqDzaS3b5soOgrf9iyEJBHkVl009y3PYy/FHChe1RJJUjCLSQiw
SSILdGrEfklIIUjEaZOEZOZNj70a0EJabZgYvmw4Z9aUxiBLSKUYJQ+1hZCKpYLoEUsV4xf3gOuW
cv5jBIYljoDQyjjaQqMtOargvfgAyJUrC5hP9jtJTp9610F5NnG2B1E6FQIZkNqdbdf8nRukui0k
fBLM+Nv/QkefiU0Et//Yf+yF6MwhR65jGa63pLhUmgdPyLVMlFfCW/fGzWEoEPkl9v5YtmaF01U9
DApG29ABnAb05mOgipVpjdgfjSRIKCmZIxKt4SzGvZqW2dqm70OBcldp+fy41hKQEMM9BwLOfOvq
Gq82t7K9Oz3N2ga/5G4qXFYtBpkmXc+hFbS2hfTo3H0TxxItEANOdWUhIwedbYf1U9A6qi3dLuRu
0IkNa8BGd1ZhuYcNaZ3zpejEpJgfplgNzaYwFO/icbBKejobNzB6grIRHUROHSNZmlkCnEClJSec
EBAZNN9O3/bQ1MpUBmrIbOeMTTHrCb8Bu3TrHUwPaHYFyX7ZP6Xb2Xwx7y2bVGBw7D7oGt12b3ia
MFWLU5uYd+m+BalAkOQHydgC8Ri7yug8nUnRsVBUu/yEyU+T1LwUgPajETsIwiRxnclvkBhzlOev
e5rZY7Ww+7D2+BCW+/lpRgzGJJDHUB/Ru3MmbYGAvwBiZYDnJCuhT49oGajXLNvI59idQhMTlbty
4pYYMqueQef+fUTEfo+gio9Y3FZR7TnumQv83iz7qbFH4t4kjFYBqeCC/ubMii+6Csj0r1LQkC4A
Zr7UAYEj9VeeoAnOZzrHIszA4ixefFpknBkyqdlPbkojLi17m2CWtg7NZf+ZBUwrSHGOElA+hnAn
rUlDMo7m2VXgg2rjNSQk/GmQ1Vc2Fb0j73V45pkwwNpMldhUu8d9fTWeYmWhFokosmSNP8p7iy+M
v/6NGBBr7H2d30QfQv0k4esE2biJ/FB8VKK0wOWdj9MULb3uysxdsp5o/zLGMA5RUD3Tsk0W1cZc
2oXUAnjJKod+rVqoRpK/+u4jecWhsds7wAe25RjO/a17i8aU+DWM/ej2U8YwoOHXIL6+69p0Iljt
eCSollZFoD/WrETCmmI48c2M1XAcPawMpq1/aJnvcpisqwvTLqu75TaCZ2H1I5WxsHx+hr2f4anz
LMkUA6WXY4dMidPkXzANq4ZTTYkJPxh/MJ0n3ZsUZLtQAx17qu0bbKgcqDGpnKn0smd069R9WfWN
ADDhK3/DbsS9RSc3rsp6vvFp7ikrX6FG86tVSN3CglmtbotyKNnQkDc49i525K6V5DyyZyNUaYK7
30pd1U9qVMxf895pKvJ1QtjpiZRcEC9v3OZ5e5RnZ/gESBN4+rkq8WUgXXgLQsNiqFzuzPPRHJCC
vUTs7oPrH6AR8mRCgYhkeVOr7iiKwbou2tFf1e7aJExwpsWuTXwLN1u89j1DIzy2BJjwFkFW7c80
j/PUXWe2pKrn0us0i0AIK1puawcAqO9MpAd1fxq1BjD2rfVU6NKbzRV5Qx14OhK18PUmh/V66fJL
qh3zSnmSEH24nTt6K7X2Rziw3wLgFBTdLqCtdVF98muL/rgjn5mYvtWy23MSR9dPeEHH2ZLlVN2B
orb6oLErqS31rpd7/G3Yb+3DZsiVf4CIYnZxEvfGbQJ9G+PjulpvPyV1N3yR4+9xNwmmahSb/S7u
QZL4kipQMbiRYDXgKogJigAaNpI2T8cNi6DaMXl6dTU2oPavhM4G5yaOm5ilxXsrO22SP1KpPElG
myZwLjUNS/jt1CQmfHN2bGcNoSmFN1mtmxK8GJI+99DftvHKQtLxKX8XoXIQ2m8Lu0hSD6O870FH
owvgMnV+cgQZSb0lVGCGFwvOTMnzLq5XF3GjSWAc+oHYr8Cv3P+qESCbFuFOhyMiUnJvMVvtyq2+
yOuIMrKGZRVJkJGWC7TGBQ+KlEdiC1/ld812c8eBjo1O2xcOjO5BrmBt1LVB0vNk0+x0nITaMR67
oiGzoVrp20Biw1zbLu0A1pYyKzmuWHS0p85dh/p4DAUuU4bCk2dziH5r0kPXL423LEz6ic0/tAnK
Xe2qdJPU7Z6oVdOlyBv93nLD2rV0C36/FoitDqZ8ecIcdTc4mX208rPC6gTEIFy6yz62sCnZevOa
M6+RqfaU4uNVnmDe9vrWGq32HbU09HzlQDc522znjac/2c9AKhhWs2MOuCHvwqdS4h6mOCLa+p6/
SkgCc+/t3jOVyN0XJQNJx1JD7yQDPQJdnzUk22zWt9dD+ccLWRoVh2wYHDK1wgMVzkENc6clPW4H
Q5g590LcZASYcvr1tg5jjQU/eQV5rG+j3DFXqqYxZXsZ7tEI3895o1CZ54feUsiROlXo+8bxE3/K
KFPJJnyLm194nX5w+lkCZCiYekMx1O68UV/fUNiYhBT0U1JM0qeTYscOTLyFCnjx6+2IMXlCDuQF
HOP3LbVw0DF4WRhFkXEETkJX4OcEW/Hcu/I3nuEwOw0B7f/yiNbF2sg2vS8FEUZi9/YUjoAtxSCF
XIH0fQ39/8gZ9CNzyRNhBrHMGFu0npzTzKUwoKYuY3C8uGPmn9JKo6Bfr1LXeahIzYP60hYnD38Z
WwrBXw/qD2+YYxyTR/RUEeK803N39NJuL9BZ+Uyqn9zvTe7WdNF7q0wlN1d4hcxt9MeKmsrHLTQY
lzEe8JdupG7rjEv43xQvB3ldh8sn4VMoHtmWDroKJFAem6CTEmhVIqsFzfHPzOhJ8rrlC71M7gNT
HSZpWwLSI7vBC49eyELhzOHajUpo/Oo33aFfAlXx+rhVwN4fXrEo5N8WnstmZthRoR+yBQMPQGTc
fZOmkMvEmQ8RA2MLoytxsYRFgOQ261y9zkoQCeJocfjydOBv8q4TzTDxVfUill8+s3F3eXuoyMx/
3cxCt/z296a0aUz1UeTeJR4efdhbuJxt2lnIrw6AjXn5xktWZ0ap/yiS1+oXR++1xqedFF1xwb1z
7ZWZLd/yz2R4CfV0Z/rB9Rf2zsWiTxRRzF+OlfLjCkN+ATZEtvuVFHfFu701bKfBK6roqGl421IL
G1sx9iI+XPGwV5r7dpISQudl2L+Yv/dvFIwjObK9ifoqkiEzXCzVhv9D+RLefuXKYulQ8GMINH/Y
h/7NJ8Ip221i6LgWWx0e8TRIrnJvr0iDcMksS5m9EfL8svvTrCCDOaBkua98YyE444sIvuj2Wwry
FBsp4o5O9jMwCpxffVcBUZkGucqCWDiJo7/1uLhKWAVJSMvinhgtLsjb9t5D5PYBytfMbx5uX5l/
pcepgU45kFUsUD4ESbsMEkiiDrfTYRxnks4MnUp8OtaXPMVizH9eDm8SZR06UYjPPbUnGg6NDeyR
HczFRmeo0g5JozOwsPlI2hTJy8PeHTQQAxX3zpxBSZHSFbyqCZUl7SkynhUA0uCEFSzf1rBiVgsE
iBQq+yKaeWqn8HPXs/QT/SFmwbBU3YxuzgaouASvmxBAdidaWjkgwuoyDStcdZFOfLYVEWz3j0S0
36v3xbxLzIp6glpYtBetflpwIWu8Y42ND7Cvpn0chmhlTYQPwJlYXKADtUUELP7/VsYpULk4xw+C
WbKETKGlIuNSYnU8s4KSmJxpAsl5lXn42k0IIT4XEduYNJwsHnzGn52m9G1yCTUQoRdmtrXSQwOK
tnLsPaaG2LlhMsT5mJr/tE+gfIgg8B0F6CI3TA9hSrght8hyI/WxOPoQLqTKJB8+s1tMy14TGt5v
TumdzqZflMBhuhZZEp9V2q7UWcePCJzeL8gfsmziQfcTdSJV+7w1xqgHNth9jk8v0XI+aox2fMvH
5Jq5RjazoTMefjOXQI60oDoC74yaSoaBEjx6ucO24SnXIayHiaAh7oKXZIvTBeY0H/+jrCtWVL1h
h5Ph6ae8kABy/D6u9eMeT/j840MyL88YpsF1L9OKNu2+OAODSEhMq5MSTM9v+NjJngFFf1U5roMr
C6F/VeHsGN3O/86D/G78tdRDRc+nYhbkldUqXo6Ud1VES7LM/gwN2zRm9GLuT313ZpbyqLcvHu4p
2Zl4Nz0UsgIzI9pgUmhDfx0ZZz/M2KG7Lq5z+PweRVPbNc0hUKNh44Nj9T0oWk1xLSdeZ0pmOFBe
uc2TcAWWkZS9713Ls9c9NLr3FSlV/qZ1Lar+TcKkXZ3RhzZalv+Ab3tjn8sAEqyO6vmT4xN3wMUd
rIlv5Ak6o5pC8AUayr+I4KChQnPKpyQoDE1ItSvbRuUbc/CQy1N/mXk1GL6I1w7R26xHrk9cwM0J
ielYLOw8Po8e4J/55VeI9QfZjNX3aqRcTGaueHseIxRwZNPXOAhhH6o2BDTVPw18Vo7B3eeluyxF
QAxj6Mk8nqju+vDHN4rhDj0PP3yGZ4F2+Ak3/EUnxpIOK7JjiEmhtiOexbQ1hGYewo0/4+B7CH8y
gHlNlHx/uvgPVydFFQ2HOc6e+uMv2ai+gsdd/i1fbLVwHVZxorFUkXjy1yrW6TUuCYetDD/RDzcG
Yk8UVtfAO0q2YISIhYs/bvTKETXJDCfdZ9eloyJ1oHOWyaVLnazsU2gyMCS2F6uhfZDwhS2WkXFY
kxPfGpIaKunsZZujp7748GyPtW1+vYeJRqfop5TMnez8ZLj+aPzesCtKIM8mgADsQ1MdWRs8aUGc
zwopnLPd0obSouZ5LOpvp+kOh/PNyr9KnzGSOBNiWlNrjj1Gd2Lek6q/Y2fYI6LObpg8MpkbGP/5
fyr68YTVwJ2orGEShMipgeXWj62BW2NXaHXTOFseSNR1oyPWQMXYhrvqlzDo1aG5tPJcjT34zYiB
xemEaaH0y4iLUQMZ+NkIQnUrxLajxhtTg2hSdr9qpgPUcIfgSM2DjiCZtsdM/71GHpiXyVjKoDSV
SzioURnjtnb1DdoCE3xN7rYr7r4ah/JliPfOQcTe9iRbb8Yw4r2mmy9yBHipkqvwKqDMJ4rPHDtG
CUvxeuY9O7L9TuQuDHTQqyHmyjQXkkNvkUrnt29Tr3tlg6tY8Z/xQ4Z0lqybTBHBMGCNhtvBieVa
JRw8qFHROaPfdBf9C+MIm/S5sl/NIOdJemHq23+B4HgIoWu0NeUxyMEoXVkE2UFwIaGymhPPak7+
2GYws5XV/KyFsenx0DwOavWxC2uy4W+Hh8m86HmefIVyS/pxvOqGchTujCM5zusQZgstHRzB6HkP
rOy/oOjLcFFsCYq+l3YHAlKZItHj7E8EXWUE0c4PpDvK7OlZ+roPz+r6mlNF3vEJZLNx6+6EP0Ny
mhcIUbt45SUF0vs9iU/NWVEEMoZNrxVedatDA+EDED5MUIXMoU/oqxh156Fnljw6+Kuzma89wSQ3
36zCeQmLfEn59TqRnL3wmO0rpooD6m/gscZxU44Tvy/EMgN6WVihav+I0qx1r6W/wp+eDXAb/Co2
FSAUKOQ9yGC2WpfZ2GEGlEhjpE3EOTPhTgKLKCi8o6RLHcc0rukWDVKILJQLj8reaalh0JFB6el7
5FraTcXU6q2PnWtwi6IT1r5r/cEKGf/fUPCchG/G48ZGvEKK0fAGcfyhUAfc1XGfgYGQwQFrvNMB
p01whuK2WPa329DHp2qnHn3wOgREBX8dnEJpi8vgOkLkGuRl3Qb8vriHMlxbYMCMXa6+llijusdE
MXTwoSIp+0qmzgAEnNnDoFTh8tYjTHoF8/M11roysV9hQpC7/ynvUvxWZIf4FO/89ok1XIBmCYV0
a4IR8E8ImHY8wMO2Lk0YwwfaJwmGJw+DATPXG3jZaUjFvwpCaEpt/6RFVZT55usTP8nFvfjh20CE
X5perVEoyCGNPLrsLwyzgl/IDGqHLj4v9Jfoy18a3oXF2upucE34FZH355IiqTV0kG9glhW8rHHM
aEANr68uPGOkju5spZ+aTzuzDb1vZpiNclxaPpoxz9bGsutixMzLuh3MaE5BJqrgzqminno7WFts
vbJn3IjfA7RrSfRSHoF0H/WfjKXVDVvfo3xNErrJHLra+xM1J9neeIbQZlQgQyU1hDX4aX4wIYRY
JrWKM2qPU1ZsT7XpszwVCtCQEmxcPWaV8KfiNH1xaUCm+DTrVGAVPI+1dX/rE72d4mST50bt8l5j
jcsxrYF9G+cWB1gGlJnidakyv/TUaqGkAPZgAyK08eAP7LetWIRw6FJYz0kzawnCkEM5DcaiQ0aV
dIJ9kCx2sqiWHErAnEI8g+a3Nu1KlgjofaArRd2GEihfLkrCfnR9ZDBoHkB+5LspgQ8hA/rJserq
xeaA6dxIzJ4RhD/dDZDqkpSPQWZF6UC+VVrEpkAhpum6QU/wYvRVOeEyPuUMbfz+b2DFqEy6p1dc
Q0T+4rjFUycFt3RXBLrmV4rIagg/WxBgETgo/amB6NbxDiyNSQH2zxORntVMmgkJvZHYBdHEqUIu
37IAPAw2So8gPH7u5T7XUA0R9hsB2zn6gLMXt0vyokwI/TppcVk6P+AVSA6DjJHhGZ3uHQemCIPo
keyedhhfHr4N4xnKfcJtOwRtyAYA0kEgS/+0KKipWRwSz1lT58jzIqox/PRXklAoliDX77vvS/Tq
GQFO22bw3Wz+QJcjNkb1aAn0N35Gar73aY5eF9ndi2AcMBF799SFI/OThGbczMB4dlIRRdUP8P29
XdLcGh+Wa+maDthNx9+1ct+psdrif/leO7re6047LDp+qNoypa1BobnsEKDpjQhezw8kf5pDHtID
YX5vNahrgLJI2bkbQmQ1P9875HgarxBmESh+H8SrVOckVwnsCMPzt0s487TsLiio1sQKg71laboP
XzPXgdYSYsdgcGb7d1vnliJJs7XTnliKUGWna9etMgLhqy0++M2I66ZMBocqu0W0i4tmmxHJsaiv
vK+8VJ65O9bocIMNAnpzpHI5zr9/4sGOFWwVaV0X2Iaf8EDLb+0YA1vtDnwqUK4xveIIkAJE+lKP
pxC3BcvqVg/+UUVK7XjFGQJ0EjOlMo5TuUd1fjRN2q78oDnsL3kwfCC6+YGSQ6A1bSA86xb5Se51
/o0FuUOhIHmmEIkTLQgzI0o8ihyuErizLdwHOj7uw4t1yOlKCk/AVCWEAS6tmOENub9NHeEGqQlq
ssucMF4fzuhMhXoIa4IABOJyWoSOsL7qLX3TF6vr0gyhnknwBQDQSFfwQQ3CifYg1pgX4EeVzCQZ
5aDLDPRnFui2mdll2eYnE4S0Vy+MMeZ9m+Tig9fPr4iYiFprAxwBJVP+IBpMERUvgHQ8zu8/+V8U
xkeyvLH9k5ptJWB7FoMHOzIKCM9T2661uQOTx9LAe5Gw24z7wn0uFRx3+4BROqtDgurmKCguHT2T
ipMu0Gy5dQkUruEaWasueZpqO5JvbNBP+0yk6RYpntAxESoquxFLFq2g2yfOfme0iKTdmdDH6Xqc
OOphwxY4dl1jd9s917Zdserf/jKFYV5QqX8sZaLKwWVC/k6aI3ibEzRxHHXWs9steCZAPysiWaCM
AWxgAOPD0lbYLInFgESlW7IdWOoBbGNQPEC1oDBDAsR2rpFxkBllhVU2fssnGIGRO5zDzrYlOFFi
zcmfvCkJqBnHwkwQN+yBKJ9h8QXPm6KxVSA7sy4x1lzxWHkZDGYOh4VjkaAu9zunAgGtuRIGxW7Q
4Jx2e5ePBqNcWBpRz379HFtk23cu9rjj1Tj7E0QdDmBYgbe85VvtQCI5yf3x4ZwjBUaPASBweP29
jeirhHLOitZ8AsjW+pGDMEBvEAksSfuZyMGMGqDHt6BaBvauv6VvUPtv8xulhcCHS4pG+56f7GzI
50mJ/uueQBUTairhkuRODW7y6t+0ErhOPvmDuY08j9oj6aNGFbTq950R7GoRzq0BzKGM1TlBvi1+
5wWP96QO/zx4RaFqu4h83ZolG8p5eX9q5S0rk+MARSf5XaDQu9rIenp4XQvCRRWx63srz0StuGeD
wj0TDJwuTfiIjqv9IlnYDE9iTvBidf5B6kHkGZDQCGnqusUgXZr1FmA2iTtfPJ1XF2jiu/SzASZD
MdOXiLcGTVBXj5Jq2IjmCVviGlnE5wmJlviQHBJY/Sro+kem+bE71j9/VeoelWODFZsV687iTtMJ
e4MF6+oj1h2GGG9V4KlL2mmeqIRGDI/1c4i754v5SUlj86SUV8F6J0LV0fH8mKfx3qcvVXgItUZc
tR8GTxnUmMBDejADuIXsPFoo9oR6PeN4/DaTWTuBMr6Mc81AiRJKPqKymjoZObVXF3SLxWmWABI8
cnnTMTyN2PLug41G7pbE/7JNuFBAa9XYpGY2gjf61XFRmMlbEi9ehHftvmwvEy1ZUMzttfKwG3Td
C10GXnpKyH5kONSWAPIJj/yEZiHs6Cg4cnzHYluBufurh79vDsfWiIq8zv4N+YW/Bu0sjTgd6jhp
oZ9iD2bFCNIfU4VWiftdfYZie2FVuBX5Ytwm14Ij6y7i6NSLY57VqP/jkg0Sb1awHh7fwdpBTiSY
zFsxBvprNFqV+kW1HxIuNeZXS0LTbtHwR+C49nA8bFZ1poepmA71ZDfH053ndDRPhU5CkMN02xyx
oYd8nBBA/shi7lpKMSW61eAWJMNsQxaMw3p1xc5os1lo3WxfjfjbWAK0KZYB16vQsuvqV9P9Kxcg
7MZxiAsvtFzQrr6Cveyq4uCZ//7pHq9MAo0UlJWZC2tgA6O76xVfq0jiQZ9OfMT0x7zzyyDGo/S7
/TtKB1zMXW/PyENPhgpo5JZO3f4gCNHdlJukKLbSgqEC8o1bLSTz9AL3N1JGIC3ipLStKHhSidK1
9WM12wJcfcjfGgcADZi2j/eRvZHbeQg7EA+uJboIaF5t5ouhKgCuom8MMci/XsBCuJX749eQLRTa
6d6JWxmC6Hvwz7/qoPU0lkoadkgbNRkx6JQtop8VY5UbpNZF75EzsYlhp6HPO5joPa4CSPXBXFF2
HtlHloy7LEb+FqbZE7TTe4Cv0ffOPQcPnWa5wDX6uSeg/QPKayn0yor6qrpsIxvBjRJ5uWtR0R15
JLiQI8dogDC6S49OJ9DqN3rSkyDLwO+JPfut/L3wdQJMqnH5Le8f1ClztBTEl46JqxKsyb+DzNR1
0gkBjEkz2CyfLbx87BSuPXA1BsEHQjT7NekBDOZmrGUqbDAK6ODr++mVxVnUeduxeS4jNpWugyPa
EIorpkDJYZUqWge9CAAoq/TaufBkHn8+9Mi3t0Q29t1+OOCdK6/kwmwgbrZsGKfJzekvrao+OVgE
1HASfX6cMZb67AuhAgdsQ+at36FafTf0+StAJtXvAev0KGeEfBKCtFgxOp4yyYXb82Go4COD1pAG
TyYnY/4ODOz6xcSh24HzORqFd1AXUnOwFHxpD7qOw0QzAm34t15ABGdj2IKFpfHio7VpR1b1jtyD
5TZ980hHgI592CZsy9aIp9o4MYnZNu0oaz8bhv98btl+ayfyUA47sjTkEFvP+9t9AQiGLk7h0Loz
RcVjf4SxMMUY0mGYa3guMiYvFWqVCpaPm7UIsGParl6PNauNxWbTBhFiT0f4ZlJ14kMVw1wUEz1N
J+XifhbTk/j3mgvCcfkHaM7SAeb6MLuoNx+ytYpJ4lB0EyLwLBf+T47PIL7+hFhWUdhRKZ9pHJ/3
C3pdwL1cO+VcZ2xAPgstune7KyzX18+GfYGLO8zFmok57B8p90xyKq0qwd9uSNSRVVYXOMA8CSh1
ELwn1J3iP72IcxY5K3i2nhfTQcKufFiwfBDigULmWtyrhQdwOrcajSVVCltNaRSCqYYkYFm1IZzJ
d6jnckPx/S2lGMeWnqDX0KV89LK2blHtjU/IqElXMqI91815/J58GzE1aOUzXrtYdfeDX74O1tVZ
jV9lJNHCw9PWfq3AUPU4T560gpsNoKtZqS2Qdf+O2jA2D8JnK7wmYmNK93S/zb0+fGlgYMPWdSy+
EDCaE6Un45H5zJlY7MdBUsOQlfVQTy6aBTM42RTt916abq+nVbQss4U8Qn1KF1PPXB2aEPLUsDxg
It6YP5Li/WpMWY75YN80t0G8sFoMWvTvEdHmQ2S+VkefPHETYSQZ2qKPpdwGG9cgN9ao3enX63Wy
PYU0+yFP4MVGiMUoIDTAmtvGh+UaTc7j3BBB9ypYdLUbYlfX4UrzwyJ20VZ5wm1Am0D0ERsaoz3X
t57hEp0t1p3P/cAgRMknRCTVtOpM9B6KTbnUQvCdXoNP8LcqOIoqcTJU4AGIveHMHscsim/zCcQ8
DyZLSA1EinB4sFBGB6unUUe5p/xrdcn4HdXYs63R1jaZQSRKeOMdv7AMnVgLzVu3wy2biLBB1+32
Kefy98KpdOjXF5ELcPi/4AXbEhgONzIWxIVpJrv4vIOoXxYZuXMg8vEC6GUgvSozuNW1Zfcrre8Y
eO2JhAhXZMcn5vDIvrwID2Qc0FHB1/xShau31Xclc0/+7Vv4Zf24Jbw6kpvVrqx93RcyF1EADIhQ
KQJjTlvzgt/aSByQV3PJnbdyVHtJV0YBvNa8qURoCiba6+z0g2z+vt0ekQVdwYqil3u7Bds+r9Qh
oJ7exmQYbGxMApGZ/mFOUxougsxfKp1UF8Zp4YdWDzY8q7/gSjDgb2gMHmLvnQlnkJYQC/2OfUxK
EQjmOv/zVuodKGe7RbpFWLksi1UjDVX6QR+dcaAFeEV23MgiUsg+rm/hyYlkQFw5bfXZ8MZQSrCS
eLoG+H27Qgy3ChU7xrgD9iOP1+sizkNefNqrYUvg+6bUJfQm1J9uX7CSz6FjXAFQYH+V9jk1v3AS
8GigHdr3R4Y+8zMBrwrAaz978Hs0NE3OPQGA8iDofEIYfONNMt+/M0f4bJV4JjU/SjRonoqR41Eu
1L8NhpX5ADvFgQHf+qUJiewQQar4ra/6S1Yf8OuYPUM6jV5axMvILJ1bTjcD9B3qA8WluP963Eje
ji5zduly38ulTlMOLJ0+I2bWSo4xkeczZ6nYVkK3xfpeuAjGKDlNmnBDetPBRrLV8u6f2K7rfqrd
2DEueDTu9q1p2FY1EeBUnI5b3vLQ6C5sd9V8JDP685VTJi604cOyZdEwGMZKMUS0xUYa4fJsoHtX
OFPgclYI8nebVzljW0oMi7ctFJjholBYEE6inK/XnsbCQfyWSyKDCGEzY4CYDPgkSkWqhll3ctum
0eG2EbtEYGYIsKwksHijtj9aO5/pZpKqgvjxWyn2qQ3sfUet4BZ7Cg9sRear4UkoT6E+/SohacY4
8jkkcs391w/7UGPJ/jncbI8n3l8ZOgmLO/Ktrpgjfnw2nRFrZjkiIrxLEU9pXL8gwC4gwgzPd6XX
gGUtvORJtl8eoh8GZre3xU0DeMJRGLViORQ9ZyD9fgV/aDe1p8IOxiMMBiiLgX8YiwIeBi53iCCv
B4T5GlV/l+Y2mIKE4xPSdgGtcn1v3q3j09+S4mHasaNeej/DWL9BaLrlIhD9WA1v511/KX2PZ4R1
6qht6uywQLuocUt3iRcXldBUj3O3Ckg2G7AeFF00U4B0MU702IqS8+6tBF2WkQbECPo06vP+aK2E
6FVLGXV3E76wJHjWwQmb8TluGMW+jP00ZIy8hde1xhG0g464ADGieJFPjsmtiUbVhvenGGAn5p+K
UC8+L38JqNeygDgxqqaOj/PL9PcCS6WRRrWa0i4vwl17xqxL6kmNg4EPrdBG4WCVkvB8rLjpF4N8
o8zawVEBNx979YXA5H9by7gS/N391NIr9HrHafI6XgiwPGPAcaLUwoNtafsgDrFjPNY+QPakpnmX
nmdCgw0R17xnCoRD23vjSAowrph5TsHPvBEjq73A1+PoB9zXCfeuxT8/7kWoyUgBvawWOE1teiVg
7ULa77vdhy94Sx4GzGJsuNuiWZF4e5WYDqfZnOt1gRO1X8iPzUxzveUY+fN73hMMV2ylYZevgqa4
8e97S6KTqhbNgMMGsnFVd42nuiCnO7PntQVobRng3U6a/gB8lA8QgrVsfyloJLVSQg6kEp52WdCF
feusw346CQXVkR2Rbwv4WOvbgdwYzfrNFrU2iB15aS1+qTMp/D0Vui5Fyvvb2K5pRBTt0fdfnkt1
yaRTKW3vIvVouEjoXt5kB7pQkbP4dfEDb5yQgs7WhLlgIVRUNPGRzZmL3Pni+RqYRKZMfue38Roq
DEQnapYTy5rTfZxUbHu+6sZYC/2x2psPAOCm3ThhiF1rANNZbuHhGpft3Z5IXlygM5B15QxGjgZg
tRqjLR94CGW6ZDvPXkrealoocyba6eJwjrOEpwIiMDWyamW0BE1LVUVYclXpsgxGeCTKqjD5DtHJ
la4a5qNxjZh8R6VeD2BqKOE0ywHI0am9UoqmBtcGL/0TkZAkRJjNP5o5xmu02Q1i+slooEOjnax4
dXHm0NlKJEP6/Mx0GubKlzifXLSpAUY1S1iSNion9BZ+ZmfaFaGCo56UA1/ag5n2lv9t7toSITl1
UwZAXBiXck1QO0i+FYI9eHEC8ADXa9tdMvVeTqjMhlkqNVq3LX4ntmovuqh9EtUgNj8PbKP1vvPa
0+keDswfdWO+idefn4up80zSqCCU1brSlm/SdnQPz8+71Y9qiN/BPCmEBma03AY0NRUNLuIasTQS
JEkLeahj3YxasZEavYgVMEiQaZ9gkChmiWLHeO8NFZeZkbK3cUQdubsWA22YmPxAI5Jz4NN+ua4d
moLBRq9OacuXFmPWbazwlWdVPm4VOPCMGDUGcVc5IYZ5gryZzRbjZFuxwX3MrvuFzivBgyWT/ujL
bzR4nCfSRrYqbvzg+SGDxnqb3+29vNkpfY4vbC54n0mSUK3fmA/NC0oAbD4fD3zYmFpIdjZZrasg
U2p6elymn1xw6vafefQPM+HDxp1KbAq79OvxzqOfClAatyTfxeNXn1VYacFcgZP8EWNPo7Md5WWH
QaWyXtRmFDghssyDfeh3zdrckqMc6bsdQUTxEGgEnrKFsnDOMaIiOUeFaEOWx21BP0aHF3LobyuD
5ZUFU7MwfJbGX0bxZ3QrfijwkRwqDRoNsaXnGHaCY/sqy9Q8NmxfiLu1tH630wGFH59urakY5Inn
ST6gDSB8iGlqeYWtz6rDjCFAgnecwKsGExv21BV5HR4tvrp+R0xWqJsBpXyvIdZsgvwVvhhqwKj4
z0nnWK+LuZ+7Kn2i5B1OBRK7k/yeitH2QIlQe60ZYdWgbC0ikp9QMSB2Edw2ocuDHroyt9Utne7L
TqlODslB/ry8OZTQykfKvT3CO3UxY9vhRBIO1EREBLxfr3rsw0M7aKeh148q+jhO81Cgmz+pUXAE
4RGDo1Wfa79zvfZhdI0i0CJSPa4hqOo6zMncHsrfzPAkn4IQqxtlX52jcA9WcByTHBNG5QquqT9S
xYVtz1aSx4dWdYWMqxgCewz7Opyg9yS8pRERIaIR2RkxC2uWEwINqx1mYOyeLfoQ+R0utz9fH0i0
9ncROl8QIuVb9VnhlHigtDxwCSAYRdt1D0zMmwfXWbI5zQ+4o/etoaNM+opCHm21nOzH0WApn2Gc
8xxmaifSVxQ9HWun27+s6LepRFSM/Qsl7UhUQt3ReOJHwQmIpSM8o/6I1usCOwNpkF385qMFpkHs
VYFg5y2pArn08yB5P5+hp0d67vF1dRS7v+K2duE/0cVRBERcEWfZNMjEhaYdQ3+MX1JtNRPsSI1h
TwPzfJwdV5okfHvh58JtbBySOY92UrDa+YgjVd0ejEENhJW6lOnek5B640s/CqbclAz6P5shIIpb
+dnMba5T0aM3suDLsjXbQM/4v6l3UM2MzsSTGJI8aX8yyuU31mAHi1moFaK6LREaQcakRim7dBlI
VrEJCyqnrxBkFbxIVLiuPvJaCWtOrh1CnhXxLoXcgrq133fqFfkQe2YoGHyNvKXoOrzZR0e5hY+K
+o8w8oQysa7EdXGEQuIFzAgOHgRgwTHx9lSXtqRbcUJYOQL0CjfYYjNcCeaTmgqpByJ/IThGPXaB
QdGBXjGRWyZhWbcmM3NVLIDmoj94tZsJ9AMofkhjaJetkXifAB6uLBskGKMcaR9x3KX4gAIYDLqE
taCA5frIaIc5eB/tc1ODMBpJ1hBcHC4MymnPDOI5RzgUDuEzgqhY3aZwu6fcP0KsUC+pCXIBbA4Q
jArxMtTWwR642O9HgmlgoSwDpPthCkoG8vvyBCn5fO/B0AamgH8L7zcZRW16fuHMKxEqeHG7J8ND
krM1rtMdwJSTkQP+bEkdlAEFcC3pYsKOuduLHcFlP8SZ6VZXjZXu+DD8KsU94zVoeC27yYNaoqd2
E3/VCCOSNmyWvKyqgNac8L2/zfHTwjk0ExVFeqVVUohgOiWbdEknmdA5poy5MkQhQ2ORCmsV/Q2f
TphaQL0I7c7yLkgoQXGwxpNVA+JlBvZLwz8QhS8NzwJWLBPOkeX/Izr9pValRlsApfYM9RHNBqrt
PdguVp9/JdLVQ7NxhsF7Qg7c3npXg1OLnIoEf8mUfj6VjVEjK+AJIrAW8dHP4VO0Twoz0hdWYgmH
+4e/YutLP0oDxfQCr3bxBu2eg5Ub1B0JFHfmOgWnggTVSMJt1iSjoUGY/ka5EZtbHwzu9RnELjU6
sa+N84n8q7Ixd+CjtshnYtM/LEOpPqXdjzBAppjaP3lr0Mf/6WQpCqaTIjsqZYMMmLuz9dxgfbX4
vR/HOMYzJ8rODK0IAA54IcUZmMdE6ISfVdBLBPjR/WhPgklOEqOH5IekytKtmC17Lr/lxBEsbXDq
KFZXkheSvcrCSaqxJ4jAFiFMYQdfJNDJomyyoXj9Smp6SJ5yaPMUg8UVUEzTQBSMDeMT0RGco6Pa
1vVyZHPS6K1+MIpCKsMyrNd+GRUBsR+tsm8WoDLV6tG/B5Bv5l6f/CniKnP5vZBO/nCOACd7XtVe
9CHzhbBVbqEvmFjQhhlweSsjk+nGdL7oY/xBXOvORT6tuWHCf31MR4D+fnegMDiBW8bArJDQsp9N
pvE+k0ilN5Se3XZOAcz6Zdcddc5ASLAQ5Ga2ABddi4blzU1Qepqf0gyF6vtanHDWHALxn/1fAMSt
rsr25RIcPNkCLouaQIdPSlRNNWRcBy7BGWSIRMo9KyFobMQUUkSEZNmlXK5jRI3CQK13aRw11vvN
aekwKzCWt2gNUdRjfjFOJFkbysnDsCh7EaNqi2G772RtfFCS3O2czDN3UBVKdok9Kb00FlLqupta
NavAB/w1v6ZWRiM+uvHhx5Y5hkrLnEC12HqYiIhzbFkiiAEdQ8uvomdOJZfLJVUJRmflTJvDvBkf
058UbikqdUdsbu4rBLS8OsEblBrjIp5LENQGEy55L/JI5iFyCVeLAUKZYtHE+zYGK8+JBjTR5LmA
JzhAnJL8diaR/wQ97fmcW3lje0C9B1LJG8QQP+77dvW+ZrzgoYvcDtccbpcb5qnUp09airb+UxI4
e4sMmMS28oAj2SizuNrLUjLvMD28K48eS5QAJkhsDwMlCrsM4nQpxKdz3heCuPG0wJn7N6aeAXIC
M5RO4UyvRPVGYUgwvplg1Mxq2qVHRwRa5+TauSnd5YouoG9xsRvk1s5/bYB3LUoCHRGFz5/vzk43
7uc7XzfCKiXx3fR4SuDHJAo21EpjRyIReFTPEjT6eVntZlqSVmDilRJkCm+QE1cIaVgISMjsbLmB
E5r9UBfzUtCul9c/DAym6MoqqBKf5H0PhyHnUwMyYEr+r64NdzHItfFH+9bwv9jmsnNk8/M99579
pcRKhQ0qNWexvRcJJQz45La0v24izZejqkWgJ3bSJtastG4sM5WkEXGHDXY011fYNLUrvUFnaWVx
wzyFrK6lKPJ3Qz3ww7xSkDBRO2X9P6d97AzkEEzaikYWN/9jAHYZjCi9UYpGMGrzj/qEmmD8u35U
ecZ0d8HU4oK+HISAPEXExEWyiXDh+ZId/VRu4keabBAXLCIrFrQ49BUiaAz8KxY4DR61hl9yESBk
npeJjW7/5YAkWxQAUC2VUybO4qaD/myel4XJQkM6tUIxvfmCB20A6n7CIHdod5edbWF/kK9KdkID
lpENoFHWSwpiGboPJQkY/2lrdn5gL3HoGh4/fLWo9zE7JvI2iKwtRTIW9Deea1eMK6QcTTFKi3sW
Sk9p73nRA543vmlnZA6Kj+VybN5zu5Y1HC61zXT2nqV/3lqELZrViLiWQEFs6LAWG7ZlSGUhIx9d
xtRaHcimNQNjndBYjtgXcowbh2gL86BKimPkCQ/ENcYuiSTgfldmIsQKV0+/Yko5LH32R4bKqDY3
kTM6Az17sQj1rYHAVsxBVb+JCIDzTQhJRL4AOR2NYmccS9vPL1j+rk0ufvVSSYWJiS3qVXoiTBoV
0bU4bERpu+pEGVFenQZo504rcl4owfcXHg+Mo+7Z7FNUkPuW06F4EgYy3HUhKWxEWrnVEdxS6bVJ
9vG9AiqqaytvI/vjaWqH3yQUv25gZWgwdqksrSGKmZq4pP7lsZTmIkutLRKQ8zsNy3eHUgyn8bNf
9qV8wImdC+D9k2qySLOz+aJaIwplB5u/19TEXpZfSo3wcCTZThVVRUqaGcdeLPi8DzTpxZHDFzd2
Ciln3PraKi0meoad6nvdL01NEARuywK2CeVy9q10pgtz+9/83XpaBV0NnB7l6JfOa5x7BQfEhtUO
py+GTpnuM0x80l7BzRNC6wvFetDBn+YcYqIn09L80KccqEDghG6U8cgRT1s7N5O4oCiVTZEA6fIR
WwnNOrtzmuBqQQU8GY0bypph5zs7H9yAQc6gJVX/lLovc27aGFZcZmDhRpbhY4Sw98TmH6yqrS5t
Qd76sv3JWiDEPKAF1AcPxU2JIX1Te5gnnCVc1DKJcABwxN6/9YaLR4zrrXLDXBBHz7AtRwCulrzY
nM6cdNEB5YwbboInm6i90zbE4L463ylDqI8QZCgCemJMNt8+qWeesLMME/FjpCuHVho0XwpaV7YM
pRj8cDzfe94BM3eXQQXwfgOy6RQVp4OHMhualcnjexgugylSHPt1QiorkQGk6lQeU3/y8jEeuHM1
QJCLeTAqdC7/G6NpF0gu4y1VtE/YYnQrGMZdN95RESCL/QSDBryWI62e/z1OqXQW+4JaIukn+nfo
tYO8lGGW5QPTJTFGfRbTR4d6U6HccEqVo0BU3h5hJ4zmsnfakQ8mG/4xp2NBh4b564CJSWLSCFLz
rX6387WP9Mg0tfAONQJ15MoJ6/zWZpoK5ImB0x4F5UfOrFcGLO0d2g1A++eR1nEewgPrFePMvKRm
woLjUUcHyb9GQcC58XExmGVcerDglDOAvmeJSf4OJn84WM7yxx1hofxWHoUmoBJ7IjWlSTdmFTnV
LVejIcnvUJMXfFhOHrL70cgRnI2KNZLKe7UypByhxOa93VS/DSV1lVpHElWJ+t+noL/EjO7iHhOm
+IIKASfqvG24dfY59+XY14+hg2ONz/cxS24Zm3sQICI7e+p1+LBR+LqWSWQdpycWN3cCmOXdu/sC
ac7Heqza0ntm5bkq43yyHGR56brwuZW2WsgJ+1u1C1xwjqJbhE/lpePdLCF6zW1Yxl8bC8+QpcjB
gj9QpfMTIRZ5iFudXYEYAImNsRc6ZueZsWxZIqvmhfvo8mr7fyPtyiDNYuCZ+Z63kf77jqRF9Yp1
/LHleyjYRboM9ETSrN0A60WSXw9cPvgvN7AXljh0c8ji1Wu2MKL5i98zhFfQ6lyCnyKTGjBCqWL1
Rr5+Y2OHuPHuBEhl6whRhku1j1cEsYGrT9ArVi8Rwcg/l13D2b97IfRynEJRkO3Vf3DRz978Z+Me
PsIEM2UqilCKEbLTQzmlYDDZR9/79JtZJr8dY7o1UFxw/fWeAX522VUeNHVjTbBtd+0VVxt/d4xW
F2x9C9rKvQsI9o3fI5tAOld9oxPTp4oi1m94f5mfEPinj0GO17PHMQM55md89b0tDwSVO/ydAUfO
RYrDtv5wc4jplyHRfHIqc/EZf6GuLu2UUt7G0nGJaDqQ1AclvJYei/smXFS5V1N5itk4k23HVwyL
/+YgDTBGbMDbEnuYTtD/QQDoWYkLNUUA4N6C4Nxa1twN8BNIF309zv7PsB3Rt6n+OQmIvVTvDBUK
OT28DSlNQE3Z0KbcqEU8Zj7TB8uzJGasxGQng4Ai33T2bJeJwjgzj+bRLkEe2tq5+LUXNkXHUy0E
rhozT005TgfNYB4sAIw2n/VksTlQw258OoLCFKqqK3pB7aT7XKFF5+HdgIyJxza8cntT96RO9E0T
u0JMQ5BeQ9h/s3Wn/8yMFesVZr/0aJqcKZkmW9gIj6iQGb4jwfgPBoIOI2vCd4aVpmM4NDFbWAN1
vS1DZmWVR6UXOlqzV359Hor99pf/puPltVtf21SMm5Y7WldluweGT4Zdzd9oC75Du4vca1P+VR+4
b8gexMJhBN3EvzNOqLVbkCEJFaqImQNlPVAwDmj8uN5Z2RycXshf+QrL+Oa1kRs4L2RwLvlOGIsL
4yuC7Z4SEQmlGk6ku0rIWohT0IV+i0i/EYYnu3rNvidUHQCQyEc6DwclutNvVij8VXqKv6O1i/l6
RUrmZwm1y91FWAYGZccPLR6wO/j1vlhVFLmG8Iw5z6oBlzNzyOhT2qELfqw/1dRdAlEioryom97k
i9oNSGAPte7sowCGTgF0Ckqgzr6SRvg4lhltICd3ssH5HzFa8c1RkNlIwMoQNnz6qWP4MscxQwCk
Nyq4kB5xDB92Blrj66DzNNs0+6LElpMfwjtPi22+iVUKTVKC4V8SJ4j5AO+F9oIeq7hKi8a3dVib
3IV6//eJLHK8nmBaKt899HKOVHGFhGka8bNllBdJvNhKCkn7okLD8jw1eJ12i/K7OV7muUG4bx6p
ktK77ZyaAIWkZV0mLAxyFhcK4CJpU2n4CkiGoCfei3RIG4IlKxcaahFJs4LVL13VNN5100nZ0PJH
XdqhY4nWgDx2YqabC9UEfROX+iz99/5WLYK7MuGclVUybak7F8msMHTpK/kNeSBqUy+2y+91dgjc
uDoyTRncxsHA0xZ8/38Jz2QDoW//J6PRwcz+lmTsm2WEOBZg5qPJyqrKXoDkpQajfoap+I/x6ulu
pGxfzwMcQuUT5zIt7LTzafrIbiP+CWWXCdFCFGvfCrTVpWvxoK8godTTejPj/MRBUaxT7Aei6+Ns
B8w0AQ7fIdPFFuwfnGJkbGBqmRzJsuBO6eicpKNh2QfRLmfJe0JWUmoeFqtbZT9lSkLc08mFrfgO
1aE9DHtD3yB+gC1HhH7b+B6ztnFVYVo+mXvRzHiIuufEaczY4mC3LlU6hckr+eBeLbhKWmC0HCqt
UTMo/2XfvxczfZrzuZNmA8+bsjrukQnqy9X9jL3/u99ntAv+ZvZ/z5Mvl3eXByqHz8DCwcv62bXc
8Ub5PxhN5Tsj74huoaRCXkNGAZebmWiwcXGa1cknGvixHq/zPFMfmkozdJV+A8nWdZYoXxGuKvWf
wiYVrEMUPNbKhOE0CNKaJuWAILReSEnkmntB721lK5FSIt+LyyJ5uou9XhMVlgsbK60Ot/HQHT/6
TxG0yInLRkM2/AYmwzw8fmI1DylJF1D3muYrLkghwFec/5mRTZuQTnuMoVwsdA3D50G5oha5gp/l
pKiUzbxs/jfN8tV+ar5zsefr/pXQt6EBGKmaP142ep8wZH9IFtzUFyocwHrlnkSqc25iZpjIajKr
bv/6uaCrJxrv2mqwDjcEaS6xRvk048Al2lyf++poRWOd3QDsBfyR7IBGgszXoiIrBgYQ9hz+jwMW
Yc2le30frWVVAxTwCcwYBfTxbrWxcAmbEFEhu21mkeMA2mqgyI+Q11qPEvLF8qXblZx7HQCmmTMu
knU8Inb5Ewqb+sQS91In5s1sqhO0YoL5VFwSVaupNjGid6zV+r+1kNdv8DR0acKHa6oEoui53Tly
ADpy8uUV2O7oHwQ7dwYfcjQl1b7alF+6SFbHyIz0F/5mofH1bF35Vz9RQEy6i1k8dm7MIRMvG5JU
ywFS951YdZygiJZlljVg0aUHl8x/20CABQoPcvC5hJON9wy2Y647Qc0Lk4zjJ6SlW9HAAhte7gsN
4xsfSvnBai6qvi7PRbsqogiYxJDsdyONYgM1ztrwdzAJhWAtMIBSBO48N8QOeUEa0LEVcnW7mzeH
GwSNGcML57r+fBtvrEow4lnhe4Se5N822/1bIJ1M1p7QXS5+nORWhR0BZr+rTCEXHGyHguGelVl1
sMbkRDBPjcjPyUPZDNyT/HRpkFsWMp1gJ6OLzbXZXzzr/UcIGriibZ7XmxSrNdSlLxlGXHvZsbdo
bhtr4YqNxL6k+1idKDEygVZ85x/dGhw+BwBtXCSRfhY6d/kpcTj+U+aso+1m0+Pz5grGriSlUhIQ
jy8rZ3PUdIR962zCZy304GsRk/DVIibLGoSsgzmBDoFlonYf413hCC7Um8f3YP73jmQAypeCcaYn
zShB9Cl9rbjo1tB/zPSrEaozA6p10h50ojlUk9YrZCZWEC45VSB1SWPR7rX60goxnhd4appRv8zr
+07wTVaMGfTPrg1J37ryks+dIipHjI5VFsp+WNedhgDvhLW2oTdQggzAP8dahd/T+02FdgvQ63Sd
zaQqWWQsaC51G/aaPN4OZhHXQv2tJ3usBTNaFbsEZIWltFlhwPQw0WmjAQjcvMOxwu5HJHQGrE+F
4LtVPduKHUnebwYcLNgENSRb8tNS/M+82Lw4vlrwJmGsergej72mkuakCvBZ5vuRTcf5gz/pSUAp
cKcig8KbVWjFskuMNM7oyA6vMvU5Q38rtlWb3yN/Y+kA5PJB2FdMV+FhH9Cn0LIgPXuTeWxtPIMn
PaSKpduZt3fTUXRf9ypwnNql1ow2dTCStnVx8yYNiixBlliBzegRLsKOZn/Bhj24hK7sUpvM5Z4D
kR4Awtw0PXHpVh3TbpDi0MnE0qdtqGU+4Ss4pvYDSVKxVP6Cun0u1x8xnkB0C6l0iXBhKQgN8GLC
F2znw7kWQ0f10CmRKPhILrlLMpC3awqRxs8BwAq85yr6E1FiWn+t4uWeu0iD9Yn2Gwmb+vXoAL6h
AK4tbKCB8wODsyTkkNjFHGZ4+rXX+jTXOWdgh2hWyPDmemOczIFfcnYqa70zJZT5JHLd6ySLZM9/
E5yLgV+rQfGDaPRSFejKW5+drSNQTkVJ1v142PH/B3VXs6v5taBs+Uwzel+xcyFEwkxWizpbg2tV
J104gWM195DRg2BVifCRxyGxMA5kpGlJ/65Sw7So1JRigDWk2Zv+Wkx4cKIzOdGZYNFE5yJvuwmJ
Er0HSI5y8ZvDmJPI4/kKKxMw+xTanG0lXE1f0MOOH1hzgmbS85aQMY+twdDu34QPQELu6fRnH7i1
1yTv6N7bZUw5CWdsHA2PjcPsfACoAfI44yLIV2YuBIzSy/+UcLogkBoD0DNSUzQnY1jT5ApCS3Ey
vt9sYEoBVZSRGljDuF2joo+QX07G2qdQLiKqkruWgOEfz4vJ9fxJnuSgfMRCGaQuEjRW+aCtRcva
UnISwpz3ez8HuvI+SI8nqBj3LCZBrmLjhPEnRnUdR6iD3fhRJHsPcILmlXyJbt2wQlq6XOojAWk1
qVBBPZTkqs9iNbqwKy5m52oAUnwGbD85ry8s0JNTuO3AYhVfJFllmfD9KlIu9sdewyDW97Q7zL0D
QCf9uJHAinFGm+rZ8WTuXRpRsWwWm/EWDn2cNPdz61klS4IpRTIitYSvzcqGUZ24MRAOXmrDc+Cx
gznIOiWUxw5CGAfaXRmowvzHTRWiFx0hYB0qQRp8tUKlzV4OVbi5hMzFoRRSqO3JBAQNy59XA2w3
LHBCH4oTmrw302981QSl36qDtQ58J5yJfn+ffUuaQ4AKHLeAtbVceRUqWhO15h94PbPtTN6ItFFj
bYIk9Oal4LzFu6TFJfv35VEwYE0zFbdhPV5DN5892KTtFTfOIn8anAdxbNB7TT0h/yN6tBi6JlVW
uxSMdTVcIJ9tcsYiNtEXUUx75FnVq+M4GBHKQVgwEguo+7CuXQ739SM2Zq9z/2zbxW45Jj83OV+U
/mAKCU8yOtxIEHDqQW3yFuPmeJFMuZdZcK3u3CmK1KKm+weH8KaDStpzfv0Z+Xqp908E/xgmLnc5
FNzVOttNSQZeNYq3MfcBmbxSGcp7/XdXXbu2mfaY3Z/Hd6sVgBqwKCejuzr91p3b0GAFhVzKtRF6
N6DCK1GINZtIWRj7bRME796uF2jHZ2YUuKTM7IuMaa7VOkEI785FlChqdGxCH9/MugA0du4jQ0Uw
TsOU4fKvL+pY5648qDoiDoiJeqqgjlUW/EWD9OwJh+AxAbO54l47vmSCqq4C0+jRbv1bj6t+Aogv
vQ682MEhZnc4ae47yhLoFWVkqLJson5zinHm3rNV2T5/D4P4LWmLBzgyIpCtOw/IgcDRG2H4576s
LZLk7hubrEXBaus+YR6EiVFmviPiv2dbq3PW5zS5lz2ECc3UBjK51JvdccfuwzYxfxpIqhLTpDdx
AckopH+dFaFQnHn7D6EMyaD8vADkYIgx0Ll8vjTkJAJyzqvFhTfed5Mdl2lLwL15cfJdi32c+Yhf
LrX1XumbR1IlHQlsOCwrDI5X5D/224+jrYt4bHn4wGvgfPk4JV06fA+6xEYpnNelSl6tPvoFp58C
ZlRex1/NlG3Q6hU0j1r8J8WGc94Q6GRj7Di8Nd0yb/H+4WkQ/bQHKOpLWCMOLZ0TFPVO3H+gwlD6
6HvwXP1/QBje1faq5skDUWho6/VS5aaaDsMfUElAZG9UhSa/bD4ExKak7miP22RQZxv+muFr+heA
7SoBBILYx9AAa3/w0vU1ozUYlbQNpU2HtDrHjgFSlyV+zObifsVdnMO03D0PkiJxow1L76JPAQo2
Do9yar4o3wrbHbMkqcpgJz11iRwfNuMyFDeITjJ7wuBwGCOQvFRlEQKutgJeH9d0JKqdQ+TmKd1H
m+7ST3zYaKRUN8Pvu0E8N7wR7F4mNXIzsIgDIVYxDo4Ogi6gB+SZ6jVj7yS0JGONamUQB5Jl60pS
vHpOMbOGi7fIU9+Gxb9JDg3c14lUeShfmFi0DuuwH/vHPsgpoCZrkHRnRugf2DOGx5Fykum6CZzL
VnqYmJYXoenJkCd9ish9tM5O3e5qx36hs37y07jxW3w4QrkwBqfXIKMKt0fJfYM4Rr89A6SpkLN5
s3WXSYACikh5CcO9cggcCBnSoO1Aw9NiKCNF9RAVbP2znQgYAAlCpWg/Wn0Z0dHPWBIJdFFgfZVs
wyGCIOqAh58us+RDO6w/ZaN2zlDZQQ24/CLEMN0jCqDudY2xak0nwFnUOa9qfgbOt9TtNG6iEG4E
obS6qDS3rj2+UKPG7w4IpIxt5/GST2OYbq5e8SQv4yxW6NO/1wPnqL2e2e8SOCPHkdhPCmL1Hj4U
QVLqMITHaiGq+Jb0Zvsw5UGEEDa9T80Qj25GeTI56Wiqqz6BeSCIvqCwC9hZTWrop0FdRL5H0Gh1
yUwWOWnEZ2YiMgZQveQaLOWPp2Bym+EJRn/G5BR6Ec/oXPd8Ae9Ef4CTEitNJWT4oNfS4M1WvT8y
9vnCXuXC5FFFUmplnGD5fpGc9gWa4oN0lmBXq/AAp33XIUYgNcsgKchpPT7tCPRXvtalEsOdjjvr
m7pXwnc9imPbVIkONBvNd1avOrxTyI8P+j4/FUXtcOV43NOn700nhvg+O3Tm44xLApHDmtoptJC+
X5gyrVfAFKrnDcTS2je7RfpOhfezEyeGBuCuDwW9NH/qGnQ8/ns+qvOGF5DSgwRi7sEk9SHLbc8m
TQzT6iF+IESVg5F73dLTDaTTipEoE4nL59S69+rXOVuEwrykGQVpz8h+IISGwz2nRCsUdW76tBqD
B1v+7Hf9PXVc7q6QaFesMwsAHnZ6fFMvGCnSXjcv6wslnUhxEa8nYeqrsynyh89/7BjVm6njPHCY
FzYzdL5x6yQNzoF5XA9czEawR+8RX0r02Gktf/92qjmmPZZbgnSgedCBD45N9+f4v2/5a2EwWlD4
OU30u6kGpgt9FvT9FvOZD51s+lcT447cLxCQx/E4J6hHnn/Fm8IKDHtWJutkbzaRNKgFOCrDIjmA
IF5wwr4B/uPfqKdsHH1ge7ZEq91b87leC4mz2BV3nVbWeKOTjiChiGdoTYla6fKKJCy+gOvrzjQB
pjj2SLMF2lOEr/FDzK1ED31eVCWpoDASPb9D4sUOpXYzxNHyWzhRhPxt/GeoD5wk7kvnPXBwcgAQ
posrKrqMNwpoHrUT9FW0aaHuK+xx24MjQpuXBfMKLWYW1WfoAR7BjfyZ3dxOIa8VrGJZ88dAJWah
v/TU7NVtCTwFp1mJK1d6fRNGDh6647kcHO5llyZKJefDJ/bhDafxyMA85Q6ZvzccDyRelwXLhbKM
pNjmJvNckwVxHMA5IsWP4p1oHo/G9ycoKLa/sgZys41AqEAhVsbgsTdr3MQt3KQCRcNAggBQr8x0
bmG7m7ZUO1yE5O+hnH7ISe8YKrnPM8wDqGW4XPsQSaB1nBahEI4C7rhs+oWva+aQMG4nZzXZr+jT
AaZhJwIEGLs7xNlcBiYOKMjdQKuOJGttYQdRiDm0mHktI4qKfaUyBiFF70+ZfdazckBqflcne+JR
+znMoAFLgbda1pminXF68XhYnHzkzmy5O7sup468AJjQ/J2mnndngYgsXItEAr6l9AdDp+bF3389
PpfQ1g80cQ2iNKOqMFpEeFjPCdx7w4GtYh0kEBm9h0IUj2cROY/eB2oaNHCkngibGIYmtgUpvLTM
92AloBHTO0gVpPTXyYig9ih4aJmVWwzLYJ9bKsn+VpJR/7j5QfuVZi2FeN0we5XgymeVLAXAQVJU
6lrhv8wSzWKbzXqJp5nV9DH1cUXsbVyGq3VoJvTXpRI2Eq7kaexsbJu+Ab7VtUQhwb6bXSvmB7p4
tsfpfCDNAY2GEjbFgnm7Ti52LB6/HvWJiNLnNonJIOoucpQCkbXX3T/LllM+pLqMpKkSgyZUjere
YqXVkIv9R5rC50R7JEQV+/NnlsfMYdh1hMs50dKwm8ZoZam2wzuLlIjbYnMZ+FAa5HvfjYtZ8TW3
x4swpJAMshLgJ8r+eFEG4BFxomLDbG4HMO+vaVYVPjEdMLwqi2DAXHgC8pic7dR4FzJ5TmTWh3Q0
oPh2Uu8R1TTu6HPEle9yZh0VhUQrLUBQRkiHYVvBz80y9BceDrEtEoIoCwlINCkAxhUUJr/XnYRP
aSWSdYIHpBe8sGUbIq4s1ECNxARwGPWrG1crvlgeyQrz8SRV0i2hChdW0JMq8upMcP6qDFKHr4zZ
HW/Nn7bOhZa84BeMidoboco44ua5YKMx5lNas2qSW4xhF7uT9DuqtbZyJuIupjeARugwC2AUDInL
dykObvC0RVrJMqcDtzrCzu3/cWlYgAnQRn0oZUuFxFNCAR56cCUvSd+qAe9mywzJhB/CPgzVsV2D
zL1GV1ZRBhAOcNc7I4c+f3G7pkjgTKe/6abKq7sF0u9nibpYpAiaAjz+FO9tPNj7noo+v8J+5poo
naOBe7gio8esqA/OU1TKr8PiRUlmNf2W7eaz2rkLYN+ooNrLyqN3vwzri3IUAYio3WAT62b0eaTr
SmUvxxw1LhM9p1ncT9WDPabZt1myBB9Qy4xWQxE7tKColbNghoh97NJ0v7RRGi1H6WfUZAQzCX3K
cahCG3RoU9fHOOK+rVT5LjNwygYu8UQqVoCDkqeVhZM9J5WUcc3X2qNcBgSDtHzE2hWvz6KFEpt0
ii+e7jGE6qeGd4gpXDGlwREdgtez62wQo8ODuGMwyCu+Idj2AaqrwaWp+pPkDA2c122v84hsumSN
h3UA2zhCu60dOi4TBLwA6aPc9cZ+Pbh0JO62q66uYLuwNdzDnZAr6978EPYSE/NMZp60c7ciy1uh
VmOShGO8e910COS78kUf1miHXeF7cGCy5lBH26yraXnZj7fxMLOaPKFbOJ0p/UMvTRUQIPpKUP8T
Yf87qvoMwOY5VZ5MR3WozfSdQg2bY8ssFQUI6jkO5MLERh3i+qYr82m6RV3+3XVZ7eMYkMoPisVb
hmVVXyDNxAh7vqyU1nNXhtLlgb0ZDDhUbN067dN5GflPFghW5d46MLmw3WEj+zS73J2P+2G28Ts2
iz+Zr5d1sGeof1YAF/owU4boqyLSPVeRRMukWw09ZC2Pu5bpGxZqZIEjT68TTKf/yBArfxQp1cRp
1ep57iTDYQgdXZyS8Fv0a4qZfJ/gOYnf2THS0okW5urunw7YXtIWdfgQNYVbAKshQh7eEAOEfP6k
4OuB0XHchxvHKPaL5YPeXq/OCMFI8X6Bo9MGBfHRgKA+VugG3UIVvhDFGMhouE2UKIOXSszzJ+of
zYObQKSSgnsgjthFxNEEgq7IEVDrAnY7NBD5AwrsV8AMIaT8z32z5fMD5tlxzoNFx55KXvIPHZBy
BibfHu0p70YCJmLYB0Tex55O2QOUjgplruzJyEdDN+KKKYoIHlnOB8YxR9lsgDYiZSAzN8/rU3WH
A4kShVBZSvkCW+n51bVO9H0ssnkve/58PvBk7uShO56h9jBsjDeXJ920TgJDpvF8M3c/LGxs4Q5q
w2egBWMojCO30mpvXwu5GLTCdV1w2AOG42iZooADV+k53egNntKVN/Fueh5J6zz9173TaB7Q0PR4
DDyIvz6RR7kTOgftW+l17nLpuV+stbQdpfEjPFmhdlYsIi9lMm9yenVcLO4lAzMM+Cidpuh+zY0w
STKhef163tQGkrTnir6iiCMKy9f3w5AYBs6nZzuPlmhxyuMiRWXeqq/AWPrbGQFmXdAe6RnTWyzN
9SBqlqW52bp47dtJ0/BsAiobe/2XXyA43DwcFZ4HEJw+SXnBlszFAytukARI7NvGI4YSsJkAc6vj
OeDGADlRqvlWja6IvNARgF1j41IkLg+NVPM405U/1emfptEOriToesT0hTqrJhPgVWkzTM1UfH0b
d7uFqx0J4DRUyPE/Ht2W3enxjJSNqGDKwmEE50rMS12R4XI4/Q3Zz9ichpTM4CWagEqT8oW3QCC3
dYL3yV2z9YGsQ0KMb0GWGRVdR2xRp7OXJDZbiLfbtr6zf7NDYW+DQUtBDF8KzGWhsxIqg507nI9R
MLQEp956nvIeg2y7YIQ7oW0ToJdfinHsstTMvJdOib+BhURhhKVI9lb8NRkID0vvI794YUG9z5br
taHMofi5buppyfTZBjeMg90JG18vcCcR6IYHDWYLy05p6A6VS+e/0YlGayRgX1A73gD6N0AQOcVQ
Et5TAd1ABjZKGud9aLJUGCcW/r6QhCEmqtfRF+08vJY7mfDHMx2Y1pZeig4rK8NbsxAno6tSD44c
mqNL317Dn8X4u2seGNzVC1KT1lukkN4qsSSWFDzF0pOV4zoTh9JOkc3NgaVEBHxGOR6SZQmTevqQ
TApWyeF0NOmUu49zyR1wxjgZKsnc0A222Bn2suHpan2rviBn9/vault27cF7WyS/wdWDAv7GDMbq
82jjZ4kiuL8jDm5JZqdNJBzC3axuF5MsmI3VfZ+7bV6yk8ze1Kj6xguchCrSmPkkCiAIBxWCAmjI
jyYipjUZ2imaS7dghjCR5lknREdo/ACJk7oMbs1UTAGptzUbbREnG3yKsvsyXhWyIOqJx+8sqUgf
1Q3SblwbYldWzLEAZ4jyicxzzT+JiwA1yBwKuTm6a1dv1/RCG3FsPM80oLqvRF7zwUtIhKctcTlg
s4YlA7riLTkLJ/vKmGEvdBAuM0R/ATBY+xyh1j8j+4wAsfAaBgcyUJIoE8cu18dl5rvst90vdSZn
YZSwC7Y0fT/tm+0ksgVVfvQvGtVJqfz8j60k/TkyygF8v7LqFDQe3bXpfEw0VTcvYlu/Rp+m2YBn
tJVpmHOWR2+YZr0Ak/OYlOHwx7Nz2jwm7RarjyUROzpmW4LD6viS3tRbEyEjQGHfosu+Ovrqw8HF
CrKfT4AKwnRS0OnBiH4fUQtB0MIyviY7w1fhU7Ku/Uikme1x+vAtSU+HCkBQ09z6ARn86JWFFLpP
InUkrWeY8uF4ulZ5aRMYU0+GjHSlS/yuzOBXOcyrImqILfNwXFHe7c5n7M821ojvBwCmOmTEzD2q
dvH+6MdoOawjTUhWCw7wVX9LLoqVEUC3fxxzZ3FnlzvwIePZHCoLeMUixNnjoS/lEwLGxvxBuRDZ
vmfxtCvZPB46Xse4u2jzVNukuCpMiEjTr/ml6s76fyo/jfLA/GNzYJL7lyOaPWqf90kyzG7F3xxF
L9c7Svd3+zWJFh7FHxlMVfsvMB3+El3r4YsLjFxjWF4znUyJgQ6/4IsVBdK5ra2mcd+anhZxp9A+
PWyq9nhPEBvAknaRsdTHg/+iJQ2CUG5su3IBFCCS6cDFg9FK/RF6O7uW7Z2nwycqu9+YCjVDKOdh
khFBCRcxb+QuVrPxWYM7vfcKZyXHRejQhlB6KmHb2xklONgebY1mHw8Unqt9e1HcEHIKJS//Jvqq
WEPkvRcezG+aJqDVSfLwDby9eYEpkhUFyvxMcUE4kbWRIjG1ghsjCMYnRjna0mfik2uKJJuc59Yh
i0t737dDr8NQ6ylonNo+77hHCF04X33MeGunRQlaYJkwpH/HiD6kHYhufNtQ2gxR1IAk0PeuBYR0
mlgDsz4VAYMjFyZLfxvinhtreUc4VdRj/wWbmKgdf2qll3flNdUmrwpqz2us/m++hGvlD6fJC/Fe
4jY0DhBAb36+XjB2vR5NtatvMTLrdjcVT/sfgyNROKdJbQuttomNOSaQWtE83VpMNAVx9B0wgcw4
dsxc3znr0NZRrRy8lqXlxnnS0DuLYKv5RSRgaLNaSimwUKOQMQtU2784sITfuEHRILs98BVcJMjL
NI8Q6I02DEZn3NX3m7KL/DY3obOXzhWRcGie0c3k0XZV2yVsE+xaDyZy61OwHqU8W9Bi+pTy9+FE
c05bqtpUJ2ZHLe2ZbCcg40TB2+qLt2oBPLmgcg27V4bLyz4wVsS9JfI66Hg3kTZFiY4Zs6+0Vg2H
TA+3ez/MEEFB4p/aGkduuihyAgGAk+pa1Jgw2TPQ6YeuTT+l8YKU0YzdjWTe6BcRz3eSNyc7DNXn
hN/gUt+Ce5UsTo8j3hV5kC9vGPs516SjFmsjfbDuRleL78ao3ywP2RjdNc+vTiCxysaeqW5IVBL+
7BosXZ2N96FAY5Oige1gtlO4HbZuIgkj0rJjVDAsYoMWJ7zhRBc2ixsMeBM7Kdcj9k/vDhVDAAQO
BPqtgYT0QoVP5j/EmFWgDbgqt2dwlbqmvjXpTwL439Q3PMBt1BwLoxEo5pUVimk2Jh35IF4kMi93
/muZwT0eO38dkt/JZrN4TcnBYXMvcO1+wtm4kxAPJb76WMr7L1VVRkF24mJUDAmu35rWMdHLbo/m
sW1tLesLQmz6/w1jX4DwtsZ5wJxO1vnM7IT+G5XOKxo5cmhNe9JKqTlBgiwrL+NgytjKJmLCCt5K
NPGCssa/V0XpO7oq9TWmLBiACJnYP/yUcqYx8OiqGugRAQMw8MbPAhSzbxuWnldDO/w5gx2TtTqJ
eANOaZPHnJbBw2+lqsvu3WLdCahikV7U4IaxkhSoE8QuBRY9JUgFvfQ0bGwoS1xQG2U2uiP3xmfx
kVVwwMxPG0EqmE1TY3LH+7J9U7qpwarTVGOSVjbSEXcciCWdHYZNujD3gugXl6mTXWhYz4BKeMME
EZvTdsUEID/8lULqrxZp2A889ZCubeM1nk0KHud/aSfADqL+EJB3vWLjT5LGq2cEMiMXffrUltDX
Z3KIVOqoWz/Nd/s8AqydN2H5k9lP8vzAHILj242S6IjZ24TL0FxY4txqKZKtsivUM6zmbp9w88+1
8/KdZlk2juWMOuKYh0W5Oc7QCLBjYlvpV50hpsciY99nwcptSLo35QPFLsCVxsm75g9yYlqqmhL1
JjQGdaNoAwUax1bQexgy7TIvmB3uRiwi6ojgiNEvE992Le6bh5o3hpOGNIbAk8P8PtyjgR1BpAX1
RFvx4qPrXJpod4SiCRdrpZC5yjs77ZmKQc54+6MgHvWJcQmCsUEq9VbsLwAQie5U69u8j4FrEvkb
PatoGlgKxmdtBDTUWKorlNLSUT6Tk4M+LOogvUypl5Phrl95/12jfd0b+4BRMimPHZpVnG2a5FSd
1grpv9DR7n+Aa1ei1BBLRlNxNw7E9NbIW/BWNKLwjlFzSYzhxLjk5HbKMp6OiCLE/2oUDE9eB/7W
nv1s1PvvOqW0xcgi9jaLfysCFjZWxWBzr61mrGWvAjci+Hp6BNNftwdODn4NdIL3KKPAGSHl8h3Q
ENjIY/k+ycZ04zThaIsqMX9zY3vBXvX+roNrmr9RkPyBQCxQ6CmqOPoyOxQJWRy8Gwj/QEGDKEoW
DDRoCWIUvZPpRNYTHgK+hIxuaWEt2sxL2wh1xwDTSVz02GoOawOvS0KtVZL9E4Bq85Yyg6OX717V
/Pp6nG29stGY5+GLTv/XFElqMlVFD7oXByUv2pliPnaGAEgxjf7LY6oeY+LQIdd32/y+bmrLKaXF
js5C+aD3+ydfwMAtVIvBS0rZ6L+Yn+NCPfzfhIO9IOrTLhDVwiy209V1/jlC8tQUqInjJheQrJj3
QhsiyI6n66mufy2Xsk35mb6eTksQKsm8JUs+gM18U2VezvraCCWI3OSK2XrGR5WCcmyD8YZmAYSl
xwmMWydacDoDlUXI8vUpRmBk39DuhkroR7i+UJZtkiotAwWsurb34X4C6cut9Qe/chnfJvxbS5gJ
2aMWOPcNz8GGxvyfE+doUqg6jfqPK3OwqRHDmDZ9MQZllkP+qDlieIdaD3PF7ahU5v4pWJTF3KZW
7PxgYcBPhmCcmIagEZFapbmWpuYbGy2G5K3FIO5BN4uBQ7gpC4wFcE4h/CpziW4w8Hs3a5oerbzm
TLCz91pguOup9XY0ahAYFTL1IuxBJd+7MHjj6HMPW880zWoYLXq7aovYQSEchKEuIkb9w551ILIs
ZOmJnFgy7QuG6eEx/+Si+cFJIoUsd0DuS42uuMV3wQtp3V0FWDPYJJiXy3Yqlr8nz+pG5ajouFyX
FJmQDRbQUgukF4mkM3iK4OXpWvJ8NuvOswPFA3PC+e/FPtNoK3NLqXOM0TSwwv9Ruj7cP6D8W0+a
vYiG3ZN9wyel6VB+qmvIX06Zwfnk2E6JY6dvLV8hLo92DDjk0ex+MG523CuyUdxO3PusbBipI8nr
GafGFS8FCtsCJ4j9OvgcRvbMGlShqaYyOridSffatuLVri3GjWeatPYCjAcBH9N0WDv31digN5bH
gQ1yI4dcy5h5VsYmEag6xIkMtYkBsO2myL9UtJJl7mGwJxtClnPivVPDovZTH2tZuhgWJ7TVHFO7
YKdt6RAXAEvI/evGaW6+tUO3DLz+ZANZU5eO6yVpqweyMfRf1AXpvmhzUsCHXGAvGroMyy3op4hZ
9rKRzF2a+AnIXCrengXjI3lLmDbsSYwWCvqhtR9aeXdi6SMzGbcZaJV7++GmJbdhI3VzB7KhFMa3
f5MZeknx2BToUZU0gwj3yiUnALjBuAxiU7gApXOJ+iDypsfYvpbO8halL5jxJ7IMd9nkbbCuDZtb
H2nq4fGaJMqg3e2xvdfOdSZ2OsyHd/dvFKY13qY2yDEyiB9tLXTlbpvMDs15OgAY/18+YtKliR5f
8eLJ+4l9/A2EXJVRPuw0JaYq0+xIhV/k5kJjcnPDtArWSjncRo/LTp52EmEmL6i7s79QJwzeZP2M
Tjn+hQMCex2Io3/zUwrZvK0ZVYOHxl+9Uc50EaphT8oLJabB2fmp/SUcjoFL2T3RhbF+FtQswVXB
F/0E27yVT9UVotvGbJmyyaBm6XOdnVKzXcCpJa4f39+P3wYrXIoODgAwTWBMfA4fFMAFno7wJma3
SDC4sBi2PgdVa0ZUdf3BL9DdNIvhnm7ZoETY0/2KBfLIzH0gEeVMdjQ5maUg0H8i3YsIsu+E2cGV
VXNrYH0D78bbiMyWRxvCOQkhqt7SQxdSBYE7Z8pLSu+mzPbyuRZcs0V1BVNSLI2nFD6UA1rhn5kG
0Q/v504ZCQd1CnRkP1+tC5v+kcyjReyvr2alDbrRG5vDhjV/ErTRp6cKMR94JLysXFDxaWbxF+Hc
CLOHCbrbh3v7zUUJRXk/V1g/2iNUPoRRi5BxXfuz04nbYFjWcUdYqi5gnRbOuR5nr8/2edcYvcmw
MawJKd7y3GMGaFSqJgeqBJA1kMYaSauTpZh6Y4s0amfXPW2j3tBGuZy0wAS8CvWClQu4qBAsZq5f
naY7NGcI1Kt2XY8dcyjU8DPsf54FJieI3Jaj2t9sBSSDMB16w9hDAeUXemnZVpYqB/h/Z+9NRut9
4I5pCTg7zv4er8/+RhgomJ20qr0nOxe1jU97TIi1GZwOVOI+RBYwebTmamfCxYU3ZWojeotVSV+5
mGxrTd2POIKxVeBr1ywhW39x9VUIqA6SAAinfT+dMAAZLsxZIYW+E0XaGzP9cNASIem7kHhaSTyO
udZx3taJFxbyF11Y3q/inawiF2+q748jTWTUD00W06YhkZy7AidcxOIuXqekV8RTjlxUt+ZDTtwl
s4jKw4IkfMWm+cCJoRBvIXzD1Xsg498azzCcpgd7mgsVZxWIsVuChRdEmBgyQRaIuU97o1aJh5z7
L8XEm7EdflExCbZZ8O8ql14/VNLpRYW1Hx48SH3XwlaYPaOF1my62PqClme5VNpjSzH2eLDm1Yb6
6tn6beZyWARjJJH13W5EvWdJRHSUn6Lh1tl91lx1zKuZ/aMNoxG1eJQFzH44E5E7fnawUq5ShX18
SEuAIwZCsUJy/QrpNhKZbVYkeLZsKuS8ON0aulDiI7sWaqMBzvA7Fzngrl5RHzOPND7YMAAb9hlg
bDp1oNxVfgof0O/jgntE94f6pYCdjjoYC9fZjTpGyNaf/YIFpKRyrwNUIvpOLrHPMuhrgi0FADjz
oFSptbVRYEzJqitlUQ7zU9by2ppLiD0aQQQZBk//zzfg++5bOBWeGLmgcDe0PZ4Gi/jXlpAI17RY
IEMCzUXO7tplsRPsHza0PAzygG3zZizQCrKQ/p2JKQCg9x9Y/BDIiZ3wGAoTL3l9PLXCWk4gosFz
W+FOcQzZJbdZ2bMQ4NcixpwqAHt7dzQL29bh/dzOePGtIgkzoiZ9OpXZXSZwMv9DyHr7QK4lWoUx
/NxeQAl3ep2Uqod2igKDbgEfQ3yD6pBnw0JJf5Fs3MkUUVYrG8sVc0Cu00BywYiLrtvOkPq6ltUF
9Rt3Y5lbHvL77uTU0k2hxwuxwYx0wWR8oYRgMzuhAJSKHTRK/efUOaDyZkDQ8XpVb0fhakz+pMxU
vB6q1x0O47MwWB+MyCnlvazhTZcvtN66/zRvyD0Gq7fm0vmvPlqpDbcyNwCRNQN5+GVBi88JDzqy
K1TP5kAXpGkDsqvumsEKRQaL3FK0ApjKwAu8GHtiPFglOEg81qsDq+bQoLMeY+Vcjh/E/CB1AGid
ZEtMQ0gBtdDfPQep7ChEfRE9Na1Vo2mUqTRXqXIGYOYz8Nf6dsjhcXjXueehL81QZFi6M6yHUPgo
PMh9TVuFuKouC6Vrp994zfKZuz5poGBKjPqxcpOhL7VdRQBvKzERm0s9xPDMnQHCBegq5VRRPD6o
zIDnJeKVQjiQNVT9yYvwQtzsDxYR7zZsaLyJH0BNs9fu043CoCw3pWgRo0vJBtBnTIcytv3XABDK
wGHrKpkmINSzi2RHNYg4lnC/p2QSKLmdtIrkMyYnVf67nQr41MjeLILjFUDDXtRlINCfac86vEoB
0Wrr2WIZeupLDRbpbv5sK2pdjelIVZ0o1hO4R8TG1nevctjYdFwW/On+TN/XPc3EDzur8bAsFNLP
EN1qFwx1Dw7MrXwVM2E45aP1bVihrvKURj26MWuD+G1HcmJGm5ia4Ia1rdk8sQYVuxLwz9M5Pv9K
AcWaAgDyS9TjzGqrA5ZHHfB8AbgB+crEqMjanEQpzuPrxuTJQCzNYfiKdHzw81f9isdmqwXcaYnh
qXPNVrffvjHwck0p7cZFB9ehW08vhNA4tfxjIwL3FZaQhuMcKHIV+u2Bk/NKEKj9KwB0eGf+Q992
SdThQR5GfRn29ZA/ZxejsHZiCLPxBQN8z1qFex4vC4mGIivT5Ju5W+2RK2k/xUHu1yEcygM4DwUu
4b1NELobykmh2Yqaefjz86Qlvqq7lJ6/yHkRP0JdeDEgYfsHXSrM5/kGJTSO2gUp1Vlz2ffrcakQ
ZpaRQycvLeOsTROlWEt+AxSiPO3xn6yMGH8GuAvqyhR/sVWDosEPaWuYg/NEr9L9eyayOkEZeTNx
sczDfQ4dCrih48ohyybJr6HzY5ERomnfRhMi06y3iujKnUPCjW/qskXQszghRxhF5E/bht6gMAs9
IEyZWlasq7n3cQKHizNoNOjxcQL7QL3coYJL2642/EBD21PRQFINanca5Bf1YwgKYcQEkkF1sidt
EALmwdHShurEdjGu6DQ+MyV6qxy496encZY0Ahh3Xoq9MngHqpT6BF8oXZE02UzTp38IoNFl9RZn
8bIntq7du2iTi6WpGmRf/q5Jqw++ypW7MjFeBTuR1V/0vd9HqtUutSOcV5Lh1F+jQvaZzaThTRBk
5MxyBFN3v6oulFejPOikVxfdMXwvhhlnlfgzZwFEP/Vxk4gXvMssQroDqsp7NlcoeeXw114yWMNB
vPBUHlylyfbOSEUESuCEOX65Z3VgWSX/+WiL8xUzqeg/Ptow2tUB6zyJi4PJI377uka1VCyeiMzr
gTJiQqq+CDTJpgSRbDlPXMkgfJLiz0dbStYAlYeePMJaPpI1x8n/tzDBydc+gfiA6DVwlccGuUil
epiKcYuMtLzgLQeMx7+fSCgkheX3cKrbWWaM6UuljsehGw26Vtuty+y7e3EsUOuQUxj+AQqZMlYv
36enIkpJ+BAyj2/hr8/fyMoxWYxRAvMp5VFdwctfXjwQjRAkSWhWGPOYLcs/d1rL4i8yi1jqC0ro
nwZKFda9G9KEcDMrMsaq9HXO0iSK1OBJQczi78MCqJYMVQHBHixgdEHfHbb5iuFpQPe9fCva8oU5
SB8aFHtEdjrqnykBH/6D2g43J4KJblZINglU9oy+Mwp9Op0J6wuFY1l6hejQ5ZRULluf+iFz3IKf
iUPrd4Muk5hyblztJCicfiCAekBr00KDULt3b4q6VFheHLauVSv12o7WUsyzGo5oH01qakudZ5Vb
hQXsQ6ud0PcpR+dF0wAKGMX20hfy12Tl+UVBNcr804VVv53uNzFIA6gTPeYt6J//BSoaznhDRBJc
eiCBuIy1K8BEb6p81i6VSdLuKzZG2PItriT+dnyaNwDPY/ioub/M+XheNSC8u5HOwS/Jf1/s8YMR
4fVy24gAw/hTndGqUhMQM2IHfHkjzqBF0tkKrqYMQc4uLZmHnmJxWJro40K5CehjHlWvueS61Hbu
pH46dLIM4uj67sK53T6JnyKeitoEnELZrJzhDVGNw58dlxZSUpiT4LF0zfPEF+HhvzbcT/nX0H+j
NjQlnaFwvNhP4gkrYpcneKW6STHzxEEaXYTBHRTJIBWrCAym/2UmkhAQWWU4eo+hJIM27EzyVG0G
VSSxEFOb+lv3eI2ot//0Nm3O2/JHu9s0qbXVgEftzam6uATUfh41z7nDgBJYFKNFpxQoFQnCbVzq
TGDgA1PHcRplq4APrjA8APHriPGr4QBebB05XFuq57QCoOhYp5UQuhtYaJCGtwhOkBaGrWREYXL1
VqVWEcPTcgypuBrgZ2+cXCWLP5crfwKCWaC34rJ5yTbkwuaxvk+6gkuRNaXjiFsAiIc1Kw11R3SF
CfZzKKTeYnzpOvPyWTv8EykCAZLS1iZ644k4qJM0WTS+tDJ9SzirJRDqnsUaCiRaCFTz+tSApcs3
N0CIGRHWKQbdbhYGMHU7ZnUPGdyuSaKYTbGeqU6vaHPtsoSgEz02e/D3Lj+yuMqeAgXsjEkvgB/X
wqE2SKab7oCTk16c86eGvUbNWU6KFuLIPbEaaucAi4WfcTo5bT1oUJdRd3e12zcS9TlKEun9aYFx
3K9C06fcr8GtsPq5x7H4cBv7MKBfZx54iYWR3n8V+DDkl7eE8VLyKP1MHMSeEHh9PRcN6psPHgjc
rmJdVSyLEU0ekwJ455RvNa6tco2DfTj/acvcKenlnxkit1ipXbsSxbq8nW3Xfziv2wOyzfwx/K5H
N62HrCep0TWn8yEIEqHZuMWMVJaQxzc8EO9TjQgexHfDTcfmy00GnFtVkDbsJEWL3O2c0rbfLyaD
EE3zEN5ivcl0JHSx6S2mdDHJGb+Rg0PWEb/mtKWOSeTSuj/FNp0wJZb9fwCuZOx1TPDdbiNQDsUW
uwfhIDX6kA/BLpMKn0M3/qRMwwcUF69qTJxgu0ednVX9AA88c8mKnOG+yOHnuWUyOvVqZu+GAa5K
jxv3u9V4Fznrlf2HKsPEYGVNkrKXcQa7vf1rqW/Zbg8rOQIjxt7K9/N9WaKFXjo6DgbmAt6c0VFZ
cLkimCd8y8POYO50ERZEJyhIHFZx+7U1U00LfwAQTC7oCXk0XHeK5x7eV3wZZHJt2Kdk/tTnnza/
fT0CKYKcX9PYqc9kixUnJEcfjU3fJ5d6x6bsnCnwPnemyoplV7gAsuj1lr5FZ3MwCfZm0U+Sf2Fh
3zIVPU0Wrubx3zd5Fi1w4ayYVmjUEtL0xqWfRCYNd1KnXrINq+2xB7HFy/TJ9Ur/63sVgKOICTgr
GBKEA5sSMIGQnnKYpVhspeU+RL7+D2raj0XXlAMKLuq5Ux5T0DH6437iMq7Nv/8dgsTYeKbEQI8F
GDjT7Ag1A8rDaYRGQyiNZ09HaNRf4VHgI5oqGaJ4nzlCGiochK702nSY68hn/2GBeLcsopj+M3BC
xPLVXXbG1eR/ThzAtBleSBr8ZJJ8g4qhl4LkBK4/Tkg5bZFAMPH4PgFG97YNrEFjASmktbeJJMOA
eOM9RAwgciYod9htTiONnQJhwt4xpjpUrhVHg8538JuRfs+s8420UWWpYnvg0krzgkO0GOgq/TI0
doWg5uZZNh7UyHp0xfPL2AfSImfRX2SY2LA31HNBiFGAZLQtqcDBXXMjSfAFgWul7MTOqzb6YIxm
QxR2Dy9bEe9hUlpJ9zwW6oUVyLbRYOKo+WEQeHqUvFoR/Z4rpHymYoDpDpwXs2yRLngJHzaU8QLz
focRVSDYm/fSVRW8P6WmBdzjCoOZa+/OJLw+8MRoidD0hnEZ2BIQD8jmSoLuBaG7JX3uyNwVvTaB
9fwXKNm/IHtqenWpAhLVhhPEhzDyHaEcHnmdUfqTIUr7DypiWiWCyCNLbEaCyia7HkDdi5iOG1gX
L4+tcAn1Hknd71rFEsY8LXIvrNqgn5iVRLwgPtlNvMXtCNscRPnung6MK4c04tovju7PBegTWeuL
ZGzEgNRJdB5JCNo3pXrKaN4ljjWd+e5vgD3nmh5LTZuaZ2/zJxJR76hTyYJKr4CcEUdAx7dKuzJx
buq7TXAxMi7TYU12QggjFF5Itb0W72SMNWqC8kikuerw2ilkCNwb5jVT3Pe93deBsz5Saaozlx/Y
QiMIwofrgzS/pa6LJhqFQZ+1zlBYaxPnLuK9yFHbwKC6YC0i1W+r3On22oPYd8i8Y2E+5e/f5bxy
bxwfQRCPAb7Lk/eWUbvpq0kcU7mzatjHZndTlBhEkj81OGS/omyPt3+sj8DAJN6xK3jNLV3Skvb+
KE3Piq5fBhWPKqVh4qQgSO724y3q3B2PwPSqWsFJiWSmNI1S03UF5NnlSGuVCnRR6ZeyLrc0ddlD
CQW0mPiuLV0xNuzFR4TeFojWRAYwulaTr/0gkTRZ18bG9ELSdxwp/KMHYm+JJ5b0UkGz3GCn3+bx
kXfJg0Y4EXZILklXzAhFl2yg0Ma8O49pbkueRicE34GFx7M7x5esQwz6SQKolA9CDbKBw4hpP2QD
l7XP2TsFV+uRHM8zISi68cNtnPgj/RxchBzsih2vBKPRg+OM1kFYeNXnhNjozM1Ick7170poVKBt
WHVgVfm2IWxK2l4iG4UCKffaGiWioWuQZY6eWvvezaQCZKm00EJJfVs1Gj+U0npGQkN1FASaZ/mG
reyMS2rJWVHXxJleMbghczU26cVkAQLGwhSugl9++Yk8cY1NXOoQed9IGSxHEiOanimU/YP5lBwf
6DFA+gnqKKSFWxcS43sBbREm+fjJ189HeVTWPsTy2vgVImHAG7uTU9YXJkvba72H4V84EXRg9QuH
Ktosiu+PzH+/xZ2RTr15Xskl/CIYdN08jS276+Qy1HYWmKxEhq7vzS4inZDFZHFQVIZduDDyNxCk
CvRmbud2VZTCmiV7HU9D3BjGT0fFFADGLik2STfqmwm2N3SpC/LNW5+PbVu1rnG7DelEPOqboNxF
VVeNeF2L0rBHedwLrHLhC+J/DXXLvIO3djKg8Tz4BaMfq9xMCon+Ao5NSPnLtaKGJ17enR5vuf7O
NHWtH6OgN7fVf0WNUVntYBthAOHYmzhC2jrvR77kV8TS44aEeoGgsXN1ytJzmWpCno6dneRDWsrr
1uNUKIztmbCcSmdFV0XLNaW+oRh1FNZPUktl/wdWke5PCwhSrM1OJL63C3QBJtA6E4dBGFsaXeKR
AktEDrcPPndSzhineYi99DzL578BpGj+NpWmXiHf7SsUAYxHAhJRaDdkU0TZzs0TiE27rfM6frq9
8plwVfDN26NesazmaTqgEW1ydY04p735bL35mJjMf1DRID40XD3tI2a726xkgE3pZssN1rYJLlRw
dTdo1k2Vk0vF1Oa1tmbAtLc/l14EiQdIWGeYFQdwOk+Bqd0jMzDlHchQWPuztleEodaGSyTTQDOc
NsQBa7JMedrPtRfl3Q3mPhou4byjd3tu2lKC4TPsjuWKIUAcMpXdUwuu7UwwSeF9JI5gDJdUHMMe
qMpY59tdqlAYPDoVHdGfSwVzvCdKuyZkqqeR/kaJiOYDS0Kw6Y0wnG8cQOLNwZYa8VihCmZr8yTG
hgEHY6IDYSrOXGOUi2ohueJZAHjUAh06zHqe9CJLs/kzI4cHALbEplBcFD0wRnDprsvTVkuMHuE+
Jc9ZpCT1DTkhEFXADpqkzwiolyAlJB/CwUewfQgRkzMuhmAHX/wK5Qp0s0hp/0RgSsNkXv4T2Jj4
g8jKzp49k+La9dIP+bFI4xhd5ZZtJc5HYlECnu9ZG5EPlwCSDPKnqVL++CMQrH0tJKtEUaKYzJgN
gGfi7BwiURJvU4m36lZLO8tHmWwsqboiOgpuDOIjuPMZCggLhQ26f1n4FpvQyTPuA6G34zZPxw7w
eqE+5uol+cuooEXfHJkyOVEjT+kf3bHdBaEJ4PqNT+7eCNj+nTLruBTd0wkdeymzWQFLFAgfEVg0
4t0PJMRni8IqGGNzjHcgV0xKTlL6qVXiRweTiW4L4Vd4euGdmgnIhNJGR+kf1TT5F/Un7xACDtmk
4IKDc68lbz7fVMFzGv/hGnUmEQpzm7Gt9pyrhW83MyEAsEHhObPbGJ3CIDNLJQ5E8DFuo+3sP5MP
hTXb349BydAV8lZUh5GD/1cdVf8kQ7MD3Ur1bHaT8RTPlOvWg0ZBVNYbzx/2uJAlqPJLwQ87besU
OkvxorRRfe3d6Nh7b2DArvotOohHVLN1HQMwEBjpYXVCIPF4AshnwcNqKX2ROdzAZnr+CEnx4sLD
1vRiZZx2lpBPCeR+gNgOpcra8x0QoMeADt5r7E/fnm0WxwYlFd3CLlI89gnI58CFlOSN2FgWus74
3L87X0zwbwgxnnZmDc5Sp/TJBrQvTdxv5wxIEDOq50JXwZcBYE8VNhBiNhMKQNjBFy0LuZKvRGmB
HwMrrMwlTghJnLy4wmQbMKjmppnvtARU0GFrAHatwFXOIw/tJ0cG+uIo7F3ylXkckM8VkVDSUAcz
Eb/V0OwWnBKrLhm4LSdrgFLJMS4ZdVecdhfluSOpWQUv6K4PYkZDW1ZDmo9N4AdIO4VoLGCR35C4
p9JZVofIJhzZTbzw8rGLaO3y6sxnMSUZg2DBaswi1DNAXWj0UvqnoAEFvQMqr4Ek5HB8GS3mXql7
AjXtJNXHq5LAqTWrmPD7LAaJjo6cKsadwUsg8trsY+SSxBUc4v0o2kdarB/cSuYwYE+7yC1KtGz2
/yFDtgTFsqYG7LIP9V8S/5xIfcJzrNConr/LbLxblCrDdhjVRdhO14x77gXbfod1Xmh0OIOLp9Q6
pqNOh0w1gzWopvnyix8FeMdgZE4rJXZyAS1TXp8ONSWt76ewYnIyvio6tsoJ3oys7oCANHA9fyDW
OUAXO8JsBK5AALfmYd0ACwtb0qk4uLZfRWrW5Ek8w48sdEQ/eqMdVSJfld7rj8sIkGO27QCyItlg
PMyJUWVgll0QotYa+wPAk8Q6n7zTnsSbc1HyjG34rxA5upa+3rl8fFKR9N+JkUYPsRZGRnYgxv/r
tQQrqaPjFrNL6f+OckZGuuGsItEK9kaFZllwe16zV6HSlz4AdoRV0X+lr1HxlKRkWNUm1xFGfAbq
tlOQJnaiYESCzT+dnS8TNJu9g93d/5RMEOws+4CNZCl7RoLkApkLHhuyESf7oN+7jHIQC79nig20
HHTwV142H2vzBN9v1BiTgV8mYonuq3wsfmtp1P1Zvt0VdBxM3hJ37oEwh3Fty4dX496UVeEHchkD
ompv80DDglSeOxf3+DoxVYhbRKjNClc0geI1lo9bQQSj3F49Lk87AY1i84S53YUfflFW2O7NY7y0
3FXvrKge09j0T2gf9gBDCnOY+SZPFgxbrtcDrSyM6S8aeSNcUnFN8fSq9tGEHSWAUTW5qrTSSo0A
7ln3thAsuMUqahkXvdBlfQ9Dq5EI7S7WYjrLhzxC5fG0ZBxA8IkH+iKRKVMywwlmrtx3SrkO4zx6
znou3v6GBavQWqVUA00GrSlJsi7Zj8jlxBF22t/bfL5eXas/IIvK4cesuzVqZ0SUYh3rtVyTf5r+
XrgJd82elJn0uDn+kri7Pjp69sH/XJ0U94gpAwY8Jq2+PC1K8srCk8cES5na9nHIGqBiowePUlNr
HT0nQHoexBNIYkUH/9VM7vm6OO+HmEYye7Do0xNXkKN7nEGmwW72N9xtwcXh4NthU5ILNaFQcUeb
jIBRtJD5iIk+emBIL8PcOcIszgrtpV8oBpIdrZqE5QPxLAPtJ7yaAmcghF6vo04UFtzDIahxVjG+
Sd/Gs95vmI01nF4wdhVRDbsGbpnPNe2joVrBoyKmRGQyeaB3ScwBPge1Z5GboAc9/9QiuVZJJFRx
5QRQdsww7ziurfVWUfYnFGudGiweT+P2AGp+roZptn1LZXnPuxL7V2nSMk85zYzGukBZccA3pvbI
5qeH8PES8aEuMAOrmTuVI6XJ0u3TkfFJZnZ2mQAugAstS/2N4abMKhd1y40cqPseoY980IKjGNVZ
roicfVESAMA3x4U4YFxjRPqQBOMhx/yGw3O2RkT0GjekhPGwbYBkWiHKyt+vu4w46DPcGObdbO0q
HwMwb4LZmW/441u/luOO6p3ovs195weKFxPjO8Xkre9XOQvPIMytxvxAGZZ7l66jFdkFyGX7lKl/
gBJhGcxG1GHM3dyVVGGIUzGMY2vGNUMUC+xMeENcS9LIPj/TnlXrSjOdDZ2K29+Xyu4jiILlgLyc
zwNOxwmQ9/UQWB0pRYpfZ6jWHrpWUW/S2ZiD4vADmUqn9qcMqV6o4kKKj1CMk9ATnvTHMYXMRzXs
wLY6r4tTjtuI9UdXAQWf5NaZQ45x2SbmF5ainZEgJAd0eiSWKlToQ+oT46B2HUY/msJJjK05W4YW
pkze0chGJYHelRnaSqLh3xYHXB6QkqSkreIV6I+77XIiNAbKRifUrMwoqCPS4Y/q0aB1qu4ExoJW
S8CONeD+rDe7LJFF+7iw2ircgBQK5tm2XXc6zsznl9vGLB28Na2D+Nig7amB5hrU8NTweAvLomy6
xH0z0x041F6diIVqKs+ICj4v4u+kTzLYoWJgVBXG9CpiXZuZobzSpbGLgJneDqttI11KHMo4ii/e
gQEXFH7OMXBnkE9ekye94oWvoxG5Bi7P4ZYz75DCK7+NoqtJaFINRE0PL8pzD0NHZo08d0Ze2cNE
mzTn+2HNGg2eRjvaG1JzITRbgLb2WI2oMwGJPCouehaDX4lH85YQUBo8HxhDd/o1nGP4tsDXcP3n
KRhKoR/WJh6z5SiapNUBqC11f0FO/iTYbkybsPPeXxABxPL7gCuiWVmHK1LLdcv0CrI91stFGdg7
t1ZZDspo0RGgqOtluvYKRO4lTDD2/Kfq4Qfr+LlA5eeW8BE2lD0ZLqfjNoZYywd9P4Rx3aj2gn4I
qozXFxQduGBPWkbFTAQfVmyEa2FwJkE5YkhaNR3dvMlEpYsN3JTlvNTOnCO3ZITkK9N/j+MBfcDB
h9ciqSRL8S5WJywZbMKjWYXXRQlsXxHMMIHHFfGMNApH8sMq7a+ZTKY1LsrQRUCTo+oxrFtzC1bD
a5lORsc7cikhRvVbdGdJhNg8veZcrvAC08wQ5UTvtHtDdXl6Qn7bSfMGKyO9DSFn+utpfSSLnfxH
84jbu9AmjlKzdZagbIaFUWMmnN1l4l7nTdKa+42721nc3bUh3v5/xHFxTabUDTyZEyQHdWZ8J7bc
9QM7/KEIYmR8RlfHP25OPpNLHuM6uwLXc14Otu7KcUWNO4sqezGTEXS/Hc56sDUbL4wp5XEUfRPI
Pf5WF18UkdizLtMpxugEDOftvrlPMQiUQC3zg3JyJ2yA65Pf7l0SaQOE/b4I+qd19oZnS0h4URrr
mmYYrQ9fgkdaJE99quwEQFQVXFuNjH6+busPDVIB/3rhpiLSF6Kg3kkERgf/mEZbYpm1O7tmCKPg
Pq/KrrvhfIj1kQOBuAEIWy4TLJA+76PVozOmXOQi1jqbyg1WVq2WTZqFJbD8Fmk2jXzn1FV05Inz
dGwBCZ5roL7gErw5ZrhQldT5EUPlkVOMdJT1MRDkLuptt5t7Xx3xIRCmaO7kRRUldnrQAPsuCwCF
B8YBKpCsZ7+w/KPAfEW4G5mcbxK6IO1VsRuqsHuRGZcyZZ3E8dxLlpP45Umv94AAxBNy8hnqDeBY
kfp45xBSrYsc7w2bsXImJPuTk1owh4SvRqO7knGGmx1WOw9GFNN19ydi/RmexjmVi6wBYEWknj39
2tuD/3e+VdtuA0Kp1ApidKCiw6Ri5+tKxLXlJ7ldj17uin1NuFvUGK5NBKk5VQHMcWk/QbM8IbO/
boh7XoQau3nwVmkJwjJLWk/a8jjZER8/24c0ppYjvo1X9we9ibC3qAt9mFRGwto8EwkFkz36tH0y
NcUO/c9wLEPxUsCTH0WqS8CFZTaDKtWB+OGURGYMzlEJiWzzvwDvCWQW1aAKlPz4SmXDWemvtjoz
77cfYT9MAU9zv6CzIRJYjBMaHep+8JzsIYbjpOOWxFv1h2VpsqzhYbEvb3QxiaprfWq5eD0m3xrI
d+51z4y1AlYEz/R7Ifc75AEzTl1hGX6wMzmWjLfVCbLXbt5/NqOU70yga0C7qeiBiIc/POfe94Sx
dTY4uJsLcFlUEHs0GRGVECSWz9Em7H6CYqZYQBWeRmfnTPkWLRVmAz/Lq3JbvYkauhqu9j2bBsS0
tQSm++JL85ocmzN91MyipUlWzX57m6TwuekG74mQqeGhYYfntFN0bxrbkt2FXymMqGfywEhjD2Ju
G4GYnDVls70UPu2KeBD13tUxfUC+TuZTTMgZfaLO932cjvhGH8tg9nw5FlY1MPSgPfo/JeGMb8hv
UGQIfON+RfB5ZQzMjSqS7tmVmzkDk4aQ9MV2tm9AlpA64P8KAh/NljuhSCU4ZYu57O0mka0nAj00
iuzmhp88GLyOEJ9IkS+WOQZZQQ/PyHRljFrTDxfBQ/GKBG8qnc44Qv1VBXF1bbYIFtAauR1etD8t
QJ5GFRx6pepmXDXbh3RGYr+VX6+p2y/wxh8hyNYAU4LQZ8yvgVMccIX6LHeAGzT2xy05nzQCZoDA
wh2SXv/PxVuGcnlzEIy/6bpww1xOe9m0XDCPMnLpxvLqFHJ5Ydtx2xhNE3t3MljFzX7jPjqeqyMn
6o+s4ULBwLgVAv4l7kXLoI3+w+hDJ8ND67vBLltyoJOGCWgcIn+w/+8jy76SrP4LhVI7qApPQNWM
iOIXEDVZ9Ay6I5JxyhuYsou33E0N4cKKIel32/fhlpIvviMNO4BqCvaHzPtywv61108607I79fnB
GEEKAUp1MFu+sFxZZmpOYd5w0AQntlY6vSG5iT/8AbLl7SLkfiUV3ALO0W4Tm5btGEJTheTF1JGD
dX8q8qrtzaE7THp1LEqG6BGtOoACjA/QWb4iM3ycs4xA+TXOU1s0idDKitXXvkmSeKS4NqwNPSEu
gboyMfmNmCafh4qrpjHoFKymyCF9WvgCbcYJ+gGb+TcUQ7c+DcyCtxkaVoiR+pZncIoQU/lps0PL
9qlG65gWlrzHHdm+5gdzzrsVeTgSl4ooWzxzR3If9XqNDEzSE42AgNucEXh7QL4z2dsJF/qFsrGO
fT7ZAJdEAYrRoAxoPYs0njJ3za8n113HfON6a2ncrsU1jIy8tTNQHI0ESdAMfTBad/MVyDfL19nb
r004Ie2KdWGk51YdlSqRxC4+j/rbhO/1Z19LTyhyCIvJ4US1RzG/SR1F7cHjkN+ff/8PhKL2URh+
xO4yNjWMO0b7QKeEUo3WXEvgrAnZhNulq7It2PxgoGTaRhhnbSyW0syjGlFAdkPSyHmN1uz32ac4
uj/IW5ShgAc6KeKtR3cwBXK6onHk//4Dl09DT0SAXrdhjWrVzTavbpxfZeUu0wy1OPRwN0/lLZM6
+Jt4hpsBMBX1wBGiVKztDyrIGq417PSxnz0G2JMJxaPHTLU2Dr2uindJxbxsNcPoprb215RiQ+aX
XMgBdfBgR4Hlkhn+3/S7J+wW277hhUkeSnrhF5Jyg4u0wn+ft6IUm/l9epxrNIyu46G6n9Fsl4Ne
QIze8TNixdVlXuNET4KsPFvXW9qU6i7zVmUwoT9RZ7b5zMpEj401DKYkHkFvy89gDBS+0QTcJjiS
pxQBaEo7YMmjhyhQBHGeWJUsq/3Rll7M+MM8WoloPdfzVCkCXI4y30AnnhZI0b7x00yCw/wWo9w2
xhMrpOKY58w2dNhkOmCVr+lGWTBb9ZJbROxHlKO6/9NMi+h9A+48zrjAfx5UG2UXXULqPQtDC+M4
XYmcvDpwCO9dC1SCN3Uu6Q6zsqNVsYTc17dstbmRrLLJTE0HrWrcyomLZXEWzMWnU4X7f7j8pdoj
+F2nFwzMRm0Env+NBtt5C2JpajZV+UYf/5WyE8NYeRb6SNkFa/yWKNmqQq7gOKujHf85l3dU8pHQ
5OXBbjdXbBxkgDL8Zdjc9y0+ym1q6F5uiGPsQdLrrcAtbERexBppgbzx49jZ4AmnU4FkcgoD3tha
OGdUDjQ/60oqjL0+k6SbwjOSdSBB1KVnVzeCyFFoJMFFygOWjNyGcPL3MusUcanJWUgXQD9zpdff
PwyqUNN1tLroo4UPPNMAFkjZFz0jCRVrZpcOfgicMRPLbfJVBa9wgd6SEcrVeWjN0oVwCBeNs2/y
oy4lAJxUe9qxDwLEqT4DMlOpWaf1C2q/dSd7p+tgRfYQ91dXf6LSrtR5EIQiOeDyK+OC9IfwUT0w
/0EXdw2ONki9Qz1miK9zvexWQgbgGca/1oxhBeRyB9ZcKFP/JwJiRpcINkfI9zlCV98Gad4YVZZs
xSqjjdN3gbSJAH3EOgUB+rKQxixmOkuhPBAIeYwK10PRJL5leNnxX7qlhLb25dr7Nsbxz1B0HZ2z
NOP7n9vW42uQqiqGk/EHcL7NzGvPXNnZzZlPSm7LJ8ykfSJmFrQXoRO+CpO78FGdStBkzjLAL/z5
ZPQk/nS8Nz0OkRnU/EWq37KCUevnzRKYSf01ty988m/CKK7duMDJGHGsCvs6YYQAJfJiUjsN2mfB
IzutxLjiQE4L7AflHpBTGZ2aV7xDd04lPn7rIO+ZA5CG40Lr4FWRDXBWeGDmsMhIasBlnWcEnJNk
oBirLdGO4I2PtuGJApj/6JyWB8pv4hYE0HDannObz4uX1MffalI6kRgeVm8YOrILmsSo2Fq2MHGG
K5HUgexX7PMDtbdIaI3Amlb0NdH29GvPmhII+aQviZSRO87D6GxvMsaexYQtgZFcXF8U7GyZY0o3
Xefn6aHPXO+ehMNa9+V6biE0Yejen2XzNPEfrNK/EzHOZIUddmh8miE6PM0YNf8f9RMwb7lehaPR
xlShbey3M47sPpaOX51OfBsDwybbu/qv2R2dI3zwS40WzLN2N6UyCMIl59ilop5gR2hn7Na0Z4y5
zj+TwFGL7X/FfH5ZP8Zz5HTw3kuSodyspZZwlDxnzbmRLk5/dsJvgSpkzUbrobH9I9rGIs9OFd3g
W/xz/dpdis9jNFL005icqIkPMNHcTXbscAJsyYYIU72a9bQ/sv+xsTB2223pPIBWOMqicRl2+lJs
emCKRJlpmpwXfB5xQRcPAV6bfSLIZ1VNqFQdyaFZ+ZCBmxyzC46IpubCuIuGPYPAekreBHZ3p+nQ
H8hi+r9u7LFL2zFdGEGvgyYArGlaCHkz7+sX7i33PhVdBD+LqU3xOlzJGcBtDb8JwHFU0oj7dc+W
qJUI9NDCLOyPs8bbU3s+YzGheaNSmWHQCP3JlFqtqS+Lj/JKHZyTqH6SP5x424eJTjSezrqEOUsv
r27hTHZhp0wPFh9WpaH4kIbgKaMlrg1/kcEc7N+1382OGzIMp0qX70a5x6lIGJgGDaGyLGhq+mOJ
T15vZLs3SLZDSoU3GCZvcZvTbBu2J1umLCwSghhgWGI71a7pFdgR88YHNth3EmE9l6l6Rp2xySaK
0ZrCmB9vn0yaNAMP7YW2sSPOd5phdLbe7M99C+EtUViwr6dvR4kj+pw2YBPTBRsfyoVOy/5TtTid
B9Fp96tNWWFSiEJvC38IoTPqbp2FZhgO3s4PgNMHTx4eDi0tJerVZuT02KrcCqrvykMLgjToCGU9
7o1yMdawZto7u3ghi9H5212paQdZbA09hh5060ut0DyOOlgNUr3lpYxw/pvJY7LlEM6Qpk0kwVgF
eIVegvxTJxpIP9/QuExVAe6KOBemFx+P2MMNq4+s4Vl9oH5YedYIA0KoHlMIKd8+ENMdBWG0WJGE
DKV2WBmWSEgYHMwqpPeQzOVehxTs5km/6CAXpKhzeghFPVyreTNp6iS3ek0bJqGJicAzwJO46kZv
cs0fYdcYmYvoMIEtCR/CKR2hWxJjY2BT0Gp062IRyrxjuOIUBFJWBwcuMvvJlI7kmJW4THmq+GLH
iAmvAb3xyLoplywG3rCK4Tybec8WWLkdHVj4aS8PXfZG4TemzhOMxa8DaCmsUS/Hco2ojQjJ7qj/
eeGKy/kLDLFDeWGdZ7uLGPeI2Ucdk/8H6DCBzygFM6wulsBNudvGew7P2CuYfoFAnrohOnICNZNN
hRmwkgh5mQooPUOpQmQbwtsz9hxQHJlTcffF2OwC5bDP4/KScI/AjsfPZ16OEICHCnvIZwF9d1Tr
caBXJq/4SjOwTdvYa9SnQcCAL/lBJzYkKouDakydqR9BlH7t/01HhE+Z6U8VeTVt8coxjEXsieEP
lwp+mPM6a3EadpT7FF8WqXmS/YqyqBKAYQ+ST6ZhriYXQi2GWId3qUnjfopA/5JhWDswMsSieHg7
ZqyL6rbwk9ZFFxA7sG99HodyMjTIE0KxigD6ZPJZna0rq8vB2FY2lQS7b+RKEmHqaiKqBNguSrGj
5sF4lu/GzZfJJHgu8NrX9bLSyF3WZ3l6DH4VORUtEDYWOwVgHTADKaJphgNbWpytYEjtTVN3nr1F
ZrCe747aUJZY20dgp8vdEOsU8I24F5F2utfXfORiehl8XYRyeV13apfojdndX0EZ4S2CFrBlb1DO
GtvqxHtYJPe89P+3IH5KndIeGb+CtMBKOq3cM/vc0OjFSUo5UyJ3bp1lPcslIokjDqvG42R7wMwt
b5DhHtN7ikookinqA1tVvjVkSXbkrnBUSgM8QbNpM/zDSQTt+T3SZdc0APao/hBYRpmnpFOCYxSu
wFJNl7haw3nWdCx7occk+map/vPzs6dsTeYioo6Mly92iACvbmvZL2jeNA6Ng69E++GT/yYVy3aY
smjOQPAaLTQBPsDrH+vuHz3lsdM9aVFcay18T5A9F5etPIgQI4jmkoW1qo/6VD6Ibx/vSEpaew8A
9fQdaBlK9JFz0WpOdc0uz5SKI3CbnuZLS/sQsCfPHMX/MOZWlpmacGk+w4nGV0ZiUoHTXjJSu1Mh
i/nAvB67mSHcUDO753CN5bCElW6iE/yR662m9uKprDik40+Xl6gz/whCafOSJQxdc2VS4X4lmbEs
6QbTLNPNpWQuEXSYEXqVVxJzkSGwgHSCWuuQSd42XzmsEVnFAe2jEvFTUt89PbPFZ2kTxEINzlu7
yUWQzZIg5zkT6e2RhpEsg/LeEOfGvkohWPo09Qwct+AIm2mmsBxoBS9d1ot9UViXrIxcqplSqVIZ
i2th25URoLV7NfGgbpkNF8fjiWeBXBueyZqarrJpAICrzWAJe5yTTJTsu7wpe+gP5WK5elt08HvO
kXftlGnTxaJeLfBIqvH4xoQHJDweIMIGxN4RmfypgtI4w0SItZr6KE8S/7yNYZ+PpNQEFKvBQ/Cl
jsvL8WTka3fQkNgMUltFkNqLWQW41sYXNBAXbX6usadLqV79E5GNVQKOb7qlq97YYgZkR+AOZ3xf
Wtxx8W93gjaITtrch2074R0eVa6KHOeGDnDlL2HLAOmlnYONwGoSdPUkfjcbKPNDdxRpXIQNIH1E
Ub2jF5z+itz2SbqKcxpHQuyvDTXTsdGbakOf7BLsKynBFNpqu6zXfokY6PPBuc+o0YUxbGXqwszI
nJKnSElTPomUwjoaUPXRp1p2y/a6Cv3Mn8aR0G6QRV25jgBvW9ITz00yW384a2SrAb/jUVw5f5ZL
cIsBRq1gPLX/KzIeSO9soZT/2d11Ldj81++N1Au71epKLCf7JYQPL0Pu+LUbSig3MkUdOjslq2VF
kYA6fII+Ev6ExCAIfw07ferJi5/aRS+o4OoojqJhDyEHjmhbHUKFG618Irk8FXUSyVSVZN69jpwj
zKsgGjZ8qEtM4Le4rZNqWyTeBM3d24uHeY2fcaavLGEWHdiA4sLZqQvK2hPDqCA5qqHAE0xULgdt
LJQ44mE1/Rg/D54kORozDLiaCNNnWsSE6f2KIkj88QvIYEiO7iYL6BeXnKmGX11k1m8bwTWeHL3Y
vZfK7itbvQgG3rmzEfTF3ICJzmcBy5QueStJSSGHZrMhiYgjGKhsfzXtvmqmgJQMO+CISnvR0cwr
AXScdYJtTwxAAFIR8ZvCTn/pT2P/MYMdsz/o62Px75UFRs4K3pM7WDrC5WSZS4S3mKsusQuVZxVG
AK4odDXs+YZMUVaEAnNVpJTjqOX8esxVJjaPnvnd7G9X0vGi7gN2CHlJawgCdcbsAu0HjfGKEYZd
MX/ir/jkVQu6WwMwvdtxe8cRU9GM/cuVWzcRzdt60V+dYuHj33rykedvS7LhaNgfnj9ZGjxcG469
Q2uVLWi/S+H59GIvHrIkpyDsL31SyKI/soWSBPOaZzdOHfN7doE47ynlUWV4fTntbP9cwA/oqN3k
7WSbeFi/aNeehEljyRZaMksvigSrdd5CBSFlPUl/cicoowkMPt4opTEgkFD4CAB5Ko3Lk2zuchpM
ZmoV3YWRVrAvR6vdeT7Jyq3ad2+TXojqR+erbdNdjTwA3RSMiJJMmO+/cqsnpVBb4LA7uOZhSBbH
6FHq1M6AhGV/ZHRDpaKxOuIOJqGW1iizhjlK423kbikeRWK5+PW3eks8p5yuZcKz3V9WKz8zM/lU
qlUfl2lCK7evIjMkNF/Vr7kRJIPv4td+ihLHMRz6y/p/zXl/+uYZk7hhS5rkqKd4GonTSdQajx6U
ByQhEdAXgUUZExOsz9nFTW39+RWrkufXwz0B+sMgrmKyN3TOAlvRfVyolFLDq0w+ehyTqq7+nmu5
+ydGrwCEajn71ENtgUdLrmOgngJT27xq3nx/ojgpab0AqU6MpM0ozuJ3oI/s9rrV1E7lEaew+wqX
mXd00rQMvPoHaEtONdb5JiH8OZ4b5M9p7n9h9HICJhXBIROyJse9bnRkdwKD75npYULFzBU792qa
fa4RwGwKnJQ6CDVG2X1s3UGJYHlr6KFFKrUbYfahYUDXxlbXrIzv2TFbCbDwuef2EE3NHyjQws9/
sSxpckyOS1deiQ/HnzFl+tba4AvbpS9ZFUdRzbGP07adworI3vSHcOlNDx+9G7dEJ9xeb+LXLsKr
tGZKxXn9UCx4dp6GFKJc39zArDizR1e/etSisvD9EiyevE/4sEl1BuJEEKEZb0luFOA42MHOyzI3
ONogVHXGUlCi0ol9EAlvSwPSwx/K2qYvM45ciNVuR3ecl1P0VtAnznL+Xv/nbOm7HFBODTK7z4io
rCoqtEbo60gb915X3gR0dgGpaeoKRmEg0ylt8VjnkekF98UZPXGvTPw5fugLKoX0rj73NqLhWpa2
u0POWwQUsghCu+hBAI9t8GIGIV9p6cDhWVEzjXbzUiNkneqvSlIo1LDfINdQmbFr6wAvs4jj85+t
MebtPxJMrw3BmntRGPLQNdzwwtoyz4THqP6lO7xhe7fLPx6CS97wXh+CZ/B9TIpn/oOzWjL9uXFy
J9NCHj60L2Utvyc94kmHwqx346v90umNT60lhh+C58+rqSvFPs1QVHK6E2DIJDPyOoaYnNKTg/SI
Yep0R3HGJehYh7uqjhz2UuOM9hVXm9mFxL6K/B45qwgPSpwc+F3Euw9RDGJVo9aQ5r9/z1Y3qJDS
EeWKtN+X+Pd+5rzoQdkw3I+jubRHVUgcowat3C6qVbFtv6t59hVc32JW5XtIqW9fd1CKbeBv3a4J
96CKotiU/sOqQTfTQekTamd3ONpG9CQnUveXVveYUWsa7bRfMnw1S/4XzSIXYroUQJrO17LdAHjC
Lh51LEdQLb+FRp8byVBX7apbYf3h6w2wJ38XyuY6t0xaBHHrSl2HngzinFGfrdwWEcFdRH+UHV9O
phLAZtI0I2DTq+qphHFU0JiGgAVYhFrwN7VRXCisqJ4BmLWSbgFLybmTIruzEC8e+wzcoSt4jx2B
htaTM1GDxdW20qafQBEZfzBOLivtfg8uwZ1G4NfD9q0B5Et6LifvgDNsKlQiXkFXyriJREFDkiMj
x9FKzErijDPfcB5W2ZjKBOBHBHNEDECrRtfIrDRUdX6cV6ulvwdx4BsiU3peX0MTxqhliXe1LrkJ
NxzXGd14f21TpLxf00DheEUu49hLSV7R8QQy0/TehtDAG9kyPFC8n9bsf3WMeSFfsHPT2FEqcIVQ
o2qdE5oLa9WTBk/xs4Qj8R8z/xoG8STZc1Ev3TbbEV5gwGl1MUVnmcfaAxgHxCPtfhz/JE7HDBDI
1c696C/NczYakRkvfkuI7/sKUoGWFJB7EESRh9KBsbL1nbj5tOBit1Q0TZocdmlKEgXmIZZYB0q0
+E1hxQad09R4aJpIGkIR/daRaHT+zJGMNh1MMmsSActCrWHU2fwQYqTLHlRN+dTQJS6lgnfA4San
waCScC/y2XTBfSMMqSgkXHn+A6ujhoOSMPMJaYNoVARbRdDN5h2cRjEmlvpVbuus2Uh1eJdE4ibz
iuhITdCVbAwd43FgBTenw/wCxn0iKV60cXYoCHUq2tgH+kmsLB62vLtE4f4c3guaIHnJAF/eh4W/
mOPJ6jpUNfG+etub0nQKLVJOBS6boOGcFLCkW6AwvrJcGx3N/dd6kRE8YzLLBpzGBsiYrxObByCv
oQGhkYRdD12lIcQ2yf1Xt1wkaLYfWZNfYmj9HsNWDZzqQwzoCxSVywI1hAr5rLCd1fhaNE7zb32H
HIEkOvkv7sJ1feJBRt6s+fRO0GfhKK2sPI46o023jCuXfrQvhDLR1/x8l4UqdxJrpxR7X66yVWyF
M8ZRtPxiDw98vsBlK8YEu3VFW8i7BmhFAfK6LehPxmO/pnYHIZKOuBeYCa6mkumhujvSqSOX4SQx
thx73JkM2aR8mKO3A115S4raNsbv3mMVqQll1MJZ5Uvr9f0HUOgR4Fs/R1b63Ji8QAeHEW4zloyo
kK9N8QRliFC2yxbx7ZC4SH3yRYv7kmxOD4/l2Tpz/qbBWh5d43BS5vhAfhSgSSTsZ4rtCzWR9HYW
NdMR5w6GOSJb4oO3N5BQ1qjHdJ6k2OqgmUrKZ3RXpXgne8M6nE3I9BQbf5ASgyu/Q/Qux+3olSQG
130CkwMIkWY5hqvfmvky3eQEzIqSYW7KiP8xbNvBcZ4BOgHXjwyGwFIpXC99Sfn3AGfwdGGcgytH
Unap8MsQ6oe/h0v4joZqaNTa63M1ByrKgT17gW7FG6gLSn3Ef4MIXUeLU4iT/3RCXBj7ZQM86APE
TsWxwTSuNs1cdjUPoYmJJLdgT7EXEnRhRUo+Nk9lOCYDARJ0q4zN9RfR2hoRMDevheJ45sjWMNg9
IW7ZQ9noAmVTf7+4JBeQ2+QFbpiK88CV+HrLF8lhM6IknZLO79izTNfJAb9F6c0hdIVzeJyFs3Xo
XeGnmqgwFaJjdUsPphJw2qGZLiPE+1oa+zZYNit2QtvWgt4LjRQj+D2nLU5cSRm9KS/MiVd2ip7B
PFfATyBOaiNtvICZqfbzxbk2TouImiBFiNap80/9Q16VjcZ0HZhEV44XRgNX//AJ/McnJWPQ9xWE
WL/X7pa0nT1uxjMAlX6bLjwUs97jLRN3dldWdFgA3/vflX96voouTd/8gDecMkFczO9VuXSSjtv+
CMQVQGdao+40G+p51DDRFdQtkwy1JBexE5Pt17IJRWOnDJKnp4m51U002tY6spixatL2Ad7Sp2xE
XbRXxSOhY1iGQe1oKIckytVLi/ZEQ0kyNKHdbXoaTi15B54b276kPa3ycLTDHQpZwzcu6uDydaZz
yqG6pj4SJbLuSN+62sZtBmzn0qRd4EET70fpaNwvUKtC28zBLC7NcsJL8YuWX/eMmikLNpBpieQ2
7QmsMZHCHvnJ+9cfI8L+KDOcNi9dUsdoj9bkMPO6RjIEDOoe4ssaBkf83cH724edRE4GZKbcNWi0
tO2BjT64543CLiRZ40zGDumx2Ovq2LwyQk8FeRaFCX9PUsqyHfurnRblufwnA935egmBK4l59CM/
yxr2SKFjfkj7UITt3vcId2VZcTAIIoHK7OiAp50dIZP/D9TiowXgCqEL5pmn0PWB4IAnjWJI4RHZ
znZeZHs7LpmiA0KtjAZgx0Axr+PcuURu5+mJ7y+6PDgzEayGWpfe5Ecx2IydU87rApcL8jGkMUks
hYivdVpzWVF69Z168PpLIxatKul9uP0JLcPlspr0DIiPqstDRa9ypoeK0PC0mXiBcvktaqeZS61h
ZHGvFrFeV9STuglUr13oXUFJCxv3hGaZ1gvkAklNUaX4dMn9O05FMzjBLu4kFOvQDTIfMegRtZL6
JZWkFIZjSF2zv/GM4HBE7AYwD9o07giPkgWgqtq85yOCTmLL+EU15VMjkmKvAXAdKgkebvVfl4qn
sQko9nR84DYazcnAk15/4KcaDGuspc1XZgtrVrWzmQuimWBUEfqMLKUi9zo7sAzTayRhrPQHvBbp
raoUvc6TmMGLJRx/CgnhJ2hz5b04d40wqVj9nnDI35vXCgbXP8xmNJXt8IVRj/YuZxlCgXeYEN6S
wR62+MvzZ3uWjYQkXxCA6XJYsYZTGPy/mXw8fPSBWpvhxHW16G4bF/zztZCzofPX8GRYYouc4Wh/
w+299BMUertgrCakMymNCsOdx915nCi2TbBn9+ksuYj5C6qnK2HuAUKAV6pQuRzq3wXNigu0FPbR
BuidgANuvrwVL9pIFptqbfWAJlgRO7rjH+DhBQzPkna1ALZ6EuUhaWkkY35JTAlSD7kqtiNPoXH8
6GGy3EvjJGqF7VicNjQ12MKt8r5rEal+zKQCNek8HcnM/NNfK5AX0m3qftWdxgVu5Ap0DKO1daRK
QAA/upVvoc7yA+LNIdVDhc4xUjcHLDFg2ZMfwOEUfHGq866leZR4Mf7JbfOn4E2C1Win9sPLQf+g
/rGR1PT6uNKf5AhDWz8BwAfVi7W/y7iCcaGZDB29zZ/5ZJtkRDBkztgqtWI+9M5Qwm1mU6JcmtZB
7fFsaTgAUMjqIu1vVMPIs+Xqy8DJRRhstJ36JUuWlDsoM3k4SYsLmdeqcOkeda577i8I/mBDRUEH
57wD94roUIV02+ebwkRH4YR7Rh4lcgzs3oQ+FIlSZIv4qeIme41IUwzNyvpWG5e8vUASFz/afmH9
Hk9QdXktW4DfTLCXRLDNtZZ2TY6N1uV55xrDfyIU49kAcVzbTqxpwAH+WZEAGqfPjaelc3VNdyzV
s50KTnaqBX38s8RvKI3B8Oc4CVMfEAIU/ikX0hDbEeP4RnjPaDKg/AYhOUPG8yc4CcYdEqJ/goEQ
rFrBgmPBnRUgbGygu4kC4vN5QU+TtvSQtrDPx0z163hNzecY01WKSYVIH3QDPy/gW3mlWrcdw4bm
OB/XF4asuTgsBglDbbY++uO1t0QVjDbsbcAtmhs7dDcmNHlRsmCW310L8dt4DWl8087NysFCbOSW
L3ugbzTBujyBh/adgvGfw4dtGKGq95iUhMEoRmNxYRJRMSAOGwK468Z0kPL9kcaXl7uR7/iqksWT
CGRh4RHT3UpQxPkROgfq4CvAxrxmMn3/exnXqw8WXOrg8OrsuPdU6zL2FAAoH6Y2FXJoNQtz8Wx7
ib/AU8c3tT7M4FVSmJ3FsbDyApHnX8FN3yF/IuO0/Rx2+cL6UDe6SPJAB9AS1ntOHcCIYbsIDwmm
TNB5+dcuBDBvZqrOAW4+/fuf4pHZlbPk2jHeM40qBrVpU6qX1TTpa5hsIoE/S7ZdfrwRLyT2vSI7
JeYhRp/SiP6QP1jMy4iWfM/akKmhGmfbpalLJj9+R8m8RB9+mosLAfZzVRzYOj9fbJVodk1VdQVz
oXJX2+qMrJAw90NwVfiyffc5d/69MX2CsnR1oxzJ1y1qpCCaB25Rh++7Zd+sEcOWZM51ZMbJpqn/
mU5plRCM+PAyGrl4IMqiCZOOxkfb8hSM/lWVX3SWURb/MDUTpQZwlX9noWsL/XPbJThpCq+TTR8+
lig7XnvYyh5fdJMmHyl4/jCxSRX6llqGP5PusCHtUA18HIuHq8FaS9ep4xk1PgQeJblE+WwBgmYs
05FajG2yS+6U/tn3W9rXKyaHeAZGHX6OtWFaEjcsei3mYSg7k67f7Oi698m26Bab+mfOFq841TEM
EZUDVb2wFyxwe1m0AlMsAnH8okZHIQ+H+in0IBowD3+IIolRSKlgRBxs+YaYB3xNaU7ipbg8FHbw
bqAxHkRHNjvdL3eS70dt83EUv9gett0f4uSshxX3a8rrNGuUGS5jsbbiXuWgVCAAmvBpX4DoVz+I
krvYLlSS+voTU2exw/uNq0blz4vh3Dx0Y7i7603R9zE7wme1hC62a82rOuHh6JhBQIHkQNuIoMdW
pZaC7dCKcNlWdmstgYON5nW/ptOEXVCi38BBg+x+rNg5ez29jstYECFTmAgN+roxZNBqIQyPm6Yl
aHsav209osHjxHSfHXCRpIO+5RVDHV7AMWymjKC/qAfvZKqwnhLvw2ZphjA0EZZBt/2y3zwzGIkg
xcWbtlFeMcqIZwqFL2IBZ/ehHf1xvE+3Ln/4w+/TWYn8JG3ZfGIupe173AqXL5C22jg2D01ecv5U
q9HUqtNxfbMZf4b6CUEk8MRvNAiSPTg2KvtFlu0KU1KPnSl+dgYs1M2h5WS4kGMSVXignQ8jr9FP
Sk+9+MmUgA0nRQ/i0DPnY/HTpf8bDHlq2ehSArObTVp88MJ46Ooli5WhoyYGb04Ff8jka7Fe1btm
G7h09Qy5pPcEwatujE0PxID1b3QKAo8e9vNfwwWl8NLCdaRdoskWcFQz1SCikwvKAE9t1g6aGDXI
flr8okTqVJYL6ItiEkSai9Vuiqvq0nOqyeXtVJ11OaTN0pHU27R1+3CgBV8Jft/krg+dl6rfclhK
z722636KlJ49HtkH7GMeTWxIhKAR8xc52yf4lJHIFY2eBUIj7jpPZwbbAB5eOX27pXi4c9NCEKS+
rS658VZT0jHZPRQDq4HGdUuyUzilJM/EeBP8XbRQX+3XCTQhSppZjINvuWJOYZ0FvmevwEwyi6R5
0LW651aisebEcLlk7/3QaRE7DzMyCa0VJxwSqozAVXtUVa86dQ8CEXyEQvaW2sYB3NWopatzhIon
N7U7zpYH3SgC1zGmoPOPXca2fEoYTB5d/TXdijTXZEmsDrs5KBe661z+v+tcj+3Spp3YLJht5SLl
/o+FaugeNPd5MsOfcmvEuqxpwkxZlp35ZsxA4vblxiLHhHmWg8yBGKGuqoMsc9tfPY8NLBETcR98
G5O8xgBHNwxm1QXw3gAF9oqK63aH+K/ipUzA8gaA4Z9fuzbxNKp//XGV5XDM4rk8Id6IFyoR5NBH
Q3aq9pOnoaiThJsndqVp3sVRRf1yrhFyOyAm+9cugRxOgUUhhJhNhJ+drcRIdSoB2xswV+PYOcFW
Rz70sSnAoCS8qbYBCXie4ynlEpuHeFVgnV0rgztONUFfqPDsHAUdHUIYe9kf13dDgmB+E/RDLF9E
8YFRg9FgFz/rQbfFuLgWN0VMLnK9hmZar30RZgso1gEcMfo/4aFQEztpxPgLlep1EsJ5+soVD0/h
BOPv1jO3GsLuWx26zm5M9Eo5HgVceYdTy0WClUI1semkw4L5ZuuGvu8Lf1npqCQx4uCx+l4mH/qP
5S3aQce7dPY76RQZVW5o2gIyIdls7BRDuKdcaklbmdFeHoQZpC+P7fULs57y2vCe+HTwdkcQxgRd
ZNF3LCpXa+U451GLtVA+y4ZoQ8QMAvsjihVFY0CT9cd3iOsjsy9kZNzBHm1wB0uRuiZawDbs6ZPE
s0N5lCiIw9qsEi5XtwI9wRfAqvb4+G57sBoZTh63VZF0MyrNDqeGIApdYXHImk9geboB+eSigEky
R1leF49ja6k9GE9W0xjQvUrgiGeF+sf8kQk/oms4hbq6ZU1mf8lCOyQ/Otgfx6yKxewqc/LJXlLp
75lJurKyqM1yOVbKmHSD6dPVdprhqKIW90hn4KAQLFUNUgC2Xs9yfi8JFupSy5MbJgdmuuu4SyWA
myn05r7s7/FsJS6AUy+XmGp+Im7/OmpfevPjm6Mug7V7tqr1g1CI+ZPV48Z6+l99XfVgKq8Qy2Ss
Ov7VythAXaqvN81kU8j/TDqVhHDElszAP3DkR2wjhH4gkK+7QF9wV1M3IygPfH+YvCcUpwhsRWUl
Yuo30aVTs5ck6mfseOwtN9502ve14HehiFEHDuRLKFqCSq1QYIVSEX9TgO/fKJ2RYj8DwP1SjQrx
9VUoxPigld66I1DUvzcEQqjJvUL42pfW+TfI+upNYw2FCcEdT4cx1oLc68zeIPBAc2dnR8YPgm7e
Ny7bhgZKrglxV570ulh+3R2DxWTD+7iLg/k6CKdbkGzc0hcgf4LFkjNHbb83CTegAxYogYVDm5oy
rpp5LFxie9Y0Sybbo9veeO0r72e75TZPUet0V0j+S3IimFGmimu7DwaCW7WzKxAT5fOJeu5VwiM/
e5UuPQnlcGXooRQKstQ/At9EUKQKwV3WjwshGh1uNtH6bdMArT0cU+mAy0tjlxILBEMBM+NgqLQF
E4uxtdUhz48n2zo9W+zd826TLz1zSWzk7pIxe+lamAggWO0hGnSgvk6od+QeHjIYJ6n1hoqJpDmT
xAeZ/I5X+MRJ316ijYQbuZMw+i78QrnRbgoQebljygOmVA3Alw38hM4/z21lq6aeqMAb+fH1O8t0
fFkvOPl+g8HFs+1OFmvpau5nfHtxVSTeDgSCOL80oeVMHMwvw7zAxXVtwGvGP//2UmvTX5RZBGZW
srFd0aBTCMc40pGznc4rNSFYNcR+72gYZbWu9Plj99Cd3voGrTq3XwLsFpRTTQNiniZWU5vsDYM4
2IWS5ckGzbg1qkEF3YL95sYtAWIH7ZzSOrBSjJrxXdWC2KpEIdP0Z3YBgeF/ylypW99P+85EMkOB
ukvXsKtryKrnrESOOmEX10OxgBcjo0RfHOk1d7zkfgCLyZ0RTXcufaEZl0emOLXuTLdAHYufQh3u
XcqSh418V3TX7TWJjeedm6KgZtAytrcNdWHqlLHSMCgeoiw7hvi5zZKnb+o2Oi66QUcBYg9ON+hX
5qR4U5BnZoUSX49vnIoTf2WPXfCgTDqu6nSVlE3YBucZchuj66Hk84I2vFj3BTZuD/pPXMyAJ6XR
TwsdB59vlwiAU3AGC/pURH5ejYeTzZXpbsA0SZ70nWW2DWAv0p95uys0fQV15Nu5Jnwrj/e843lS
ikZBLNKIk3eFVjxUdimiHAhkhwG+ogG8a9hKwtghIuktyHBJYzAXbAZgfsxLMVdv06f7KNrDZ2jk
jFsVh8hhJf0L6NDl/hjh9KHoz4cdEK8DClyhnkrTKd+ldXnhcz8rs1NShXnLWilfkW6l7fPe67Vu
uPA4jegHic+IJ46rsLZDq13rD8dX152K7dBt6u4+1p9TBJ3OEISPW6KQxPlBPyr4DrK+i1n5zPdY
G0KQwcTDeOSETZZ9vKiwNfbgnOa6vdUg1VFHE11j5Z4LqeNuhj3/9QybeaZvsEXGO6XxibOLXqNR
06A4hGzD1pw2rdaKzyurzaKuOOCs1CTA1Kpe2wUJJoGubygiXRnOMZIDnx/oTriaOTEW4tYHIWnI
y10mXJFswFN4EGQPWfxmDIPrVKH6vAWqGXdNkXWhrAdvg5CgLbtUgXILPl0O/HHMqOtdSkjQ9KRw
Z7cYMRcL1J7vQd8iQj3fU7iqjX3K376bCcNDNxMYIek6ZTxbMqb33LH3+TuZXQC/zw0YOydd5Rxq
Nkk0j7ZY/z28a2zB8Hqh0ckHWz0O4T3ZEVUAqsEpZSOQNjLcF/d4yhWqhtLHJKsJiS5Zoj1r5CHx
A70skZNGW0jDwvgPxVVlnQCFsJWN2OOeCIeJ9EtDQbOjVI26kdgHO+OqsVeqS/aaFHoJ9wl0KXpx
uD2r06zpapMeqDgS3AuSoiXE2JkmPoPWmxGNil3/u4wNidWv3jyDw4JVU4GfO6kxnoafvIwieGc5
T+4DwP4J3b3+ZWPZacNc4sAVfP5AsrnEb8r8LmQeHMqzwCd52LHCxEuwdu5dH54v1n77wSDKPPXk
3aJ1niPk6B/WDshR8SliO07xO0fQ8dZtVxf4kGoMG5nUaly7hGRk6IkGP42zJQVvRd6i9pVUgMWz
5K+lOJnPeqJlyx+4RpFk+iBAI1ofD5ih0tzO3ZU2QDy1+Egpc3dCnqolAfvlpZ2nLGPBO6xQCHsH
e1Tdzf4DBR+WKuZ/y8sbGvTkB0GF2QRohP8trWrF0220VVvJnL5qZY+WV6wTIEqkvb7ew2SHYfpE
KAsTI1kX29ckT7E/R5dvXifglk3zhip2itSM1iq3GilXLaM2DGpvEPkJKxglAR84ExCrsjeULGH1
saHE65M6cIGspaEiXlHtubcp+KtrpjAMM9tEvyEwQGHyP7S6k1IH5B4UsMK1LulrWakdojjWsK7x
ElKXLvUK7+SqvJAJh3zgUBcD39tK9IH4rb7jEEsNMKH1iKhClcg0exUXbBIR0WqUfiwAXKKWk1vU
XMY1nmCjxqQ1YdZ4tRPgPZJcOktlCWsjrNskYL0AC3RVARvqQU3N9nsqIBrKWbuzpvtxIsqGEtb7
zGLnpUzFOEiPCDgUHSM54ZNye3Y3XOsQ4UQTp6T9xCiXTJd7km+uPBZnF42WQgKUnVbwqnUtFDlz
jB+6M47zHYBEyJCdZdj5e5dKuoTcNZd9bVjnxdGoMt7a3B3trmLslyqoIsnAUgpd0mQ/0zgOQY/t
yPY7E0lYY98UBI4tYy+pLW10GXyOvYYpeflSQ+WUq2B2zmeoWxJBI9SBXrgrxez64+7zWEGXoT5s
3AcunpowYppx0bJDQXzKq+yXe0SnUZzdILZnHFlOrVm1yEHp27fCyy7GrJhJeUh8JtHQUFWyOY/H
zV+PP3u5tsPWbEqknQvwoT5mQ1oQkad6sWZvdBk0odgS9AnbrZNzPVwoYM488hR7NJTbCH6i6q7c
uwEGXzsoi0MMoBkZS5C94WMMJP8f3qdmdjU1V5mFs+ZQJD1e41OIyc2fraVvDdFs74p4DBGOzs5p
RKhOpBPloiYaG412JhfE+IWZ/I1UzeqnAGP3O5PaQMkFU4rnajInZAQr8rqcYUGDUUodMWk+j8Aa
dQUYONTTCQRysrc0yGV0rosEG2Y07+r1xE2HQmQqmnbXoBqec9NXnQ5PPBl2MKgCYbK9YNToeagX
3UBmljAE8YGmoISxyIS9qrX24Q1LFE5wmCXOT3T5aOMo31+QVSlEIEBdox/YrHII5LBto5L3lGDq
+qMSVlIXu/KVtjCdStK1Edf7r4teVvf2mtafxckGqyuHG+iBoMVSIQXQA58SNeDgj7J8WcNHstjo
akRsRxxKv9YBegp8X95yiL/1o76wKsHeqY1D2A359FAHfgYeCLvkk2NUlXRr4Dw4oVJarGFtVSMC
fWd+81NNLRulisOTPPmxcWo7doeRHcnE/8JpHZdA/P2FBqhtlZM1YVCZ3JpppxgeunEBNyXxETcG
2evshmUkgmvAAPSm5UG/BUhv6+jb8tv+Xff0iyR3FhORYT3/b5zOWTz923XA1izr8g6+m/soLOAK
klFG7DS27kOUC3MXUcXa0qLK8QalK8REbxWE7tknryJTBM9Pn/wASbe1n7cT9Yvl3cZet0vKyXGd
OWD0681ysazQ1PLyRVrjjkV08dKtIO2vJ82b/0EV5boxBJa7dH9rYrTuP9FhOnkL/aMaSRETW2h9
0nYXZIrDErLfl1gBq1hqKLTiakuxkOiEb7+/aT3hLY5fgYIwTxjS7D5aZfeqKSUlsazIaD2HEjwo
Qv1mF6uC0Owglkr0x7wRw7CzoR84B0i1f5EXI22ScpGnGQImsRxOIU+Q3rqr6T/eH1HW+hs6vu20
lEqqIldZHAbRkZBUYNOXgJfi/mF0mSnbTj+o/e+OoADodnASofQbzYXOUB7sFwB9GHdSNZg1uxPf
34rtRvn4ym0lbHqFKspqaN1ytymZEECelxXiPIr3LeAKYgzSJLr8Yynszr8XH/BJIljtgHbgUCkn
zZIreGonRuWxYAVhfN3Yalbl7R3c9+o6sS4SEO22e9b0+TShiXIHoMnc+4b4xMAOzybo0Rt6Mhb3
qE/hLApKrawqCb1dMnAB9a7qXu6GkFBDbQKcBeQBxPb+tAiD+veV6iQ5uZoKEB/aDRo8i2YOPbvq
6BE9qTfXXYFvKKjPMRc2hijyjhqw6PLD/tX2Z14CRyt89WqLlKwGELSkeIkJVI//GNkQDyegelie
yaq5YSJBJQnOrLkdIRmD0sYyw24BmeFhe0d2Qv9wgL5+nayWdebV1feMKm0O7Otg3CMZmolSprEc
P3lsXe9/io6qMJuE1YhLmkSO+RqlrZlugUNDFXx17zkY+WICMEYYS1trwd5cw/NCqUyItjyZW9jf
yTjOWh5jE5Q8WRHU8epa3U52+3xmXEcQCaI80cE8Kokshj+OVXb8PdOG3bcgFraySe+WIWoxPl4M
mOPJZrkO0y2ntAqer6/YcFehQLbnAOB91amZWfRgufAs1ra6XBvZqPKwsacNJYM18TTVI7o20y3G
W0yYvfljFV4hOuHTBbrbfowiYfZb+z2tdd/NgSGBFvVPSeu6/mrmQ4uy3XL2wtLkkGtWfBEuoiOx
w8af/I7A67Ecd/b2Un86iyzShadJqQ5CMXa8JvMzo377yd+l5JBoy5wcaI0GqZhlzagmmtlSkrf0
QCu4rig1IO22Az9VFLkXsm5eWz/Ycv37yt/fxAD68IxlfcmFhHyULKaI9wdUoT2hgVXuQuNnUcVF
xnfqB6snolvJVGAvLKH8c2/YDel3gwpk8/JTdOPCu7im3xRWXosAFxRW0N1q8bOWUu6K3uN3jpQ8
JMvJP9SRMTpM2ihNYgeb/ebFhOtGeuFSslPZlvEAa0amYqEAHO6Jskj8GqHlyDUoaI9HC00i6IRJ
KYt8xrKe4bvYOSYS5nSW2VPNYSZ6boa7f5fVVbZDu7a2TDKNFDkSAC9ppB35wyHbp3QoYG3V3C72
/5Mvhq/owDhHpzRqyrni6h1NsYJSeTarwYTES710ovWhCNItTBCHvhxqRyFS+aG1YAYG+j1zyjBu
aajeGsh1+YCp5OSvI1s2XjsNjbMulJZNiNmUtcQpgTf2Wvm2y2TztVh98F566kSkuidxslfy1Oja
Z1QYpQp49/j9QPhcBprd6hp+yf+230I76kHauBIGsy/oj4DbAwhNuICsZqK21H5j18QgYnQg7Ory
vAV3qYlf3f2ncGHWyyl36nHwAF0SkVPUrSye9cObQ83cmS5nqd3DfK2vv+vqi0OaTwhOAr0qHP0a
od4l36m3N9i1UdaYoYQBQl2QdxQArVUHfGp4AMShr0sJQ2JKxFMglw7FtxtxPLlTMcBxib/9f/2u
9ENfyN38ffu0Sv2LSIT7rzcBAg13fSm/jrIQRiMxI09HoevTCXe442Egd0Ibg+JuTMCpi/eqCexZ
hK31LHAxP9hiZPk3Ag9SHyvVQxyAQHp932ihd1sX7yOtE/dlwkpqNgoYtCh9OOfgGfFg9Fm3Utc6
pHMr7AMHJCZQ4HK6UVzsSzhFd89ZgRieVh7UtP4l6P8l0wSPBCPBgn8NiMLypOXKjxYp8dQm9/rw
dMqd2s7abn8Cr02heZxyCSw/FAKCrTG/3wSBsK4gQ9AhwgSF5okbgZQ3NG8YFvIQGsUJVpK8Niun
PZ3ZAXB8jhYW/nE2pjcqn3/gTASNjL7R3SKUsc0ryRT+qZJXhhn1yQgRFzlgPwZ5VptPe/zb4Ao1
nd9rPgty0j1ymPcrJ8BZpxaD47lU9Sa1oSnTnhCGj6utz7APxDj5kv7Ov1ZeYbK8cYDH6WSc3b/4
ilJp1v+fSj2wuNAyCMwyLwYrMjQoNquzH/YNx00RCJoTHCqQ4BH/Z+rDl0hs9WZ0M7Tsl49euVN3
dpqfgbBgk5rXjY22abGrLYDE94kwFjqbmNM/1zSbEz4+4vcjsugwuc6Ltaof5NYmrvVfdVoA20n/
RJKkOyIixk5h/cE3O0/XYZjN5i/zPk6r45oJgWprgYB7r9U4FCGroYLzSJdi7Qgfskaz+jicnrP8
ZLypwjbp2NRgNMaT0q5D8/ztRBAq0zD3peEc6yxGs0Fkpw8OjI+SeJUgjlFyOa+wfbkLQFLQjS7w
FceyihfxAwQiN5hayLwsIJfx02ngsu+eQvtpaXicMd88ObFDGYR/rrrSO50vB456zhaQY/bEO3FH
FqcTDHPHno81BVj33do0MUGjrrQKkuMWY2Jf9BxLbFMMzAo59q7gQpx7gVrAZXiTwYFHVIslxOsy
YodFOzsy+5UMXSYXXJAmTRF8Z9ZUYJcge91N7q+K/wTPQsTTcKKSzkmipEjB9esTOtdD6QLCxTHB
iabEpHd5xGbntsZm8tK7FvKMVE8a2HvVsMsK68zVlSgP4TTByDALo8P5q8grwa2/qVz7gz2lIPNr
Kv90N2Vx0OikKM8eGDDdCBv/OQCY7D31q8cJcFf4VOHtFH0z6bQ6h1yJQqYfSMvaFXSCl3P9wZNQ
7Ar73bsMb6vcKkfIWKvK9+TRUJmiap5q9uXtnYTCcdywdmF6HfSz1JMTvx5pT4W5sugWsoGS4oWK
2RCGa9Ts/CNQEnnuj3Zr/etzvfTfwJ7DWpL6ntTlBdMGGJfu8Gi3dSCd7On2ei7XwH39hIvdS4u2
bfb6fg/3QneyLHuXfnqlOkQ4MKC3JbL2y/AkDfagIQGn9ndRKkRcAAiWFdrPQ6ADXdxhl83w/RUe
nirYqEfNmnDEtwfZqqZk2393N3YcpKu5oiGa5rN1WGPebr2ftCo1aHc5VtpfnNYu87k4MQQO73ul
QroVlFBWflyfGLfEt3IuAGgCjWAHVoSRGCgxbUGzkLad2FEyDt4zc4VsE4wg+2pfYCtMakQp9Ssc
RpnFy6STTGYUJdMDX00Tk9jMhIonh8ICiNzfjyBgpUE3L0FT9TB4CPl0QyNrJErSzqIexu8x66+D
b1PSUxgp9UueO55t5nmYdyPtHqbejnakUSFc3ywNzjrCgD4sJvPpYo75Aff+MLtyVeMPDkCuebgv
z/yVbjJesFYbIwYhgVbDGUeydE++drEtk67dtdXmh1MKugjBZW1T/g8gDOLwn92koQZFGyvR8BdF
YwgvAi0Lsbfsp4H5hKS0Kig+loWK0xIK9faGekOkIXI15LtYr1ibCPDy8FPVxNo92oZFWihLDDsp
zRtkr0NXcUS9Fw8Bu7vEqAnGRIuHO/pXvGBYE6Pl6b0urYD4ALq0n2dOPqDNrqNp01D10QkkJk+g
kNPKwGIIgIG6TYhbCjAVSQUko7L8XIOI36yebUMNaJIp6ovEfBM3HDcibnqO/srGpwcOwwwJAcJG
y1ECZGfr2GDXtNUsmH/XeKVG/M9piX+z4w2dUhBiiJY2QXgbF3oKE0djzwmH0nNxisOoC3AePbck
xoyPKkCIzy0nj8yR62LUShzFbVs1GSDVVN/Vk14op8FOXPt5X/IoVABoSlXSTi8OdKLKNOcQfv3A
dQFNulr95xhtAXHMrI99fNIOKrRob3L5FRfvNAI/MjHCSyPkdU0F8HBAAbZSJ6PFp+Yvk+nU1Q6R
Cior4J/dClfw0IHfM+LsK8AI5fkQk8Of1EzZypAHYuhd/hPPwwl0hOjzRIbhWEa3uC3ADoYq6qri
mB+DdslsztzyaSb7HUAuUuucNsLoyxnVSE2/VB0v6PPfoGAgCtVWaadB1Lal65O5cZnOAcYL8LPj
iP3XzW5NJNk7IutMw5ZYFmiRbC0EkHzNiBq0X3sMfVsXqXAfp7DjVljCmKNMsrWPD6ybbvVFMJ4b
+afmtbTD6DmNyuvplFA5Ge+7hd87gGW58DS6zinjr+DRDSb7wn8qIFXQ9tz9663PkMUgVNqB+d5k
Pa8JIJar6g/Gdl5H0sIvvROi/sDVLpgCcHOKFwDhrQTarpRTcwZqb3sgrPzCPtH975ldlzYaNd+M
HEmwCztw5Sc9s4mW/5lqY+AXl6E9JWoRE2p99kNkNaZmP/bPYdJIOFxsXH24nL0n5+8g5Fnq5N+y
xcYQyPjNgByk2RN1nxlj1bjzXgoLNNr2O7eBoiuQ+WOlIIMTkmwMWh0HK5h7bGgilrSU/7fdMg7z
BdRutdwRTF4dHdqzvIL2+UBwsjm3+r9I2cJd8Pf/BvlGRD5s7ggN+twTovG5k8+wDoQyMDUPTH+N
Ezy7a6fuy1RfOcHql9/4UCDuY1oe0Yw3ClIuzfKFHQzDMlRhslWMaIskuCK/I6tDd0Vg8/VYwrfU
YNWfvUuHADkZ96Jx14bQVHzl0bPDFhY5f7y6zey8EhQRa1ex6oZhjTWMDN/l0Lg0cJfJtybJdFeb
ZikU5/JlgYGmk0aocLg7l3nzVX0Ac6bn9aqApyp0sJIFdnN6R0tap2wdi/pQHZpIkMj9E7gyT3TN
OmlKSuuzyb2t89Ft8Soe+v1agji6fPmw9hNkOiyC0ru0k0rTVcL9e+AnHEnWWx28baXqIBYJ+SBB
WG3h3OjTeec0y1gX+nJeTsBrmuPYWYkSB1fFdZVp45IYzNKjfOLTSXy4LTffBv4f2EU5qV2sPnlk
dqJR7BJ3np7OhRMTdv2eOklTgBW/LAHxZoQZ432rGp6I5TrE55cAhQBu3KKG92PqBUd3rL3pFKjV
bFfOQF2AE2C7mbnEACFqIlY2XwpHGx55U2sySAyigZEcQI1fmW35sZnBpNuxZmhiLfPH6pnVKa0u
tIANtJKox9SLDCNjmVh94jBGbjeAuXYDm1Mgck5xsF6sZNdXok4H9WIZBAYR8HOQkO0Y/KUmFQVF
sSZShkkKwSydWCPSQn5EsDQseBrmJqFDlTWyV0Qww7zC8ORwmcehylc7xJ20lsgl8InsAJ3DWhwb
T3OlbF6agRusGdHVVb2mT2Ttnq7s7pMgSw2ID/sGwYGTX7Jgn0n+oE0VAxhQZy0HltPqKMcjwPgL
IPPH+7fmknvxPmdPZwYc7SjgColeNT4ILpFsuyaDWgJrnNZvvEuhvy1GnoRp9SLzST1OgMsno+qY
/95/j7zKlmFBV9dAnh0NQD4T6tZaviLvOVhAQXPRbjo62U8E+EiULcAo0Atz5WCyspbDedDPFNpq
YSd6jGxUN9eOrEflTVm5Vdhurnl4cZz2KsW+VlA6T2ik50uP89pXfmvz6/vSkF40xg6MSPy9VXRY
tS/2G1Vejx0Ss+hqqw+k7G4Ch47dj3eSLrPU3TZxZEDlL3sY9mHyKWsVtxG12tP05eiKVFPEe2Bi
g/BH9bNJyCnKhTEv+Ax4LbOCVKGG2iBAdMAPadV/IYDYMhmYX0BScWYpJt0ZzmDEvg5bRBaDKsmO
JCRVSA1pMsv5fgTOo7qD4jx8Onqa0eijGtCfQWUeVwLFhYy/TDDwz81dgqjDIOi10o37NrLwSC8C
6/rr3KVg0yjtrAuOXVuP5ICp7o6NAxDLyj6UhnRc3IgpLshx2g92Xl50OKQlp2VirOMtBAs6ZQrK
3yTmpY/ctfsdhJ7Nn2nZJ3EBIdl7KS/Q3cjKqcfWtEmtGzURUz/ZOM949t1HKmOYKndCYQ8qNsXo
9M/1nTCU3zP6pXWm1kRR671EV7SnFP21tjQkg6a96jv6vLKhZuu92DbuFMTqI5Zj+BQK9IWifhjm
j8cRT3OdEFty4Sennbi0W8QJseVJBG7CR+lS7TGFE90wmmdkBcsXs97J1akjrS8RHdJXJyFqEg7L
D/5eu3kj7GjCm9ShjhNHvH1BJ5eezD4gsoQG5IN2sbCAnjNu8gyd1fjoZp10+LCUA4t5Guk53aVI
cSI+rqhkGV0WXLDutW4pluLAuJ7s+l/0AO2I0zy9LdlZagVmm20y5WLS3/59VO72NiNj2RyngMm9
AtO0NxUO9dLin9HL+3W8Ua0o0c00oY2ijzNPpRcwbIl6wA1HyMT9LSIavOUhGbvO6PLOo6ortxPl
CI7Zhr0ru6t5m9SjMAEwD8DOn1ShPYQ9PXp1+o5RTMuz4bTYe4VkOeq2FizkejTkDr5GlgO87j90
5ESA4AG2FefzliROj4W+u8gbQCQih3FRXsfJJDAQOyDQ0Sgfiqu9NalHKxBZSnrWmrke4WcrqUUX
6lIHANCnwoiDQ42ovHX5I5/DYg5X8eYL4X4RGgeu8gxa6NmSJslqb8/Fvz0MQ+65I55eM/FPWCnt
JclfXrlKoEUmefJNOi1RC6peCAhikMcd9Wh6ohIDOp1RiSSMDEAdqY4KZ8cDSqc/7c1THgXcUhKm
xphSQW/0CoIhDPPOaPOoyyedujd1pJaiV5rbnHSnaVljDhGrjIwTjDlPXyDdQRqwIWx4JjMkoPWO
Vnm2IcgdsaP+Fs9oZEAXvY2dQKsMpu2LNJl2m+93loo8zNnlQrCKLk6vy3kcoDedaI8/Wrou6rE5
efiyMZ6VW5BsnwcXc/EcJnQpd2tsQjN1Zrmfe0ly8FLZCJ/toiI61bTX3doIrrHKdALAJFS3y2x1
8DIUnsllEbUS9WVK4HMSVQD95tL0EKfVxTqvHJefEXuCQFOrJ/a2GUxuQMgpzjOoxdOrRHH0PYeR
9TPQFMIv12cCRc44W2SvnXt57ZFj4v/m3Vu8a9z9lxYUuRJZYWUDkpvqb1zTeAEtCBf3rm12bvPL
j9/i8WNAdppGoyKeMemCrnNONPNvkdOC/HwJjHrrXhq2VtgAvPSOS4lrKFgNBgKsXgTuKZwfmDGE
BTaC0SapwGwDz79cmUqn99dTQMg8pUcUjsktuy6esQ/sl7ymcHe2nwCRqDRP1Xc+CzkBfkZT3EZ0
U7Y/3M7cvB8Rz9rtSqE3q+56VdHgDtim2PORQxAtJqF+LFaBN+6fel2JVLt0zdLgJrYnUTzyvIxl
iLS9x9jtJz0V8iChSVHdZlWb6RgsRha+zD7Ps/Z+qPkk8WWltIOi8uEAC4WaaSSjr4LAGZ80ONuz
HfkSTyVbDNvrdg+3k+1Ph2JDIYYXbakldhflDeSZHXW0U4CV2HiPNGNmVm6BjxKeeBMwuSc4L7y8
EWN9fYeKOkGeSjOVxu4tkPfjXwTgsNZEDBfFVLglnwNX6A0lzREgdNnphIwNNT4oD3n2z8Yk9elV
G7VQ/Efqe5H3FEiQr4VokFA9y32u5Qlu/mLgHtFM+scUuCXy/WKX2B11PsTmxAMDgTSkhpMmsKaW
BFzSS/3igl1O142/Tb5CQTdni4X/YqR0tWWb8He9glean2dSnTaLmUZTmnrgox6dT4XRXGaxifkU
z1z/bSHw/hDpq9kyFY9mIQ3icjA16Bs/eV6nf3MNwH1PrzY0KFkbZamb8IfaOOepUStqfTVet0E8
m7jRCb/ocSGglgYbYGAK7gdeHNOvFMMUVRGss2fYcYa4bCyQb7+TKZSHzMTd/oGrA9Atyj1Xs2ig
o+lXVPtNEk++vXYB5pqfbWs3actpIiUVrIkCpA8KPqIWLuf5oRcf6qFZhq9uZ3mWbJsgwDNXCluy
pl181CoJL8QF7LLJXK37xrittm3g082XzpIO/Ln29jam2sh9nDzGdnLpVy0SEUsTy2uwfRFiAH/8
NkYySZoYufDTlKUeVvOokoHc8emgnYjEWFe6dvVoDfDR04uQprcemI9rLWWvzSCyPdHBbOl/177g
5Z0Vphpf89nlCLyKgvA7ZRniBNAKDxy0w/zIZy7kvNY5WIVsIfR/PaCx1SfeZx9orFMOw4wlRIk5
wh/VumIeprng8aq8cKx7/u+2TVKqaq7E6hElld7AEQm6HuRzbEeOGWgiozDFA3QMOYdgAr93U3xN
9kd2YMO+cE3EXqB7VzLOtPdXK/N+C38UpWDkLz82lS0IPQmjd1lw2TOWTgTC+s9Rr+NcUnpnsBUh
SfFBgSCHQLvhLj6m1p9Y9SoTEqtUgatS8jKZq/CXTB8DLOQiVL2Yj+JkKMaZ/dku8lT4fdyt0j3B
QXhVqp2kG4LsBfpa3zEmPqPA/jeq34YAlY6zJNS8h/fPBLqvo/IwC1PubL/ZwWBIvm5ut/zKihl/
yZR7aG2wpdyVJhnnYcYgQOk48MoGtD5O6jMKsxhoL2EO9f3pvUCVZAuIHlbNMNYzjVRHKD30BrOe
YhD3jJr6QTdJXJMbOa0E4T1Gw0C+q/c0XtOgb3sXnf8SaiX9DuRezoXNYf2nLe+tfa10eRYHZFAs
/IoyRjf+N/amryZbJXHajjd7gY1LBF8fgbCnYalpzWcfGn4DsVylj3MYUyxjmCzfQI9vzxEXC4di
A+HRgakSnMi4Sq1VIXApzreQ/QHNK8+5uVdezoRDHU4PGwRRbXZHSxul6QW4kNH31izcH/S4MIkM
c095G4ciML+C0pc7RkoZG7AuPfyN72OOXbXuB/hEvdu+8wBuQGRiqGF9BsPbbLY9BiyJypd82XdP
n2y9AXshBNOx9m1EgudJTLiAF0piI7FH/SCu21tOMMOcVZAHlp0k5a7bP3Pp/UR/zQw8vMrbqJLV
fyJH50xjGhHCTU/Mm8oF1pkWa/9ghbMRBSGSAbgE7TiMYlmRBkiQLu0/4+S9btokmDtT9g1KPIZM
ftrsb/oj7oWwjraaPO1e0e31tyIgw6d51KOVSBd7/vA4PDoCoBqv57mhfOBuZhTsg46JRUisqK8q
gx69YYdVpoODraznfBdWefU333B/L1qH0GsWRSg52QN4mgsUfqeYEfGD+g9rTE4goQ7hipErksxc
+gqUGy6arg9A0xcErEF8PMyV9EqC8mrzWDztsz3Afx7dr61l+h32rP412Pb/v0fJ/JqJ6vdgv5Jh
Ql4kB8PBDONC14yRG++HAWEs8rAhpWm7GLV9fLPqxOHye2dyNufg5v6/Z8uPwfeWvX9uvKKu+BCj
vTg5uMMWeyaxtUeBnvLGrov4/hM2x3uM563L3sm6DYcaNk/hWfvHN7AWgkvRttXvT5rrv3CsveCt
mzY4uHGEiuvVHqKrF4umX+iLCxAuzs7A8LoYUfsW6tJs2RLNai1Ab/LSJm2gqrOStN2L4VZKHbNl
hBd04O0vjTmpiPqvE3rf9+lW1fDLS6Q5Ooy7Un+6ukxIDKhPGr0mxlDGTyTwxSguXv4w9NKqWbWo
MkEkvqKFzebz8ia5ighTOXTcLtfu/6KRha9wWMouDhiYYzwao/2rRG/V10b1MGH4PvPJTdhvNS9M
kb92s1bXfujqCKddf1ld7CyiFZIuBGBwbttlSfZlwxIg8SI93tVJ/z4JXZ5uzotOmzWbr/OzpRLv
wHhuHraWgyv9DJnSatb9IcH4rAfn4do9SKkKldh53kxmb0cXmk+hVzzYb6cL2btbXWGNQn39fI0t
Gh2N30vgngeHA4hU0lybOd942+wioZFog0ZFF6mQ9wng40yC7rxxE/vMaWff/YN+OcLbKfH9VbeP
Qlgb98UX9uTdhjU0bxj/hDMnq+7AEJe/kHJFZkB3hxm8DxkgRggZ8zsE+ulWyDw5bc1lkKnU/bu7
YMlrLEm7oNjFTsqG611SO6HkdsLcS1O1GQuEK9NlAM+nn83m1HNALyDWnWfbiVm8rKFuKSCzTlUz
MUb8W+ujYsE3nePHgjqt72o791fcpXmnVxo0asLmC5B79PoEhZH9mhkUSo2Snu+BkokEQsdqdvxa
I399dYIqfBtheX3ZoV51adM5OFLhNakS/938zdCtrPij0roqheV9aT0c12g9cdPwPfidyeN/ExeS
n6KSLI+BujGJTvxyHBDQTLg+DyeX0QavX8z0iZW26z4tMxKD+cmc7egHuiVvpTgLGf3eQdSssf9c
xTzxMpyhjwtWCqt5yJ/KRcbiNaSHBfk3LAoVphvzQQPdnh/YfQEDS9+m+pU6YM4B26pNWBVPoJZf
B2UgC9VMtU6/YI0lmrBgx9eh+KJmU5YF0ezOXN8yh1RF8YYLwdS+b6Goyq11fWPCfD6+7J0Wrwjw
EzjSkOiLl4WqmlbLwQLvW6D8GqtrGTKsG1EFsr07L9Ye3eSgYIu3+SIzpE/KypFS2JGxT1JzHp/7
Bz0fN9om0KHIEHSLblDXabdWu8B5tCcxMnvwBiNxPGAUr0lwsEDx/mg8zVdGd4Lr6+JimZVRvspv
QWQQh9QcqlU/OD3RzS0RJbiRyCdZ0kRBsS2VPspEp29eb5CK+PSuxd008mhy0eUgN+Xbwl9dgbWp
D4uQOehy2y21VZgIiidCHcfs08Ul4RxuPS3+2pk6gI/+oOgUjrq6+IxcxiGgWFQYORXOirUEk5xQ
X59BCfFdt2TzFDYqz07gUXt7t80M70eilVxv0e2FrAMyO9JcYGj1d8yFALYpE6EBd3blHoclQiJZ
KL2FnbnqFd0BgCmD98mQ1lUlLRwO6YZ2RHy7CeMKeITTq8DHMzXT6AF5vdNr3F0tMllAMDeQ1bC0
vatQH1QrfAlzgtocf8x++MsHbcC0BTCtgrQ5MCDsWbNx1PRy3HBaxevkiFde0eY+DPy3C47nVdHc
bd3dXAYgjX2cN//nwoGPPPU8PyDpe364xN5F3Q6YxOeMuvC2YF6fTkYfC6Pwu63Ko1Vu0jgSexlc
ZVjMlIwC0MYP3rc96MIqGkHFgWz6zfWumOHmWi8ZkQjQHg9ymr4ciANgmtIoepE4n7RmWVVudMKC
T8nOnbjbqI/5oJoBQY6+z95KBOZsD9f2vSGe7W147jK/VKRsPxxLRNAwAMsBVCHZ23dXVvswZtWV
w4qF5rY0yrlByQ3at5Vt9qDRKMibokW5Og1DWUhKMxVijgmEt9xApZ8ba0R/VwwsFFwJ83NL3BMW
J4QxL/uk/OB3bp9zZy2Zxx69+SVzYo8Pwwbctnr/vTAIWxcuHFiHve8xhL0GnB5P4ktpr0sCH3+U
HV3ODaxB1fJkcH7EOgBulh6tgjpqYx+RaJDFMO8ysHrtUKPq0nUNX9lH5UN3TwJ8Uga+5G3lBu39
+bHWQC/bzkZ5ltTzR5XorivkvpnMTQh3durOC2BC+9/glJF4u/TU2lD7O0WpEQVJ+PdZvBfhS5KZ
sUltM4Vp4qTIk+xRXLFb/TlSdcEkkwcBf4qnzbQrPp5t2tpjTFK5OjfCpmAy+uWiDzlhmtcB7qMo
ToR5WdbTsPcXLY+Ez1uoY4gv9MHP1++dZlvJX1c8OMyKAGYttifl7DetX0r6NttbkkL1A6ccUvCb
qY+ZFHP6DIP3tDvMCzWxkTCV+BUoU8WY0q74Ywf0/sIh+hYvOZPrlAfDbyqUHr2/vmO3QUD3oxeg
KVlHPVgpjObN+AnhqMJj7ftOa2EQE9pOHCkmbWCIMlO2iCedDLdI84qzQCKQBkOkW4VQHI8GesMw
nLkDX8pQFfbLEY6PrFKgY7paCPZ0tO9KeE9ADUEw1vUc98AIuM3yMc4Zwg9W/WkDP0AM6erYiHUY
wWPCFTpMueYsoXgGG3orO0aWMyFeEntJ0V+tX6mFTM5nfUuR1ezX471bjyfUCkio5Df6n7pWAXsv
e6wo4eh0G+hK9/hbSRr6bB4tax/V6c/e1pBYMEJAjSmY+QCDzvKOHJrpqnPcSY4Ud7HrJ6N1H+S1
QuEIa7ju1tG55SAhgsyODJRAaRcZ7apCghoe+zP5YBP8QJknKdDpZhnrWIjYmrZp5gSTH7irwQJM
4uypmY4pEPuCZBuUw+KWPZNloxbx4RECl8/oZtQXOwhLh/IDiZMV1Kl+5seoqLF3duNOgniq+VVc
4oxGOfyITfTt+EELZz9v13momNHl7oFyHIn3fNrf0gQ0BJYqHVlKexK9I2fNERq+g0g+d6Cl3P+B
38+9MwHpAqRnCLwEs3zWpyh1TEXgxsj7SwqiN+WIRAd+O6LCFWXgDRz1Kxy8C7FGcMSWfA3+iTiE
QBmhXH3LG1WfQNpQqbiCzLDjncKyAlOdUzOoTsMv5/BzxMZ6j+A+UuO53WzIA7yEXBbYLMgU4DKz
GuHrjsm39rdOLAHIbG2OVyjFu7A2GipireDVpWFBu5wyxZ7U4MznFXJogwmbkx9zAAEx1fAHUXiR
kqpayKyWj/YuvNtXL+mFB8VS0JBRz6c1YCpm9kk6Ln1WOSCXTBlfbOZ1iSWE8jzWNDt0VFotBaGX
GcHwt8a1v2vVnWihbkU2zINNlvFbXgw6qxffHUGQ6vwbut3/BAywqTmZY1kO385ARTI7zJUBy8jo
Xfma9gD9/Icry4696j9Mf8ac8rLceIz5RGCHy4/IFg4uP4TCSxNHMeDmxEbRTRk7k7OoFe11cVi4
tapIHCXBhu3r9qpH5/zjuhQnhoWNwH7p9iiUlzUUCetD8y8cbJUD5twjfKYnywJaQpxlg2ZEedwT
2BphlXGtwoiwxQsEyxRBup5dfMPtpzJCRa4zcOOr9YdNQmiEl7SfaHkzLQ5mTd4aw9UP5xgO9jsn
jKujgccbMqYYPydTC38w+NUCTxiin6hfpcfUV9fxP5q4kpcpr6yDU1F561nnm0iEcKD8Jbj1Hztm
NfHG4vOo7DP7Z4eyYLSsdMWNc2/WNvH4awmkKmGq1kfwGfifPeMUQYr2AIoHnJbTShEHrnQ/y5El
UiQxHSowD4uZX0fwu0JN3qNK79d6gcK3lEclgWiK8+kh6xGpFfWqrf3OmEdferOBh+zbLTGWE6O3
/nDtn18pJ0DdVEzOb0T/+lls1QRx4hK8bpG4ucoIAkjyKj6Ev9ho/yDkI6HDhtndsE/CyGnktIlq
WCFvcri0JKZP82TNU5oKrGNGdJ2JTYbTlX/F4LZvBaUUrtFC722BzYxejZcF4LZv1MNESmJtHJ7V
skEVEYq3w1zhFtFhQgvG8uYnKNAO9XQG5PIIvPu1sqA7gmQddORTrMErKuZO7uKdsEyqygFksue9
C3gC2oWB4Xy1UaV05n6prgYNKjb1OHxp8I89KH9U8hmiCbDx51LKOj/NEP+Wa5Ug2k9geDcyZajD
RWyU7W6BiCcE8q1+UDeszWJ9Ott55kdPlF7xUC+c9Xy2vAlLrtHJcGZPKXyBBDzRvfNc96yVcLgK
T8LcLNfI6QZaB2xtyeYaNjIci5/gVpOFHOR6ixuJiCS9Il3YYzRUtTkkLfxarhjEoaR9wd1ASuXv
FMTI04WGhKSZ7yCu6GA88x6SkDthIt+bJyfMxry9Kkt6THNfnQms0dmAJU4s5VR1Q8f61U3xPhRg
zWCHxbcgbaKv422WI/meiL2dW0hogsy9sKDIVs59okCm0LRSSgB4giougXv4R/7D0K0ceed6MNlX
8g5GNrJSLV6oV47VMr+jHLwLKDNyo6Z6U/crdI+N7t9YJWJWw4yxhXFRQadlJLbIC2XZPyWIATrU
rpCUkP3V+8R0fi2qyb65CCHT4FsX0/oKCJoRSZkqDWWp8y6IMpyZdeh8XaxlN/uHYQjKtRbmEiQb
5NPc15dv3GUnU1kO2Q1BkwURGsEGPTvdaasiGWVBbMuvz2X4O7vnoTdod46OMq768JKvtZUardqw
XAuoEQWwhc177eIGrTg5rLDsDp1bSBotGfwVnexS9bxAkBwclmqOaxVGp4lxt5W2zVIF5tFcxoPa
yxiu8ttpE9jVz7PSI22N2yNDZd8D04xgeFauaC+SUoBz+td3/9YbRsa5odoufX5B2A92201HqBYS
69FeD8LbpH1c9H84tdMeb9bFZYFVKpGHETWuthEq1e8jhtgVVB4zGNxY2km85A2NRqcACnb9HYol
P1+kaeJhK4PvlGgUJKPeiphRZdZLmMJloIimHEefJbnkOex5fYVC5hOKbAoH9i4IDcMxcFVQcQ7O
NeR0o4qmr7yy41LIhDVeiYmtVjsTyXout7QZJG2vw9AA2hv0rpnLzVvUa7QF95soL5vbFG0P7cYJ
DF/kMfekj14HfDQkKsIM+SsU+wdtxiQErWIbgNT5MMn3tAhfTwcmO5CkdX9cYJ8l9/Wh8Tzszf0a
Z3QN8uWJKlTV7VYvROGzQ3dZQCqg8vO1sGJwOC/7QXKtroKsJWYAsn9dod6SOIVNYUhwpIFE06lK
502Ved+7+fAYLtV96bzCxTsTNs2Hbq6rCAKYtj7pHsx2t20QL597fDgHWJx5JBrEIdtUe1swhvWw
MSwlu93Zmvi3GSRDSSVg6L+5v//E79h4Wm4iRRTUlZ5yh3Q+nugmKlmBhT1/tt7nQjea9/7jXhMw
VmodxVUU9cz/ADWWqhmNQNctDlcwGXJSs0HrKaFNnJkK0zDnszK10q2/rnFlI3QbAAMT34prFDNY
YxINKdNxoHg2L3SQhpKKQHG/3GZMQuJlTeAKlPvIgTkqnKfcukGRAwgm14l47kqm+StkyQmQctSg
Qzfn5F+F6zsLJJZCaJx6gY1fBXcTIkcwmBHLEgjiMPQlqHOZDbAh6GTxyEW6EJqqK4jeAf7jPPER
5pAVMJ0N9hh1iM8AcuMgTkUFY8bY4s4Goq+FhSasgZeywxINBPXOW7z8bhKg3B8Zxzhy494JN06B
NbCvmQ8BHi9ZW1hlnFa6O572wCyrIHWAxT+msL2dez1A8qN51/hVKX3LHxVkQwHAAztULE6aDWH9
pIAZ6qBmiVB0D4nAFjOLiak10rIe7+FLMTSZdyVu74GPazOVNIPdqV7aHKcwxbdilFTDU6JT+8ys
bEqPAMiNYg5CBi/PKIvZ4oUXOe2KjPbrhY06V1tpHITXbXCfQ+RoC+qUihWOPVK2w5HHIvq6sG01
EOUeyp/ob1eEnPnzRlkc6hGcPg9fq+EdWBKzVH9O8asmdqTuNvbXyplCRAxbbiJs/OJWjNzOXnAq
zS/ME9AYtWF00b0zHWYiVbudclkmz8UJ8+m3OtKrNpZqGObWQV2SdYogOzrCaOXQyMSYNY0qKYM3
kfapMf2UHhkt9MoRfTCjdL0lfK+yC1W+Bq7QXfNB+sCOteId9y6H/ZzHBQVRA8n3szBUfcuBakje
Fu3B2tHEThsAJyYEZJoilU43ggoanxpc3icioDWLiJZ3N31y0ffcJ1O3FLLwMwc+vf1u+BLo1en9
5jkr3EbelzeshTEGNCvSeZ9YskPRYOyxyZ/3UIxF/vU+FZj/tbrXgGhRGWmCR8Lun28dBCHi7KWP
kiH2wtZZrTYnsxcOxDB3t00gHzNOWSv9J7cmYIpIURR6wRiuFKe+w6K86ClmZJXTaUUbVB5i3SyY
yJxviY9SsCBniuNELbZohgT/QbgPP5bAADrYtpMkGyHqIHSBwpovbHz+deYTPoCG0BWDWr2NUjka
1i3Oc10Emc8wX2179KJoA3r9H45iOFMgw3aLqg3funXuKznzV33nzhzrnmv1p3asGnI0ik3Gd0hJ
t9tYTZkQXor5yqF4CYozklY+u/hT6Ls1gjbOkn8RnhhONN+RPFF7dpNh86asdafotup0qsugwHMk
4ljldd/FxJ7sOkjS6M8ZgCy6zYQ+iZ6BvHrSUG4JT5+Gxe5OdAD/ha2PECbW2Fie5V9Z2mJ4Jxo9
g3J9YFzKhHE93YX6nbKQypvkD/sFgPXqMVThv2X8J1sSWV4qs/fp7NVPNjy5qvL1zOlhzXk1xi/d
yf5Lz2/C04yxmOXP1jgvhGDeJ7VVMAW8dVBI/o45t6mNbxnUu5lTjODbrm7tmmx7lVXxfEgNmiux
3j72QUTQviFR9G99M0Bgq2DOVGhO1LyUlJLaiwV7oFmvZiD8Y6WOPdB6ubKD95G5II7BTG+P7358
0/CbyO1qfQ7vbUS0Rfzwnjunz+7IGiL1u2YKEAvsdXvuYIRXfPbjcmmZJosnThM4ACom3wviAI7g
dp0ml52/5nak40TcFsjlQfJxSZZpAfUhCA6FRx368B9QTOvwNSxjmJjlGf8M54Mq+fNoYGtcpOfz
GQAaWl0Pft2RiTgKh3HYe81F8DVyI6uEjGHP+cpLLzZkdRuyHQ+1t25eSy0EsniK3slh7TxWMXIh
WvG94bXQt8diYZs15dLXmpk9809xF8X/d4JtBLSDJAhzGvhnuv4x4wzYJmEc8e2hIVDwbAm8tJWI
FLQuDDhcH38ZR6CcgP+2zujCCZID70npNKeDfrrsNh/1c1PCOJ7X7RjCd+Db+sISKbavSyinm8Dg
M0W+fSkdVtKh7/B/6BLu1sd0up06nREcztNqvqSLDumbsu4Qy5TBwxZi65pHYD7ys/7z12bK32Fl
7SCt5a92M/B+Iae/6xM65GK36fImI6cJjYuiDbbQQxG7laDbvSL53zhD6p0IaDAXTODnseO3MdwL
KBplZ8VoMHBF2DsysyLrUWx7mZxkCZcfLwKhuvN3O7V3Ju7jcHIs1ZQcICWxbxKZQedV80GUPzCj
PwmM+8ZgeeIYP9AvXxM0dZ4NLNG43TUSX6DLuedaDbH+Py+I4qczo4KeA5WpYkgw777teE40W5yx
9ajAgmBkt6UDBRWHAcWHgYsRONB84k+3tVsb/vxk+G98CiLydvR6cFqxupWJubvbC84b3Rq72Eyi
4omnjMFQrS1Kni6AfN5BRCsn1PmCMcdtnoulF331NMCoRYaTKMyutg8hMzfuuTytPhk5h5zhUPKj
Iq6jSlznqd22X3NM/i3xdtKQ1YbsuVNPfIi6kLkRJiLigsHZ1OqVyQZvc11Txn1M3oA7Zcdwi3LC
gV+4oPHaYKxBu1zlif6TVDIq1Ph1P7CqJ+cTxU02gh5WJD8r8ooWYOmWbaO8f6nZ8pblHgW0LB3N
OydfejLjoGfHwlOF7LvC+fMEyMHd0+MzsCUqrw32U9a4YQuRwEFPhnXAXYT7cJsyNVa9vjwzfSbi
giZu2djVV/sJtU5Ok7WQNcLFDDPqxG3H39MU5pk6Ha41q2Nl3IcjMkl+L3pYYyMScfcCXJmtkea+
FYvCtysEWcxO0lZ7GVAGU7FNII9ssX8zyggQPEfPfdeoDmZTOrNtTRdih5UfG4Zr/LltyYmc2vrc
NkwzcFhMKiajfYhiUXYOhArOrdE4yW5FAbFASWZHIyaHbPJpQl5Wf/M7zAUs3Cz1VLDRYfh1WsZV
Me2T/brrHiM71ds7R+pKbNx7T35By4flyvWP8t9V8V8cC4owyaUhtnLfLq0kJOZuyiiB3cNaX1B7
37jijCq6d+Np8WvgAnezvSuj5Bw9iPoBWwc/QmpDbYVNq/wtJgsdUnb/RPFrUJi78moJPic1zcSC
YFV2AlpYEe+QEroz4dD9ubfnKqTAn6MqNIBYhHNaPI+VXDlXvfMAELy+UGXOufgQrtrWVaX7SpHH
1MKu5UwAHv7kgR8EZF18CCZaeBeWjkXiX6HKmSapY0DWhuC/ah5E+5gty8IRR0MNqN77CaDgxA76
gyxG38M/6Q0620s+8iUnHYOrxQjYnBi8BDtD3zoD6QkQTCfEgZn4Jhcf9LU8ArcRSENjhV43oLU3
UnuC1craAzNoxY74xwkgcEVKR1G7MOlqlQCyE1drcLbmQVN1Bq7cQoHdPUsqbWnLd9BiKyd3XxxF
wgeLy45Vn70eA6Dr8ab7UFFCRcBzsGqqyLk6qbjCtpffCWGJdG2UuScFFJdS+s92BadNgyIykgjB
RlJhppFEyw24aes8UyZnmPeU+fgvXIfFHYuceo3K3i2xcR0uGCmn+5UgrcPbc9A/h+Fbqzftagvu
aYSJ4O/clvjStGcIhkmxuHkweXey8nldmbwVMsw9Ht7mUpV5Fve5X8yvGcLhV3VMk6kDFfPgFVAN
XSAkU5WD8yB6m1jhDwdjpwD3yILqaVYwWiQ0N8ZdFqE5gVC+fz5KiebN6J0Td9PCeVDRKOx+OlcC
Rog5D/hybnoTSHNRawMRUwt86zzA3R0YgPc9EfEwlSIfhXsyr1mXwTysscj2LGFakTdvSNQIC8pu
GAcFulZSrNsy5/mp/nTnoL5LlsL+EPtR4WrQlsfP8MnMQXJB2b5LReVkS1fr+yNw2NOw8YZ6jW+J
UnyfS+vP4WTLo1a9jtoIJUhucUowFtEtPWr+OpHtZFc1F+KxO5stpLf/o0xPBubHMwBHEvtNVEJ+
qMhVBiXJgstyVD28lYDWJ72/9eXos1OL32kfSD8ze9Q9nYtNLogOT+u87nveNoz+b9UZfwUS5PYR
ERpOE++IU/B51PCHtBqdMHPq+gesHbyWX1OJljDMYFLW2hbAS9O7yY4fuZ5HelJpVD9REBy6DZKO
3hbAOsB09ad7/qcGG7gCV71pWsOD20cV7/8NYQB3idu7gYX2QWBa7Ht0uSa23lLCJxoV2uU5XkBQ
1a+MDj5NSEyv6lLYCxf0K5Djqg3EIEHZGeJRoU5wvzlwj3/J6G88NAggFRCKuL96IevBC2h0g8cG
G59ZcFQR90pM9UgiGzWw3/7tctg9pyAxr2+1WFC7lbNR/qJhXp0Du5HhpGwDQIcRWO5DwPgjHeE+
5HkTkDBiZ2CfttKS2Deok/TVOT2VxhhaSkwHPiph51yUflhfwlRlAbfrVKmLyH2oTI+nCvGDMXco
eP5UPHLml0z3S5xwsiVkFm8A9JQZrTJKAQpOpuqw6H8Y1H/xZV/HGBgKvJw7QYAVROTahp6EYa5Z
BMiAFOGl4Epn6iulG9eX20asg+QZ9b+DRWuHneQxAKtcaNUCho+tNafeGC6J3p205V2FDNV/Trm2
zMe3e7OjHmw6MlbavuujA0pKQt0vQx1iyp57Op33yKscS2aFVZGr7VGm94h/6UwRiX2zX2jvRDxF
eofDdjBD428/RHy56mJyu2K+T2DPfNObd1igzwrz6mIyhuYv6fZrNVGNeKRrzdllKUrtf2q6Xx5k
LcX0hxjiIookJPJQa8Hgy+KQt2GE3LiMHUy8D4cJzyWsURBO0teme5aSlWTPPSCzsj0WbTPRalft
hvzB/xXJfNT7SazyhNyqIhu1GprB/9tRBZoqwfYUxxjfxblRB9tv33IrcdjAXvPTXs/BdCEAMO4b
KSSQDJ2yIkSlnDTdvKImVxDi4ZQrpZLxVHIeVoogctZrOuD8S7qKtpDN6a3gMWat0fJz1ejhR6Ba
B5CEEEJtnyELm5DBGlFg2wb7vUG7l/N3uaR1sZ4/3BTLen+fST9DJ8KBsEYteEoXhIZa2L1rwp49
hin+lkx7tPMOZGiaNDMxXm7WGksC/Zq1/nxPKevyd6aW1nkYheROJgDTy+x+RawZXBHqU7dMdsI+
mAQ3zlLN8jGKEtvV0OMGNJZxWIsKaZaA6x5uOEIo/ymMP/WyL3eTONqjy8pHDi5vuaDjXSYQO996
ZjgYdT3j77+ceCA4O64fjSnEzS0ahaHH0vtjrs3ucjKUnPwP+UaEdenpz0pieo0Id8vtWJbUPzgY
SSZDPhRVJBN4dHZMtQeOQmm54TInT7R8b5PeoG5s5/ZV9zMCsu4/Me0DZwZp4prn0HfU+3wuAGK3
e2F1032K1iAuQh714f+32rYHLU+biqijCumTZJq21JDRFqwEbxbeKgewMKjWQeSYa8M2x1POldfs
J+E95qcucjr5++Vh/C6yPbNE+PiXoNWf0kIfiD/XCZ6zo902dLyW31tHwvuqtR2E0wvRwSkeDKBc
LK6b8DA7T42WnMnNgySNSAD0fRlw5WH+lqIIqIx3zG6wYizpkHckkmUnAdeFlbgulmycH62fm6HX
zuapk/l+gWELhSshwQUQL1Nid07xDQvq4Gv6YRj2T1vIp2/uNuQ17oXBHNDFTKRgmxUjXYKVOcyl
B9GCAxVxkfMtkZKEDeZka+1R8kMktlxrDMiigvgeacqtO7YhfSf6ugtZqQdggKse694sWzezZngd
UcPEwoFtWyvRtCXRSXy2+dKKF2eNJ0mZ28j4KEPeEM4jo+/fmnZweshQ1qGXC484nrTdLKmudxq/
6Nj7uyvEqWimXzs6yRAfGlTuJiW9A87OzQciPPKUsaBN0SE4zJsXcdJcEtuiM7QA7X+h15qNcfCf
P7PWGZ/a0GIbPbk5/7KxsXrYAWKRDnWQdlY1jtf8rVglyP1ikB6foyx5Cf7w/CVFcANUsWMfQe72
Hhj4KDt4J1emlyWh/qoy0K2xkrFEqRWziQHEms2O/IXSPm9RpQP9a2snX8odLdfn7u3+hYYzRoGD
0N9oFhxFwaT0e4K+iQgnIqVpP3zM5VudWvtkUR2FYcvkW0277pVS+mvVPSLImzQHjwqrDdC5ULu/
UWWxPgAgOB+ui3oJ3/D8peUPbxWBnK2nWlE99GWcoGMJfOX+N1K0CsIAZSN82eFOHCOQNIy8qLI2
reea1Ny7/4AEJoFTFMdypGA+u87MDUH5emOZg5Z/7/fW6n19FdQgYnJxxOQknoUILGXNr1/Nbs7A
uvdXUl0XBXCMrw5fI0XOdxu9iNLoXaNqaSM5iLqihBcmIb6xln0A1+hTzU1GcnOFGaFyvBfRvUay
hnIrDvnlXcAgQ/8p0gbsi20r1rQqLy04rWHdehCj0HTvNDcL1yx0VE4dErCGr/lX1irvCqROkMD4
OpKTZ5P80Wnnuuhoe3e2qjzzTxmPR53o7Pg/JGVFZYLaMR030AzSTTPSrLqd1lnwks1Q8bfsu6Kc
2VyFgvU/hmNQVVxMqwLqpGk7SlRO41G+3n6VRXvqcUgZn7/E/nfIas9baLHchHVbJjj2c3Ro7h9t
4p0d6l8kLdYbAHRQh+k+a00TUID7a0ygk0u9r0GDOAA2yAFvrkNc6nWbJz6lnnrUEAfYmdJKaR4n
8/CzGGAAGJMNDEGVrgCGldQMky/nV3m5ovdIgxGsYQ9wmU1y7Zk4A31S9BIO9KBCFuf58FuO6o/D
R80N8j0ph/TlgmLtZB5M0dJVM0mjxhcVWsQn9YvHYb0qc4geMnfnj/SjY6L1XJgPyyvxE+yLLMiK
33Wz9XYiNcO8hK9HyIMfCtSdWm2ZTLilBve3oK/dqHqozJtZ1OvrVd5sJ6uX+DN2Rt1lQnuhZyCY
AiCdTXqKo0y0hbSS9VVq7avtxSj711h79MTrTPp0OvXizlTiVHk0WVTQMunnIbBvIP9K6gVpVJOJ
cPXquXUAPbJu5Q4AbXILJ/cp1vZNeVD3tPOvjgzu6C8bV785urER1x06itWQoMzokOPhZJFdZeAS
RROMcPUWecBTeUzQdmo6+7KlEsm1TtivewBEClV44HJCneOayj6purjnPBe79SbAUyXcok6JZP/D
geCd9HhQcsyihqvkfEi0D2ao8HaxDWlisEo6o9dlDMkosAe4biaYctI59afARPJfwQow2p1G9dEh
RxZNOoNCs4bPmLfqLEJ7UhcKA7S1p72YG51mkTRZnnjl6TsGwb8Sb5shYLVUXahI8uKA9pTBZDkY
Yq1wuiOCjhFojcnN2l/PT6IzD+wc3Qe4cpKvpgc/gjIpBk34f11JRxajpN4kFN8awvfFJivyF4Zx
JYUFDDM0Zb5UM7n5v1MpzaiqYJHsc3g3EfnPWpi16e1IA1W2FyTY5ALgaqggU2k7FxLTKg4y9YdQ
59qYlr7Fn85Eli6FbPw6NA6OVabpDBWyIebMqEhD1pNsQ4Uj/YSrnkowc3OgcK3uMSV7QvbvE8Vi
duUw25o3RSLfB5PSQo9ZXB2SqzVNNBs7jTWajOdAJXy4PHlMnfZEnBevv0IZmQPCADN+RbjQGjgC
bzT9NabvsofycDIOlQDWiEXsp8ChtHajE8GEPm2MYK+WyhMfFeg3d7eicQrbZv+8pbcGy+7qcCqT
hDdFNAbYQy01A+Olfg8xlUgap8xTQBBCfisab3iw91HoQUwbKXHegmtszn/fhRMQzg+eQUnJRFrR
D5KtoQbfwg4b6AAcL0VU2gARK+/JUtDc+Tuv/y0guoeaZPnaviACafdQlCmLNN6o5OWaWeyoUuj3
FQvQVf2DMusTWnHiZx+qgwCpet+XLxyzs7NdThALjYh2NpKLTGr9nG86f34jQMjPnia61ekpJ4xW
BQptvz4UeCx30ELWn0GBJOs+Fwsng0Oj9AjEO4SarcRqC53ciY2IF10QDN97UR78rlDsfVJDB4VH
aSi5j1uHshlKDkr1jMvasLlMMGiqNkcaNjOzB2WBfCkgcrRqX67cgagzprNrv0GrBdrLuH8i2y7Q
d59KmRsnZh+dcGg0SfuZRW5sjkYZ+fT47tTu2iFsHPPmNROHknybVMZMR2R2S97czulHWJ1x0cn2
Xbqt5iWZ4thtyL0WjIwMWnbhPWyHGcrvJE2y+bXykvbkO5Dk6p8CQfFtU5fKOxYuvYm1eNAfl3mS
YhjWfX3KmWMpSjBMiDT2rBRVi/ygsQhwtH+Wt6HFQG/xLUnnU8XbUedVaZ22B4puGniB8aqxl7EF
51n/m0SO0iMg73hbfJ5rjoNGQmyz9kLWUaQdmtxTiCf+yLbiGtXRW0XjhFX48UVHoc9FKjPKD6Xc
vu4zkXBiQyKuKTG+GlgAL9l3PFl0yicZ7j0mBYsqTx6DjyZY5QLqs5yWKdi7Ighl3PzjYICWdsGG
MWErGIR8t2fNd8fGEcXYN+zzwmAPbFoOcxSC6HFWYhyon4ZVeY47q87Xrca9ZUol98oO1IUP2tJZ
LyIIrSe2caA+opvVpfiWmx6sH//J5Ls+OpbZc5LwnV7EjvsZkykPDeD3NCitx7iH/4ygPslvyds2
arKsYnw0x+uALNq01ULPiGJcQEJTAha/argnizeqR5tnkw+oQIbl6ViNoVMH2A791ltd4X4OYrLM
SJWZsywZVp91rjfh9nuDpQjf4uuw7+ytGVETSnrEstIDP6wJpB2Oh5ocAmtom5JQqC1wKGrnbc2y
Mcp0su2jlv3/O6cWXlc8U+AS+mqeIav/EZC+aSDcOerwJ3hAv9P4sTeR5bgtCYXtFeYiVCAPjw4K
Y3AKGViJwKdq/KUa8st5Dpspz3gnKL5Rf6ZvxswppeE9If33zyurchGFmIBfG+R3InLKUeYmJ0uw
qXw8zO6+Rq1+zEJoAQkcveskEOAd3xBT196jbLOnetYnJthD/SYoYPIwKAYFS6xnGTn2Pag0ak5+
XA2id58uZBZhy5dIMbcDZTkt2MieutLWBu6BlRkascrprouY4270rzITPQMoDx0WVDZh2tzsY1l4
wwpI8MUI1vrkJUCiMAoQB5+olZNme70vomzGtG4f6m4UqoQjm6ZpTTl0eI+6SlzusH0AvlYTVSts
dtiQWTTMtsUiB/lYDm5SbTfoS4YFm3uRbYkBGEUqvosYNeiN8SslqBIH4QwQZW4kePXBcVsRrEN+
k/dWRof86KBLQSFDkZXX+LZ3rxgJ/vtQJyUkff0L92aPzqIBtsXIrq+T7pqqHqwOvlk7l+KMR2zZ
wnmYGbOnwvQddQwIVivFCGKYJTE2AU8rza3Hf3OMbsWnfyBlMkBVXpPqgsoVA5BH305Euyg4DTzf
y17jU3gJUcjG27oSEYJaxMr7WYPq7+4N94i6ZFXnGdFeTOBy+787HGMxkxb0YJzbywEbr1BtHNV1
PVAEaL/28GVbiwvYmfLgCyP7XKLlRiHW4cxoulTPDFYFDX5UAVwf4ebTuuyUTjNIBmF+hHsd9GMV
1AwZR8VEtMNqQ7KO5HfkjjeeHkOQWrUwxkuQsnescYebKEioa4EQjRq258UkWWUL48CCfmWhluU/
F0+c8cR69NooU+FOT7Z4GQB/bir//we0Ji2pb76BdAREKwYuPiveX0MYwEvjk2Vln+GFPYH6kUh2
lpIU9fwRhmISFymKfF6wXvow3Tz6R2wmupIn3YjbvX1OR+gTYxxzg0dxgnYAtgvylcWCaZlcvf9h
9kDwfqVoZM66ZeGcJ19ZZDMi9tOYc0J4pjm4h0nOOAb9Vpojeeb3lfk+wsGV2ErbPLXkphxYMI4O
R6fH/9/Ul2/wubacpczD1M741tJipDo+4ZXYoJHnmSd6PbYggpZr92secxxRwKgY2GFCzfYFrGGk
cHMQIzYPGiUKxgMaNKbafM+wT47dz3R2O7y+BEp7qjW0lOt+GG819gjHcD5shCYop2bY67l730im
tCAKjQ6x1fbOt+oUBSSUCn39p66oarnCwAzpFbN2p6N9ajtGu+8P4kd80dg7YQIcDjz+i6h7YIyn
QagD7RnA4MeHOys3PpIj8CZydbvF4ZWXaIoZUTYLTOadveSL/tr5TKYLWBgEU2rWCBQZb7Umko6f
k9gFlngRlTiwGVhsXs0Ex2DxbaPx3pR3Y0IGZh6FMitLa/IVDszc9MEcQL8Tu4d7fWcwbLVy68rf
Hs2VZvZB0i1DiY3RoQ+ssBIdXi9NhhxtKoNUs4iF5S66C2LuOgkukkARDywbfzLw6ikVj10fF2Gr
ebvzltG5utZm1cRP70gM0xr5KPy8lcnD3OkYmUvCRgMsaUjxnHziMEgS1AWeHyGRUI+YeoTTz89u
fDVN/BV5DnlNuPow69iyBeoZXhoZQe9NiTh1RogCIgkyeb4j6I0gqy3cKNlW91pDeajc7zJzT7fS
tLGAIk1/pmOfMDw5s/z9rB8JZlEWlt/FM+N5vjC9/Xp1yRd7FY+467bmWCIxfd9A/vxv4mp0ZHQs
zNsTRG8emKbd210aLaRH1uuXkNRXY3aXuLLs/k6wIGAFzSjGGAIEjVMrZ5SdabHOt9E3Q58Qt6Zn
EWAiRZxS/YvAkAxUIVT0JBsoAbCZFw/DcqizHCHIpioT8FUDavxdf1ft0fzQWxQyFbLBQl42djZ6
4G3eoXUy8q4AM5v4nXMFTwXr1x8YrAQMhflNAENx2zICjLOqbD92oo4NuGTKQCE5arfYfP+NfbWz
NHKW7+WJp/JxM1NFSdU2NIzFcDTUheZ7WUK3rHlJyR3FdqnRC+tHuzI/mRJk/+tYxXetpyoiSm0y
t0raceMJ1oM0R94mzMJAHOUdgohyM76veq9fT4VVZFvhInN7R+MU0QIPrA/1fWiIK2//2PRb7FWo
uRdnWERc/nKaCUezuUy0MQ38t7PxE3t4ymgAVHOr4i8w5XWnK6Jypodm610UHA6N6VBAKcBhHT1t
vkezg9nyBKe18giFS5uA3S2MuhjkjnUqhr14XrQ1d+Qfjgo0NVP7UNRME9owt7t0/vc5waKhE4+x
EDnv/YBtMAmLxKPLiwaLX6WbsfT5ISiuBUQv+RqfyRvafOTUdRho/R2pcih6qML3CbbxoOxWZ+EO
bIEmkOIdNxRdTjhI03/Hr4KBVYocTu/PPiCe8aJsBwPwY378B/gRekW67AQ/jGRIeXwWltou8+gU
zk2XSw7KS0t+NdOuAHDmgtWzAj+dE1qrxfUWfEjH8ax8IVUyfY9neeF9832B39eZfXTG094wqVPU
MxFHt9hg8qOrNjoa7csmOlQR58VEqsbmZe5KPOziGYOxyLRqWsTnAajuBKO+bfMcabGCc9JfPEPF
5Iu5gj/jvkGIQoKDQorbXIOgO2oQaHs8t7nXeIvrs6loQoSMNXNzvceZzClIiMCeHI6AqAx12LUd
Fobyo5e856mHq3Ni0wSpabz+pS1lokqiNC0C9PZVkRFW2ralwb1xscK6SbGvOleWTgP9o5YGcjyK
kFMwQ+wc9TduaHQVJPvqSB1r1C1CVMtk2ox6w7jtrmrgQ6uZ4bxQGgW1DZTdgVlmuhksreRC+YM3
f/wZ/WrQeZDNEdrNlaMg4s5fvaOS50ABfemacWBezX7o/gornPFh2wX9r514WnwgZYTnGcFenCZn
fVbYLMC2zXFuPo9ucgAOaPUwWgt5zCF0srigCN6JaVqYcEjukF0HWz9UAAr/Tm4fW4omvL3K6u09
HuRb5rOvw9yhRatO6mRib5qS5Mx3ifnl1ckHkTfEnmt1jtRDIm736EKlaa9LWi2d/jr/80uhZCKe
GCRO9MinarR72V4ZEarE/ALSjVPn7vO+EgK+vGCC5cKTRbd90CC/uRdhn8Qj4eZg0JJGdOXYxFhu
VoqGpFxBE2uf72m0M0P7UDMQy321+/PzptA9ZOZRgtvSQjwfTb5P4zD2fVr8uPQEI0JaYqoJhfCW
zIwAlouq0tVrcWrtA3H2lCBZkNmlB2KOymaGGv8nNkl5X2JDQjTIeeZwQk6I9+QcqNtXQINAQTXH
viSlVUM+TOHk3CPeFexpck29hoQCAOp9ZllxPnYRkrCQ9o3eOQpj63HC+g29ZVeI1v+zAc1IymKh
12RVPue8jXREWbazPx7WXPwxa4R8AHZdQscRch2MUrjhzQ6fHiwKasMw0MQmBGNEPdY+Pai7CpIj
PWQf2Tct0DhORd2TrrgD0f5/PYiO+YAerUYFijuET5NGiU2V4uvjfkaEljybGZCoQsZ2kgygXuwg
lEkmix6rCf1gbNGTj8Cf0235h32NiKdzdWGDacllQQk8zBMno4Hj2W560fHec4BCPnqsHSePwQR9
IwaVh1gUxoCvZgu7K/9RfH3S2ZHHx0Lc+ZA1ywRzT0p97Bc8b7ONi6me9tXIRS82CwlH3WO3cCRn
UIZ2dwRPizm2W4SdUnbm1Am8oVLhfs+CPrEP89R5nLSeqkz2Iv5OFnunccL/B6FO4C20JGxmjBjc
QIdmzEKaGV83pgl/9/ikFIbcYRe9fjNcXpnDayA2Yk07fwNWnSZ/rtcnOA6SnhZ0/rMCg15N43dv
O4m7AIq5RK3JvghdibCtOwFke8M00XQEEt3+RjhzsLeCaacGLcyX8aj6ntsYe7u0V9LVctjockA9
LWKyukLRxVkVW9IA4tGkpkKIRrtznsOfRWaW9IKuJEdDDF3Lbay8UPpuSC7j7Bq4qa9AdRTFs6N0
aQqAt4NaMWM5YSxd7EWBqbO7g3udpKLCW4yK9y8nnqWJ9RdMvwSgFkzAdmGM2olIIgFsmWrmtN9+
iF1vRV5EGQpAELxb+nPIH/j+ZO0NpXPUwHWB/JrHs1MfGG7Ds4jm4L66mk1/r5FY2giEHe8Z74uK
xCyz9WtYSfYUO9J6OOq6VFZ3UflFb+Cy36uK36Gy6xF7H1Xb0hBud0CjsW5+GPTANwwBScA79R5K
yA8fb0ubdG2dMmqkEYY8JRaR8WQAjqa/40XA1sxvHI+Fv7mW2JBtF2wzRHuVWlxKuSYj6tBcEbJ8
7mdV25fBpBTX4Z0B9iHdhygIoLpL0P0j2yriXO//b0TTHdhq2Ra2/MoahITPOASZAHXTh734+cnf
Nt9SGqF1c6VkNSFvfk+GYcxwjFHZA4Fewvstknf1XYQH2e62pMPryF5v7hn0gu65GTlyI6xOtX0V
JzPux9koiaALp+S0ibPckOpJGJ+sDpXFgdJCdbGXDHw/9+uvZbJO+12JzINR0lDy5JDTIZdA+i4F
xVSUMqGiY7b1Yc+DmLCPX6RHebDsZ9YODO7NeyzA7na9rRwa9sHKZ9kA0qFxTJC9ulZHHojmGNk4
HYUMzAL1HeiuMYcQbZ5/svgHW+ImnqF1+LbucFFpGDV6oXUr4KDZyINMrR4kIxjlF/vznTs9R5yW
9D8IfTl+edS99Ox1Q/IhSScl1ilnQBgzcXlAJwrkjJ82/0s+Rj8pRCvFp3WNvh5qtQ0b9HuKmQzl
5i+hwa7cViCq5NaaZxapT8jRHyoWcYyksVkpgz/+fEoLupIct5GJOldsMgse3BdoxiORp3hffzux
ONMhrhlpfZlDPOsO34MPMRX4tuFI28lTvtfVrRMlEOdcSWV6tdGdakiinymMhhXEV7Bsdz4qo/m8
Hnw+dP6hszeQHUj81RUgeSn0UZF1/dj2pnOM5uzQpSvmoRf6RpzMqtCgkr8joC93NrPoPCq9GPT4
48cCSv1ao9T7N2/1Delycz9+2KWZZpkfXDa2r+KeadN/JXCFJnw35cyJ9BBHjadZGHx0ExdRNvEi
Ig1P0uHJE1HFvAKdOEx+P5bWbG34P8Jc6PgCSBFl4nN4xWssmvNxNXps3yYI06vsNNgo+kc/gsZ/
5RuxICszXaXmXM37vDG6aXaV/eAfrJ4X5eJdZ6dIJyx3GBj3iMILhtedRmE2FBmaP3yPxsxckkR1
p4xKP8Wh9jSoIbPA/eq/ZKFka3SOhfj8ntg4+lEdUltOt/sQ+IM868Kucvm+Rhp6jkmNgXVb/tCv
6iEhyUYvH1RqHYv/iD3jy1ko+HBhF+ItbzyxaGmFV9RnoiJmQse+Pe4Jb7jXOYulXUc3JK4MNZHA
KmGo/1l6coW4Tin+1c1XxS7kKTNdw5qZXZvtXnGBI9ygTOaN2/eX/K9N3cHlZaR1EFzvDuUlHYET
3UKvABozgCHdzTd7GBE+Q7e01UAiLIqlEuRnOf/Z/QN8+fmXJVyXDqsxKzuqu/RE2WAxo8tr9kom
K+2XOSCBWoYNQ1I8fdV4poJ569sg2Z0rJHiQo9G60VPdAlcg9e6lNY/ArzGzpvRFjvo0zUvHKqkM
TOxy4whU3dzQ5ICDD9qGjYwOpW7zSOOqH35pkuCcxVZaNaC/U1tWxa0Hc/ugc3w2a0CiNZCLdZu5
KIgJ0zFwlQfRdF9KW1yxspLErIdDzZGOlHB00ia6mSA/WWsJ8CfZYrUmokNrKsdR2x0tCk6pcgCw
ano2VE0kr/j3REmnH1McHSzpc7Aj0rHtYdHp+wDrU5n2rlBrPVzp6/ezoILTlQwvn1O1ZCq7+RlW
6e878qXQ2S26KFbJJXTcJ0peu3g2S/r4rUNIxxEn9HfaB4dqbCwWjFcwJVwZwhvHAZL6NI6Zgx2o
b1Dbx4W8cZrAL5cbxpDJWT5xHZRNchgmCmM6E+WXoX+vgLCbDXJI95kPbpho8EN8/z3e8BFdRZYY
zbpugBHHS57LgXKup0Jrw1ZeEmVT2YSF3pWlZEgz9o4YNb/KIC6drLRo8phnsutZQOKBUlKRD7aK
2FEp8E+sMmmTCrfftayiG+5FZYFVmapo5iFO/i49P7vU1H6LLfRMDavKZX6YO19QrCvarwiE2SRr
dynNVaIyL+/r8dNypAYpeQHhby/CDho70CwtoHcK4BISLB0gwXWqLVm0mfXntOrQmSpZlOqWEcWA
1/GJ7WULHDGjJE3H8adUj1wTKjqhucQc/7tLlCU7KIcxCnof+apVIXr5usJZpODlrYxgRohz+e8S
uQZ3ddvWD5yaMKRknxtr0uxO7ucZoqK4BOdMVVnvutDfClvMN6OUqpY2Hl56c7RnQXl0GKyxFMA9
ncCQ94iK+YGBwRY6IQYZyh8HfGDrwNwQz5MhyRQnKhupQU2K0XT3K2kvztAc8j8ZNKGPGHFPJnhv
AxUOxK6McptiflcnBUxEiWgi1D48yNRmBRFP9gZXzthnjX/VqVGse907HFrPRu7Z7vGd7EB91Ond
Hynehs8D1UjRJ6BkbZh/b/J2ZbNAn/yswvbLiCZ7AXfRE3OlWHSIKEs67SUDAodmcdyPawJfT+eC
FKquME3llOuHGM+zn+xrzYok5NXjN6xYf3SzpFPfCZaDWpKPGGErJTF/IJhcA8PW/QCNNFMbxTLp
Lgxkhr/Kv+Jh6Yxtd1OjYHBNh8Sw8HgFgFzeGz9Y78Y/d8tqjGhR8iiqYsspLDL9iBzn7ArpHBA1
5uFKebH4AalWSgTlgWvhP2kMdXNb79SAlvjaV0pEDTNynpYV7ZZtB1dCRG10RdWXUVMWDkc0hDSF
wxdsR3VARbvPophx1TOiMPgDFo1qmXP8vxPh8lLyrmsq6m12n9GhFx+5b9gc7bv9pm96xCCT5emm
10ecQKcurY+kH8YV6Iz9dT6MlMYoHz4DlToF3aru6Z1tpYKdxfO3UILuagvoqPBpT4HF/l/Y7t2v
Acle10iGJUB2jft0axgBa5I93CPJ1BZhPW2hUL5U12Z1+48MOzW6WDjnXymRPMnts8A5x4wFCK52
fSPeJUV+EI5WSY16rxl9UuQDtA4gNiX99CVNRpGXpwoO9JIFEY29QNtc1JY/rDKAg3NYtlCA7CRR
rHwuQHqH+5EMzDslVjlAkFSf2/BuY7kP2rb09rrFCxqxKuTlOLQsvvP5WqL7kxKBAyDhOpCcRJyF
eutj3yROvQ/8iLAieujC7XDf5Jf7lDqUqjSilPglHSwb5AgeYEkilghhIK0fUqP+m/exDTgsntIs
nv307MJXgpn8fkzQcq+I3RPnzp8eDksZrjQWip3hXKTMWPWJ/9JXjeHVeM7xnhqc/2I8t8LRIOVt
yJyeiWXroz8lXyV63NN1QTtL7c4BunVxfLUrjKqFt3HqzES9G2ZqaF1atmQ1E2AsXZQOLjBiHZgO
BfcyUyxJochz3loVytOvP6N+HFjYsHL1umqQE4vsIRJvom4CJMVkbFyZdDogCaF1d45h5n/92I+b
IGEbJiqKzPIi72/hEuXe6MztT3btMJi+4ai3s6mPtZ6dL1i5MeSkNTgkgNwkx6I3mfUAZUj6JrE2
lTrLY2FZCJWTsIaiXyVGseE6p2S2t3290S3oBlvv3WzFSiShwCq6Cq9woFYCO7Xdk64WDk99llWK
jgc5+8m6jGhP4pRwK1IPAe6pCWVZQ+YMOKPt4EXE4jnsJaOgMc1k8A1c1lBX1j4RrYAqr4vjf13N
aLI6kQphtlYTL7N5AEAdByvwpmbWbt1n0Kag7AkFL4guDvG2RYzGxUVQRt1pvSYyKUq/c/XbQ1u1
dwYk9yNB60ztoSjNj5bc5s28+eBpwIbiUwZhqsP7l9Nocsb9JHW8H2kwYIwuIhgQff7F7nm6Mlvl
AoWuX/ohlRiVHyA7UrYWBpXfHJtNn81JfSMzo4DHshdc8xRC6/LH0qaU8tov5zE60IwqJHe3f1go
n6SHb6cwG+HcX0c6PeffJOBh6Z6tj2RaYqqxIizVMne7M4ooyvUyev035+oyprzM0gsHG0tmMiei
mba2uFXsjh1363xUzedEP3QSG1a6drWoHIJwv/4+AHa2jo+fnneTU4e0GIu7gbZRY2fiSZeynYzk
w4PLRQkM4cRt2Wq+qdVMhrW6XMW1MAoPmdKqMms0BiWcZMWyRA8utxvPHnXyEVR704UIxJLQGtDd
GpidIFDC58qruOR6lApvuJhUf/NAUP7aUs9gIy4BK2aiOxzn94HcHp0jK0EaD9q0n+jIeD1an/cg
vdWI5R7QRaV/YVjnU/BxeE7W+t9fCnxdCGlPJLfaAV1xgZcC/1ocN8Yi69ZF3T64Mw+5NWAgkAYy
gA1kaLzNDl+JeR8aN7UwjAQ+zEAgGlwXF9rxJoYPwLFluyfSzwMtDzw3owXGPFQOA81BRfXi/Fqg
fVSpOwsnTF6LvIl/XTUCID5jjn96GM7UMkcYa4fIfMFydZXnkHIRdeNp+sSKiMAh3vJ/iSevwhpi
JjcWkj84j3Z6jRTt2FD4B12UNV/EEfxbLKj9E+D6HfXU7nuy9nrRJu2vBCnp7uBIVrIN4xq9Gprl
AzNfkqsrkNPoZAHK614Wcu3XGXgyfhxp2ajMK3Ry68uGuW5kY+ShXmb0Igp/rLoEMv4K+t23/l0f
YB1txJDBKZIN+wQcq8H0gtNnquKOB1DprN1mHs7/ig8P9Qy+9Di3SnqywjYJ13PGJeFNoZjQIhEl
yZUSKrtSaAZfYRpGJJawVOzRNfxy9YIl8dPqjUhoOXQLHNo4ZfQ0x0RiuPn6Yd9GfxNrWCxnevra
1pzwns4no7qBugUBPaqyeJzm8ycazh4NIDwM2A4vInzNUpCRNGcRnh5TKcsCqbJdAu8dfwV3vPPy
+HuoAi26XBjuk4tRxQby2Rt5D22/kXJWfKcD9tRasfPq1Si1pCi55/E6yHQr5kKedo5Xyrkno0Z7
Z3OwcOWQ/La0+5NZl7yNOPfzSra7a9NHTI8ILukGWQZZpJGB8vU+p4TD4g9g4aAMjMhRWimETTcw
unnyZmiIgyMvJNv5HrnHEO7ucgzO/qrxU0MpRUVtPPrDbuPjp1D66/L1dDmcrzURFdnsckrk18v0
yBbUDYStVtTyFEjz9Vk+5PPx159jGbDziue0JXhetSwUwCR5esluVU1+xstdESAaKoko14RQ+OK9
iG2CbCwpiXDrSaceamZ1Upb1bdNgxyCG/A4oakv1ieuLpkDotcUnk50MBpZjl6TcKe9mHDoqdVie
I22bt/gZcfHKajojw+aojW9Pis8Xk9hzWywFMfvBXbCuLomptPjlrqE8AB8nRnG+C3K1iWtPcr36
SLQb8+7RLcxswFkFkzouXBY2dGWPwIxOX3KjC0IstWgeT5YOvc7KMah4HmMVQ4oJAIfSzc2qYNp4
uHHn1kCXCPTBnhjgAPZV226ZWL8m7IZb74SUubjfGoswiPRFecxOxODOycK5bACjSoR/vThusX7O
3TEG9mJS9+DAWCFXPVLZ9/ajg8FTIbtp4IvxDtoF/95jIOhKiyYuQd4hsA3uf15XtOTYiC2WgGkn
KjCLYQ3ZtPP8svnabfPtPhCfID5ErDGh8a+wOxIy0va+dusKaKddNRwzLDJFs1OQxYNzdJc8AjXr
yiyF7iYtYAOLipF5sZFR8fTFe1cD4aYG2Y/jR/92l7XnmkEQh5nJhIjsgoVVAxX1JzUO+nNO+1MM
g8Grx2u1FwyYk3dY3IesMbzf8R1t0VtLuqzyB+5rCp+Yl2BacPBfnG3UGQXgnSKHo+FH2gaWA51y
PA6v1nrECeDizv6Lm/U+Ok0LPCMIWR1yH9z4XuOkT+AD/chavH/DX0hta3jwI1bOBiZhWtc6RW72
/IVArrxMGd0utbrqg327aWzBs0a2IbhKb3mK4ERBubMzEk6WGQ7zQN+L6g9Iyz8vCZ2mHoV1qfDd
h5KX+KhcQ4BNXI3jLQRDyXRlUPSAd00WlKGdHtfQMqRltkruZgIGQ1gJUK6mWUyfRRwdB064Xwnv
CU6u80kDfs7xqqRRC/4lr01xbse876wZlNiI35k3zfuuN23UUoO8tSYEACuavkuPqg9rVj24enLx
dG6ajorwDFWIueV4vwtZ9erXyjMQG4bwMESxXyVRk7fGksXuBXnK+aj6iZSyRZmih4u24HqrHXuN
lJVEZFE605K9oqkWdr7u5L2QTllx9PrqZAyEmLFNj7FR9EgIp1aGMcJfVmJzsz+iPGFdXXAQFY2/
/qKGMXqo/WHLCZblXmDkczbLZrB85gjcx0ACzr/Qf8j1DYPd15Av7kI5oQlgYyXiDCSzJrQE2rtt
ZJzuT1o5OAVOdT21VPTfyT4lpLkOcjiHLXRC00r5ep8az7/mZ7wq+sEuLvzWRStF/DnLpij4x9XU
8mur1NBFo1NHuIzHUvX6WCwOU4IugHE597soxcIJKnXsGc2gaguwaiNUQ6kpFeymiGb5fAlFHwHg
DlFKuh8cJjh4ZS6RVxqyFkHljA08FH+xnSAcooS0K+OwT+097BoMtBxmEjjzMvb13mfkMoCG9Cgk
vJ5j1oPrQei7qDMoG5LorrU30xf9LCrdro5tgO51+DT2wbfEiF+wq4cFO8QGpv4b1KdkMdAhdAYE
f6/q9Nj04lgd4+8z+hIyVDMDQSX6HM0XZAyajLNwkj+569WaTuMoN3jSetJFZUlDQcYmvk11+lxn
ONVG/6S0IMGAyLS675obhVG3LE35b5u8/2Osd/XFYRMcLOOpMOcX8g9z5A2hv3YPZ8WHvwlOwE5B
4gtb9AIKzZfyi+VPQILJB3eY9pfel+ad+nqWJU4X97kHHbUcS5zKeiZRXoLRwC3WYY0uhx3LhVx6
abIhhzTk8R2kmLU40K7V5c+Z0TU29n1lD3gSh4BWOpBhsifTbmNutDNOr9mu3X7G2n04dhWJFsPN
5itGSHsURR0RyYTcVDdKzMIUKscO7pLgrkKb7BpLG0j4F5E8BdTMh0qg6N8Q/EfKsVU334T6kcRO
T0VRYNMa5FJtHZ/Ls2bvXaP/zprDZhJC1X+RnAUj/KFAijFD1puqc7hYdaFNR3o0G0gk4gJGEPEE
7oTVZl+pRPHOTHMl8iVXOVTn34+Lit5f6AuThpMmQU6SvY5phpznltdjPp5BCRV7W+Lfy9HObh6A
FkqGoTfKaAUyfY8do/DU1dL7MJlpSDVs8N8wdD+Tv+jG7kFRxTXU5SP9upcuEj/mfgT5sn52AgZr
XLn1ALzd8IQ+qMF1YfY2JrBiYv+5Gx4td/8WeGd+jmcZNT6pvquraiyyesAiI2at7mDCP8M0C5um
5OnOyM4jk8FpWv89zsb7tDgtwSt7vhNQZv+6UBwclfzpDHmad9/uzVFBuv3zjLdoEgl2WNCOp411
1cFbDf19HbVyd9PCT/Of/qN8fpEFFaxyXKO7y1fN2HnBP+Ook68yF3P7AgmdX08TPr30NRtaQ17U
qbYOtFRjt6r/V5rffBLyNfg/zghZBy9qY6C3r5kuujDf/3tXMPEl/V3wr7kvH0UeNjyJUDwzE24w
9HvbwCe/Yqe3/F6sKQ5+hLQelXFz82NDg1XXpiRjFzt+imMedLcHvpFz0qa9fJAm/PXMDKKr4dLR
ncuzzNDJaeSluxL6+7bpsftGNtmkPLl8mP1kyZ0XoCVzvMaPz23oltgo8+LWRIKTFOXTP8Z8Ilwf
JXp6OBCTVSzTPphAVTpM91mz179dEV/+J9dKflFRZ76OHZLf7+9NKsDSwK/EhM1M5qAnlgc2EI/J
p18O/4C+O2UgrZ8HbuMqUGUq3/vOkGj5k9PIXRYu5dKx9+ZBjoszott5110pscYL+lP9Cp8Sewcg
6iiuWD/Qk+KQzsQiV2gXhArVnB054QcvA3EJzwgIOLG3/cyoiXOx6YGiSssnf6/1NgN9Uj/NZmL9
n2/6ZbMRDI+JRaLZzx8LQ74QOPrOAX9k6G7MYrbMdWr9V+iXMyV5MtpuN3TMvV6SwRp4fOKl7Gha
gQWzo+u5GFQjUG7NlDDUvWSP6fHqdQ/dD/gyWiUksX6V6KcJEm+DwdT8tZ8Y+v4uWPy0bTzyq1ca
FCeZMHtJ1p9Y/o7QT4KjwA+fSXyTj9wdsq5w8FEC7MGDI+AjhP/9sbuKtQH4waZ+UlNr7pMJ+bDt
oX7Z4Ox2J1fN8JOXoSn6/dUxYZpcyZdtPuYUGH23Gj2sdnF10tRU6w9fO2z7Ft0etZKdSS3LLNEw
dusX/AK0ppwX3dnbbl5NG2mC5X3gdJWEcOgTwbr0KCZ8njw2Pd5vjqqz+FJkpeW+IxDMKeo1HYKw
wAajFEcmkXtRpJKSuRLcjxWI2LbFeJtDAksA/F1BYRTWs8qIUYBVpoEhVt0awtxVlwcleewnRBnF
+NI7vSqKsKqrXhKvr0eeXcbnNQTAccVWZLzNdFNS5NgpTUb3znRjC2r6OLp1xBcnYtb24oEuU3hJ
/Fnrzz8RRI0V8t+zYV/+kCHXwr9Cgj5VpN7knr/kNr9yqTxTPnEuPpReNnSe6jLQO4x+pn3QLkvr
AUHntaH3u0yZhWyeV+ixxoz0xmj8IjVAol0RcYuZd94R5BbhGehcCIdN/QbgS6j4jyPbow7ejM/v
5qGrgWw749NtgdhNr6tT4lT8TbVOLn9NyK6SuhPYJ1/ralHKdJrvmZ1vHnjfXkP4hzL6UrFrDmHJ
xhOpZZCh23DvBWkJB5wNQBVdlYsE0pq/t+4bxi07xFuLXR3xVMmX9Jm2iJRLObd2dqoonMcv3dak
GxQQ+zQf3DHJpOL1NLEtveDny33vdmVtWXocOcvmTFC81fopwzTDKqFicBdZqTSl8UqFZs1ywpL9
iz/+M2RI+klJF5VRab48rCwcsr8T6pxs+zS8aFk1gI+QZl0eCSB7kC7N43dwb1w+hDwjlRHsI1ko
OcG20orznKRtP/keckCPl218+aGAM6iKJI/K/ABiWXucDpAR4wD1lqAbLw6BPzPjkpRU5wM/XYKn
eSgpP/nRpg2phJRTZewo3URK8qfH+DnDMJVB8RBChUg2R9x9IFoCiysVXjN0dFhSWWFBRH5Q/kOy
jPSFp+0aJgahmQ6gHnTvjbHlqxo7LKAUbRCIm/efi16qPZjyO7XRyxADiNXyLIWjMQaY//XKetrU
nhUV3yUbJYsR/pfKN9RNCdWvi1QQWN5G4o8uUAGGPSG1bEMuWHZfGC+BIGKBga0ldd4RzLmMBJiU
SaslOu6MBvna6wkEFs9wrHMDOT1arzQYUz8DDoIdqzb47Qtf5TdxVKfXQ4lKvDMwUfhouxyv/riz
EDIIK+QGpU1AlNDzUQe4ZTGGexv0LHUT+gUOZkLaq/5FgGJadJluMyMesK3UK/FJesHQ8IfEjsVM
OHFIyWvCzFTPJGBPP7rdDkskr5K5uHjBvSQ9fJiugry5nkoSI3H210cqF7DRtfN0eCvc5f1BbjAP
RM2KlHA+frhigZr3rfwOvOez9Ih57ugDLbvVCw394R93fGBR5IhHPV2m4EvpytqZsGrUtEDPTbC2
zAEZk8uGVylunKkfmVnThFGgStgrr0yolFkbuWMwgpnON8rZc9sxJ9fOEz0YUuf/3NGnE+e0yNuj
hHYYRuqzJlD8iMaBqs10zFviJ+fiJgmrik1M60Hg3jfzf/yeiEGvtmmVcdBT903WaUR0eNnqAa3t
CfHMxNlU6e3YiQnOt4hincffbKHotDezS2A55/gHxh08ekvCVGta1/YL1a9QE0f3FiPAHUl0lBEb
uH7yk8FKmNew4jUdKBToeLUUXbD4blgUq5J3ma69b/4iJrOZ0Bu/RcYBe4JXweWL6IgYtI7AP/6k
2t8c+ER6qbCc7164Tvnikuh+TpOUVlkRlTNasWNd2wuZR2TDEO5vv/oDVo3wnUCSsr2cxLg7wvy8
5WJjEWUg9qDlz5KJEtmnxquCSA4F7CxKe7agqVWDkFMyuN2HbjwlfcqdwM/Ksmqk7okGLhqPu4nZ
kH2Sb/hf+KTAVP5QCq/WjCDNsARFQEP4uEzrmWG4BD10UALBbzD8SUoXbCND3XLVogUWKcnN1C2L
6y8LQRGVZW3whAx6m6P4Bq8krG/WXMu4peIu/bNFFCen5+vEwOPOxqVsqvuYDox1A0hIzX14s4Qk
gYf1sQJB350MNURlWymCELPJWvJzWLsShv18UMuCK7YusQ9Zm55Mkj7P4BXIEr4pYvKHTZ7UA/Xi
V8HVQSZuf5NI9CfRl+g/1zJ5qBHaMRwZ0fKxUOJgGGdxQk/52CzIN0iBMmKSyYx9z9mE17fTk7iz
0kyBF5+TX2aYSb9xpxnC9h0kUmK7TNjC2m99+HMtPAFvinQnlWrYwomrVqeNBatyVDV/Iu1nm+F6
KnTeCuUFyXVAMG7dYtPXVNKkuuxKpRLA1IgfdLEtkxw5bOu+dy3f51f20fDAE2ViieyoHbemMfCh
BaIHesO3vtBQriePaPTT7g1mHhkWMpSO06euwEIYi62vrHQO+umMp7la5OwJe5shp1cXuwSYmGcI
pm+H8ZCfVa1ktrYNAVPW7s76tPfnAuESIhNF6qIOeCUo595qwrJNrpU5d0vOX39BpAq9s5p7MoWD
SNQlc/AuP9N5Eq7TOD5YodV86YyWUzxLibRYRqPEUaDvLlUL2xdEvGQJSujRZYAExh7vEw/AQzTN
ocuhCsyhe3LHjFRyr2my6dCPsjUI9BOLvCKaiiRE2BEjZvpHHl4NaFUbZsJM1hQxr6BMwWFcjw1L
6/r3VkSFnGQU0kZ+kZ+7LbD77KHk9PT0v/ad6/GsG4g1pPKIq764ELSXUm0HN7/4AgWh6iNuulkJ
Ita+mC/SVT0EG1OFeS/NcHfvQL9Qgd0oB1MnpGWrhFubrVssRHpabY773n6pFOEBofUtqxj6iYIF
Nri+mVyQR/wIBDCzOvsMNH32glgxMOCeejUduDmkhavafDE4sObYd1hNhS71MGjSLFGz1jTfEnm3
BU5PRjvd/3XYrjS8BNkD8GuDmn+9B4ecKX0uYyT8xtPSkgoi/gcOllf4YiWDdsLxWn/BN+nJC6/K
/3y2U1WfJx+sLUl9v7lrGlJWuycgo1i2bvsXh/GgYR6+YMZ86srLR6pTQqkDdDC6fsciJ0bQDAOq
H6x0XGGa/e8fLH1TwH+FmjZsJYrsDd5Wkn/wqc5GK635jvDJ8icfiBMJIo2ktfdWxTJa213hHV8U
8BwP/T0yO7HchVonCHmGHISqV+ho/2sWvrN/SUGHusK7FDzsEGzNAkZREy79bjLVQxgsILpeWAn1
iEAp7ablD44Vxgg4nhCZoAYZBF+vUG8mh+5WPPCi+nBXz89TLNy1klgAuNt1mbqGdA9AAWy1347/
5VB0G0LV2N4jmdr7uJbaONTpAK0aO7E9rzUBsiWX8QWJ5jK84S0BwwgUAMAS9pIUVc75n1MosORF
1kBF6q8yUH2M5CyPBXX3Ccz72OYHa7Be4Wq1N5pisO3I3VE4VKGaP9Mul67TaL7Qcgi/ePSGCNO1
OuWEcxqPuL3mPeLw7Ky404NVM4mo2izZC7ZA8DvTbtk3DYMWcteyzMc5vN4GcUQBeMsUqK5BHsI8
X2IkXeDgPkPN+6nyhP/krRITGo+WAyuxlcEn8dY6t54i3lx+Ijnl1BYeLM1mQ1PO0G4ChrkwvBOI
2ntbvk7hwdpKCf2cMlfE4BbEJiOYTw9VacfK7ZtwtPVdHL747hVfloBTKILP/Due1LW0b5UBSoJc
Sv3FF+1XUvEFwr342vZV4v3wTkVgYhTFN6ERq+CO4GwYBzLcDAMHY5QzzcjUHvhrRc7YNqIurvJk
0nLcoNxcw6n0B6nymYmdFGaO2aMzG6X4jk1D/w3fVyM1n9K0IB23Ku76W5djQ0GBqVNwWfvRP34H
IS6DDuVUUGsHObav3KCxqQ177msCrAuM/UHqnFQCBHTF1n3EKSNna+Zert2d8AzD8jdHVZNdN4Qo
HJIpYIIuppBNwWnOandLmtTKo1a/Y+gBE4uElPOvDOA36iV14gOT/02iSWqHNTwFScIRsDp0D1vJ
hkDDDPZGM7lY6xanSOsYD9/O1NiqCRA740oQon0BHScy0yk9aBxAniSwbKllRrh6jenj5PUdZmAl
m3hH6NRc7js00ShIXnVb/pZC1U9v2TWmfMCtgFCO5PgQ96PDaOvBAfxoVz8U0EJCXadW4nEUYCL9
5atYUy/QTUDtPptQjSweD1DUIIIzix1W8fv3duKkkjvX8knb+eUwh+SzHn7WmOS14Dy2nxqWpGFO
eVuiuuFK1+RgDAQft3Ez+aPTOjTfOu6jpyuOG9Q/P3WNYiLz4g+FpgvfITYpgcOCveJwXiqbddi9
GNfYRMMqDpAb+O9OobnGJBFcujdXvJ6Be0TsqWVU99K0OBCsYGcKBFgBP98Fa72wCLg2Uwq37oOd
9n8tLwJEbEymMhUpeTDSRTRrBLsLVu4590QHQ0ElpCPdAFwxMdrGNn2+R/nEeoHOOx7Dzt1pncNC
+VH06TsDAzU0tGVFA2LpkauLSYK86Fas0DI6cDjovW3vdrZchpbXbtMSXcN/y0dAHtRJOwZlWTAp
DlVlyRxqC7oL+xWxCLXnvorp9l3+UeFPiE/+uApDhj1F6s8j7EK9DNAJDzgOGtbzCtHy6e73iBok
j80m3ofWIXSk6in2ibqww5/5J6W6dxTmx+7HAoNl72lz/IgFcFuGWX/e1Zw5PRhYMNQXqWT9vPGI
Vh6S32FVYOlDUlPkYZGLCkOJLBS7Jzeo01l7Rl0uIPC+jv2j6gLtJYDBoDbjBsT3bqqXXdGzI6Gw
QP+NJ5b0S9TJA1yBQBUfBHm9UPduuiMFzO8zvrlgTUFXBiiau/dz7yb0d7vSQn/ujAILlIk0Yiy5
hODonDjlsaAglM/OBdvvgA6YMg6yniAARaSpyOszWG0hg8H4CAscuuTK9VRYqSe0pSYYd5riZazk
+D37gzGdt99MVadNsVXGovTaGgVXR35PG78LQHVCVudv0JTrDxIMkP2Xcg9KWUaeUBvzpo29IMd6
3AVU7OE8v232lPQpDZRXauX49jEA5820A42rCYIc4pwP5TVywKFomnu4LKmE3plodud+6YdHHLw9
akmfkRgoMoOURcqw84OCiWDq5TaBN2Ax1WU9hc5UziDWAT6Q879eLp3raXjU9QJg1uXGn+2Q+gsn
QyCG9JiKusdiE1S3CsBaEwqDx4tiz409qpf/VBzer9Pru9wEIrpnnIYcj58jNnhYktu05tk5Xv6t
5u3UUUJIK2oJaCpOaCbzaNP/ZWLcZCPjNKqZc09yvXCzMWvDknmXTUEicH/m8iL1qz9juaZNetgN
9A116cICu0M215bTQomNsiHzpFoZEiZiX2FJgEb+RECox1/peuRjQS4NW1qLrKGtfeCjJ3pDH8wQ
BCZdVl2t5jYn2qcENfD2PFRwA6h2FdBTH6wv93pILGjOyYQGVqUv92D1nahMUREXb8fn5F3hUArt
xN/14pwYf+jY72th5Xh7RUIN3RTBNaXWEfjO2+7RZhaWW0jFONJKKOrw+mOTsf/lAu1uHSaIVTww
rUGSAZOWQAoaPzH4rXPwS75LtBeoUMKq7+VEx+mrE2VTj3i7PTGpdTGRKaHN4ByMF3XSQhCoo3IX
n08VHigL60oz3Pm4ycTUQlK1KOsfMBheTJp6vUWTusav+NvA2mleWKqSZi6b4pOmSJGYQUDKqP6r
j0nN/DqA0Ho4npy5hwO8R849vdx098wHv9lmXrbpsTAe5KqYeloAaw6ZafuGfdoHrBvrLdDq53WU
qK+rZRmzvlxLDf6bGErex/+aVxKN57jKlUingkxQJlLC4qoXe6nZfNcTvlYzNviY8B7/qWttEBW1
J1sfrqM2Ng+a1DK+3jbnCyZmlDdY9g2mYBH/PFGuVnGum6BC6quS19igGdJZMn/wrLfnFsEYfsEr
LiLaPtlWeE1/wGe2j4ojkeU5urVmtPkK0MziA8EWSwPnCSIVEg7ALZ1J5Y8LIsdpO8HR/Wu3vkO3
khaRIjmz4rMe4PLm86v0hOVXNUWeYosF5OnxzI19u0+puhDdWQ8uFZdTMaUsNvV1Y2FHPf5ELVPs
95uiJdo2jvq4xnKnUbAJ2zJopnIvET12PM1Pbio4as2wCFmhH9XsRLxZRec+eLmOsz0Cx1kUQiHv
TKGuo1LiMfaAP9RbcV/Wv6JxHAg2qQKZ6LOdONNJF6x8+iFf4T4ZKflnSvhLWIeKq0n4aoeGsHTP
usghgMvI2Js3L4BKEqOKX+8M6RAeP0j9eX6I6ysIHDBgGpwpa/ELo8LafgzKQvEihQQxTJx8m4i4
WaYlXcARY2KBQG0750DofZZqZ0NOrrGij+WmgT78S+mAZJ3nFbJ7ise1O2KrtPwMC0Wt3G09bjIY
m2XE+KMd5NEHaO1o/5x6vquL5PiQCwekpZWTpx1GA84o1m2mYup4r2W+U0T3SsVnEZEKHE+489FG
9/lSZiIaGCWtG5T3bNShpC2gyPn0NKFZQiJdRoPZ7xdlPHd3EiGerFzt+tuEJXOyYPQ/F1jqAgZ+
R3pRKFRGj6WGaXhygWdrI2m69WXGROK7v63Wxwu7Cgri8LlXGPQBliPPdN+AsPkEWnM+HNYMrCKF
FsmdvHctomEULJ718bUnvJQ2Ep0WsLHAiS8BGw4Mw/o+hM8YYIFyiilAuHxYqCdWsvb1sgmu6TMu
oyvXioV12wL8naKNxTZAcPio1xrCcZxIyq8YFxjKIIjrRK6yYYeFiMM3DECy9i7r804EbMFLpcJW
aR9n20bDbjFj1IO3Ez7DjGKBOLc3KiUqayncII/ULFtrbfnFfKtOD9AjhBIkQYa9qsAHndDFfyX7
Ukc57TzlKPLR6h8/NMd0xQ9Ms+bLGUJnu04XmN/nKxaZwTcQSHmHKLvCDCeoC7TuYl3OyK5RIHIw
g2qFd+MgJeETJH71S+Wacbk5gm/AMfu3VE1juH9nwlcQNsRg4O7Ms/MiVffZJSPv6z2NJMI+8SuP
kBHQ43dompQMl7ozwvg4aySE3mphkgxLO8ZjwxMCoyxREjsOASK0UVVwj2v/99f630Ic796NFNvk
4P881DWTpA4vjM0iRV2hd+1Rhx2NF+cz9qZRez9ufYRMx8/1mVNxPWoa6F9DoyC8fClqKAhnY0g9
gxH4uURsnrBDelR80Hvb9QShFYmcFIcbx3snTTLfKwWqC5wO8nHzG1Gnu5Ur3BzwPgyA2GnqPXCo
y0SdhJb4vwezyOUU04dVNHWFVK5Fg9p9+B3ADXKOY3ESqRqjtVxydZpopSaiAE6CRy3Xpk+aH5Vz
aQ18+uu5dYwcPhCA4FRjPgmWmkspd6ALwcIW7sVCOjYR7PTjoAZmNxd9dlTK22Eb17QXEKQYja5n
WoACrf6g8TkfTEPE+8YepL6ZKya/WbvI/W4AQBEcPHzdD4VH80hg+9dc8I9RgZgtvPFkvPvN9QxD
DdJazqnYzS/oIkr6wCgyw+hO0T7ZA6uT+VrZOf14RNGbQ9x7Df3BRotStGSmXZvTpKWwoM7SEOC5
u0SoAxeagC6KIsS/FBuU/aTAtHXS3O17QE967axsS6KDK9tLYsxttAEtrhn+Jex7PDtjOrAy0vL1
ft/DjPz/gxsmuiQ5j1wJx4+rkpFgULGCnnYjPw6RefgTIwcH9VNnDLPz5z3Cmwoz1Qqq3yV8/hxj
kdkCUAGJ+K52nQoN9548ekGzx3ltvpLBoDDqWfyQYWtvaX/22FOwe7aLhiqXr0C+AqEsBmXrsLbv
27Lvw0ltEOQHCE58dTXXEljI4JTbbUX7mA6n05g0ufPHwofdaG52Lgx+r9k4RpxfghpNaOEa1eDr
Z/yinyCjWzwcTg0CW9BRYEnbHofR6QLXeaXv4yJMuSTHsvgl98BSyTToiU/lMlk7HCkdyAquDsz1
jZfIrM/1tmKebR0vtL737/thJtVEuQkIhpf2EU9loWNXVSYk6MyhEhqbFVRtRypuOx8tSkcGkRaT
y3j66Z+Lt6jv7DfD6rpHcrVlKE5CtmdbOP1r9n+5JnllnHoOUYuhlp7RGR2nATwv9eGrM1dOOElN
Obgejma5ilTAuMRVnqyr3Bg7QrMLDX+M5iGKLX4kdQZfoOEAxDb2egJcutEbTAq070da+g+O5Qij
YSVGKTQ/y9QP03zjKqD73KLAPnjnWBMtJSdA+J93B7QaqGj4s+3WEKWnHxv5YtjS+u9zRJ6TkelB
EyLSssL6z7iv/O6gJ2WXLcSMW91seNaMSn7NbxTgieSWwk+baY93TWejhthgzD5gdRszWtaUJ8fC
AXGk1nbeyFhoCE2H/Yc0g1ZjFPcCq2f5GJE2dE9EsBfa5tCVg5CnaVd1eowLFy3rrFY4qYnJdIaj
UB0754Z3rHVKdsN7r/4Ee1Nguo2oj/IJxkZ/7cBvzJr2Ofl8n1qvhnNYTGEOglod7EDNYFrmJJ/C
8XU1oN/uTmPIacEVQ3TmVxPeBYAj2L7e5qs/U6XZHTQWNIdMg8A6KEe9cdVgGHDXWTmG/tHD2nfQ
p1v32R7yI3+t31kXd4hAEjmgFDB5A5Y1HNK7YWxDrBTJepf36wd3X0sqeogwxBKQ8uldYvz/2+D4
5uuoMRKZJhGE8PlCY3Wz9mQnZvlty1e9AilKMZyDcgTy6sEO2ujoN5X1qcleT8BmPRRMeIR769FD
oH2/Qi+4FJZ7dHATcgV+NAeegngzJAZLK4mJdWq0szB2DhCb0nb6YZ0t64n+OqR4f2ljJZWv1TEJ
dcfUN0PlimCtSUB88NOahOgrM6lk0+dNQSv2ZkEo50kEUYLoqDrl3RSGrru6nsXZtUFTbjyRflqQ
l0uSS0k6kVWtnb8v66UiYKGzWmj0AwJa3fDI7pX8N02qKv1lap3Ow47ZOMv06S9nOouaOmuvLAup
t03qFp0dYoOowBqaNPrM61m2pwS+miGFGN71Um7LSHw0acDcbZCywtCnTA+LwLE7kzQjd4VdhZIC
boL30NLG3MQkx3x+Wk7+DH75VbE7Hwhdnv0bO8DalZoG/eE/uw1BYkMox2dQ8F5ovu7GDajDmD3I
VjmSo+jrTyLqZLfOT2MwJyoZLHju0EW3cyfrqlWgedzta2H/t/ezDuI5Yw63CN0PznEJHky6tESw
da6goGl3U/8qolhnY0c8Hv/kYd8ZlYfCE72nkli90Ygfe1VpnL/Y427SO7GpqeB+E3wOzr48ez+9
gp1DH82iVt73NE//MAWdqF3qSANhsf/nLj1jzJZfIV+72LM2vayF6QvuYBEFeU71YSDeMo2Ob939
f1eMTMvZaLYVBWY0MGs/5qw2acoMRy7ONGaYM/TVjNWu989DMKNXg87OEfaxl7wwuM/QCzn5ZPGx
3kyKStVzFvlYKZvKbtp1i0J/++pReLn3TfoGUp6XGbqlfsIV2+LeQNNDK0arT2QJY6Ln6bKZohO6
tWKLn1bIOqEpkYq9icsPSw7h8e9sD68lSgzGkkDSVGH9jW04zAHxybG3Y4UX8wCWhMszdbqxSNLk
8QBqaEat2i3kG3u9cUooN12sahKHltY4pfJQ3cRUQvK8PbiuW0Mv83s6dqVLNpM47D0yjGgklLwK
cQ6jSIkONJ+Whkw9dFEzCGrK1JiJ3QlIH65wollEgjxPLp3s1Pbx0uW2VR8kovoRwt+owFm4mq4Y
gw9sKxuGFg5WQaB5SO2LO7/ns7u0HoYgMn+PNNjV4G9UD90pr7CUZWshSs4Zo/Uvgd2Ts3jYAmCk
J9YzTFo4SyxDVizGDbmKgMujwtaRPr99MardqwSb8jPHrub150BJuB60qVE6ECGTQV197Qeo6Duo
rs7uL9OGcODEdSitfMoVQaFUbeZqZPn7fuwIqq9WwF1a+OT0cdzDsJtYxw5/9PfnTJmcqjC+39V0
7YRRX+r+hf9aneUB+7fiD2yp7AFKbWmWbyxYIZl22mBZQXkZ6YuTOGnipIKKVg00zQXYYDaG3nwh
5rF7rJ0SIyOjbUq9VDbBxOC7f1lJiCGEo6tyo9G8TZr+PDIxNXw2tehQYYcOeJkJVO9+j9gAhBuf
7hUnuegoTXvJFVevid1gS6Zawh5t6oPZZR7Dyuqzk4DSmUF9gToCdCkHdZDFWdit+6HEh6rXOf0U
hoyRaiG4+ul6ugr8Lp8suRmZT9PFIifkFm5ATm6GgryJVOp5YLFKrkC4sFeBuUnGrmdCyZ3kPWOP
yfPJP+XtVqYO7GlhGa/kK2Ki5YGTO+Jr4nTmfTrEuQkr8hj9F8adFgbfpuNsPyE42QI0fyXAeoCp
RIa97RsmVju0ZmMH6GiB3aas8is6XFMmFhVbABcEa6cDAgGy4K+PKEuHlivmagEOHOy8LcNY7z2l
hCPojCMzICJGioK+wihDAPndX1Nb0nWPecSf6JUkkF8cgUd1NvsLrPkxx9go4a8ZLt72GcrghWhZ
2ordrULMwii43w9E/DDxbPMYfUBfLxa10guqRYXaPDL3dfKyCIPfpq9e3tAJYOCI3k+t6EZFQPJe
BJtjAc8EiunYPl2nRk9zK0P+d6vVhauTBu7TkWdOAGpxOdssOiIS8zsEaUgEJezdhNrbP+ekW7KV
qDFbDJdHqMNlcC9TCe4Pwdm4fboIBBqk2cU/Yn6UQtJEbOOGmseX0Sy9L+gDUNSroYwKoAhswgwp
xbdMx0XghgHmTK3JKuqXGlsnPXMUsT340exi2L+aahGfY345GbS63ibvrtyDFuBZExJ+yvJHWp4a
CWDGcf8ijrCfygRNhRTV0bPzVZbctbwUnSROr101dVK3DrMXuMLqJBRgDUxt6yubYqghtUCzK24a
7RRh+ejJmIQD22JJzUYorBLItntL85pP1lfL7zokcwMCLciyjH9+l/db3Avwb8FidIgpj/Ea350u
SqajGFQ26tVKeHkyvE66XpVuVIEgp7rxiuRmGNKZqpEEEasGqLq/2Zw2HPJAtiIpC59riNwnelTi
vogMRVC74PR7769YufeQshh7yfOERM924N8nEC0NR2Uu5nJ6awTaPK3Z7QTSDsRhPeVXZCiCCy4J
HhJqcT91lWB7PDifQoR5QSPKY1QFjacfbGEPJDJiZLXMf4qTKNJ4XQ4OZvJNrp85sF+NmHqozVWF
lbsKbhnWrHnBp6GnzgoVCYOl6CpVt5LP2vN95Ln5nPTzxO7hRfEF29jMXEpfuX9ENk8POSK0uuE1
fwL7yS3C0lA/upJjMM1nXo7miX4Gt0MPbcvdN/B/htlT0uVPBOehEUVQqClWlolieudwqVvEaVTJ
+geUgkOgj2QFcc3NiNr6/lOkvyGJ9v6Du/5hXQC6fIk4y0AxjAh6LpYKImFY960rTQVcqSm8GkVD
CgYOEzDeBY2d5aZdIJzVvG/4wlkfEFFxZGbrSxApb/QK7O2lYW0Mb15rLykFHf2KEusy3BTbpTX5
d9RrGf5yEs2i1GPIY56g+U2j/KGxlGw5B9rB31NCORKRK6w52l0K8kQeyo3fSoN3GB+6RyIVHgt8
LNw+nGLzsX9wKI75JO03V4SXJ+w6iJNzzHQ1Jt3YCVLDz1FjCrbFBO6C1MaK+V0b+1O9qh9R2qAa
uNdJPfp4HiRfoFIETd9zj1+fZ91nwKNzgEL0tNNZb/pWs1eIUHh70NOPPu9isHI+wjwF3Wn+zbdZ
BgADR4Mx35ezLsdH5C16fwx24Itb2IW6gj1/6mNSz0MtqT1hTDMY2VTquyPy4/YtAkaWIoVMSGuR
33Oj8KKDyoD/LSP2OTVkn8ijp5cF/MYmJdh2ygdbcBfRT/2lU/yVCAAgDwgAlnQ1e4a5Btwj3zQz
fN+nQdDfg0bOwAXvoM2qhDD1Dps1Jb8eYjAUoxp29f7ZyOFC3cMO3uZS1CbIoT9m28iPDbxKOO4K
Qi5m82TOEthhfWUdorRiNWegyt53KseXdvJb2SDwtaQlAtO1D5hxuNQL25zXENSxt3yyPWj3DlAM
UleF3dZ4gnIf7jiY5NueGb0YGpnHKvnA0rU/P60CePeCk7UJ9QJTBqnyQlp0ZeVR2IjjBxx1kcKd
q0sTuj27eUjZ9HV6c4U22NBFCaNY4kNxRFHsH8mRjaNnGuit5WPFqWfch7hSj9Kx05oVeXiL1Zq2
3FPzdrmpujA4XB4yIeq3nn84OZOP0R//pUOZ37+Fe/IKH2tGcljX7nnip9gJ+PHFWnqrdyXb0s4o
1AnS5DXPAHmcvBpnAkHV0cv+xqng7BgubZ1gMV5d4buhTtkJwPmzfLiNz4NPxtrcBtgFHbVILi/b
l8t7QntR0WUJ4GJ2Ha8wrueMKcDbckpewhag7bKKM8uRkQN0P+cmFQmhvNzrjG3S3Fqxdpi+RUoQ
jtBozcxaw8jnoqCE1m+pQ77dkmBWEql2EA1j0Pkyu/RPZnnSr5IPtriPYlIjmusYa7m7slX/+mnx
H/lk67bQ7PM4+bqg8rwN4LACOmwVli+duu5DQEBR+7sZ/dcGfh3Wtzvw7hICxPyOHMkoNcMPPiIG
XKPsIO1WyqEXbKJOlfPU/aAD4o5nFnetNH8Qcy8hjS3nVphKvdtpabSs05jgPNrdGe1mZF2ivCWg
vbPfbPEcE1Tck+/YEkSfS5yZIumJk57+VKjwno0FRXbeBQM2wDbhcNM10a9GN22cjJkvYda1j6hf
dDMAFDPlPUsDfr/cRMtKO/Z0NBvMfAdzEaAh9ZSgsFatLdgFAJh8dY2Q9mqt9UfEwEziXIaAwv2T
rtMe/wlmh+GfT4LSqNr5VfFxd1fGT33/+Zia6a6jR8l5kjcAEA7/lASM7xBufnAEUHI1MSMxxn32
LElH2xlI0by4k1wdjhyg/DL03ocWe+9edV9NekqVDO8a507+9JNn21JzfOqkMeyJmSfyDIB4TX2U
7sc5zCYvDhZJjuLwUF+rlu3oWFvv8DlYdo6NT/fN1xs/DKa3eMWlkWBF7K6WFbePxY7AuCHFL637
cmtXnzMxMjLrzNfFUaOLMfJ/28ak8qXe5TRBag/ucVW0M4hIHhJNP33yHd5XVVCpsvmzPDQpRh8G
5f08hV9p9eqW1tfFQaytdOY/g+52e/1ZS6Il5GiXQTul8+GT++CL/FI/guSoE83apogqS4MqVnE/
HcQbKzWnLhpGSgEU2lPJwr6gPR7QWG2M4wDOhVK6q/gjjAcni5LSPY1iA3u3pllOom0A7cqbY5id
mlezZ+WcdVWiGDdGsbsICmoyF8v3Xp54JBBGo/JCcmbSWbDoSci4H7l8LUvAIT7Xt4frsgGci5R3
lNe/iKXooGsNIc3Pflff6cloQ7TdlwonFGceXCftFh+s4e2waMf4Vdo/P/aYWprFISPnluH2Q//u
cn7mq3Yg77bIiCAqAHeTBswT8OEGc2iqEGCzr81h1ZWhQ8FsTLdzAuBJiB/qmIN0tRoefpd9EolC
fyeOFzyUPT6ErwB9dDa1zBLsDAlBBNX7pYeGwdZxXNeVCGJs8KGu+id91bTtbrh8obFkfZSN5iLk
wwXr0p9pD1f4kRv1eD+cpiFLgjBUgKdc8KHlJIHQmwoLbmjwRuiZNye1+GTHPS2cBRhoRrLI85yN
HZmjvICM+AGf5RA0unmWzhCh+nN5FKHZZDe7E6q35zmikZyxBqKsp3rTxcHcaGpL5Xx9u8N7SYT+
S77Vy4BLfIOUL9H4QThXkM088dXZcktC+BliUp7Zvl5B1ky9Jn4dw2Rtx9E61GZi82EXhgctJqv3
+MCcb8o06lciQEfZwL+J0kmmgG0HbbSint1qgBPEG4WFm5ck/yT1dvIk3roxl6v/fcLMmUFIZsyx
dIoMv77P3r9nBa+OqbbPFQ9mcMEzxWppwLChDBgqgHsPpTxefQUAxM4xJfX1sMzoKvaUHc8IB0lf
7aXoYTMj8613SswohtDT56WBapBdIB92pV1kqfx93pyNKehM0romX95mZR7YKpM4tj8Td/J9UHMo
vi1hOwmDL0pyBYw0Rdr2O1KvgB22/2r1e5G+7qSiA+Dr3ykd66vvP8DReoxCKCRhGTbT2RY3tpHG
lpBD1arIJUsVWPXcvpo12fd69INhMmTcICIatMwE5NBIZDmPqTBeDA2FXx2D0+dvw8GXqqtc21MG
U/si/bC0iq8AEGWfkAuhbpBqrGdTc9FQ/t0Iv41kd4XjXVeCM70hVY4WBgipph41NX7AtKAXUZH7
EAGrnG8wgS9OaHKrYVVVaYfIaZj/qEZB6Y0KFj9I4Ym/jUQL0fS1l8of6EOlFKMFJeFeDEnSXlff
ZmqrBO2ZJhNeDAbYB8S6EfQWCA6jpRIp7r6xhm5h5a6+tvd15XNrbd849ZL+HG1ViliqrznNCxWj
5BkmwgshBr/nbA+PZVj/gdPqti7BnO0s5emp/WtY1bOZJguCcJR86iLMyTP7+JEloOp45PL1DYDf
dh1zFeeH042LeU67JCPIPbqi7zDaAYh4F0lhfd+vFbi7UXWtVpcil9ZHMsANuwdoUDugU80L6eei
zsKHD2Jzk4afqZJoRmgxT9Au4O458paQtjA/wqCIPUUWHQcz6DuVEnGp69az79vlGRtvjgVX7Cvh
IMbfXbdmXAAkHL9iLvY3yk3jl/By8m4QBKMmpnMs8kv1rDoXFlygwbqltq7tZUEiQK8MyrORQakJ
CU+qFG44HbIk06XENPw3d79ake9P+DLX0tWaKI4FdT9yi9ydiewunwddWMlNq8B3Z28/YLle43mF
BUZ7zteol3B4cs6Xaw4YXXKjGA5CYNbPkRZK1bJsiKlsqJf5xw3hjuJ8WRwxA92V2GQBmO4htgjW
3MxG6Tmv+QbBOgZS5UPP2VxfuCsgcWWCpe95uUqqwwRST90fdkrO39i2eCybpKAud1IWzhOXd5bp
+WOavMwDBVshOeJap2YgKXfTBuBVAdiUAol5bNDZPnMcQlMg7uEDdVwdili6zC8yWaUe0WeH6L3x
O0QF6L/WN08p2/6e7dHuxdrayADTeBEy1pAlLhhzywj/Q2jYSpTXIVQ5Oyycu99Rdjn5kO3At/hG
ibxaA3uyWM6Tg7+8mUG2PJXoqWgabYtKMVnRkjYIXk0L9hZWkIUH4YIfYYlTlrZBFLHc371ZE2Ua
X+OxrpEO6nJXHCM9OMEmKjC8YK0iEJuXb/PV3zhVieQM4oku+SKv/g0BU1MVs+1fZ7S3VzzYR88s
PXv0QxjUCi5QqHSpObF4pdykKnWyJyuC+O58jvHgsIdmL5lgxaV72qDZM5RbwnvVy9vZMoyAtWp5
1R4Gtx6E/2it439/ohO6Iv1vHHceLbxCaLXiKYDcFjfxUmsA7x9xLMvU2eVbSym9d7reQUsBSscE
3sj2zE2K31ad9vBxZE6l8isozAlN1OmVotv/viIqA1GVSZnyiH9wErdVe2Po/5D6ePF66OYi+NUA
tuZW4LZZCxEOF4+ck1nqtWXYMlBhnG/WLTxpLMPFbIhnmCSVWyYX4MFjwtU2MBAIc2R+hZM1whqK
JqdCxwPYWZY1oln8Witcnp+E3QyYEOyEQHToB1SxkDLxGg9Ez20BgRiMvcQz9X4fV6wKZf9HfnWE
NjxxP2MlDm7fpM476oExfjlsTysaYKo/io+CSIjs0qHggACkBytRG3exXDbfC0Stu4LznJW/a80I
MzkeITU/lYOGs/4bRqOranNyyY80lwusNxErhzty0wu9O2X+bBjZD0Ty+u0u91wzJzkAP4Kk1ywN
panU4CKQk+FFhqOLrJCUcWim9gM8sEDjqoEYIssZZzwMJKnLrW/G23VfRA8KD5dy3jPuQURnq0/h
HhvvYWUQ0WF+IBeVta3Js7hiyb8Z8gY235Wva1PT8YdPWJhApAfx2ax4Hg5YY91odSX9OHJCsJcT
OVOyX/F5yvbHNPfKcN6T+i2YEuLZPuVMzKWJUJkJPOQFQkTX3zR9djk5OwGrqq1wGITsJyHtKp1O
eUtLsA29hTa477Ivon9EOUDW2wrI3iN0E9YRWxPcLGZ6UiuzJiIm79DQ+iWMs7fJbR9CHHXjy5dP
BqQ8ATtK4UNIEvlGLyBkigO2u71bG8g3STnXfy65L+TkiK48s7KKMTdFcvwab4Z7dd7Qg2L6vqtd
a3bXlLyGtAFY0Px/EB6PnCbdw0bwr9cMOMiGx749+HV+qsFoqy89upzyEnFckAo5j6mAL9CuGzaB
e0gwQK9Jr2yzSdSl4cOkXQubNPnFxIJyJNKP2kKbsH+fTcH43RdclwcHgu6FNxrf9VJ7vZEz+GDl
JeJ/oxuV4lRFkZRAjrSnTs6udKOtJ1lIGC1pLDbPTbegnH8LsPUDGXd2khcCa0b90jrEQKB45hKt
9Ovi/27u5XZweVBrfP/+NUyFNlPYjZKqeKy1TJraeV7s94OrmMx9orhEeqVYJrpSPLB0WraibcPd
GBklTfTkPC927+JUaPlAg/nFmsM5eTmPtN2oPyRHVeuy6vFdGABCIekq9lSb8Cgd6dVFWaaEykjG
ySEmF89JgIg7NIJWGx1+uOymQCoiHx4/bqi4XWhZOizMLF8KJ1dOtK7ErelMpkP1FCpLxFuTOKwb
BJVHQKh/brEIfGUEy+C2fCoUDmMXZRr9z08+rBZNWpFYhfKbn3+HSrxEVaK4/STboPmbIDvMVijo
mi/cFPIanggdxxMS6VSiyFDzR4PMiBrbASpqy4tk7YOX2YJVyJHb7iZGczwce1KSISnc+fCogJZ8
yxS16KlJynTZOAahybkofGcSLiUbr7WBNwEbDAZlgpRvO7evF5YmlGVhn0UTnghnr5FZcUcDtkB5
mnrfd0TP4+a/7wD2DAh0I9vGIqHsNi1DJgPh8GgXgu0iMnH1J5Dr3VGogSXBo8927H+AmWTSFXxa
OFevrJjnUi6QuTgnC9wuU13qWwn5OJuStgO756AJEGg2EYw2Rm2yGRxlawZ/iABpBcNGSUbdbYAN
P2QhG9+KteZKOd0jXcpMc/e4t05JFjr0ah2pfrKcnADPFggookvkzMtqwMc4+yAOCbytFuHqc16N
BoNQ3gsNyM+p2vXEgfVNmz9ermffGngFkUr3glZdvGuzTgF7bCWBlRrxvssDOssVOxdWkPL9XcUg
PYAocin6YNr4zQ98wgUhKsLBCNQRUTp1spq1mkDkR/tu4HfSsR/OCmWYY4iCQdK0KBmMmo/W4A/J
3Df/d1BsNn3ML/2xfYoSb31vKvyff6TrMnTJK5mDoHKefykh6ksxeW+NAmSuHVzwBk3JWYDgwFY0
tmKZ0bt8hoEEfxZ/65B2BZfYXgqG1uOeysImTAVxw6E646qE1I+her4XRU0vXIyQvIhmYr87BzvM
0ZyMyIrFghTfZG0xgw/cxt/LTTf38gumxjsHqwSonvEdez665Su+cx0cUexnbN6qrUFFITEEM5xw
PeDibYNwXO3xyH+H3mEfJuQMvNRZJePgRM1TByRLyp80fRtYXoRoYeBTm4NLvt1oseZOlwKxkbmi
KvJRjcNe3jsn0gqphXhqW1gubI3JAWYzD9LPiKuKzf/tPZkquY0NEocHAZ5kJguBVv4Wtu6gMqvq
DCYBAWgQ4QejSxQ7T+hHQ9G2rst0ZD1FLX2FCl4fdRWUvAI3qN0ZJwOPxIlfvJyG4FVHTVz1mHSJ
b/ZsLGe56PiMmDW9AnyZYOhH6sZ+49ZSQQ8DgMFQesxyWVn0gWkXF9CdV5P06IbUzThGLRuMFaCY
uMCi73flEW5TSAEmqRR7TVXq3K8QFA4HXGhruJivhBHHS8s/YBFRJiCyuazTmrXzAfIa+xji09nV
kPJnearoAMdagA0rAzOrEXMVOAU8MlrTht8RX0VKWSxPG0So8H3tjFcRDf8vVUaRuqoCdjAVpbEb
m3OzhQwQy5UJo4wvSM4yOtiezw9FdMaMpG+LKWqjdrtHUVGtohzmfCzL3XOvYR1vbN5Ia6Fh/1o2
xtXGWW/IQ2JZ+5fbUgJv3cdJq9iWGNH1u3JCZhJAVBeqkxmDkdYWs5p1d2X3Ll50+S+Q8tw9Kk2x
uWrUTz+wgmkQhbjwfulGG/hYl4nPJ/z55ACfGds2cOnUXu/DqIzv407ZBrzLrABpZbnEBXXgb7K4
Nq0Gx6DQRJFUMssEsh1bSDNSZTYai8o0MUDoC8ScwIkWtSzp+mSvvZBlZgj97uJ1894HE9nKe84P
wFI7Fp4tlDUF4o/1GLALC5cBrmL84wBZg8SkIioqTJPwfkc9jPtAIORzjPFA8e2AcKuMuzFm+PPO
3pixMuxC3pI7PFkvtnMk76J8RFfxNMfkF3ALc+Yqql8AF3JKzqjqB2l+otvuO6ICl2E3auDl3ke+
7mPuJex5O47E4ELV/ygekI7xarxzira1ZerUN1mcZZJNOzl+B5rFHCXwjyq0UIDYJK7FxU71HqXZ
2Kr/RkfMSsl90BDYaYxsLFc35qpAR9X2Xryy5HZAqDm5Ueyet4h+sRn9xRurUB0JVaPG+6MO0XHG
/10hEqCU3dkw1IW8k8p3XCHRnhJN/bRsOp32K/ersEJKt7LDGWBeTArW7g8YDctsFvKJrGpPf3ko
n9Qg6yKI9VVblt7H/A18X+M3ii9y7igCreCBln+b6Ig5I8Wnnv3h/L+mtxvph9bJy/KdDesfX+J+
mOEeQ/nSuoTJyuehnDLUBgfIFINP3rVmF2pxVgBNbDzEsehbkFcGx4QCa9zTAWZgAnVkBTOfu+Th
2jChd3y0ZhyVXTfBnIOJBARPPX33j0CL81wDUJFQJnrXl8Zq62ZiKqtcuw6fyOnor+J4SGcfMQ9p
qBmLnrSeDbJ+iZZ6DUiLjJI6nPFnnACyI+2Db9dI2vtQpFAKSCnzUlIQLPTxJeRmldrrkxxXXi97
AMuCF0O1nubCfk28PBOtc3P8ZuGnqR4HoiV8sjPEBM7s4jKgqHHUGNuNhcO1+EDlsRL3CNEdDGVj
FLcVnowHXcruZjryXs1pp/S4N5Q5TsIV4vj4FIbtb7hGxPqzWaW7xrP9l6IDl9GlpP2cz0IF7XMO
Q8l5VWMuKZsN7WpYHN+HiDenrERdlsF/sA0kSn6Fj86dg4r4jSKTnzeXM6x8X/po4yJwGY198bDp
gvyJD5N5NmsgnuE2J4nNlkkPcCfydRi418MpFrk/1KksxS2Ie61sql7TDFVWJmMz6O6k8cw2LACU
/PTRJoTdpAqlx2QPbXu0RFzZVpKGCHv690uheyByT37ng+eXhP4oNEAdWv1Yb08kN3GfCz89bi0+
VUNIlgXqhpbkssYHafKCainW3Y1g6YuzANs21cLVA2kmGeqJFpuHHED24PP+u9TwjtDALAqCm0IZ
1mlTAYozFuNYiNPk8jR7g1V5SnZe8GivQUv7u7XjZF7bswIIgt2S/LbV+Tr9WvK98GzI2srUbYKH
DV2UUBeY4hFjpE6mhODuvsOpUjPyPf5jZUQAdIG50FZtG1w3oW4jT94NPa49k/i1cao2eR9Mc4uc
M40UO57F2uqSNLnb/v6lay8dxRgzwtJpfNwyI4uC3eBscG8PpVH7FdlGA3qMziPwMKX1XIq5C54e
tonj2F1MhcLrl/Rw65Ozpf4/XmN5S4XAYBgMtvJBbRO/Cyc/05ZsWgW5DfzGpRUG11zHmMVS6JsT
Yu+N6v2AYQs0cdB/wwbsFnmPod6Q9F+P3Npm7ST9BvXYncr7E2OoJFzhp2dyb/BbGO1SRtGaa2z3
NcTGicH9ZybbA7YH9KpcgTM+XXUk8adbGg3GfuYzZ7yK/bavHktj+3Lrfh0hgHq/Ci//9JyyK6Z2
ld8eWOg2rEcdjzuMfdQk0sozqUkZ8BKP2LFnW7tQVvnRR0GHIclARCh/Luz4h6LP67rFHTE306WR
ErVPGCqtM1LuinMAig13yIG3wNuLUA8mcOa42aDytb5oHGl7ZQTGYfuM1E5uWzzojpmPTcvJSUD0
UjRgwzmMJNyuEoCgT12Y4TlFNw+T8RGaBkcotY92S5Ihl62b/+ukgSDs8KKlS4E9T5Nbm3EY2qOw
SqIteHvm2APNID1tOTIPs+wvCcM8PTmc2PGvhFEDA1GOqs0iZ2duPOwy+9bI4DM7ll0cJS42zfH5
IopuxVj7q9WpbujWM8NYaxs26DaoecyFWbkqT38D++MEoNJyM9JzGEfoarjPuWm0PReGGul+MVIY
rjFYbPRFYDzMbyOs+tGrHxLraBZ23Vqj05/BoS+7X2Y4qMfoaRrRw8ccrw8M5ccnLI0B2znVnF7+
C1NucV9ePgZPwH+RcpYPOv0joc3INX+8SOLwlGMrZNbS5HmuwyLBi8P9WGrcusMZx0GKh0B1ir1y
EMCjkIozgsiY1OIvvIrB4xqKXbH87cvFp5We3uJ9yag7T+G9A1j0C+YgF/ulFM+1Oh4vyoSPVvZj
eQU5KmUvrOfkG3dNISdxlDV+pDKK+764aggjmWWbePBJ6q/whx3IkDiuqsHKVoTHRc5oXNcr37H5
ZLccO+WUo6mx2AoFYGcElGybnF5BDsZSSUFN9jBmG4tuIhD3UCcMGE9FkyNtPmG276hkcDFaJBui
D506iHqUa/dntBbqi0SSjAAsFvOIQqea5Z8l6/NfTJ8DZHeVRfORr9l9UbfPA6Mn0acsGuY0MbWd
nVzYRV5vY+QwLN8hLhSsH6kegd3Uoz/38VrzFZglZ3FFClsV/cshV/LJxeTHzNvjvlg6IV9Bku6U
Ash14xkbS8d/1V13gMNTdD6M8lYiZKM+9RqpERAd7HyXQXnUGc5K6TPBKg/87FteYmyePexowlTo
y1XQJ4NhXE6WZ+p3HlTIG3155kok8/QDzdj72YE/EpVnLZLqxKp703eSuy+dfdVR5rBHHa9uMy+D
fvJJkDHJUNGFGEVzXPCB3v954sroe7sQ/3/woGFhaknfhRy2q9f0E6V7aso1b+W6M7bvfPgIekEg
H8iXanbpT9iysuqzyzqsj2zV/qY0QEW9BV1Rw3fvbfUeMae/lwwto9DbAf7sJ/cGVsVZqRtpFBHc
+4zQTkTqaU6l6qXW434gwAMDZsSr3YiU/gKz4UW+OfuLg3CsytYU9ZQTVKjRZRWpzDapAwhlZeXz
lvJNob0+T5Jq118qCjanR/2ATbtRq3o+MKXlLGEFQsEbEl1jyLfzN5rbjkzJUzZhSfN8sRpqJQ/s
IOgFqqv2rZDXE8uUaO9ez9uddFBxn09YyMbj1L0FW15uEPSRFf7WPa9Zv1g0hVSsU/gzpi1o2wcN
k6VVe0eEqIt5B9VRVlW3iA2P9TSPBjq1nwdcuUtm2Kz4JhWczEwnFY0Ae6wYUKa3A0rdMIyF8UYp
5GkrcvTsDdgEkqSU19Bf+VPPJccMrqAHuc2hYh4BPUYbcYIsibXi7rmuk6bouKeHjMAcTdAw4cVP
9cs0uLDdzbiKS+1OoSdAnSRNi2fgtEgevsHAobeBCRu4cR8EAOsScXnX3AiApZAWuQ61xTSqi6Kg
f87HknvIs9zr1jwqNEelyx2kVie1Ud2UgypjqEZIIVoCyvBVVRVzutU/0sWdSPodQhd6eFw9OsYg
mPT99DNIEGDvewlzNeUgtrs9Lt20V4hvy/kzdW5X2VDq2muOn6E9Hk+gejucCdcoAKO5/BhYUyyk
q/21qDpYmDok7r8llEBCQSxwep8TWTuHw925ue8YU44Cz3F2GvDFgX37dN7P6gF9cQfMRVoQq6n0
uacjSoLNd30sOZubinYobEeiAxAu/Td5RPfYLUScjvp/cPkxibD1F8gem+d9gVMPceEUVvHTW/Dv
oGGYn9o3Scgmzg6Xfz58ZZGrYUv7W9vXJfLhDJqWVl6gB7o4UHjA1+XsihcmCOL8USKUL21JwGmx
QD4+eHrhoYZvqRVNDPJz2ZBZgVDSn5ZOmpN7Qf0o3WCfmdskKqCLO4wSLjIPhPVyq4/VLEpsD/NN
HHGks/8Dvd9grmuZ8T6t0W1kRqlhK54x453c/xUgsk1uW3b9qFZEfjQyv42LkQI8zTrpnNlZyDZe
E4AvKPhFfC/qsGQzzQ8d86U7spXswz4bo8/1i5GtpXG14QbisxEHx8vPJnL6XvPbXIIns1d8AwrV
KVLhC/G1nqKtXAD1QjH5G/edAou65Uf/JkRx4JEliEBzEa6CdcZRjtXU5O41kwCHTNOVwH86XzAg
97Xrd/z6yX2YvdY92VUxrMeUls1G6cGOe0mJaL1yFzpNbbc0PhISvOVSL/KikulRxChH+1qn4X4b
GpULcvOgX9KRLedT2Np6T91hmkBq4hc4BE2tFho5oawJs2F/eLYla29ql/lIelHTH6+WK9HMGUQx
/UEXXo39B25G5F2jwWiR5QbQuTx2j6vKDJOf0c3kY8lT0lCyTQLoijRWczbL2+g09bBj/QKMrmgq
lqQJfqdusSgu/ww1ndLOkTZ1RNgqoUtDuswVQXyL+QO+Ml6upCe/HiBCCcU+Bf957GlqN+KKRBt0
j/CUQAvC3svR4jAYjUaYI0MBwpEaIVRLey4/B0M9OOBEFeMl1EpxS+poLxz0jiQt+7+qt3aqEavF
4f61Bjsr8OMkTqPAMXg0R5fWB519gHIqZOq2qavMqlJPDPISr9dZqdERFM1ReaMbPamzMG/uCnZS
XkDZULl1k9nE7jp6JPW3yMmo4eIXiVJFYRi/tDQDnizWFaX/Xk6DlsoVXxzSBqTr9CETa7AGCefh
+ru4xLk8p5C17XJTeDVMmBnxX+5y4fHDgKA8MpzQ1hGkWGchj1eNEkvMC+rL4AOqddSXZe+LnOEX
fc8PObG/R/7aHNdEbz8d+Vw5hjXiTTeV07acTdO+pAUlAWsLT+QhXPgRzmPqBPWOQtCphaRVMxqC
d5gXsRj/W6HGniREQ4MZt6qwoMqJcnJsGlGFmx4wh3DltrwHzJSKQqtMvF+6k5uIXTUFUpmrMDoj
ImcV1SgZcSxH0zOA5bszgWsW5CB8CPKG6R9t43Nuublwz1J9CBqQqMYkhHeRuonhx/aRy22NlyEd
+DpX/B/Y+gjqx0T7hwRKT07bd3Y+IIijuHPMQzgOMD8Q5s9AqDiYM3BrJGupqElhjrzY1DvV1COj
xe5cnsxj5GJzER/o8NTIDYUYCYZ/gIb+MLTSDg6+kZDzvAFF+rhFIxTu57Hh6yTb7FFSU1q9Z8ow
cWQEYSMmNDnzhzWz3iJ2bVyw7/OO1l92FvxoRwtL0rA/aOYgEX8QcI5kqTN197mtnGUgGoLLyYDy
LukQLsdTzb39NZGfI12Y6C8OtHavWefx8lfJV4UXg1KVAf/pKlLV4tIh7NYF20FtB2WHTqTBBDm9
moudxQSqUXh24chiPmHcHJ6zQqLukWx+E2JApLUT0j78MOnqCfRHtEaMJ0f4ubau4i0PrSQenN/1
MpHbJE6MdRhnpWlg4pl5vG3Z2fUXiRbuCu9BgqJcLlRJyrWvGJMHGkJPnwNiMQC75vjnKjmj1zxj
cWvFizQf2Zuj1fPlfRHxKfeDo8R/TkTQ8xckSindS54HNSAypW8gDr7mlo/XTmC1c6Uv2H+/T2kz
CPWzA2vJWzDK9D+OfLusbZwAwy621etGgOjgydMmLNb592ML4jwcjJLP+GS5XFwr4fNqVL8m21jS
hbPwH/9bltCDa1dnXCukC4qd1UlQg63bdCiD2hPucmHCmssvU0CZfXPhIq9bPz5eOv0FnfNLL54O
On2fyMyEnVSLcVaQYboxbd70QUrYCTodHvMhjZigYtQhsUexlh6nmmzz01bBgA1FNANV27anQMFX
Ww8G/LdBqKfQILbE+0BWF30rmUfI1zr7NB+2XkKcm/HGEakKSUjxIovAMz/b50e9A9YrDhzwaCV/
Z6xcfFbXKdz6vYEZJMCw3Vh9sXvHglk6J/OcU/Z1NCnMiK+jGvwpfV0N3VWmzvXzvcC4l3BKg7nm
gaKWHabUNIEYhdF8qo1pxej7hkpxgCQkyZsi7yrABx0f7U/bOQM25NiBEKGilVENLrpMwGKw+r11
Zi1Faybm7hIomoI9DxA7hsOk97vBciZFKSfJy+FdUEvBvlUPJLWvQClZrpjtHNbk22jgAxbLL/E/
qWaLVSkikDR+geYf3swZzQQI5FNd+7OheT/1cTvEBCi4vDxxG9989ZCgIaX7hLI+7ekz4WrHVrzs
5FyE+atXU5Kt55mFZY0tFPWJ+l9lq/ro9iH8QlwDL0WgdwGWV5cRDrtWPejoJtqKd6eNJTSKlVWS
CEMHE0Fs2VcfJZkvs0YfBu1d2wjaqXcKXW1fD4o5p54YC8HMD7Hy4NADlNCgXz9JkaMZOk7KaOZA
LxK9wnNd3nSZBMsQMog2ddULnEZYmsv1spShjIKwDQkzLhEltiZxZ/UzMPsbGyYbz5GXo9eM6Mu7
2xi8j7dWZK04nvCLTlndM8eOsg+Upzh3dVuVSUE+8Q4HU+67+rufo+xr1kv3rdx/zZ5WsXc6UJu8
o4Rw4e4SsFCx4RbusI2/f4LpCNQj018l7ixlE3vnTqU3AML71nejOqrG3v5ljMlr5g/kQHMbhl1z
1OGVsGVLq9BZbRNw5nclWl39a0+HSi8i6LFR6XEVfWb8pYIIHu+mrUK6RQ7lGrUCtNPv4epGzoMp
9kbDbF7ZxzR16BRkryNmclZQjYl9JhA3dXaFUYlpY9DP4PYIaqcKvF6nhkVRcsjq5W1B2PVUhhcq
t7PVmEXfe5x7Nzvattd2VtPQHxP54CrjwDBceUz/UCjc5sbRSBrNRVodYsP7Idmf14M0aH0ygHQU
st0JFUVBE4APNT9Y4t4p+UymJf9IKmd5PxXfEY1Me7zn7LH5e9s87NKUi8lIhyLaJ7KD23w0aTXu
Op5wpM/jfSoGr94ROta35SajNeEUIhzAYhN8ex3FGDAmmmdX8ou69dIh6GYwW5qKU2hSQdSSlsxi
K32yT+85hx5NTeUERGYqoE7HGPYcMGddui0eQZrJTRjfKoPKq4rlFOrgg+Esfaxv7AKzFrfGZ74q
fmb9u/iOB7GOphNBt8a5uX2d08azSMIfZoaOpjn7I0F+SwSHgBJTjFsTKj3AVB88ujZ3bwfHgL0m
I7uX0ev9XJPDH9Dp4SXMzY3h7pgalMVF0J4ewAPSmHfOp43+Tl8a9RMBSOQ9kRJPDXvs7cG1v2aP
aOgSkEFUoQL2yz5VkvQCBF3KQ900ppsIYVKxwg8+1rTjM+0vIuvubZLn9t1eJHVkFG0/aHXG4cKf
82bvfvaw9SDmgZFpug07/scK3C/6keY1V1jDeXn7Oo8l4mNOqFVIYTL1OKHJt734eBFLfBVvn6QE
/I3VTyNuTeCzFoHQnogtk0YqCU0qXmQMF9yj7ukDWR+8WSnZfunEkgI6kJkeRwkZ2GsHkQUpva+N
BkhGep8ZNvPgWoB8IB7dkIt5+pHcXhhXAXHnI4CuUqG+CRfEASjkkRJmkakQ+XveNfc/aXpF859X
GkmPC2ka6qnHyCUXhsKfWfZsz72uQKVLoN34fm7jfDIVnAaFeHG/HO90eNQqmCK4GiJxLgE8MZEm
xgLOKuFUu8eScMJcQAU2nOgZIXhgxyjEO/DNOlDjIenclZkk3nTMm8TDhWXnnHGTpZ6HYynPYBGO
DUwXf4JWvtzl2PBg70Pdc3/SKanqfDTnxMlyAGIs5t2YS6g7/mdH3QpmON1yOZ9dFSiNZC7nBNP3
lLIgmaNWsrO5KElFP8lCY7VKCNrpWK5CHKdwbmy+g0zmmYw3CpyTKI+zl8+kmeLLrvS+yc/ZLOsK
nco5YNAYn+O7WBZK+NZMqXmf8pC0yhFc4IqwyK8c2mxoC1q+V1QZjdAlv5JmEFVCYRpoXJhwKwqk
ThT4trTDY7AVoa+I+HZrjEv6dYhc7gKrJLXtDmGTE4Wa9jhU9SVtj3ksE9f8iLBoxUJFuhabJjsk
q/E9NdeSvSdpJ5g3HeoFKQgO1NbRn9ZC2rTxkQU+vGXr74dGk13lKRR/bHXNxfF8AL6cP6Ellk1T
I7WdciuXhUjoKLI/p1HP5JTFe1iOJgeRHGblpaDcnV3sVZwTUsRnQ0Td5H2ZKkwOjh/XetOH4DLp
0i65Tb20ja9M2JS/sDLRdLu3vXigBUT0/IVWwrvm3n3v0SQubHUCrdbKsc2xBnnl/O9CCFuWtiSs
IoP4HmmtEyAw4Ulhhb1rpvs7L8S5WCeN/xKmDdfzBPSNhOz4AclCnmICa3RFyELiKhjRMmx+qZxx
ccWNXW3xLOz+40V70jCVgjG4YR8gR38L/72aOsD+5KiVy4WJvrbbL6tPJvHFZ3BlC0JHMV+ZTeAf
BwePOV7CiblmyEKX0I4jNvhT1PEAPIty7qhdWjLBTKivALn7d8CsTxUjX0jmlulx6ZU33Lz7CF1G
XhxslKYZJ9vxdzBJnZBqQEUqKuANg3d4tmJniRDhb9hFsNt2LRnK4+5wcXVWsiiu2wYeHvHhRBe1
LVwFX3EERdszGFBkihVgXfeqCpDsxo45cK4t9n1CwsqI1GEz+V/5yQ2jTt7Y8TIHcc5/UsXqy4dH
TS1JZl/o8ffyvZPsItjaiWxD4bGymOq1PHmiZkOyMwYlyvk6TbMtYmWRYSakMO8SUXoNfnvmpI7r
CY1M8OQpXpmU8nVgRGJF9gjFwFHRczhMilazq42vfQ7xIrlI/Lgxiz219AnBYD+/HfsZprBEoxWJ
heOH0mpPyjh4u+EvbkPjrq48XUIrwRkAhUGuA7gRaJVyNFwH8PDABWJLvFH6KCPd1vse5buKNTDN
U3dqF5JgJYdFX8uVSeoGy5cKMPMbAHEtxNRczeYK2oKYGFKYEbLAY1WDdZ43ANZ/U+6mgFNZrCbz
7yG4YwwUsKRMhlCo9E/G299bqAa41WxMsFZjM4LvYxx6rm37jr1pAkF6lB/wTSbRi9fwGE9f+Fb5
WecFIU/0RHQoI3J9u3uAVi6gGviBtroTS4c3M+tUxdVBWn3GNmhgiRNoDh78wTyR9dTaMoQNusve
ZqMfhMywZNqYOpei2W29xU9r8aQjly5WWNrJA1iZFKOFdel6gi4Hj4G00PmViwrMB87iRs+X5bYq
UhmFooV9lKfE9oxMCJ0efA+v4ObK3Y0FhJ9kbEIxs4kzfUptqV4ZQHH5OrJWyiTADKx3vyFdz0YE
/SwkEGGeYUNBj+543QKB8L/cfIr+b3QCgX1dwLz+sBEqrNEixIL36LsPzPFyI+n24Ew0zWnPzFyr
xdWGaB2PFSJ3uc4KOsRg2ecGAcSffAih8W0qa6Pv3ORsauxYJwN2ZL86h0sG+8n+ue8MRtubDBM3
19Q900ue0r8m1y2lKixHbc5n72v4dnsyTYzhPNo8PzvIrWTQqCnKxsRO9zrf7WHQ7z7QdD/c1BiH
mxCOAQtU5OKEaz1o8zFcvI1+zmDudQ8x8xWq3odTzcRSq39eOu0UzjSJU5JOXl6qND17YBy8WzON
XzamodMrAgOnpj3Rrq1Oq/qQZeo7a0RTiQf+PUPgwpHPFXzBBDZjC0icUPcjtwUjEWiRY6WWlnaj
mjtamSSMXpaP4ZBZLDpPVGYFMOL0nnTfZDxCWxl8JvtrUZAGsJ0GVWr7amz7PnVCfBm7AX9gcT+Y
ynjeSAUiiPXowbsAkaoxJa7OhVCLONY/iwWIQoSfYqKsuiuovk0sYsFzdhUN8lBgVPMSogDzfNmQ
wxU9k1HJHMngzwHPQaDTYboNpS/gq74GH8xtmpnay7Bx902QW8yJs92EUOzHC+G5VRlQsAmA0oli
yStAhHBkAVbYUSDTiUla40uzjrHg5OdtxaU2NbBHiskGPiIB4vC4tst4J8m2nMEs6a4jeoKD1cNz
C/LXbp5+1/ENq40QfB3gItZjUMRhKJ5+WT5X4JAAcSrK0185O1VV/w6WcyNOhxa0UagwAF/sE6HZ
samo0QTg0ZKdMtt6M39jxXg8+z4QWmW/2+2ZMWdo+RskvRtLQEvsLvr2BpmmMeZmyNCifxEWfLlY
hKWKgVAXGWBwP+v4zD0pjS/OKVEGqImvGBdqzOcVJ51BHEaqBJH/uFghNzVROuB0mmvX76pXZ1hz
IQiWnFPgcqOmO/31DLrNiDwIOOjD+W1KTL6dbDP+nmzqWshMx9JwWMIo7bYhormeO83/2B3v770G
PfHwb2Pxt+DyMHEihyf3DXP3mKf4HenQcQir/8DN/d6oyNHU2Uswmjze2IQmeZrRHYE6vXEcgAxu
9hMTynJcEzQRHx4vgTrtSH3zzd4kO5eCF3uH/tT8s35/ptyaEyH/jhON4yK7HMRgDgVBpOh60AJL
xIUpzF9fPOb20kHVS6Kppa9oDzjMjDLYBvkR1u7U62TSruiqrNxSBhPU+41hMQWIPIjIFIT0NcAT
O/7VreSmjHCkdVDZTba3471ZQgHvhu6RdHqpzHfn8IHQXnXS60vTqF4KwVCXdY1AkE26YsxBOddz
0Z1QotJD7Tofc8Gf76YgaAfe9N2kJpFymJlz3iMgmOagvD8cukYpAZDNzqJNfkPogVp1NtUGxZSy
5dIf4Htq3gJrp/RezETDiUiLIQ7sE5Xlt/rBD5kjU+vinUf8zf2ho5J8nyHZka8iZbuHJUYW+cs1
zD351ru/rBxjWnNBGUx08EWf/kiiqNnLYY+hicBof8pIhez35LHyCR8aeXk4zIcUShiRl7qoCm20
6y8uKe18AfqI0s8okriMUtAuGITnKhDe9TP16ZfcKJrHGz+6ZHNH0d9dW5ZaYjWqiwAkQO0UpfyO
/uDXQt0+OyjthtYHpSa9Xc9tFxqhpkY1hZfHB+PzL9xsrkFSEYzCmtkFa9YIw+R8nj5RgGz6nMFB
mKk1E7msIVpPfGauUCkjL4Mc0aNL6ih3Pp5SzkP8jnHbduT+uh/17Dl0IfC16seocF7ttyf+uwLI
MsDhPq6k9bTv7YWuALxSlT0/55JcW+HPNKJ/U8S2LHzUuUe9a07bdiAlcSupS6+lZv5cHnRehmy3
/XrBH21khrAy7eX4NY9yFu+zkHqtTyumxSl+wuEhWZEdatDtr8JP7vQ7JuSgHzKcugW8CSQwEg5t
BDofvsgG0gpOvwYAEV6Nv9WqWarWU452/ISvjeqnB+CzLg5xnaNIp6BfewOhJDeKnh0oRHsCISNG
UcHslbouVKRshSnvlmCGX4eDQwaaIOCjt8Axt3hHkTky5tTJlK2WkVuBLrUSGMkgKq8x2Lf8NitQ
6kbTLoQuajjL0gUXqKR/y+NYClVAjUS75t+h0LeKI3Z7bv1armF+m6jvK2OHyC8pmJj9QjA1uYqt
GDr7RpMiRhPee2Gtm+tylhpeN7m48B72sxoT2dka5PZnJ8MM3eoiV1ommXxqlZ6oeU4prbwg79Ve
SqGz8VNENsFof/zpEla6Kv4DQUp4Td5+FPGzib+ph2w+EnqcbEknf3CkUiLhOK6TcvO40SNDykmm
rld+MCwEGMw7ralkEST8cr4Ilxekbszf8VviA9ROn2Qdlug1VHDe495Sc+eJhDI8EWQum367bE2R
GCvxdHOP7K4NXvp/Q1hYgvXUdGp9/LG22HB6RH7cYuKDXNXrCFUHJmLdznDiKOS7tBbD+vi+YjQM
h4RRa5h+H5UET15L4EmWnOMvLqzs5gpW2aiJ1mHokPlaFFpsqxeYXwiiSpDXrHe86+f4fJgvr5oI
oUSF2faQlJRUZavGb8Q3EP65ZRtDZE0NZ73o/pdLtPZG9Fr6UQBctIENgft1a4zAd4Ic7w11HVCZ
WETrDY6+JIe76J3FYiU+eFsXoB35I5692hTuCwcDrzdoL+UeLmRSDq1tohiWdPfXluLMVCCAuOLf
XoTCCgrq62LnLyUw4tgKY+2oVk6VdVB7cgSmigfepzMF+zRWvfThEJa8uV42QALvmZQ+CGSJzlHi
42rDJtpaLLf8i1kX7oyoCeSVRRWW/usNDUO2PjSN0tIa4ixl714V7j7r4OtdrB8LmS+zTwdIE90B
KXKtARuAX5s/hIoiLVbhQdG0FXBWzpge4w/ERsIY/PjWMSwYwnd59jV/JocqeNaadYbqMbb0Qp6s
wT4pq39UG84FvleOA5TvIdxtcFxfOeZlQHbYxh/Z8pMH++dJvarfOpyRbnCbxxMxUSvVZJaeCJKY
xvZZwlB5mEpjEngCfMwDN24PQdvcexNU2san0+Sv9qOUHiN+R3tdJHCe379ILx7N9+zr/l3t1LN0
omS8vmeIwRSW+BbLfTRKM6JVXq2Z7Zm1ILrLIdrzY+e7ypKqAKqAzToklbUi30YQgIidnuLG95i8
qgzwvbXGusc+hvQl3gMPLdCo66PvmF2nS9pxu8icY+1GDBpM+e/IIXWQXPGhq1b2jGnO4JBzgq4H
CG3yYj4IcLGEgqOCOHXtqpZwwe+V5RUDBLqeieaHLD0n1sVxHpZAw1Lhqbho9leCe9jkih9y7Zab
JG2r4ASjsoY3NfNi1Jhj0u4Bi8wrLw/nZIUNwxxtHMVyI5x8P9tvg2oSQyAxaCxZwzd2Ysr6QvRr
dPj5c8l/T7QqGy1DfwYUTAbYDWhh3numrVWjMqG8ilSMCBTA7QcltY7/dl7LBN1t/9CGsikSrGzM
PJDVSkOqvxEETI2JBRSXFE2bJeWpud/VWbNmA3H1szv+iKYlPhQ+THPHltcTns+NRnF4fnLZ2ykO
Pwk/nVQRniMm+jAzm94VJqV3NZUHc7qAgBOpo+JHYuz0wi+o2k1hDyZTQsIWILqrx4z47WIQYu4W
p/r14ZDeTMAGYjM3U6e5LU9s1rQr7ae9p7QcznuFEHRsTkKOjK5PVG/URBojc6BdZ847tkSyvzcw
5l6zPP1m/f1CkiUMMuwX+MG/WYAt70zM8zW2Yv5DYqft/GK9MSlVuy+z96+g3Vh1epEPhsfZEZ5C
erucA/ma7CHkSIE/14MPPyH+HqS9GfWNm0R7D+5n1IsyNa7x5NNOk/k/axlSdao1HjEHb/kDou7j
0AsdbVfczCddgdXlIW6D8+xvwWyxKel6hNIw+zbyURF5WxlTLSRpddr8usVSRIBML4SoKjb4m+89
KrS3ThvCVVQ4o3O25fUmFU8BT4OpxgQBVYF1dF9it5zgtN0aLSHZ9SjLoB5ncawLS/PVDkr7kVb6
zVfi4mi0G1o5N2xFIbFcMvXKUj/tvzz0+dSiKLtP3ku6hGCVHQ0GoAGjAGEjc4936g3y9lk/JzI9
/Ushgb9CNVIcaNt0d7STzjJK4O0QtxEIRx2oObRLvfOwPcN1AtWjCVLlNNHSQ4iOcSnAKOyRFq2y
bFuh+2qnh6MUuiNxLtkfSI91m9LbBFA9h7R6sDdWDCnDwVVJnOvdYTJMkbAsiJh6gf7cqXVKkXGX
gC4Sx878MSq+WCEb5Zq4AFfj8R2zVaGaWMf9evrQTTJpCnaxaTUTIFTBeWiVnCIzIMVV6BlUs8Wy
0gthu6hlLuCfidVNDSv7rhmhLgX/eq/pYMD5GnEsh9hX0sNvMFAdnd/y+gjrqOWUGYO9F3OrqGdw
coPoLXejtT3TC4BPA+3m6+TB93BjzLw8gC7E4HcttASunmzYHZEeOyvxVF4PXG+6VL7ndwvRWbRZ
fIDcLenUeTh8q9ngzccR0KMx2gcxQq6crI+t6DjF3adosTKQpIpxeRlhcLYhQRPbb1J6zH5aagvG
opwr3uGcT8DD5+ywKFZHM6V3XjhQ7FYDLntEPoU6UOxViI5CSctkwb0/wr347E60Q/m0xAvbs2C6
LYRl4hgunpwtqs8T0Oe6tuhh/5Dy7aSvMfAYHt10x/DNPx/sS8D31LUCuzsgoDg4uTIlXI54pJ/o
xWuUTPQUaTs6MtygfgjHnbsbwM8waPvWWca/WefeUG3RfVdtkwL7TuRISmjCkGtOufrhH8ODJbyP
MU+YSQPMavtLMErGqNVLmDu+PjI7DMB3QWORELxB5GAU5Yo1Wu4BKCuKlJOu8aIkOuTFLv4UCDtP
mJXZHFBqF3tUDAv+YRBYk+vLBB5niTEXTWdZlZsKDyGD/N/nrkan4Q7cavnjWhhsQqBkvg8ahrih
Vnw5SG4NcM7aHBac3og2MnUBu4Rv807lDsibroulXMnHbgkc4+hMxK5MlZtiyGs8oq9ZZ4qG41pq
qqPj8Z5FpUAZW0PyvZSd2bah8e6HG7z+BiAaEMd7XXGQWYGEZic2ZPViZjmLjhtyYzUOULTk9Sgw
BYZD5i+nmDGIU4X8XG54DbiIH1tk10+7Tjwxf9lOx7oS3q/A3xW3t/3PAc6KVMzzLhnZ6SAke/lW
y3AHF1oGqklYiskftbn3Ss3srdu+zm87bW7+H2gM9yfif0uJuNFbkfuNBSRpwrn1NKD0mj7dH5C8
ArSMfgeKXHdDJ/l+sAotvISqy9MEz011ILhknjm1SV1FTrj7Gsy+t7anZBhbJJtvk09/x7bJAWUu
w4yXZI+NcLVTl4PtUcycStiX9lBuMgZdUoUvhTTpeoStiSOWB+AKweTsmv+sB353AJycBcRpYVz1
Fz5AbRbR+Q80hpdFCdJvuCQ6/qfLOHud52JzM6DobT6TAjG8xEwwzqGEHKFHNpxr5sgnM5dQCZ6H
xvdIfeMgya+0PBePkstk6A+5lkMPFp69xSt3IFrnkMCbYyO2h6cAKb3YOC04RJE+Qs1g3/s2yPWK
HSKiNrotmBVXq7uxi0odCo0Zhz17kOxanfPgqvcMQflWtC6cjzM3dFVkgH5NVZJZ3h0C1DHkU4Yg
Igycf9P35JP8gJTvkx372raxVhHlo9ryO4pVdc5dWKsgf0LJc6I5MKCKUfKrzUeD7xORBcjEL8IC
11nnKwQgx0lZR9fxUoZ5jQAjblQ8AkM3DPf9UX5H4qKz82i6JDIM+eS5h20iYrzOrxUciNa9UDVP
VpjuXywzzJeRisrUAhEl1MZZN/ZdXA3kRs2E51sVowCNzBg/RLL/3rgmz3hIII6FIsMCUreNm4Hy
Zb0aFlZMDGHbWvRbHHgjxXD6gukwC4Cxvha5N2r4Qppsq3NcHTTADa1VTitNWlYZrs5kFdU6XwB/
d1DZPTIo6XBrtHagkEB3LAxjFvZXz/yRpRiSOH4QmL8VZbUdKl/9z+cRykHIdtemd9mAzooq8Ktp
bzkmZt2N9ly8MyFUN/1zIo0pipX29bj5bpTD+xgQLdaffSGOiEYpb2yK3EeMWHaz3ZENFZpTu0MP
Aoqg7kiylOe765ovW7zXcA7vAkERW5JF37houa958qG94f8MplDDG6Kjev/4gV9kXZutRJInQWPm
qU6yyMOwts+QQDIe3XZCcy2ITRfC31QyKaS095yg+yqq8PnRXT98OATmuV5MLc1+kx7YX5Bv76Gl
mb5xS30teUrIrx0xOA9iSv+qnIzZbbYvyvF5vL0Sv+ATq0L4pz0N7wD8gyf6TnoFDv1x9IjxLbLt
k0ubYIGY9tTMBi8GqQtg3L+BhggZnepP9sBITZPLbMBuN+kIUKY59OHbtyvGgcWi5Rqm2fJo0Ls8
NGR20p1n2DvPiyzUg18YlJQdIEU8gmjP6c66btB7eQ0MtA4m0olozrCdgitikjnid+F7dDh4pVCq
5eElKmJfufeZLGSVIMG58cC+jN6gPxQ8WWCtjz5WR7tRC/bXj6Gp6gGQjDQ6/ttHK1jvCvxBAgzN
kInIpGJqYethOIl0+czcvUVSNhT3zmktwV0+XLcdVg4L/hldDNrTNghau1DIFOcpSPtwenLxhukH
stzuU5GyqKr06EKwqSOMWyWdlHZsS/957Y2TNo0LWYhiekxYpMtNkoJJ0jrt3fhbdl8OzsugjRf9
647LpC0MG9rQUsAtikyhnK08ECfdxMF2K+iYLwEsCHrmc+1DaXE72/T3TCr6WeHqP5HMMqDnf1BD
2Meswv3E5zce1s8hS2ukfBlM5Iwmbi9vx/3Dd8ImEsfIGUgEyTCTl0WVi9GWXeIDn1sIthsWWhN8
ETjnJKzJL+GGfbjUUXEkQLgN6EzxaOw6Hsru593SeMEOR1BDKqoQXQZ8RhZHcNDcq0V5CZjawAwA
1j9F8CLd57mbzUyrqAHhomHt3SJQm7NUnzr5idTKqCSBsoPqeDv0zjXEc1eNzf2nPPnFLji6WTGc
H0gTAcbeJjTEgBoz1V1ST1jxSTnfxnxgXEh2QYlXu9w+PDGuaD6jOeLKu5wjA+Hgs4/nXfryJFKh
+LlO9sKVKlyjzEvUxHBly31E1D8dsEaSQ+fJbu20S9q28s3K/hJDNKDj76cuQWrCONb8Gqc3NxC4
2u91Ixn/DfoccS68pg6I2XuPsxE7HNkoxijhVrkuKGFG0NLKlPJQ3q8zVjYAsnUvomL7kTuM6wAl
HLirttUL/R/IvGs3ASZrCCdCA5d3sdu3cPN8O3DsrVsPZrXgMi4PViY9HibfcWMi3lirWJhl6D6y
QCv442y8exf7TcLYiVnY0QRfTTBLVhySrLxkiXFdtzCF9kf3yCgXVxR5XqHhB7doh3GB8xup/vqk
KoUd68jsr5VRxO/okzexUFaJaPqKtTJ6gbB0TcdjDa0EvSIYF4aGBf4juiSta4mX/kUpjNtXuWKn
eUzjGFRgMWcmqFfTIWQQHvf+SYzTl3/lsZx5xa/c9kIAa5r4rvmmzD2N2ldHa4WOLhMOTfFh9v55
6DM4Hv/BD3owHLebXVr4GTQ16TIzNjzTX9MHAf8hZUvf7EvKhhNFfFXyD0HugDF2/PJnuDD6WPLq
/wnGwFrNpGDPN18q4678MltBw1lDcgI5c2iTQez8YNLZqrNvJHJS4ZQhj9RrRGVCeuSon6fbLd2K
aplrJ40Jr25RRgrk7uYl9reIYh1yNbZJYMW5DdoG0RB0BtFem+RWMKBgRRLs2MZ+YiPproD7n8h4
qFcuYZnoC7/zX7cvlYFFWkWuxFJOtfRWj+J360TIbZv5tGxH+k3pCXFwVDIZhc6c1zUWiwvvesHp
U1550cCqazQ3JInyJnpcY29Hc/M2oNSghzCoQ+aE8iZQ9jxyn8esYPyuTB7UziwOQLcwowdxfZoH
SBCO8f4D4uoh43I//5b7mYTKPjR7/B0261FpIgssX9MwUKrteZ//sdfs1mbfWhTr3lNKC7putLJI
+Y0EksueafRYEMMsOln3Z4dL9wh/Xqoxrecn9j6Eo9yhcFsdwWeKjyb12h7gZR2CBQ015zr5bGre
e/6MIDawjX1+MqkUoYYK17WrGPJpzTJwR1x9XBEg4cfufFIgLciPNtGj8kSfo1VubO3G7O5zsAeO
qmJ5HlY7mkINt5kBA8Gew1e4G5gzGbEH4R4ER+sGhOZuN8172KfXS0QoVx70cbf+ar2onFs8Jbm6
SkGDznvAvDE2bkLWBPp2s/8bt6H97zr5AaetvHC6AMfvbHhbnGHHmMREHO/XaeAki7IKjJMM4drN
4LXUrvG7RS2+U46SmblS8+2q/bNTfPSp3+mNYbFZ+E7hLo3drr6S3buqxn6C0CvLupsdXWG47nsa
fI+5BmYKLGMmVE/kjUjcnk39RG0ylNdSgRyQ6VM8oPSmS5Eh3JpQSNArWUlfBqg9nKApG9TkShEB
aKHKzFxX8MrKHLQov19FPuPAf8po7ehNZ7iHeBx5xo74SulWUVQ9seAmX1+IVLxyrlT8IYIaUcNi
2HbGyOMM05E8imB8rHr8CUOVHJX/KV6Mc5TJVjSsaDzhK5VAjsIWWhlUVBd/6UCW/B8xA8LNWP75
ZFu7QIS7VCCbRbEjoyrik7syIBZ1GBND/3/dn2lzcLESkFt9NOSeF/Qu8YyinusZ2WZcv/BdqDJk
j5dtC+SQu5RKQ06Og2FA8CP7A+KFhCr5mv7/jTMUi8iAAxZ2FJ0ZEOSQ951zElGtbuDHVVtFYzhO
zu5Nhbr1GzWA7HlyYCxmp9f8K0XJayDtP+nrNrdgiWuxkuW6F9p1wLK2VkOnB7sASI0mx/68t4Uy
AIbDyu2eTXejG//WcAIcI7zNw9nyDw9eogrea0ZTUYkrgDpUgbhI4dm0wdSejYSLNM4yYPnw3VAn
Z6npOpfl7PM5Sg8zkkpVdN4aUnEnK/bAggPkTZ4JXUa8n1SIa8bQUzTrGa7tWfZTPqp4jxeoeo2C
HYv+fRGUcAu/DlcJ6su7Le0y7z1fDY4YMWUxN+huB6PLis8pg3FhFC8zLqInms4eyrPxyDUxWo9q
bNXqoZhDibqoV8hRbktdt3pfSHI94R0YJgY+t3J0EuEXG8wvuA/Au9dA1DnzERZn1stj0qebioug
bKWNSHoGL/PFykOv00ZctfTY/bKh9YRXrBt4yaJa0uHS7ta6mdQk4fxYNQ+cYn7E7GAZlMhTs5N6
YfY/pPvcOLMKbB4wpOvtT9XgaEoQWlAORfkFgW959JyxZrU56HUF6cO3v+YWUdeyNtfM47m1sAw5
9GMfXqcft6fOw4b//fVluBdX1AMInrXTSDnldp9643SQJ73QKrwtXH0Mn335s2fcH5ycWFCzS8eg
NsaymD+2K9OiIBui8adIPVy4o2ul+9tON4caR8bqxepQzBLDL6OEMjvCpYuKLo9X2I//XR9PqzcD
P1Tr6jWkc+TyvyKy/iSe5PfC+Xx5X6jtr4Y8/zS9OjbhOLkP/AgcQy1+M+ZIvtC93K4tLcSZ9RK2
YErq2ldYZPxHne2NT+WOUqasd01PqQU+D/Bn2HodTJZC4idupkzlmbkZbij0jN7iLR5qBxnK3TMb
py0OlrdY0AWiuL1LvjqZwkevqxSyVM1n8ZunK4ZwZcRopE39jI5ch+eXVMRuurLdl4u+4057zbU3
S637lh42rM+miNIepDhUzUamBuYKYn6QJ/x4dkZOyGcAniISX1DA5fdVIiTuCFBJMGdlsoLZTFL2
utyx7uMO+GLSsN9Pd32Zp8t2d8Cy8mJNGASoTnzf6PDfMxOooAVvQel/Rg+aDrh+YgQhng2toIqr
5GW8ArAd8yg/eXg1SGmTrRa803Z13JDLiXievBX4BZsHCh5cQ9uYVMRQi+A6a9DCY5uNOW8Fk7Rv
ZNbcqff9WoPCiLYFoS0wMoDs0oOcaOdhaULRg34Kku9U/o4+3F4xQLs8dEGELbJ3bdqdEBxN2ETN
aMKpYi3wiCmCkPfVnwe0UlfWpx7DsW/b49C3ANGOL9TvKZaxHVEQjsose/MGKgFEFI7poAYwHisX
APIqFuAT9Zz8g/XuGaVsUF3UsleI+qzmoiR1qYaXasOco7fiWsMKkwBnku1nDz3kEnL48bxxVW8P
ChHo8jWkZrLpdSqshIk0r6CayfOzvy2CbihlLP4HUd+OEooDHVpOWvFarw73eZRVXeMFlArPINPo
Re2fz1n6uA5lnAbm18sykyrssIhYfkXUhxNcGXlLJjjACP+xx+YdiOY2lKGZEm7eiqLPEns/O6A/
H2ZFofkDYrKDDHzh72y3SuY0ja9CwH4GFJTmGkr2yVD1+YnXylpxB22cJDvQtV716Pc7v7tS77IV
BF9vpneqYr1U1/xskxL+zoubOhVRmdmr+0wHpGuB1CnQ7zGEboD4BCtS77Y5GDK88W2VByq4G54k
eSB+1Mo4tAS5AEXlpUaCGzLJmQT+XfpuKVOyXZJUHaQC9shhHrF8sT/ww2nR+icpI/HIAQqEeHYc
8buKNNGwJ4Wr0pHClWjylv79tLbvaCwoRpcQ3psmOMvFmoGWfhSbLSwGOhWnzAKVVbOPGn4XM12i
cqSkR3HEEpSTK4vB4jEmDs5wY5u9klPaY2INoIEGPqb9x0n0HQdMMfdNaXJ1GcgdvRf56vJeWUBG
xGtOLQGIKt67mU2yjOg5B2iuGHt0oIl+Wmgd0UNpYepOnAybTcmQdhoJ4RHwxmS2KJzPHh1OVgpi
XbnOQo8VXTYXqEB7R6AhRqIptCjX5BPm4vN+/+mUIqWqxTjYVbaURfg8AK3AYpbaJIBqWtA10BqV
iGoN+dVnKXaRzcrJ/xappvhd8dqEH4FPmDDn+8uC5wb9nhYKQm5gGub7R/qKlSBWDlwn1YX45UHf
BrVXSPrz87ev2NDQ4erOCUwXkqWQig2Dh2ErLq3u3Fp09QA/DA0+LPLt5BGyLXRqhSRqPTozLj4J
Ag03Ucx8oZmK0N+NoUSsh2z31GtdBi6AnLBMBEltk4Kp0DOv11XjBTeRhw8xDALt4uZD0HSwW4NI
JzdVuNibnekn0ahZVlKLoMn29Lf6PfoPmdsMFzf5wpe6UlLy2e4r/mhkI0i4Ksmv7z948gOfyU7P
vA4/KN5DdZiu0AA5HZolX67/Fw1GAaq8eOphpGd0VLbS7ugYpx+i4PafBavLKoUpe8SZ7Xe2NO5m
CfUkWw91ao7jdimKVWVUC5JnbYu8eKbD4xoij2hVuo1qUjrMe0xZWE8NRb7f7efTDd03dmlk81Ra
FtAk2mKo3MbpVTRXETTX5k1FI3KGkBqlv8xbsz+vw6FwZc7USuRVwDHCmUnG5Qqo+5bi3FWcH8cQ
T8fswsK1qlEDbHamNYY1MTmjzTAFJYHsbS77JVZa7YnFFMJvOn7nmwJZ54qDqzLAjQP31jhM9E3j
+VE1CTSRcO9cgHUpWsvYN+nT+TOnu//7yHizYIIZ70FcPYtGBm/rI2I/KceGVHKEYjlVaHvCeoLV
ZNcamDwHgFw5XVdHSZDuUnzzpXN38BDSb+E4fmysMpG5nwzSAf5P8WpLuZW2K9RXmqfFf385v0lz
x616+0USTp9DFXMbiC/FXCsEiRxp2gNz9DohD0mHxVy7ScbBerFXqUq5/YlG4uSqrS9KFtq0ZGpE
6dO3tH2hX1CIS7yULkyOo5TPSEX3XgG1lBaKJ4SKASXOM5e7xfsStPyU5wDUIp4nRtpGkiJFYeRR
ZOHeGFhXf4TOzY8s3s4gte8+h6H/nenfr56SMEv3XE04b+FUpe5K/pJQjCDOQuSUJqT5o0DTtlfb
0AW5KC6SoBlBjuM9xpGTX5OyAfarOa3v9Yr9ctVfbAyHoC6tVmE95dK1DXUENmyxWu5ZyFPMrn6g
EmxoJv3c/hil2DieOo4bRD8+kgl4Ctz1ETt/ynSivxR5d4HRvkOtWe3R5ukCyUlkY+MG22k0F7FP
EriQrmYZIfAxhcTBQnN9fHGa2hE6BmkAC8hK4xUFiloMkepuArAZD6AjciCZwESzLgrxcV1cAZNV
JlZR/7aAKpMLBFFRyz0/dO8C2+ikxZEwAz9NW0o/H6h4ZGcZyDLYdOHwSPaTtZ5g/FH7I9wf0jqn
gC/FYrwKk0+yzJuXWrf7GJuYFuVrJ9Ki3X7OpsapS4BeHhWaSne0GXSzQM7l+UDKEE2TfXArwKak
UWVRDZEu5UFb3rIEIXdDGqqwnZV8i+Vw1EyXNZiP2YipxgykJH2Ayaj3Jz/yI39guOFG2KzoXwiH
hEser1uE/WLD7fp1bEGvpi9Zm7758UDiQzQatxskcpYLhS2TkpYnRvmEP6BihLXwsPc1W5HmhoLL
lgp0T1BKxWJw6neBFHBon6yIwIIYd2s3bUPqGT3tryLiBC12C74wATx/5GNAIMDWYROZh2rkKi7X
Ony1eRiYba+OZbwlEO/OTTdJp4P3UGAi7+OkiPo1gHZrp/9yUYbVzg1/VjueXZlu5X7OhHF1NjGB
xoqFhZD+40gRAWphY0jA8IQfou+wJaf3rDfwfEq9UMZd4bB6OE9beNFV2wkLTIv8a9/NQP/fJru9
GlJPOBjCeqrwcmmJkeMOknIu9pfaGxXaTHJEoKws2mdkFYm57w6P3WwoVQJJO2t4SGzNXRVabp8g
vmdJ4CBbxhiMJPcs33oMhDPvYzc1lhCDGfbV/wTAIsUZozK49+opgob0/vbikxuTS7NbWuVw2mCJ
daW+ZdcSfBw64Uk53CYQuCA4N1so+ejhhB570KthklwrP9AEAxZQwIVgRIhReF6BAbAAkUvO4Zxr
FCwQmkugj9xW0tIPPWgn4yhYfBOV5FIWhf7FpelBFVW5v7B4NMeW1OTLO1n7y12+AqMlrJmzMVtk
vWmbPG73ALBO+OuLxLbVJI34YCOjxI8FMfwSgCKM5KfYPlA6HFXj8Pcv6smYVHZxKUzpReSiNgfR
Zbi01+Wkfm/gPaDbcgAgLajVhbMnBgGM0REnzstFP5HrQJH7IP/OClluGFW1/DEMN3752dtxRsYY
S8ubmH84Hl+O0uN1EhfVjnNKiIsjtbD1MuMOOHQHZv/O6H76QHfZ7hIR4bTcldW4zypbjgE4pwp7
LB4Rk5bRalNjzbzkpOSdXb7T6C5DZhQFYNu1R8Ixg1h1ShlX+VFZb5aWyqPXhYuKcAckCOTHoWyd
GM3LWBwPUJBgIW8+1LO0FPIBwFJCzKImomTiVIvgsEUWlJZqHat/3pkgB9C4AP/ivH7MPvJRDeRc
B67LbnR7X3B9JJhK2EJihO0VVvG6NNZBNpkoffNYwEAK+fxiL7KK9dtqKFdKs5GjTncpQU2RyuDf
/+AfV1VZIl3iE0D9L/yUglNXaQDWBK1oJ3lPjCyWoLBZUrnIzai3EN+9AVe306SxZSHoN71cRx4z
LhulJFdV23h/9ZYFeuhq110fKTPLNv2d2v2wvoPywDkT6SS12eV6FOasdte8dxLsFMHnv4DRLlBC
PCRSD+51m/veA/v0e+BH49bxvmIGw4m11Xd8L5LLKvcShjjnRyi7UN7gJ0M9fqT3f3bPqlW2xB66
td3eWPU8QEVUESS+i4g9LFMMczI/cMfuTZhTMz5bNHFD01rDd4JlFhWgC9gw3L/pwD9MH3/MUVCS
Hs+HfD8Wb2zGlD3YNBnUnzXh+GRaigYcvmz8t/09HS1JQT9M0Ty8HNwL07netIlGALsZoqMLNqpp
Ne/7y5aN2m0GX7RHWeUT9zUkomU2/Ud2PkA5aVT/F0RAGK+rCMK4OBsdqUkBSyoBKRQP8KT38i7u
N5qIg6arfT3rbzAqu+CV5OJrl4ot6KTRlSosm02KdrbwZ35dK/qH9lQ9ka96LlL5dMg4aLfWPrqU
VC6o2XnykMQOPbdn+Gnpp5/sCwlu4pv8HK3tsLO+FUQaeRod0VIMfweIFO7bY95TSmmPYmSOif0J
n/1m/HYKdsOljt3sb7yU6s9C3O6ZAiDJYsY9R1Tj3/2PmnfejWiw+8rBq/euRZ105r2JXVJC2JoV
i+zcnfxyT63VAeQSZhQroopNdU8tZeNQlA+p8ZlXoISWoi68lQ9qsXd3QkPtkAqNvmYt3JKI0zyo
hxPf7D15UcPO/e/vn/5uPl30mrk9+jLYcI8IaDh31Basb16eXRfpo+bUjMYSb8ECCutkG+odA6VK
jntrTMpeqhJT6RZJuSeNe5v6jQgAQxNfweMw4WZuVUBPgqNvI0ZOLSMtY76f8qA7OvxmGE6iYuE6
phAbIg9Jzo6xPoiUO5ZRg6sYdDX9zrtDqcZSht3XyDSh/uU/VIShu7cd5tcT4rQojERAQEorWCk/
10uTcFeseEDXnPM0judRTAUX63sno4Bgf5xeLCU9JURromAeECbbXOnJB9ZPmYknLb2qIynVoi2P
O9aKk5yew/gHtkAB6u8PB+5lIo2AdTtG4DG4jxHsztqcCAFDw3gMU0HRb7Mq2wmAxmqo9OPlvk0/
znbuQWhsZZnC44hMzSMcO+5ugh+nTTaY6grCMlmqXzp1kPjHZFlXFAEhYlQXRjj94SKtDmQ310eV
I4EShkBLUkgS7A+QiLVw3SW9aqL+2ECRnqzBlw+vw0rwWJ8gtY5h5TU7hNvyCHmsdDCwdwnsnaUg
LJan7FwfQ049AmGNnBeQNtS7KvaaATkwYe+lQAcpTfnkxqc1gAVRoi08PNEiRSUehr8D8j/dVKg2
VtnrhGe3gVV2EUvqtDcM41KZ0wkOQvOsr9M8Fbr8EK4ReXF2ime+TmE6qdEoWdXmTUhdMcH9wNVI
NO+SW/GdM2K21SBME/9GigOGsWYa4/yd9RAKHUEgLroC5HcJVVmhmFZz7qhRlk42pfZf2D4lAip4
HPdGX1zA99LjbhnOI1aCxa/PQJLIH0+3aYG38qtXO2qD7zhlASOm0FsCg+6u9U8OCUX9apE8t+rX
iXn8xEPZ3sIQRE16hYochEufcZMmDT+0Gp6WY+KvQtRTFS1wDLVXngHh62FSq/Qs9QMKpvuCwS25
qOF/OzS9u7kJSTNLjRMo/Impt7GM8BhioBDyvMh9hbVJpFrBZIosioPnXWNyj6Deb4vStOaIUC1v
W1BuxidZhLK0OxQlbpWo8UtJ0GjbtMuGzUI2Q35/5LGcNFxz50A3oJZHvIx3xc0k1Ppsp5+b1HCw
R9C7SX0cLd5bZW0zSPXb+2RCcXX3evDgSMD2G9MvQU2YGByD+NoAT+6MKXKI4qGbWzS6jIOvLfJ5
3MO68LSOnPCt84DUX9P4Sdu60+HyRDcbpMb+bVtmB8/CdUhwyamk5DrTAfmeXFZQE1qmh/Bc/S/1
oyJIyuZzSiksNZFhQnb7c/q3TUpFBAj6DqfCRqI3grFRy2kHkq90SznaZcgut0Lp3cX17sPbYfpM
biZWAqULVDUbnXRmGLmaUVqe39k7CLrUKvhHuQl8fED1qawxwLtk3cVV5KEO6x4rTKFLkqoX+/T+
aO+F1RYNJpRFnxATWCutuS9H7oseauWNSUlgvNhZZJVy9cWBvDNfQM1+qTVMedT8ooUxBoa9XcGg
X6n9qgwR5s4b+vzzNzJfhNjooWvQZN/em+t9nPNWYLiflzolDKd+HUUS9Gogi2Zv8X3KHaAqPRXR
gCOMFbN/zTTuf4gTAHN6pIoEHGZKAWzoHCQz3u0eWwuPDvllXllQREtSmv/cixf14Rnf0LXxIdr+
gBGO05x9YSbPSw40yPgrqnzqXXMuwOgNZpwsQvHBMZe5mYce1j/hMd4CXYzw6nHlmYbInsxpmwk2
l/S6C4HC24armkfXh1HFGFNOlU1fof6qfYNQ6RCOpjU5Fuh+BbC9NPHljCO2hNPN46NbgiYnSe12
eCwMvI+N5DvRBv3rNg3K8sX1gwf8xVs1P19lZeYupVgKqtL1phZo6txpA5nW+jErNRLuWWAa9enZ
Wi/ZYbyUWUvz7evCLlU7U4K57F5zyGzUlwx3cFoA/0qGoPozI76rsdq6iCWed5l2n8h60e1PRCUN
6Xemhd/8B5cEyuNq+jQvf/wFhZEWJG7cs9+GZ7LUvDKw4d9+q9qELNdCs9Qw49aWFiYnXWvUcyFL
X8Mpasc0KgiDyDvRe98SNntMp30uhL1WgJbAvebGcHABQfgfi1A0DA9QGtRodh3CwH6/aXHQSULM
zasx+P5LT8hv7E/Mqx0qB/w6OYs018ZW4OJFi1jW1nUZd/psjki+zj7cQION8ncsyjQHJz1VbHYx
PXPSg66nyGDcqtD2uFrR4BWBtPHe5ncwqyuvgjMmmeiBVYulnqB0SV/2YpZYfob9AVRkunVHYE22
CXRPbM/e3XX2SEziWTt9zkTncBvlLkmHfHXw+3RKBih8mcMeaTw36cY/gU1qC6KS+AhEOTv0RvcU
71hWAPS45BhtVtNOb8wTQGsqyxIaQJY3jB4hxcAy4cSGzNFgRKrqwRXbxCUZVpFYJE3O5yOMYxKe
QFe5b4njFXCEt6UIYP+Cp8udOTvJa4zOg1RcgRIemKoT0hd2VSPm++hgjIjs8Zio0XwjAyXIlxvv
zX1fuYLXVmEgXl59Z2tXQShS9dkGArXnM+gkBvLMAm+8eCS8TzPWFs2RsUVP3Z78+3vOyzx6fy8q
07xJmiPbUbM5JjBJijZdY7Vv6uzyo0TO1Qgu7N0T/scliADcxbMs+cuTe1ovUpI6DFqUos/xf3/Q
5ocTzQ9OAqfEbpEEx8AwDRSYhSz/CbGR6CBALY8lPQjox+0X/bmvMQ4NFdzu0mvgQRyh/Pemv869
R0V4hP8d5GLBqvvKEmT7Waw3gPKdAL9NTeIn1PmW1D5ntEaumKH4yYIml2d94ah/5Fd8VmnJiOdA
rstUglnf4P6X4uyGmDarW4cXMz+g62TYfPKm0WkDAqWvtu32sQbcIWDEWV+Wam6XA2vgx6XL91gz
+DkoGK8j/HMMut5XDNdYmd0s0k22vhUQOHf9zSD7ED1wb00hzHXrTh9/+5wYks8k7vBozsyDGe8d
fw0+1ijS78ETn/84E0BmMqhhOczEaLVXEica5XRM/V3iuED12+H2VA0J86KmvUt5kOBn/yTXkJtD
KUff7v7jYsFpnd+/CAq/27qlUtKpyVp7HwB5Zo+4F/IxQ1pPOEcoZz4lhRwvzqkizXl2m1QUdXTc
HXn06CavD/TtPVm0T54S/eSmSuFWincaSKwj3ZE+F+wwb99hNLMRLnh/LMuPo5rc5IjnsC1qFXb9
p6FE5mH1IyNsvKdFdW075/WazblVlncnqiJUKKaA6IBlAXNkG0yRCNhEndzubHKKTNml1RcXT9kg
0GIeZHksTWdIiTRqVMEalAie3TylyItZBZjvHq8IC0EqvTG114DuamSqDzDaRwwl2VbidQUNIXFB
R0fwoFus9fuLlx7T05kz09T9/zXbJdtm4vNNJAOcAHuzrGJEiAdXG4IJBgBrZfeMTyVkr1XNAbH1
b3qrEQ7V5Jhh51U42EXbfL93JqzqiSjMQ700Ysm5Zaj17SK9QPcrrIpm2s5QfPja7dkDp5l/0W/p
7X4fIThQOqqJokEjRpEuNQIk4Di7UYvd6U68bXO5bCihPGCDpQWKs0YqXIx8GfoXHGLQRC0kClxx
Qzn8ZAjGpUnSgoM7HxOOWuAt0eZ+3h6RUS6h7PVQ/rlxvAhtQE3QW9fxloO1obpjPRWpk/wLdHEO
vzh9/vUJdGnsDk8JI90+GYsng2K4zOS/XctEslmt+54d2FIzx2HY1/1KCBG6SJu3IhUwxrPV2Ku+
49cYHxog/pe+b0SxWM/SezKIjVIce38RpJXIt6qusaZcJ7TUTmU384bWfUhn19bnxRFbW4ciXaiu
0xeAuTn6Xwjyvpoc3wBlgpmsx3TP5bx5a90eYYTYN2LEgKqYJxKB4eGkfC0hzllHKYeDVfaxfbcS
bTDDTOYUTfJXoQ0Jh1XVnYXcRAFyv/BY+EAjN3272L4K9VmtcdbB6el+tyq2GyRIHUFih606C216
D3gWu5sCgkGWD/ko66I5bUnvBICZEt8yd/MmosnkLYR+AKoMGnX6K/PHsJyUUxXv10njPZ1m506y
KOLxfbyt5JzXiewq4ooaKK7sIth+suuH/R8PIDSnPyQAT0J/Ho0PUVGwHbgA+C6cnIjEM3Lr5hEq
gIFwlXvtHRkEQV/SDOBPXvv0Gj6PPujyG6qWYCVHyrOJZbGjv4r98wERF+EyQJd5ZIMf0Mc1+20E
xZ3IHCzZNQyJQ//+/G5yAGCYeyztzbYfIkWw2kuAfcTh2dMVQyCHPJdf023o1wcgHGetItbq0kNz
i+1V5vrV6+7mNN1Yz+i7ob40DRlx1+WdC0QKjDas9YYLU683JmmSBeONUa+mWF4ytEOSx37Tqz/3
CRObjINORfPjHR8k7nGwdrSycMM8d5I6SAEVEelJG2KbdqKaaR+HMsc9uFdLBwl9N4YVqn6VH4PS
ZZPDHQmcLPonRRl1wjwtwZ6dKWGYVSZbbSPyRMHjRphIKCm9naWsH9Vb1vD8txrnEuwQXRtcxWF5
mrTyljQohwyR7VgHjxyRRL2lFlitdZTwLx7bhjZcvBTRn6DxP9lAl7zwzvBO/z8YAWy8f9VZopHj
DW8e1jVJ/cH8JHk1w7ndZVbapu0JTmjDmzyPNK0avtQOqUR8M3vdMZw5Fugq8dQ79Lkbvyk1Zh2E
zPgYooKpPRMzoqFzhSgWqm0lp4n2Pyb2g/5CfvABKAfFBQgrBhpR3o2uandvna+x1LFKMILKLFhc
fI4f2KScRxKtcyZBsSoSC+DAKL7ECVkOcofTRIbILc5uRhlodlNTeNRZQTPziFEldVCudRJngZmN
7ABRWjeeT7GpW1iVCs0xI/0Nt6L1AvId+vihChvM4sd+wkDJ/vVfhhN7G8D2CZ/bZhwjd+rHx5f3
iJnRtGAIhEo4cn+eOV7BfgE6N0FXcWBd1qR4fWDSjCnpq6TBrl9xq1BgappULja6w2IOBzTNwRz7
HF5jk7QkxbwGAC1aj+hsISOME8bDRjFrXqxcbRBhwI+9/21tJf8GHwGiKX5kwoKmn42oswroK8v5
SJLpZkvC0AJLhPQtJsZ3WoK3xVZBcZR+CNKwilygHJCEo9F88voxL2eg/jxGFIVj+08svvfgF4HC
lRW77UHDMnEKZoEKrNGWGq1oIT/9pWkUzyIYJLf4IXTOVGMbQCFKrNhOPQbDHKsFu/9utFVUX39P
shXLh2F2swZU5/7xjPKL+zQgm7u8GW7tL/p9ri3dvIwv331eX0FRCAiQFu5zgjRPZUbKvbAvnFCS
H+QkOzvPq6TOv5XTNl/U9b2px99aTd7yyLWmT2NxWTvjvEn0D/g0QyltMXi/PZlFmrvEY7qArOcm
9hKgZHsKT2tt/t8qceck22lE/J9XbmwhsXXQCf9jTyznYFfbtze/xeF3dVx6Bz2bZe5AWP/aCNg0
nu+iOgaoYsL+UQdVbqVJ1pirDnWTolU7KjuFUNSf673aoEItgHI49Qob+ekNZ/bqotpimhByxvXi
Bu0gsK2r/8IXaIIXuRLb73R0i9pjb3ac40EdyFg7O9+vs5Dv5QfXfBcTpx1qf6x6nX/Y41C+bERM
9/WKIqzUEwm8mVuTYG21JcNvzBkBZJsO6bMFSerk2DC0Rf9BymRuYfVTz3sTpsI1llAmu4MaHXkv
g0+UeQWQtUNOclS7fu8bMXxpP5nuJ/2hV+Q5gIRqpHrgAwSmhDpcI9y2FdyVkzXRAWwUdbRjjhW+
U12467jh4fU1nzIVoQmnPR99yK+fK/VDlX8XnY520/c6Yv5uo6LR47aozBz3Ep2fy+zj/J66QqCQ
CJHmbu/+gYFuibAa8+69cLRvKfnYfU9lVPp+fWddxXAsd3UL74A9ZDhbVUJa/OFx47w2jscyC530
3TaTTCLwVvexmek3oGTiD1SH9JhYzT3xwEX/WWS0PpD1AnERy/MLd61H99rXN2qGa9eDvo9YBJbA
0kAZUXqXLZaFLEdCBgDWNtvdMm9BhJvH6ooFt1A6T0+r9eHg2wEODzPlKSXcpBo2fJLhyC8TGDkT
f7Jtop1+2ANTI/cnEKT8b1JXTR/yMQhr/3QXAAmE9xNGP+hgSjL9bMaRvMLRgx82Uuuomhu/IOk2
64IF34VenV/nHedm8xXMKsjxYURK8C6Rzjlx/LilLD0pQl9/6BR/CFZzXVdZ1UAFPeBa1Z4Doo48
vlA1YRr2dvz9zEbdK+dh9Hl8fbr/fBNK01vQEBJEob0Lmz93O65imkHisjELXY67JPIAB6o70IoT
jVoITIM13mUBHg6D9Vm7X7GWXhaR3vzEGihziot5xLTlS1A6wBN3D7ULXscnFYtALkJ+s13R4rRt
KcFSattHK947Zx8sV5PZsuOUR1d1/KFR7jgNRj3hg9907LDqOlsgRNkfy13Tx78XeJ0W/5vfgFwD
Tx/JHNn6APwm4K0ekwYbf2DW2Tma7Qe4iRCU8U9RSTif+ai72WVh2CmRKNIKkwQO7EuVt/932TTN
C2UPvJnzG5lNKJfqyG5/PkM4tbASg6uYlRc7kZCJmlwjWFL/xX8pCUCxiQ0WCJUqPv28bq27XGIs
jDaSHBLLoQyQcXVa60T+d4cjDHS6bvY+E63fSb2wcLRJ/hn90Ig3ZR2BMOv3tUPppVLVSIxaET88
YW+kt2UWFvdsDoPHrNZmrk8B9Vl47cURbIMxLyaj0kwjy0XV6AkypW0uJXj0FwItvmmV1Q3wgpSr
x4PqhfytNZwOCxXEWncCztFcfO2aJY2BAC8AjJAkhU3PBmbaCMnd2epzNltUsuewww9vwMj/p5Dw
0XzX0lpf+iYGB8nDvZaohu6oOi7zmJzUkcWVQCaycoZxCBQs7U9dBhVaTCRdv0MekgQUqbrZ4ciw
Di9dt47ER2xVKV4/fsPrNwafHONcvWLs6Gq4Ofvdg5hOeBazk7x0aqdFcsmosrIhs9ensSTgLa8P
NxkZF/yu9hECEjdsLYp6AlcdGoh5qFsmngqj9dmm0D7ZKfpjIT7m0Wck8UeX5sxOaEDUX9tg+eCs
QANmWhs4R/repI7+RWSyb/biNb43GOeM7kMYJHsASpzYA61i1mch2fyQxXV03EiRTPr86jGubVsz
A7wpBA6beI3XZ3EN/rDUM4u4YJ7knWIWCQjwBTWdDYLwODBmmdBkpbF2B8gIags8hlnp5YsQf53R
t65FjpUbPBtkC4pFUeUsUJ2h5iD2haxV5i8ij6unZvh1n2eAbiO5vuO8WDb6arfiHK0YNh64Uh2u
6iqS5fkPxKJr4fkgSEtFFaVzixGM/y6wCa+y1k28TDIVk48+QH1Kk90dHfOiv5vw2OxRN1pB3RD6
chtMcrDEMgsYliQa1WAKNcdJez9NF8MMUdlnpzKlV1g2Ie2o+24tK2jLa7XxpCvkehLElW5gpewD
+jLYucc0pSEKUB8SyEZsZKj58r1r3y1zCLaPFzEC8G7ex/i2I7mdXEEzFjFYjsTp8QYCNKp1JT66
ODD3XeTWJzWEIY0vnGUxfoYqlf5LqWnAZAcbfOc1+DzYRuilZ2oSviWrONeB43Gs8jpMHyhTRy6p
pjsmiijJDIWWGHvOkmJNkKlUAqj8UpWtTNM91rLI2qy1XJqwLpSmV0bnyGoBZJabP+1IDj457J6K
bPxXc32/xVBksn/FathjJJ8Z+S7T9VKlN0KzRWpGX+sWhXAZJaZlCZwwVLNnVikjB/i3Tc2tlfam
k+cTFLJdXWfPuCnySdzOkF4fwX2pDkLOBONFGwMTtezyUoguyn9ATijI02/XmmG4wUrfWFev/9M4
gBTl9rEsd/YPaJxCntMBkciEA20dDdgH3HDQliWgLxNAApISMv33WReRvK3hNo9AL97oiYiXY/gG
i3c0jnjKRYx14Uy24bczi0CwM08yRWIRA7tF85P+LSfHBn852+xdSW6FqV66Z0e2sO+emvDOapMp
HItGhx2oB1cGou74cjrrBLdjmgtxYtjqPErDXchpKWs6hc5AzDCYEEt97eVCtbqtmPojEu/zl7nu
0qzfBIQiB1IpHNdTcsh/uG79x40KE0ys8uLqZaMzA2OCR325xO4MtsdmZJxuG7WsuZnacg8ghEMx
hQ0ge6NQDv9rxu0qSP25YjENm5QGX2OsCv0Q12LI3bT/hvK5NUITwtUOpr3H3xDaJg4rc9KcBeA5
OAM8xsW5rt5RNhPWO2APPJw40RDvKpJfkVJpya0+ye3Khrz+m5JAPufKrzautikLogDo5P5z2JhW
OgZiMUomyZdH2yzmOiCXzCrWFEp4IsbCDLR9TcsZYl0bmxVZC+4NHUZ1eYCSOlfOmvyDlo4Tt02W
aFfWatzP85QIg1XQt/9YX2h6bwSXXQvnintF9nl8EEH8TYgxX0GjoFRKTGOWKv6RV0AIjXeWlGxA
nTczppN2fII5qC6CuSWE90iyWfDnM22xwYsWa3ZXmErolPI9wFKYc0UK4wYBGx2rMZYjNFOhYlqZ
5mDjRkad5f8+e7Dzc4Af3t71SQyIJG3ADNDsYd4VDUlIEEEJtyMeOA9Ap7RVdTCVINm7DNmOgJxd
y+4eSjkIBenhS5K3u9XzUU6O50P/vYM5xLzYeg0ZlpSp/fbsxHZ/R5ZLmmb2GWDMBHxtD00g6H9b
Ka+65TpDblNrDN3i7qVuuH/JI+MnZpTnum2fTmnQ4KUzmXwEuNOXl2Olt6Xx8t/ENP250v9bqkmH
VAfaLYthU90KqkE3l3YPM47I82SkWe9bDVHRBu7fehXkIzGFx/+ghQw5NQq4M/HYMqCZ4pm8bE9V
vFT2VBid9SkdrvSgoYD9GuPlGQy4UbCumt6zw90Uqt8EVVW7oUQ8/fcFF6ua3m2rVFFK0kDtX1r9
jCjf/1xxOwCjJWQ12+cQ5qiGxo2Ff51Q3jN+w1h6KdokCtGFZVhRGYygge9eji2HNiiOA/JHweyo
+lKELh7omc2hiCE67k5UWtsLEhVMhl17mZWcrW/dAsjNWW7ssUFScwYPM7Z2vApsGoXT36fueT3o
v+7/brjnDKtfnwu4ZPzh1+8yJTYa9e2Rdpol8iOdoGT5hP0IMgZWYoQSjRyYiXyvuKDHoqHaNtPC
yfZNtWKJ12SKT5ABkZARbVJs2KRDDKBjVZCAhqPQmmxQ5oMzJdenzP3/S9jgl5GS3TE9kFoeMa0w
oGuOCS6RnlSk48hSJYAeznG9b4ieC7zGvXcPsZ1iNHNsHkkZoJqdIKSljMa7RXOdYAQWyaxg7r5H
fcSVdS1rKDsG6wWYB5h9eNGo9/9cKgYNNw8/48E2SUKSfwCnw7PuRjqzwLGrIhPH5G+KKX8EGj+2
k3yeqHUEkgRuAFNu9M+guiCVBK0BapPU2jRLkdObo4d9mH7VSLqv/QjDVCJ4s5E8NQvJSzp4Kux0
JfiA5afBVmz/wIe97gL0apSoNLrq8ibrdL15L+9u61fpSkhbK4n2iq6IDuE3qKwuUDb2YbuXBiXq
wZf9LgNaqRmKS1qCoVxs4nnnhXCvR2SV9a0q2dcl8ZO0Q3VsdMKmKlrrQo5u9NlUr1/Sbre/lNP7
1M6J6OB3hHt5zGkfL6ghqLO3NE8W1C4aan3ajYqIpWnXoq+U6O1qqA/jDr6Y6wB/7bvPw7RV96Mw
XQly06fI4mtDtbHYoUgMO7tIjx6u/IZKzduLGG0OigNLpXxUB3L7WufKwZcfbEV4033p5ur5DdBK
QQl+cpytWfBl/gNAqEYDkGgm01l3lIs5g5Q4/LnUeyJMQzps4VRQZu1AfK3qL6jY/NKM8eg8U6Zs
Zq87mpcl53z6wP15H8yfUjXxCDD5m8JLkvAY+qKhJw+FRwHolfyyHCGwgSUM+dXq/hdiJ4dYSluT
e/rUjx8CAM3fNqzgUPTfS7cKNCiC0j+qfPAkH0/wTISi2/UPsIu7dgVwhp65SBvsGwcfVvAm2QLx
ltiARNYuhRDYflKjkF8mA+rj6sH+4ECz8YVs697cwQaANE1E8Asd+/BoQb7hunaJrpjCtJ0W5aZu
nZse7NsRlZVFN4A2ET362RQ1Qc5qamPYfC7kmu3ZkB4OsMaTwy1GalKoqpqmyXevawprPwNGYK7j
ea/y7jgTIijdSLQTJq4ILDao1pKHLCaOIwj4GUiaUMIG6HUllngLx8eiod66J5BTkFQEv7FD5sp5
1DC0WoxNu0s2JAy72gy4USRouFCZ+eDPAfQuM3YCIxBqS+zgnkH2n0s841pnwbi1ytWVUTlMTYsk
cR1Ce6ojqDUMXypowhqKWmR63x0OoKE8ABSFUa+EmOeaoOA+kCWb6AZRIc1YhQpaMm5/H6/X7CEr
BjKGMiY4UTYirkZ7n4rw1b/D80XAXSiH8TmiaYbwQIV2A68jn4+sMu79mvw8ixHVp4G0eQD1ZwUU
Z3myiw74/4WJGHTIUW1azbvvMLMlXSWzjebXOK+VbxnOMx2ZQ/WzLTlNQ2ivZmcopVqLp/7MFyb0
DDuDch+jZ1sVkUwhkRYQstAERq2v1v9NSZ5FNdbV2zHSb7Rfq+C+Gzy1t7ic/o0dwr6yu34lQzLP
3LyZwH/UfKWfPeTiuH/zrJDc8ncOy5zEwNZIGo7zbccM4DkZEP/3fzxs7ZT7TRLztxWqFHZ//SkC
HLIsBB06SAiOrQAws+Y9BSVqQPsAvNMhizqrhorDfFoLTDTJ5MvDVr7sxaCEpNjOuFkwzmJT1rF2
5lvnxRuTEPX9oAgYMK43KZ6ZcHlZOPkv6UOtFVhWchLSoly9ShGdkD/1XfWgwWUjqdAjSim1JBwt
zhJTB+3HhWfmYnbz6msQ+OoncgJVwfXdjVu4rX1akbIZQyZUPDPevDV7Wj7Ip0iTjTHAUx/op3Tv
WQX/8S1wMJSPW7cQZhcUdhIMp8DIW2EKHB7wVMT6CRYwKAqlmMy4EMZ0q5Qq1AGIR47a5O6bAWb+
0Hat2OAe0Cy0qqeijqo7RH4zHwvKY4Qc3r7Ga1lmNmTB4gKSjd1rlm+XW0qy/ro0dX2hDuvIdZ4B
RQ+yHbzpMJ2CQmupaGLmvkJ8Qk4FJwwl+wS6Qn1biEkr9XNwTR81v8uCx3Xr6bAIoeHpXVd1CIFr
LtHiJhCIApoO7NsaeAnNhGH9N5BIH04bieXFfA52RfvRrtrHUhcoRrqL4dKZ/v7QIeF7HTX1f4lT
iYGbzuLlchNHs0EEqj3rfOgfFo+clKwv7bgWu/FspVHGprinKKMwK7IG+8yIdSp/fKvmD4PwOIbY
b8KyaLufSfLA3MUIfre9/gfU4I7Fp7fH/F1GbqaJmdEyR3WEt8L0M4DMpnqwXxpQo1pre8bquwzg
7uvtkCWa5sifm2MY37A9gqogX/Jf95IcOT/vLXyEMKjk94rWqAoqE/ematjgIm9gIkoSGwtjWVJm
xxILYkCnnxaLT/9QCfqrNheUxRYM2niRETuXqJ9LZcnJ47jCKI8iPwFzN06mHX4nsQ8lu2MUWzT8
Khzwrsi2BmSNWkPIFpzJAnjME8SXc0WRwBUojAy5mkfwqoatSDPQ7mjYod0A1LLMyMq4SlBTAQBN
VI1MGSrTmJnXE/TQfu3VyhyJg5P8xUuiJLshpWK/vnPj29nHFHcgCYsy3arqtan7PvsW7WsiZUZ3
WADGl2Q2AiQbOtd6CQNwv8V2w4YL27X1kFXtvprD1xnQI+uty4chFy1x3Je8aq/YmrJY2176nKUr
HEO3loBp5Am/YGeL6IJF92Du+nNTRe+rGlMkoTyt6LhTWuLUIKGHRmrbKmH+p3rk7G6g0/oBotNl
lwjtVB0/paYYSZhpv39FPahXFt2w7zF4s/9XFsDsDgeO7aGAj9hDRBuL9bOMxNOzPf88Rbesmtzg
MXL+UINwcK5syQSRdhUQ6sFNIz3tL7jqOMxto/zUNCyasfUCMnL+zVMBcMc9eR83bw3TER83dz1S
4wysn1lDt/SwxAZoLMX3BtSJ1L1S6M/RaEuPiQFS39ZzWEC4U5/9e4flknyOOAfdVamKvQB80NXw
+AniTpKdkvTVU/WABNIRWUzj/FkuEjacDTROV+nWN5XcCiLa/zyGkF+r1k5OGcaqxagMTIHYwwBV
WYbsdHnk0UJyZ9+lvs8BLYnxJNz6fBMhRb5tXuYitFMu6eIdmDnFXPC+e9uJhT3cn6V2cLjS1s/V
eQctGMD0kSDvV/SjId4P88rxBE2CBrTVzldMuK5v3OKQuoQerPPdXZLTHJwGhAujURAJ+gNv0MTg
F66AgnTbP/IJQ/EmsP4AlDZy4UgdHVhDW1LdwE3yWpvokE3z7AADtTWpbldpCBNNfoeZySxFh5pS
CUz4+tNRwsbJb+77ApQGnksvub28nGovVnz+SLrNT1no5HZPBH300xkP2gQt3oqy8y8Z67Dr+wST
6wzMeijwSoNyUjEK4dBX3CBFd5Aff6pE2OBA4J1pRuw5Ksilmajr+P3D9kQWkf7Fdq5o6/nMVDWg
ClIiXU4ykSMtIOaQ1oLVP1mHjVqee2960hPDpf71nfupdn1t0pRQsH4v8iLlzW+PraG2qVIYeUjJ
uIWEox5CPqeAQVcGFAU3KIJE3GbvMO892xwXLlLi5/UJ9NjZWhekCmcCIPPEx7wnZABM5Ir5jk4v
eUBnkaDoqefRXiJYlPO05N1wQkct53LHjzPF0qxjiFnfjnkWulIhVJQoRu3Jje6LK8eDdjXH/F+C
yHRI77qiGW6gd5x4GxHXrR6wqQRX+lNLUJPbGK2+EpvHW/jZ6OVotqlC9Dm3paAvtoJoit7WE9Na
GbnJ+6/WNOnrJSvy/pMLH97waVrB/Nwian9wSy3Ldcp4ETl6Jt6YNLyeixsamUpyaJ/vG5WKuv5Y
GMC4ciz/O2CpnVEhyhYvAKhbRcTMW9ut2K1fQ844QB8ddg//tVOKUiJLPGiTtG8pMcCpmVQNSkqE
HqmQ+j7lctPGxExzuejmlmf/Bi744PuHPBP8Mxt+9CUB/Qw5fZ7goQgWxBBp/QhwbJi6ha6I61wx
Mbe6ELxXiG/EKdBAEukQTwrSObAy0OW4iB2V5a14tLup32oqRkPdBoI0WAL9ACN1YsGH9o/bqlgP
XH2m4TA1S+zB0Mhdne65z2USOcOw2O8BAjPB1XbeXCcHCgSC6fyfJxOBjF8341Xhy2IfXDnYA3QO
u0XehSMjExuZVpKrXpbMZ8teoblQJS6gdF7NpiaeHVsGhbpWAcEXh83kr0do8HDtOT3QTQDZrs0f
IIoMqnquw4FgFvl+ElXJ82fl0qwmU7xp65+24thUXvQrZREVNjrKPHeSuIZer25e7EOBPvBUuWHl
mQ8GnvFqbW6f0wAChi1OMePoAY/Xpuhq3abweV08v0DYNbTafXKN856sXT8cz3SScrEf2Kd0qNr1
Ir7TebBTwmbY2prFiQnYOfrVhK5FXsnxt+JiGhUzdfwOIHhuEeJgIfiWfLYXBU/ZPqxUvCXuut/b
9AWTZ8186TvF2g5eBCHj7qnQVriiaaS4WGCuHvhLfb4VD9lynnToV/27jda02Kr8SguwR8DCkovF
b1HjOoxLZu1MGqsiHIO9FSDhsv0NhsmHPA6XwVBb41nnQaSGgp6EH1BbYYJ+AnEGCuvBfPF43fvY
Ncj+6AUDPTtan+5+wqrVuHpFwloDCkmwwHppvoczq4kgupBK+Fc71CnjZhEclbdwayQ6JlllYyn2
od1Ddn317woH+HLjXF4bAIvJdbU14XVfd01sQ4E0kOLlbSfY2CIk/9Ej6mDbBr2KrdKk9tYJDDel
UJekL++cJZ26+WvDDH76UXDHC/9dpnRcXVi6lZgDRGdLMIuPlAW3iURc4kX9wwJh0T8EezXyHTdi
s+cjxjcAcj2kJ4op+G5Ha7ia1lzxwrbTStNUk4+ypMzQvvUGiNt0B8cCm2mG4N55QZuxWZgIk1Da
vCq4rwdhKb7EXJoI+2cvDbcrIyuCrfLTKfAFe7yua1PWcNUQh2MunpY54bKw9sApMZ6OCl7i+gWE
c2N5W73rkJy6oI9aGpKua9eL0DynDLc5q2uLpN50x1H6uGpA6Oa3CXevotTUmDhxIGMVQSrDmsJk
vqoiKZm2VyQrUeN4DTvv+Eg2lNTpHv6Twtzn8B/Ju2LFY+hdhsGMb9afz6Kg7Qi6KYVIEx/RmzFe
NbJqqpvMP83KgReRzWkslZhoWvCNSNjC9aVSSwOGU+Dc4RLhi2G3UF0N2ERQDPpmH12XuV1BIXdT
FcmVtCBtS+60Pr2rD1lSu6MtjD6FN6/2dTKjOLCykr3XOO8Clx2VUOuoR0s7KGUZ8TSMHU94ORVL
9Z9e+Zj7eAw4N735Z20D/IW9lrVOaBnvKwSny4LFnUh8Pt7U0ZRtpflASiK8Kg/TQ0Bp/7ZLKBUB
8G7lbf/pw50k96iQu2p8QvARDbOJOwJMiP0kUOcUsCQZF0sjL+HlaSI7E6bin9emrshzx167HpR8
TX6bR3TGTPNqdhxVvgaQFnZoEvioFJULlgMrRCYAsB/BjGSlxYdjvKZoj+2fUj8n6RdTk+P3SHVa
UTVOVVtWiXU8IoglgL6dohDTTUwcl0aS8U8I3+lQdP2rDze4XOWVaM0CDlwn34SRWsaH186Ov+NC
9mi2v9gYWnY6WQ0ozjcYRxKpYlMrB5M5IhOXBvF4MHO5Uus7jAADh9z3lh+DckANyN2YOYBcTBkL
SGIkjXqJ3qDAnClNXfIWak4zuEM+3fS6bxndQ5wZiVAskROpCyZJ6gF1uS+LXd7Pxeefxgr1s5ug
emiiRJbO9+MNKywOTEAdU+BFyRIBfPElCHjbh29F3ZV5ilfFr2OmaXqQIhlI2zBXhBizV1ec2UVj
soHyQo4HkQpaZRFsrfvmiVs6D9YzJUsMz5WXdeT6gRSdXfObqk7p7CFVx9Yc4e1cQCgmgLUZEetP
tHE789mynbBviafIGvjDcyYkl57UPlS1nmJY4iv7N4oPP5a/fm3AMJRaqff+theLait43oqW+uXF
ZogAXwWAzX5E5Ro8nqMPNQ5emEX5tQSN9JyypL+BB0btgxDuigqWTWAKfuHgaUIIvsTAFYAqqMsi
ohW6PJS7nWZt3Ji97ys6hDfWKtuupj77DepjvZLX0dm45FK6aARrFnxL48D9tyhDadDpOf6BqxIq
PLm6erRlm04MszPCUzMJHrmypYy7wwHVpK9TABYF5mE2DWL1tlGXpu0hqu1trIlqnxUiitCQlnl7
fPQ0jgXeWsifgcxeyyUelic4DgEEXCfXs1XZ8S35jPdzRDKwluJxsYJAJ34xOM+4ON8W+Q6PoxEo
0+hqxL0MkaKfHrt36ron3vctyJ6Pfcwuf5umyF2H8eB9KvyfMbY+5AOrSvbE/FA2XHdHXQXG5R3E
pDV3AeDcV9E59/UE77oiMWNV4hYlRsvAPPB2a6W08RrCULQHOt6+VLPma0kaSljSLUHS34wLKk1C
I616XN476AufjsH57LujVFYXc3MXfuGQxJSL4gDE2ifO//kDvy1fuBJ6vQQIAOQwv9FVYiss77NJ
mntxRpoM/WZN7+P8UPZ8eEEurv8qOV+Q1NBC+POQeNpLCfFITLxZ+QvWXQJIFNBQ0TkVrbawyJoK
KWuXfN+8VMc78z808+ENb2gpXuhbKuFN+O3+tWwmaNEIYJuAc5/MraN7fn/FmT4QvHnjZYa68sQS
9UJ0QBgcWSNvEMQhw8/IYOAcEY1Bf4dSNr9f9YWBpTdME4JsRyh5Vn58UN3pj0B4fkdJDbN2TkJf
kKQIjnu1TAS2n1Aj16uy1rbhZEcXCHb36IF6IKGKAODKdf/4tDCPJB3piCaFXuJ9IZKHbwCL5cPV
tScYo0oV0wlO2Q7MCDgGCSKeHgBJnkCppRlePy1hiOvFCgu+RunLsu+pGCBIOpUVEpE+QiBBNUdC
RR+L9IuXKHOvJPCwF7FjOYfeTkQHeL/N6dk7Ay+PvgP+8GMrIldJ8dxB7It8Wd1pWNIuZKYoG/cP
r6UwL8tlwqWHbziTR+DZRbtepC1X3u82Jyd362FvnOJt8BPH6wHbv+hd6bWcf99W/kv4IuItXuKc
+sBNOGmo8jpoNci0BdPx3XyCXl3eXzlNdblUUIgbh+7bAH5ARqLdJtXnbHlB8RV1Uo90PHDYEQBU
g70cqf87It1L6mvhGZ1TClZzfuYOH1OEpvJZX5pMFHfyvUyjRNJ7R7xtlQFgqsUpZ0lc52we5m/I
j/D2HLYcAZ1UjvDYIEpAsh5Wp4RoohYn0d7xNUV7eaStcmzrDK/YZBAQgvY2lpbN7ezZ+vy+KtVt
KEFy3f+OM2ab/jRZfq5yMsjWoSmt9GhKcaZMiOX+ys2s+RQq35hhXlkJOESN1VykbEdXoYCF1r/8
kHDdx7ZFob0e7wsy4BCWJydLXe3eN9Qpz1YnrNi90vRZbN4CHkupgd1YB7kdX3d8gNHLdJ40/Vw4
2KjMXSDKjh8pKEjsVV8plwwRUCSwBuT7HenpERRIKNmp8nzUSOUKBMnr5eo4TI5bGezVEI/nGZYl
Fvr+/oO1q13sOSI/Kyr+qb7KDwkm2a6woELilYMVoxMd6nYx1d6vaOtD3v82RuP6TL/stpZjHhXT
jnpnYW2bJU6HCx0xaO2zHIY3US58V8SgQZXPMgGmqe09e5PTE7ec/cB23U6Zxnod584q6TvPC5hx
IgjURy3RkdduKOIkGCRCiO8Dks0jLjRuguRK8ux6M64yYQlz4a6rWDU6uXdtS1/r8uCdHbfRMw84
idehEMNyFhnmC6zr61C2c/5BZPhfoSNjJtJ+rdXX9bd0NHGVhTDreVk2uuyBYxCRrd9bfnYrS2Sq
+bkljg4DWkVhfkuMSWQdhb08GsfmswT7uNgySrxIdD5jzbkfYuqYH+VpFgUD12c46gOEjOFZ726H
sc0P/ny2ZvwxcDWbld805+qZvICq7FLX80Jhh7isGZ9LD4kxlEx4v+jtiSaNl4HfdmrLZioK0TPC
OGXZkyx9KZAnRC4Nk3+f6IEsgeH8a9fUDUZ1KG6tGRgICIrKtlQEjaI7J2icVrRsX9WbCkR8dojx
BY0QwDzS8YDZekNF2tZqY6ushNazj28MrocSR7Ww6iOVOI4ZeMwiS0lxQWQYVGOeDWMzmsI7Ha4p
cIdSbfYtscyhtUc/u6icFJHpbUKAIuzJ29WngDc003mMt3LlHY0NyHbfwemK6jDLDqaBmPcRqzMW
OsIefIK4F92r4uy7JtpB/sUOpc6MD3dwzLsFomOzlT6KkZdD+1GXn4vbF8n46Qh/nKBVV6gtQ1af
ATSmFqvspBKO6LxxH0zgibEMwHuQ7+iTmTZjkR5leulYRJ274XqCpeZuIIx2bBg4TXEonZ+5X+Gb
Z/Jx37zOaYEJgtuII+69sVHUAwH5hK2FGZ57kgcCwY9W2CJW/OsWK/ELq3zAmseAWQ5J4MDstfOS
Zato0abTy1L0/Ud4gu58L3alNut1xdZdVOEu/0Jm/9Ojy1G1qf1QxlSFH/eckaPFv1OWXb8DVutA
hNTHJPF/Bp6kTrXmLYV5Q4Fe6vWRq6CVN29Tudd6XAdUjzeXKhNiyj/ASaJhxeCA3vMPMQVQ332l
GhU2sq/ENqZDcLGpeS5smRVatVcmUMjmvPUi4cQBzHaCb10Z/0WcacgUoPYukLuQ1Mi3qIkPM9ZN
EPLFhHyZdYVzafL3+sIRB8WRbbx5Ybr3uDPSJ/fr15Jp435uGiU+J/zoD4Z4fCE0qVPGLUJpxkP/
8blQpJ1mWAJhsFCEHZ7pfJNzBjy6rlDtQMpnlMFBUuOZ1GheUSUBNrdkBYbWiX5Qy2qO9u/xlJqI
zNMjwvkB/aoJeg0CGWELDx6BzJYR2rObxJwY2SHcE2V9bdrCyi2w4RjN9PnLrG4Ps+bJRV9wwzv2
jNMfpUP8hHXmUNTZac6EKl8d+ecypKW6ZehhOzCKBSAvCCrLPAnUFsotJl3U/ROHqMKvLGeUuYCL
sHBJrbvJStEElTxMx1N16d8xiZL6x5HXoZjgwt6fue9sUtbWQAOZCsLJlITLP9nsyAKZUAWklxkO
tQlmVx/O0KfDSwwx4JzQSUEf1GyUflMePyHQT2Wm7KmNoxnTvSFw/izZ9kiZ6bN+A3RG8xDDMlli
pPLD3C7dXTyXYV803698ttMWnJKLpRv+RxSfCk3xhLA3S7vSGfJXBNXPZ4+oyYQddRwVTnZZ3iay
kXcYb+tHV0S/udQmTG6UTEn1ESwS0ijc/VA6ekt41mSs2IvvnkTxMYw3Sk9pnRSkEq6DcVEa9ybz
EDDHA9IuzGF94ZXKeDhgmFlu+T0sioaDiCCm3sOhHe7fR/jLWieCU/qVcN0lWrhSD+me6hQfOU+/
/XViOLIkWT2ji05oybTsAboWSmMh11l5rtKGgV98Rv0DF7Cz2vM6XeoXF3rjyFwwgdHtlSuT0k5t
AY06F2LrVhaejGMMSRqgaW36hoETMzm/NtgVmiO6T/2i8VwrX+rWYCnikWwkxOTIOCcTnLzjh6Bj
Y17xQjfegIQC/9LAVAFRYoNWOsm9kw2QGnm+EK18KIpgviEM0vY9t543nMQlDox42kb9bK7eRet3
Gm9wDbk6K19kZ8p/9FJrAjCGjPEnkryixZvGSZ4/WfdR02/c8LJgyVn92Fca6ncXlrOFGouEhsrb
9AUp5x839IMEvLvWc3rY9wPPBFYkHBfe4QTXImx0igWW7uMpPbB3pz6riFLn2A9aZjNoIDKTvosy
FmG4FaTYkV67ANWAYWzbNfUxgcT9RJnnSwYF+LGzor2soVpwVgNml2onAZhHR3+2Asq8kCrJXPcZ
eIBiHK1Weh0CFrZxEKU27XbgHjTjF/9PU0i2YKzw9RRKWmLmrTIj39/71yn4V7Pi4Zuzo44S1uuj
44hzESGP1R+KDOmUZENhzQLnLwsBDARK9JxEkYFsnJw3uvLVFeaAyGUIJx3zBaQAdoWgFguu6nB1
qDHEDjwbkYbMBRWMQQW52oJcDwdr3hXTMWndydq2rQrgKOed3a0phiK4e2ZeyWPpAI04e9N9GRCk
vF63/GqpE0fY6kNep0fVq0CEzIaq98xCrlkI8WE7Dad8wzs7aVUgmdInfG3R+4D+Gtk8C3aOX/N1
jYd74DQcrZKFy5ABRpJtfgci3Jnn9nqqYcHhCBzZ8CpPajOcqtlDTUEBaZun8f2UD2dUxs5ykAWR
M5Xf2surZgoPVC0PlyZ2QC3hY+tCwwbCxTo3h+PJ3QJZ3OLFpkEaDB58mqGJMZivKNDfH3C5TKJz
8UbvZoZcaypmeggXplTRq3XFv/yRCUSowNMKFf5Z0gzP+HIPwQ1AgsNrBMJg3HxcDSPsckt+nrXV
ccVeunPy119ikinu/pwTDe6jpHeVmJFNghE7k3kAcM7xVK7J8AxMUdHwxLx91mNEO5PzoWqrfgSE
tgGbSiTh4wJBEYNYZf/yFcbEKoG7QpdCxWGbno9fhP08sIyFpdPzT4InMSeVYmEh3WwLhS2Z0x0t
qGdKqM7JOwGXurn5T0Cg/BWlFkCoajoY6gV8N0iHJNLIoAisMO8p08CJGzZtB1HxuVoNawn4cttD
OuKe7LOrkTktno8Y3/t0qUEEEiGjPPUQd25oxwIIDR664l4EAR5jcxzGNkbNjdK//p9jtzGR7eHC
MTZPb9JvUvt3GokMJ8ziXVauPCvrQHtU4UA08Cx1BC37Ehm9kuRUGRd/ZVsjvVNxo05T2UNaLwXn
7yLTAwpzmlaoJ8kdnMEwp6nsArIOI5scfTNGnYx1xYVamQsaLj35i6/aUuUBT/EneVsllesytCgS
j1XIdGziHbb8uF9jAkz65KgA+kivXksVdcmZt1qAnQW8QNRj3W4dJWWcmiTswqRKm1EnwbsNo7fJ
/J/dAmEOtUOO6oF3xNklWqWb3NLULYqrQi4Fmxcdo6gNFBP+vKkat4Velt4WYNklVtL9igACcwaK
DYKUnn4y7LT73tb+fgXjuMdUricBKlG/WtilFcUu0kkO7qALAXi/CFRYSLQl8ToD3NUSqzkZBlYy
WyGRdg4obpXWZA8PqOlGNu84t7LTDBqpbFRWGcjfulvU8GrqOnbounAtqJXSo/yNsMU4Xyxspr+W
aL6YGDlyhOsj75ywJr7CgWBHlDdtiTjQj6Og9i4jJ3Oyd+2PN7Sv5OLztA2+jzew4I28XYiEAa9H
tf4q87Tpy0p1s45u14/Xob2FmqVNuKAnW23EE8rAYZYxRtGlQRMXp7ih77NCH91enYXOIjS34VUr
eswgN8m/WdT1ilYrgQOFKVf63knol2yiScR1ZQY0mRwMVh8PuzKrqIJK70SIIXxJGtkh3dqIIGvu
UHbX6y0JLMZYtKr4G7fptbGNko0Dc6qqqatN4qJ3fA0J/AZgl4eNYol2COwVUvOg441W+TfUBEvV
9HJCs+Jxly/K+I2Zz0IkhfTw82+T/1rTymyy5ERU/7doh/hM5HlZW1KFcN18kAVqDrweOGHiEbFj
sJyA3rt5v4sEu1DYL8W6YnSFnpP2SD+Q5h4hAQ0393sx1mOf5bvEa1i/oC1af2DhtM1wXle5zf2u
JaoSvx3FUIn9PWvMMoRMB7yvqwOlq9hPkm8731eUoKEanM4+rqTqG+a1MIA8eB7zUMm+JnSoDULU
SE/Z/XIAOo+SY44SSp4C2aWwBMzg44hHr7tYVU1IlJ3ECuyFYMJUTqeBybMFRaPvY145khdzTtKy
LAhs3jMbcWhjV0eXd53rIDY36/SKI/iApFHjBQQ6d+8M+phTEhY+6bsA7lfNMATX35fMTPaFwEhY
5iKmJVuAiTuyMlYQre0YgmDLwl54c2xl/od8QeLoFCM2NIbl4lv51tBVSjesZ+fEwBMy0MxvGqhb
SgpT70KOhiMH8ZWlBGAjmvQOBz59UDluLLgCqSjIA43JQXIKcTzdAeJ1EbcccBkuLPLBVUcFNEh7
uiwqKM5ihsjlDcaZXiKhaXbEqaEdazau/Si7OVHtUKdpUtoNT0ve8KpRG8P+ZFGRQXJc2eNFDVLH
+mcIO5R4YkJPLJRuDbY/RWDVhON7FkPiizw95Q32pW++F5iPmDbTup5UDxogqejpwxugC1SmM//a
ie66BkJXxqI61KoRfWn3+wUQPTiLgSHvd045mTGuzElxH/gkChTujPvzq8s/Bf6nVZ+h8Rj/FFqK
sVMeofkFRo41jemmuuGf/npZf0RNrdkyrKWfEszTCJe2CgOGISR+nONnDEskJ/cM8vz0Jr4oWoQU
R6k6O2kIXk4b1qLmsFN0lXmCgQrU90ZtzmxJsdDoV4oUe9Mhtd5qk4CNL3XCtN6k5ZeTnECW/p7T
mbV5GpdkEm0oi5mfi2OmfoVsn8BAwOcb//PQyi2YLqnsGnp2apAsawBbJRosaM7zOy51oW40Stwb
3Nu9+6iG//ndbBwVs9An+mVdp3ino2GcfaQYNtQe5csjZfCZqJw2osIJ8MdELucSsSMgAgLxnYHJ
vl0WoS4nlmEhIMxGP3OlhKAsz/QuggQtoT5NwpFB7zD2T8zm+QK6m1QRp38LuQXLEKzKwzzpCAU5
zf6RGpD1d1rTDWm1UkIOFLyUocej1s75cZLDUHayXVZDEuWn0HZGpNmajK5Ybq+19LBQOEZKyrSA
B7pM6L0spNTWkIaiPJsSXhH1+9oGC1eNVKRVOhZOyDiIbh8KK3NBZvvAeHhwLIzPcWb6OLb4UIgT
+pf6e3hRtWVYaLzb709oGnct6GVnoPp2pIy8UOafU9954wZbwo6D48THgjJYYR8XG2VoVJUzVgg7
3FHQx194n8mNsSUSOK/a+4oCJ1P7LzslNE0yFRJYYWAfX0Y2jflcRuM/Hcv+e8yV3hu1pcWDNN/x
H3mXm4DwLF4FbMtmD1pkz33lCYGSN3CBb83wfAuLFHljhq3dUnef4ivsn9vWGaeJT8w192O+++yr
bnnK0214ofb5VSKcLLq4S537qeSonVIewWSTzBLgaItFoux8St87kopsGQyacf5MjfVGvGW8AxMA
2f8P6xEcDL1vOGc/u6QGYtT8gaWeoLUldB9qLJ7Izgub6wz8aCnS2q3sok6FeoNHiSdgjbFgYYKJ
IhhXim4BgU2XHRiw7LfhsCyJKreKODzj2t8lhpHLcpQbRMyNFc790IR18CTmmeQPy4Np4PlApHuW
5S5tGllPf3Eu/IrEqZPrdzTyxHR5bT4UKPlBDi3tmF/duyetI7S8tD/n7roouQ6CvwO9sW3d8CY1
NUooluDeiObOX6wrBA2pRD59uftEUjSBb15wP0DFwiNZxNjsyGauWaefWMxvHL1CbsHNnKOMyu7O
Ukve2xugGyGC89hNl0svB4XwglZCqeHgQXVYAd7nny1CkHR0D9KAgjw3e/+mzEjSgjGO6eilCwU4
te+1uQVdi9wIaX+hzMJKHyzg0me5CSBV5gxo4GM1XmRRavn+L+Ai7m7vC5ONa/q5cNOTEtvxWiLO
YtVK02DHlX1zf6r/sQz+Mo7z+rnh13YlNEmUuL6cwqcxBAbGyeARwP5Hd7Oljn7YNOdHqywvx3yK
PbHqjS9eEKhfugb1nR4i2Een860fyr8vFYQEK8E9p5vIOzLYelNMliHCOxnLU9DhR9/pUQb/p2h6
2ZTKfp/3aassuX2cWfRy8ioBSg91h+f/M3H5rKVcngl50hw24C26e1AXKDXt7sbpIhZilXanmtcg
7lv03TIPtmi04QR/e9ZOygCj/7SMnoo+771F908dsziIfj4B/JrkEFk2ABmfRIcunQMCjwg9L7ya
riVJPyvqQQ7syw1ipvPUQFG07D3wwYlORIUSvIHeUSPi6Qp7cnE6uwzpTEc+weQ7/Sz1N/1ZKbgl
09FlwOpSokzKQhy0DdoQrHVCSwNda4qEG1tANjfy4ZKtY0y7bcIMkUCelC1O7FxD6y/0/yjAism9
69P6HMKHj8LoeBB7ehqbv916Y1l1mHCrmdrTOwLjmgURbo8uQ/K8cKP0L/hHCJHIXRkR/pt5NXXo
Ok7kDEg/yHcJ23KzTSkmUaaGtA4bJ9vV6gEjxfo7PyDnehehjQx/WF+NLwZiH1RmTyT3T/qXMma7
Nxp96oA3rs8qZPO9BZV6t/3mth2bhe0hosPYiEQH/OWBd8KbwtNDpXJClfjGyiLkMpajqKxwDmhE
Ad8TEu2UXcBTsE78on+fTytWtdM1Ytl67htPp9IT0OrH82u2vg+uiSjgylyeJ26Gxa8LpLZSKSK+
mBmAU6SrLchwl8Ez3lLOKdIEKm4yd9AvvcDlyUrfiPKN1zQUSReadz45Ah9NY9kfz9qcvYoieSXo
AcwU9EP23pjob5B8dLqV75PWislGJREg5TFyxwcKSd9s1WQl+WUCZHbi2bq5T/KwMfDORooP8AKw
t02DOQwvBDuFZecOhRRmdUkAGEDbQ5QR0G/3oyHVly1CPML3YIKL3boCE/G9JIgutMQOkKDh0dXw
WvPhNyg86NCkTs9sKOS2tYb46jb99O1SsYpV+evOOBK8D13+A9wSBn8/lsdyZmKwIB4tRbvlKUWj
hmn8mIldO6gGFKDJmF5cHHSZYJVGOpaBfPr/2Eeu231Hxa1F9i5bvJIT5wDKWQKCF918EORB6Mp0
0jhkakpFt33yz86eZYhkSydsThBRa23gpFesLQVLPkiJfFGJAlgvxZ3rjeN5cRBYr2l9x0+BhzjP
/l94wjvqtkoMZKDGcYS2AxOEJR0Nc3hAdlH/UoiMHO0F2hYswkADfUTc9K5O2KHlw0YXQpxEfMQ0
OSyjEuDQQ/ZJrtOGt7ey0QPCKUuH1A3YnoE/p9C8xBSqrL2CIBQ24z/HmYHNJGrU1SAC4N8X3jEC
aYA3lvnPbtClXmEsGQCGUNCQ77pH2zZpNjmxfCujcajdDpHYl4Y5rAZMMd/OAbM2yVXFsFZhD9Nx
4ZNA6AsMuvtqVKs+bizGnArdmPLwn6hOYV/cEr7jRtnSo+sd9OCkY8LzwUUbTxeFF1w59MpEk1O4
EJOqiSS0Ed781kN466HVeh2ly6yFRIA5hZ0ARcY/1y1m+3k+6qL8JlrgDhY+t5tD0Mrfo21qfxrg
ryEJXsVG4EP0iNLCvPv0Q3ytUT0X6quMw8MMAVo/EJMq75pZ2ZD1LtDA/o2URrSzUeLcx2P6sfcz
jhaxikPfMDQF0pmhiZ/+M14/XkE0R2jq9OX9BaNBGeFW7lf4eHwUXif6DmjBZKL8Dahzs+Sqyhmc
YAiklC5ME8JaSvACs/k3k1amoJjvhR8e6jEN3NxSdWix/JpdS6E3OvgfLMe9ZWccqxTMssununUw
wjDqwxKxIBcy8kuI17NQzY1Si2nz5hvXiw6bPiJYnYQ8Glp4V+A8je865GVV5weuMJbhyyBWbD4b
TuKOGvIwZ8aNMt+V66zboJJVMwpJUXWQtklLoOixHqdv5Rgm24+UHBk3t2X8482o8g/PHhxSgu7l
997WDIrFx8DM2p5wTAPupMXX3NJvoc7RtCPa5li5kf4d/vzbEZH+uJBqVvx3rbgfwIE6P3PHlpyL
t7Q0KHXNJwfEgJ9Hz6LiLwmxMge3A+RNipoll2sAaSZxf6dDX6rPrhg5+Kf6263lOFboYOs8LSKT
7SgeUHSXzDf5Mtqc6mHsKGIVaP5zW5Lvc3YaezpKwbphOrRjdMwNjLtutoB4YC5nbYj9z+Oxf1YQ
xgt8SGw3ukbZBVT2nZw7xVh+nomIAqjkp+CWqWPGbhxFXhIhJ3NHLrJRfj1i/Q2wUC5xhkd25LpI
AXb0dbUyRBPMz3RkWAp/A7B1VZoym4ZksCruK3W3e6hVE/WKuMyKMcQaNr1v/lIQH8oIkScMjLn5
TWmmHBQE4D8FzNx2AwYs9kbGojwjAdamBUxl08N4aoyhSkScMoipLvXfGIzoFCxb033caYHxiAxv
jydHKXFf3Og0K4PcRVHWtwzjxmmehcTVPIIEib/xBuktcLkYkqyW95ViqQVF5UsPWRaqInisraQb
eI+1eBLODXvnKJLQapBJmCsSdViC4xCZbkSIbO8auneDnb4Jr6Z8xYE/RijZHJRFx6pfPWrc2/4M
I4nDz1Ul2Kgm701UAr8HSMD/1q7JAIc2s8eTUU1nLJuLmnbvrcjUrEJeo4zHzgC1rFxJ6sIVSKsh
TA+0B+dQRdnighaSE/XciRIYSZKLBvQPdmXTUuyffOueLtnj7X93aIAjC9WBK2xOSmja5pWOEQD9
U+GBbD972XuJitF2+X3CizMVT49CqlduGNVsUOhiH+k1Jpo36yak79xR4ZmX09w1d5iNC4K2bruO
zEQC7wjKGQ9cBuLSxSoD3PInQ0ECPUw7tnkYB/qbPFTqI+ujZbfW1+cPDgyX+c6Jder2JhR4Ho8W
98u/L8T2HW8qUjPczfBwjmMDRWHKvXeceOS4rFnnzNrbu3Fe3O9Zo5aufVXiR5qVFjEGTH4075Eo
PuAH5DJXJjoD49FHnFBlSINZKFbTBlpOLF4GviOJ1Ruv7n+OvWA+kL4aINXWbimXloZbeLeFkMz/
ztXBZ/WTWML9FooPeW57QeuTREFy7Bt7dZ9P8UaWvQT6Wjp5/yZjAGReRiDEDRBlumyfuAbvUfnI
HKI8ZgNTIrYW3Tyt1ljKx/2Md4mETDC7VM1EAOSTToLVEjsj7eEvRRs3QJ9ezJbxc+eZw+mEKFTM
uXcjGTOHgZyOlBFux4p3mJxhYLVkJEABX6GTBFvtbFIqht3RjQdJIZQzm+mLg4CXeSJqqJgm1mEy
m5H8fLeWpm8suu4E1n0Pl0bBgVFNR4XRv+foMu+FISwyhT3xecGoYED3Epwy9tpUEPy474SdrZX9
MAtzjE9B7j5yedDiAeBbqPM+swy3uKuWvIn9/JCeSeIazktqmVC2YQyUgrMFd63HvITkiL5Rdk6r
AZ+sy3i/XIRqx0AIMCUw2DafaGIBHVU6Haus/Yd2gO8VKftxX5rtgO6AlPjiID4cX76sPVXs/sIB
fy5RQjdvEDUVDMCwfUfJdoP4BGYisrbEGqIPVFq9tGT/3sMii2+AC+EkWLMhy4iq5z5nzRKc7AjX
UQHwoglOiCL+xgNLR6BNJCbfy6hotNOK2daMguBLuYiWvkg1OK+5cOf20Roi7ka7hEs2EJ1qSNHS
zi45g+OUgGN0Kx7U+ckRY91OCZAPQbLjyNG1wjNRV9bOY16ppKNlcz2PrK5gJkMzNUzgzwmJCl/f
sun9X5xf5KjlkOVOim5PnlVEiVqiY1lCOLXx4qC9ACmtPspl/d+OaEUsrICLFCVjSS/2ttYy4mS9
+nGKrisK8OJKegp/Oi03tbzLeoAL+2BeeNw8f9bjgAA0CAZp00OA+uzavycoIJHTz839AAGwWbxF
6xVxf5K4WqLlK3L9wOGzWLlfnjLwSKq8IBey9XCOgjKkidpJyDrMut5qR7f+bngvBgYjfMlgCTAb
qEUFCxLsRR9AIO0jXNckxMefXeBDmO1iox5f9Z+qU3d4yAsfOrfeXX5zRqM6JGs0O106FykdW+zq
PQ8VuDabhPRYu0G9CosmZhew0xVFTT1lGevCD2QKVUDWfYtd3zXE+1hfnHxU45PgcMBoGLVTGx63
FZ3LxTr2ZBsKbIwXqtmh/4mULwY6V46MUKQDQ7N+fsrRJ6X6kdoLq+VFED7q6dQA5Qd8Po+dBu0T
OBJmbL6Yi4q4nrLMne4WxuEfIj3OP3Rp8FxcHpv/yUsoKLveBmAmHBOIpsx571HDpP/UzSKOMadA
idZpg7mhR49RVQyYDM/JE5RSKYK/nDbeO6kso8TeFgqSPkR5iA7V12X2/LVhSho8tXknwSSVwslu
0xBepN5sD3+Id10vQlRePVz74hE2L6TKU3IjHs8+f2yEJsWBTXuyHc86eVCdc5Jlk48jAsu9oJLw
0cTXi8r16cK5VlIgDwR4JrcfNIEdddeYJS+neKdsLQfP8/0QbUCZRCkeZ/pXLPF9vNVoj2sMKSlo
eYzuY7SObUBs+pt6tjsBBVXqHMBhxdwd2UarwkG2mKhQoQ84sSoDRD1gQHzdRoCeqTzJghWSKev3
SUdAWw4cGmJfLWwuxkruZ9BH2qeJ9JJ/lrKz2NLEefo10eoZuUvlnM3x7nMnqA2x9HszmRFNq4E+
0k5cvYQ7rE0lAg/qoiDoXuJ+DvHQ0zCNrC765VUJR3cavuynK+chOwK7Rl+2vBr6XUWzlN4XEkSC
B2LcYv0t39zX5jqsJbpZfcFW3RNptNRQER5ogaGQFHPJ5kvn+AQ2xeKbz4zfGrlO+WkNZmwONGi0
gINTfNv9/IeVrZd3m+driE7Ot5whg66O+PX4kjkaFA2TEg9B85UIoL4b/AtVG9f3clBAk58de7AL
9RVVoA8pXptHeVbGpXNPCo+yEm5cNQAUuNjeYJniqh6dcOV7ezilSAEgxZYFsK6ooBGAJ72uyPQZ
HQyqhM9I4q/UqJxT7mcxJIYUcIHjd9E9ug1lEwd6HIkTWLDJUJIosCfeGmmQ29AxaG5EKj6HlbdR
AN37ZsLMWEiq9C7Aq8QNOF6YrZKq9hbN3qXRMXq+mlj7IrKoelPFxGvuXNcMYRzV13ljRnnNS6jL
7vm9nmciYQfzCBJk0J6XCfAJp8zkoHrsvaY7jbw6OKxFgEj1d9JL+8W1UE+1flMOQjDEgDdQdSCk
eE998OmcBhBjHtS8CdBRPJx6f3BIIP9igpXSxT2GT0nqhGAnT2A18VA0QjXebUepVcPHYM8AH3jM
aIof0VSlhFr6d3Worz5rRzlZd+glsJT97qsXW+kxDQH5usFDd7XQOQcq8RNzrtzPjUTxDXxaLei+
gHv2MT1BbBP5EcKtwO92iTFL6wmRhhX9Hdc6XECabsWkWnHmyU8D8e13uhB5pnciUQprq21TE7Kg
HZw/BnX1QAczer7ARwJ9xUrik26qpPkA+KkQ1RBEyscIT/EVyk5TBvHNv1ZHD4vG3EPTinGTq26f
8nsr9qh5PRJ+yrc9g1kaGOsE3U0skvctPE6FXpTwX1WHwAEumqT15P9VimcIV7A0Fz++2cEPSilp
J8r9h58LQCIs4mmxmvtuYpwFIPIU+2GuXx32XGaxCuNiwTbJbTT6Cmh+ENyRWjc86Hp2XNqZinZM
2k6LJ26j/ndClFTsaiYLzyyW5Vw3deS67Jj6apQx7vl/0dXcCZVruC9kzI17dfTVAkDN6DXiDIbh
M9gCvsPikXxo/t6UmFC5L3KRr0gnllpGnzqOtvGyzDw6Z8ukQIRb9AZX0H/H1kGL7Ou8wLs/NkdS
fSJtV5IVs39M0QmBTBt8SGNoc1ohMZ7APXeNeh+0TvCyg/ve51CAr2m/LiKah0qxoALl2UlhSix0
dUraUm83jujNv9sGnBlZp6vZVBaKsQaq30Hkz4GgGuvbfdjhNW3LrZHb+Fa3lN0mBaQgAs/f+17R
5Qb7elyROMaOHlezB8BMCr0XJMoq8GrO2eM+crKi9aEjWGEo8dtW2CcuzwywOR+2AUpxSu4D1Lvn
P0L6DB0JEw/UYSVKiWqEHTtiz5NpOuPlQ3V20vpkVlV0tTVLd97ivjHErF1IxUL6sGfCz1C/LTmF
YohCkkNRqb9R4LTiC3MhQpWS1qSiZJddieDsVLZ2zB0Gx8bMKvmAW4YMPezaRjQPsirfK/49LkEw
2ow89PGChSiFZv5xOrCJ1roEgsqysVYArQN+AOKLajfjyQFZ6B6KYIrOTY5zJ6ksmC8WBxS4nL1p
EeYfDHphL/TXbPUyPRj3Sb802OMzUF7b4BTrThMu71UF/Qbsn4TNzmj1fvnGgtBjwFIV9tS+R1nu
SUzJG1TS+2ei984p1f/rF870RuRhnFdcKDa4YEC+WRrRJk7dhEZXu03FtoSRoCVFZgI19q4I5K/G
rXA/dz449GF668IXkbbOa0EQtodVX9xwLfu/AH+05CZYI+mW9S1Hdsg31P6RV6d3RouojtW38cGy
W3PuOJN10f4ajNZCRrMg/HUJBK4kuVXsaUO1yGrGpADhWQbbJviUPtWl1PxyVCq2oHkC5+58dTvl
oThf/u86zrJzF124OlpKtpjuAz8tO8pi5zdr1PBS3aKVqZAukCG4KPawjBTkOKS3HXV6Heb3qHLM
NZlgnzqZHJINvNu/yzeJtIo16LOULNezAinuvMQGlN4ahyg/dfB2kfJydITmN9eoOM4EFaT9ZfQ+
4s7Q/zmf4Xg4ZwimmFh2jrLVTqFfFc+A07S4QgmKQQ+UKmdNxgVfZYbAAvSwSOhMxUAWA5MFhIx0
2Hyj90VyaP7O09W/jmtkPnPI6DPtRnomIT7yT5+t8y7bk4du3YXmGvk32b7OWV8AFcE8wcNks10m
CodZ25T5SizgUf/LtRNuUoZsLNA1eobzyOhp/96E/cyxzPSaNe9fHyLnBz8O+qqjZiKEq64dS5LM
eqWmfonUvE2DFNMrrjnZ8/j7moiyDhoUeWQeM4eLTO1JFC5iFQRlSWD8JOvN8nl28RyluplFtJbC
gsWNUduAr7RyIFG4gogWptZrikRbIkSmPA8KFzEU5s4XFR1NEeIPwxqfmrDywLLk4vgYP39irHIR
wlbOz/PYvr74OMIYSp1LPO+fGerYLXGrT4BamOYYIwZ9M0+0HtoMvMYdUUyvwn5SmvLI5XE9Pd4+
MjcqYZ/JjsZ6euB+lBszxOTzTJ9kED5LL8/Pek4+GVDVn99pXDsYEd1TEvwc/e4R0tscbd7e7Rgb
nH0G6U3JkIujRLz9gdSwnfWdy0EoSdZ9pU5MVlATS7Z7Kqlgp6AqMjpXe0+QPOiRwz9OmIzFuYN5
/WJ+5vr6YaxEMeCNcXh09qvUvs00JRQ0bc/xSKVRFnA/oZ/uet4HuoO57mDkr1K8XZj67DFK4pbt
rcN32N4QUB2y5WAz8bEN9eOxSvS1PCF8aRcFP4+sgzx+1Yk3oPfKG9DldQqrGkbdbMrGAgg75b5y
2KZdzY/G1iWpYCK5iKE6XgBWwTqB+YjzxkulAeFu3IOdGZ4/aDfGL8qdrJy4sU8Aoa7V02mq8/HA
9/se92PLJKD5FJRPNMs/Q1r4QMfAWAJrVciqGjsFtpP5DhgcYhpG8ktrpXUauRtEwS8YIYgBliOT
LmtbwUcJ2q8MvrcnZ8AyQLM5F0Epk6WahfK7FSsK2b03a2ZjRKj3v32e1+sTmK8HjrAWVg49BYOs
VK+XSRNMOj8OKsnNXskTHRhX2I3W5KffLFrO8NCNkZulo8gMjtBgbQMsBmKkF2iwTXBd+3twOLnj
R27JcZCeaNatrHHw7Mq4z6jq9mnq3i4jkikRX5UNnrwFoHQndCD2L0ruVnKI4efilmSMb77oSOH8
fMjfB36xpH8ZYSXsbJ+pwHoaeTEYDC2u+lxY/3ZnGUEOfTr6TicLyQqaZOIQ10UIGt8MyaZsTz88
NpGeh/7q8rFv86Sq0nU/6BNRGBw+82GDAzNoQG2Qzu5/e5CNdl4tginaYCa8s+OZmtufDQkKb6qm
rUhYpd0pCRQJt5/XOzFyUEbqdldIMTqD0hPZ74lFXldtJ+rWULeGF3kzsH3ILxymviXEj9dB3G//
66mYzpZ0OrRUPSwj3TeSaw0eCFlvf310/+keOEvWAJgHzsd81qfAC/l5lL/0i7YpLTWLjAIFsv1P
DZfwuR8MhGqqnXSBLLkurnpUs3uZ6mbRytHPFlzCh8w/ICI2fNjgVUoHxDZ/NyMsB6DYznzM/Cdn
+chQE8pPCPaBw48qNnY4ceDp0/yJRDP8KOx2MXbPthsDD+etm8+lgGbkLWqVGdMP4pWCJcpvqnpm
c4I64m4anlxuooYE0A4Ya4sIT3VfkbHL3rhF15Mxfk9+rSQBFT56dm7N+/8K4B37gc+Wo6QT+KvL
PBqXgEgRxQVRrrQ/oUSEFJetDUlwXuCqUhDgWaG63eS+bCu0tO4i4jcmnOKY0Jb3dV5fzC7McMMc
fUxNj+ekOsBRFF4pBxFP9iwoN1d6/I3OupzXEPzvRQbTjv3v3/idioeFl7plEsoncpiLzOwS2a3S
wexuQqmaUMccPLWUJLATT9uTU4hL2NViYhZULdQPHSLom+QO9Py0FtZJGG1G5yDFxWHFBGjDnz6I
x8kpLRKTBdw6IMGZd4ovcqasNdYCm4Gy3knzCruqrUS9aLx9RsZqGL0UKNa1EXVfSHEl5hV9gFYv
+xTyIdff5GwW0agAAfEa3UptajBrxw5D79xGho7I9JoZEtB6JJsWYxZs35XLPow9ndtGc6L8vQ1j
ktZFPwXzXu/MWoaSqwNESUVb0/HBMtKJEYPKwI2adHU7ZBsP58mprOQewkIWeaFehl1KbTpPXZc1
4m+Nv4f85LD8ekSWS5z8haTtTWZjBx2vvJaYUcmuuCb7R8Xt287jUQVpThxA91kB9JLEKKfd4J3e
qWsiDALugFWxRBvDmJTAsHx92ge+hRlENBfpblGeVE5I4zQzqExiESboB9iRbGY7K+n0/iMyicRq
lW8wHc4HxEBmijmDQ3XNyu/3OofUdRbQaYhCrHbbvFHmEOLA+kPz/e69Bt+Qz3Gznr1iYAtYhZw1
giLGsdKQuDOaa+UzgmkNPfx1Ej0I3xFIVZz4osjTNGnIL8ZNYMf+NE4hDG/GcewEw7h8ZY/MTBoD
kSET9vemyz72+g6XV3GduLNun1Ag2sMneTlTMIlL3TYvgxM/LXFoR23BW26qgELsp+PMTEQY7BL+
T09CsRcJHzdMMDjPG0jyf0jJg2EtLVCw8Pr61gPOJONNMNwA67bXUYvk74ecGSigCxuM8PO1SEmz
rlV0wwQOqzXIyv/MjNDC2Y2CyI61zQtn5+EVHuJb/D3qqTLPNYEPUBD9SaWyEdfi/A2y+Y8JCyq4
dNcojgu1/JUWjcd+4vDw85WDswASRjuL6FfFF8RJNszoFuB4+xNxViCyI/m4NxuvAWtmYikCn9dE
LBm8Ch5Mt3bJ7Huadsa3FC2cegi7wg4X4NPN8dadB+AItL5IKrgZwaDk43Ndpk2rVFXZYCh8AmyR
5tFI0CioXbG1lCFli8APMTf+PK7XyIpI03mKdjo2TMfSp5ouZ61IyUJF0SAOuMazEA3r7RUdZBWX
6sV3/JUX5hoQzhAeEfBAQBa5UrHopNPh4wEcT6MZabLq6danSTx398ZIeokeiPHodkDFjq36qY4B
wPGLl7DEo8v9oXOV+6EFpKuSM660kCgqMrtcz4zSP0CdgzVxZCcYkg6MP8xC1bHRqMsNfAlwycXF
C2VaiPZiY5N0mxS/UTpglqzz1oLCvjeAksArUKTGV4dsPwAGm1QKhTr+ymTvKFsWnJSToDdrbu5X
F7qKUSl7qzaEuHVjY0x+6rqEAC7SloYVhxV05wvPmZgYF90OGD4JzDx6jZ6yET/Os02UlNe9lG5S
ul4xGgK1jYD76yXuVwlQrB02t3A3SkB7SSHl/O91JPItUti7YTfCfQARPTSvqfPxxFgIN6J1vzUB
RDy+DiQwxvbz7YvdfVAvloZTeO59qw6UHfKt7j2DEtRJ5fjRqlgfrEE4iEo/FNDqKqXslqTz966Q
ai8OHFpapKqrhO7YG/KsEXxEwqCDgzh7/Ch8L3fZQf8Hm0KynjVqXC6EQDmHhS/TsZNbkdb+aSsT
Y/1CcNMLA1nFXH6jZ3LChoZ3XNjZqkv/rYXi30DGCUM/yxdTNOQAqX0jhFhKU4Evb62KmBlNv3R1
gD1kXEmc7ELhrwmuPaKlaRQ64j0a2CtwyHGcZaE4QVhV4C2ELfj/ANWapioROtWsXp8WMWodPtYj
QLYsORN6Z1rMtr2ZCVxMdSzHXn01GgKj3a9WWIfjwOVLrl+SMNqslfszIU5xOjsXmzxilSgBn0j6
WFHly2FyZQPoeMqLpv8doMtnrhLMtutbSeqLYYS0v22cN3gq43MtsXKF0SfBtjsdydp0sQdGNHIf
6Xy65Ll24ECDT5WCM7sbNY7gaz5jxtS38KjRHXkgqsivpH/jyHP3r4eq5eny3wWrAZQ7w3TCXk1p
tdJjf8teal9sHFl1LE7YQMUu2C+NYC1VWXZ0czv+88aLsjbcr2rBhQ9lj3dRWquXBg9ii2O1G+LJ
yOVugVXR1TRJHhNGQmnZV0uayUZ8/2E8ITcHNAdP1B5Z6zmaF918w4tGDY1cGzZCs7DY4d5VuNhN
+bYuJF1bvvrHhboYdgUXgGk78FmjziKd1DfxaXFUi47oyM9Z1bPWWP0b2wjLIK8BGkfgxRaehNwC
jx/SfPglZEtmUj+2g+kSGqs2fkjn13neaAzPkeyvKermn3OD/m7aO+/e8LjBTJdz86OopuRceLgL
jn+JG7VyUShBdFkQtruLPRvSNBBwF+RIPT2bMtApIfxsCxjoLPjU+R9Ii1ik5rbMlm0iXqAwYrQv
qnZ/bUCQt7PfanjytTCszfpm6CCUt9yH5Y9g/pacCp0iAuN9XWLI+TxP6iaGINEOPwNG4i5kFwYt
V3Dtp1WC7qm2F2Rd0+ycdecA0K8xr5aDt5NQS7oScvcObXRxQ55YXAMxs9ybJYck3DrzPH4L3hQ5
rcdLQNUE81K14Yn1oO0yfVsBli1xWdOTx+/qEnBtSymoYvm9IQXIOA/amgLCj/I9j6eQJepaBR1O
kkBiopWQXeiiX5hzzvOGzqhe47bMTmqI8EC2GaWjvhzrcv3SgA2sf+AyEVWmAJuCYk06SsI5GVtH
QDcPy61bcqFZuG6QVdnyhwXaXvbHmnye+Ah5cspMvElssy8xt3UCnFtBBcnXpj3H8OArCrNa8vEw
P7NE1iZDGRpXCCVg8lKpMFYCA1pDCRxSs+37DIByAz3BDHu4UsIDR6W/7Eq7GqHLCP335aK0NCC3
orSMfLl3OBIkX5tk10CnAwJyH1FFk7bnTXzG2bCtdB2BNvNQDB/nKe5B7rYn6yC1Yrr0zRa5WuEw
3G6yYXXr8hgCH3PXmASJUtMWH187+xE4I8PXRGv6mNLvgjW/pF1/vMGrYyDG+m0QTOeXnc6EmlNz
hNzUX1acUsYZok1/NEXKjv5VE1s/KEZlO1m6iTz7XWVlbncqmtUVtM5fBxhRT/eecTBI5IoXe2Bu
lPS5nu8VLWaubA/dPfMZHYQkYKLjXX8Z+HwUBpyL9QTH/sPauFQmEHnC2Mz5cXHfbHCTsLiEfcrZ
hrGASOTIUATnQA42JVKl8mhdA+NZej1cNBGyJT/bykxEB0xz22RV7gixWF2eytmH9x+9xvOe3Oa4
uDeTl4zJoqA8KjXWj77zEKav0DxFAMsOtvtu0m4D8ndDmjzohjj6wgNV2wtnj106B71pfyWLLiA7
PyJB94hlMFQLdNZdxWMdGMDfJdhhbJoYLE1FUbtjxb3Czg0XFm9mXx9qKbDkoX4FD8A2AUp5EpSa
euYF1Lwtxn5JLJSHZk7/NgqwZH2HzqeeXso2VGXHepdDs3kckJRo6mP9SRtDJNHv4qUprNLQmoOT
r6mV+Y/WHOC19IAllNE9Qrn5NwVkWzaN0nwD1y4gX1JtVv26JW8LCAjAuWcRYmJ8q6sj1cvntJfi
6BCj6krJWq+IzY41ChVx/W4N1JNS0cu+/ZH51RvFbQuqM4Zc/1HuH0OXI4f09CblN3DDY/MPrtyt
5PZVyeXDQhiXthVvLezrQxhqaE0ueZHy5OvustHahyXISxfhhJrC0iF08zX/ZkDlvh1bUFSqpiAB
9kl6ugIcv9GVFUiNfeFdedc7LkeHTmodcX8mTMoWZPjvRvLrHP6II5/qWcOE1HAH/lPMRuzadrKk
RY2npP6R+JdbzGPSvtLlWXvvSbURE+qDoxTNlc3ixTlC0eJWzyxNpX5p9yr+t7jmYbIoN/pFiQ75
NZcIH8mFljh945GxzsOb22WLy2mfHxDEi2BJ2RxBC+yzVuDuurpECripBOpmKXZFZ++JGwxgb6C8
20VeTUAWzpoRmcmZImiViR89v8bmZZP7kU8gKc3UHO/haydmmKTvilcteylm4IkmNYxlY1oV++D4
ww8yTmWGP7jDZtBzJmHpN1si9QeuiOlEZ6hGtCEtX+A5qzTwLYXVrsBR9iRECs3onGUQnjiVAUgE
q+KOPYIHpRy42XpgKJhDfl8SavlIB/QPWOkcxeMkuH4v4RZ6ZxvJCT2aYxkQ7UQaFHLmjLp76VCG
6ZH6kqdaTvtJ9rPOdZYjBvtunjVKwFW4fxNtRkdMEOLaYBr692IKD4LVVtWqAuKHJ4YCODus3+Xb
k0hXTmf5opae7o9xur3w/R34D/rUtC4P4MbxnlIGjO5c9q6+EtqIrpSe+pY0r5z4/G1rnTb4+x04
07eJnYUQwuA8L33lNdmYzgAkxiA9PTx343hqX0ScgIyUXEBtwoA1J3ZNh6VqpUYHEccRl0TlnkUZ
zXrtN6ldZsXchxajF7zDZoPrsFYf9oaGnVPTPaNAoMOXrK6ZaVGWMXvUjQBRpiILp+hsQZ2hD6Hb
gqs1Tf+cLRzYMGWhYmxv4U0sesOjwXPYp17s+q0uoJFv1OMh9c5e68ii4L7pGR/91TdKN+dtaOQ1
BGUj5pYN8gkAiIOD/qSOPzF+TikBgLdQkfX8HB8gPOYm00GaP6/+mr59mIDUOCX3OGZ3NXLTrSnq
hy0sDNVMxOPobMkLo2CGWJmhs0Civ0OGPutw8t1S4XvXiOwvtjefTrQ29Mnu28wkcEY3ctijtQqe
nESIInBCcSmt0Pxr+V8kbDz+hO/vF9yENr+pF0vp3QWWdUsxfYiKwrAFLi3rH5/W84/HKJKbERFp
o4MZKDTu5Z3RSqoJU49ljRwmSYAiO0wNE+/h3V8vsKryrmPq316qOCEDEC4R3iDoP1ZYIe9p53Rp
TBJyeWAKUryfngwutAqFxzWO27q6NVya7PFv4FOGIv9zkdA/cF6MWgtkpWODXVGKfPkfOM3IPmHK
mdzc0QST/OAUsLGGDuqnL66galpffkyG4jKx13h2oRlpI0oAYW5j0ZZLnXOaJeDawXZcC+1bwDI/
NmfCVmStURs6v+fUIY8/kgq3lovP/VARo2nWqBiAEGs7XJQS/nMUlk+/ydCdngaUyb86T+foSIvD
1Dz6IjwjrIxdd+u2RhcX4afhY+U+wXdUTgBnxDIrFtJbKjwSOAjJ4O387aQdRD5EKrTHLky+UdiG
THSebTBPG16IjleHbWTYZS4cDNg9lMnuvZE4kcPEuc9IKE3liwvHlTH8gfdpqHfNTrNGUl7UsToT
g2g4nFBRQIzIFjaUz2ShCEuGdTlojwrtF6hsxYu4Q3XpWHT5GXN6Z7ZYYE4x9Q+5LewUS6OUqFv0
2I5pGGVGPdtP3uvXjX0DSF5rjaWdfJfA/f24SLRtMwK8GzHYMjRIqjR7nq4QpYbJrQcbLHVEhVJL
K0fwaYa0Gle4yGLNfS5+t8svs6SHBWSmJL609X28eL8O3uBgtYTN5KTaRs7x4enuMKQwP5RWyFQI
h5EMkYlHdRcdQj1YFKzEGIY5wEfOgsHGcjSubTZWuIq0D5/rKOqf1lUY3NeVC704iN2K1ccksO1h
Qc6rF7cu9LogOv/FMxSpiPuhMjSB3nfmgLJfT/oQZSoNgLk9hl6xzq1vKsmTUc4gbPrPPUtjqaJg
ICrPhU1+zvPN9QL7ao/t1veGhytucPG/vT3n0k7HSRsx7E5bq1auwQwt5opgq0J/VF5fdbbU+3Ij
uGMs+JJPU4R57pTPoIQ7f+Cn+aGYYJ4lnYPhJ0RCacEL0me2qD3p3wB6ccrvHcq4bNcJ2waIMcgP
Zoe/qhk4vx0h2E3URzxoLquFpMQBx/RHjoCsosOVMHJHucSRjrExfa0qdTpri300th3rJnRJi2Oz
zLV8x93j29svq2ub+kzDENmf+QrbvVUX/QLsWuoDetKYfcLJ6Iho5P+p5+k8xNpgrtNDOsDILmrR
ST7ch9pvEz+GhDgs/e2c9+by6LkfFPkAsFIT4AvjK2lQNHwQL+mlsw+EFp8HkVK17JBQdEb1GO3U
eaUivKQ7/+K5GTopOIuKcXCz6IdUo+MIXVZL5TK/gP2SK2Llz6ySYUU9eRgup5Lmc5IViRhDPSH3
fHyitrLXqCCIIl2rHu6qRS5bEJQGz83O5nDm9Eb4BakdRYOaZrjDxgeqr9mkmI5CgqUTrf+Ifop1
V1nDvMvCzKdsqps9HvZOhFf2VkJqay7Wjlmz/YLKBR1m4NdmKskEtaX9pRTVL+9DrHk7rNql+j2w
poL4uYQaqT/rTgD7GDRx7Hthin+TvzawZxfkrlBTJD0946nZcjJ6DB4PA74x+Q5WYisT2ktlNZpC
tkQsrZgFtoPh7p1c4KRj2M2ceW9Vp8iv6KkJByX53apjhtDqaXc4wYr+VjWdzjVf1JfsufDJU3T1
gun/mcZYu3A/sMyb5BjEKy2Cd2eXSZBnKPMzfxB8k/CEq8dHSJRYc/YEPk9y+kz6eELeeKe25S9B
RkJX2+93etkk8L7omhs/WaqZh14baLtHtth3ejqAqcj67u4FxOw86Ld/ZUnTtPb8ZJsHttbsMGip
CxokGsoF/QBSql6fIjPsDYDgsC3WvUa6r1HPIF4Xf8qJb6BmgOBlRQ+e6D9T+gOfCjTi2p4UZymH
/p97UOb6azh3mEa24MUBEg/8hq2uiR8WNIa60+clkhDhYhIbtrC3YeHfrMMRxT0YHPqm2S9gdGOB
//w+jjRcOmeF1tAGntlAjvgfQLRNZlCfmrlA+5YnYOwLrGLh62KpgiLImq5AIVvedO//dm5UONzJ
QeZw0+fTnfdVI/YznAYOU17ruSd9NYoJLx5lyVrTm15A64phFYspiGKCylp6yV8gBYzGvjbg4NF+
ytBy/XECy4MiLPpnCu1PK+zBoWRgu4VxEIIeQOVjgW0/aDTXZB59lgU5ipl7u9sGusL5LKwxKjs8
Ez0faRhNLmkPFbzDK/2Nc9i863BIrUUNYQf/AIGsU6JaJXvJ2Rd2hCKdPJiX8gbsxc6pe9OGRxqg
StvOlvhyaew5xrVq2jvds15rO6Pmf+T3BcjrQg/s0okVKlnMbPcBSuN1fObeB2Im3WZLaX/zZh3T
n33DheBkn2d8/QHf5yQCzoaUg3+o22918pfF+mGRNACyHsXNhsxM89WKRhARoaLlAQ2zIU/+EwHQ
Jw90nWd9JEz786ppGijXnNvK8yVVWF+clMfhKtBcaWtnZcb69bMocGgTrEbM3Y42PSsFq97OCyvq
Y/TM0AM4n4p7e6mOdwqNDmH0w/M59YU8sBSztOoanXaf0u04d0kt1BjF0nL/T9yXxD10JzmIAN7c
6BsbXOmFl9nZJbDrFkOG/kyY5oshz8/HOmgyVZsOKPvugGbfHrLI6CDA9n8ZxwJ1DMzuHv2bgS2n
4qNMMlEZMw4iKbBHH6Zl8QOX/1A/UtvlUtSzP8/0/QUrHsj/4/lYLClxgxAf9c49JSNw0K0inonc
Udt9fqhXDxm0eSGLA8pQPYMJmgw3lcNWDuHf52gHVkJYQZGEsyVXrZ/W4yhj1BkKN1StGtJJHl8N
yr0ImWojNtlouLV+os2hwLtGGx1Mhl8O6gB0cojlVsmATKbGODDbq33NUWpM9UlwI1PZu/3aupWv
DfYCLuFTziqx1Pybaz9pmGLaMUB3/u1IyGp+uWvyO3ATkPnuPxxvrsaoiUHzi8gzAeo2t/OhaTTH
7m9CZrzcZ+qkYedxdxpx+aMNFHtrnYhv4t+27OfyK48UE9FJjDr8USIjXtXOg/YqrxYxwY7rDIkg
TOuRojDlEtiAHpo+FITqzbj7up3VUzj6xaxnfwZgTI5QlPdm2+vH+uC750ETrC8Qwgfz8zdpqJ4t
WgwczWHEo/j5M4yHhjwaa5dtqXhTZu9fboVE6eYnBOlRXnW8BLU82/RrOPhDT6NAPFj+MMJMzj5u
j3ckIh3k3IJ9FpFm6+pi6VXxQVVL0dmvHs42AxWbmSu8KMMlB3yUW0/4NSSjJPAPuXH1l087ZAsw
CrKHZl6TaScJY/Gi9ssyA5od2/uJlGe1fVvDRd4AIgDYCbhnRB+UbnEVWLJLaADXGKqlDozYMCmV
khk02GBmoMU4BUJFRjDRSzx17eR42mHQDyC0Y5ywvxgtvlyZid5/bSbRMUplEkLecY6eDOsgcxLo
PoLsIFEcxE9idlI81ECV2G/kwgLHX5hjOSV9FhL/JaxE9NWtfx35KyQcROjVlCqxAyZslwXIEED2
eL0fr3pjHJWFToLqPXqJ/1Dg1Dff8s7sBim/YcnyYHD4OMRyqtZUlBDUIHyQVYZlmwaf8mdSxVvl
K6FzPHG1GuvCXp7aQvAuL9wNsX/Un5h2HkNT+vKly0MVODfiEMHtras3G6/JKQa4qyFGoRir7xS1
vGcGeUPRsl0O2ZuCobGL6JT2O34UMyGM1jtqtYb+N5ZqzZg8yiuZYhRYMFoP5vjSsT/SW0wGQoKr
w+Fv5zcbcuEbX3Yr9qhhDHGIRlQ2wzQCpGUc4xHVYiS7DnoOofVOSTLFQzWw0ZBSVdJmp19a2ayO
lKG3hpTvYqVVViimoBPCv4Fm/W/tLDOWlx70z9nNyuKkpext1Wb0jbooRr4MUTE5yPpTp1zxm3Xf
LoV5AyXjvEOHgsk+E9ZshxN8NiOA2fiFu6YBJmFsJEtl91znw4NR0QSlKUZWAdbR/Y+oThPgoJdf
YMkxLVoHw8nIn3/sIFmG7ax7agBIMuwZ05pmuwuLBk4WsxtV+Sm5JnnV/GvqT5iQvRm0mWrFa8tG
cOnHzAi1OolZSYmODFqH369l9j17HluW7qr4WN1KWTcSmKJrKP+pWbpx+Rx9bbIe559iqUIssMLX
F6QKNqlmwCpoInmYzo8jcX9B2z0Ktq/Abg2yrF8a23Igj68gDpMOhGwyeznVUdnyg+yXMw4xbWDw
gFYRqitr8ekspAN43kzk4oVGEAq8s1ZNl+RDYgpv+7WCgYZE9sUtmq1+JepIc7aVIwboQIWgcAy8
+D0x44wn2ogNaLBb/XCv1RwC1ZmWjH1pPHbRpLPk0UXP6l6Aws3OMAptYMwhCzJPcGXNdQLIK9gp
wc20B+2A0HPsctHPopD8oRzld68BFo33vZirQ7JMfCYAbDYv33erbSmA6vKMlrsNOVMdWxNf3UC8
/7xyJ7TUjkplk4AfuYS2aSwHg0M/nxmZgh6WkEucem8yGWmnOpMargHvPVl8txXa3PX4sft6djEX
eAisoQE3cfMiHADZuQfZGMQmQavrEGJjcgn9T2xuzufvetpUMAoGVTsMBXBX/m6u6Bg8DEQICGHj
NAhsK/Y1lGE68ZkMkyvMeMQciUio73WrvQUfQ+4m9l4gqpi2MbDT3Ah8sOf2NemH3jXYnAHuSSXi
ElbPD3gjrxufVO5byG5LG4YoLaB6Kwau4NhyeimmCSvQnjO9qPyn3OiRfc3QYiDEuSHmcPXU6I0k
L4PiUfiaUG18SiRSeOqdvlaBvJjSAz8NdSblkkswveYbPL8wKO6wg3h6SUtACqWVIMnwAwy6fqhq
03jLqbm8hnJbu7JXJ2GOykh1sHM/HduzoaXgxdiyWPqJaRkgcOwHNxsqSDRF/TDdGGgFTRnjkC9z
CyMAW+t3QYzIJSKDWrURMIeUzNW2hFk5mUi+ugAPvzKRPmiABRhO0eqZZB3468fh4JHvML/3mt2t
j2GOdB1SrVSOdvQNbjAJ4C864uYo1wB1gMAKIytUq/r4Lq8VfCGfwpvA6ziJ12u4P22K+IRC7uku
ybowhZJ6WAYL17BV9abFUq17Z66/T5SlLXQUqu579U1lcQOzpVLN92+LbligSo7o4a/b1WXijR7v
49fqrpwB/bmf7D4AckdohASgzRhyJyIKeLw8DTCUTHv7H2pxhLuw4EE6On+OMECx4lQgUPFqjHOr
S1NNG9fEkqBgy3vNvPIrMGxn8LzrnXd05xqFqXOfn0BpK9huOOdnceMWtZsmr4x7p3zB/KE/kgJi
KZV+UxUJMFauMjVjtt/kupKDM322dq3/a8KJMlXK57SbQYGOwW0vBNE1Szg7Z5uvrujonsUj8SCo
T9GHrniFQRCL4p36CT5OG8KEti5uwQj2Rhdj56bJfg0Lw4jH4ee2423xen56PiDnRWU/mBgGI+WZ
vdQ0Y+mhcyPdAePwrxCWTXEOZrXuvELpzDWb2f+xGr7hzWLgpQtpEB/1VcJUWzucwpbrl2UbMDd1
7CKGwo1SBCnFFsi/+u4YSc125OZfsd5DVBwZRt2H+MN2iufyQzXf38fv9JN0PqxnBxr187k9stGL
NFcSftpKr6vpEZo8dNTAe4bXsekPZX/bSKu7DS3H9BA57l6Aknq++l8mm9nWMSGVo++eOx1/jJMo
/6IYGNCmBicCpB3Wgp9DNla637AfV2cqcbnUsq477j51vEEFS58tpqNSd8DUlbkiopSxXotMIUdS
NuPPyezkMG4S8qUw4wa45/SjXruuRcUDJjrjBaH2x3hEQNcpy3gO8AEdXgKFbpeV+gj+Rby6lO+h
t3PehmTCUczvQDMMA5l2ESZjAQIPMZ2oyDvWxnDbrz0Y3bG4SeYOqjtDACLrjyhaEySlDzA+mN8d
ZNFl6nvOVT3aDU0t4o8GgONkAAuOizQQAzVUuYRXUh2KUX3QK7JmOdwLZ2Km4PrIfZ9CM1nXU37B
HNeLX7DSIgvb+XZ6dsr6K/+vjFKcORSMkcJ26WSvAoxcQts14n+k8cepPRi3IgnGvrQCWMrIv2Ca
U00y3xs0fsROSV0n9b8K57B3ynMJPaDcBROtwkq94BtdsuDCfhCzI3p1A1rCvYy6NLbmpiM1W4g+
Qfkpo+nYJnvFXZHBIK9fdk5czFO3kCCLdJf1C+Slczd2ih62ACfcEeU84xFSiixD65cpIWYjy0xm
5df3cog2ns5/aWLxwTxGzyhpYvTgF87IblVNG2zU/86R70dfvwtEXzVgWCBGNvsbvwtKjveDrBVx
P7wS22bLjCjc52Zi+fFtfKsd6WKiGFuUaLDWQxBMk5roiSw3+tl15K28iRnEaK5BYgl2mXjHE9bM
lSQBzrNnpaLvc9ND7GX+kvnsUxdqGs74eqzp/pWx3K8Sf2/ogWGHp9eprleNrPaySuKlDwyGEcZq
4leC/sRKpxGtkMyz5zm5Ml3Ln40/5sLa7d25mPSFHFIh1H5BgxMBh9bAdUNaath78iy/mGkpLQMe
6+jUB8T2AAV2s9W7rWqF2pxmZqoPz869CGN4cGM5X13OzbegQlkureo4GBAuwXOvUEL8S/9aYMkZ
A172UFwDNEtmx+QkOm5Vc8HoLJrMEWICRQPdQaQEk8gwsMAd2lVOTQJc7snFRM5Jdq+z35g/c4md
hBPsJAnFzeZZDqOvj/vOl6lhhlY+Rq0l5byGahJzlOp+8jtD8vcXobthL6XWVS1fNk0i0nwLGql5
oJyQs2uIYzA6iaJ8iEmaQ0f/qkXJA0OoJ6j2V7uIyGMgzzVK9nw5G2/BVZmjcWlaKYbeeNaASl3I
fv5VxoSgrooh0SnQUCzLBFfjw/x4sgdlXxltqKITOas7XQhhMQy3ZF/6+4iB0bOl/DjXUTOHD5MT
iF3DmYnVIPF0rpQRmph/Cl9sgre5i4ezNPYCz5lg2XyGrhG23/w+pe/JXtJSpQH2TT0+9WQv0vqM
940S2VBjdl5SCWu8YkvZWM9ZwegoCvviRTYANg/TJX0M8DGnYkbgS22ZoXbLEPtPAD5/hab4kI6+
q06A2vIBRSW/oeNg098s7QLG/4MqyuyogTuK7QXBm+SgHkuSkvnnLNICIqvGDmF0Veb/8D7m6Cdk
kGD62JJy4uFlP+Bg1Qo2rETDJYmM/fUtua2fjvRgjCDsvIwJA4HV8Pft82wpvsX0sU95NhllYh2v
0Jp3QM/5JS9Irtoh+I5NQJerH0EV3SdxKdJCTHYTm4VUHyX39qhNRsyMIDvNmLZ/kusFx6V088Xj
3FI5948L+m27T8dSOy171FkZU0Laxz+sVKsj725JjZ1HmZfPlyyO+gQwQJO/05az0HbaT9H9Rn6+
jjJkg/5WkNzq8qHyZXDKP+/XzCpCCCsf/S05LXS3jFjIpdZgp6Y4RK8CXdde74Ec27VFd+hQU6SH
S/kUJmnYluI6dqlQ1pNm8zZW54z5N379OAswMtIQ6PCma8/5eTmfqp+614lz8Dd+lYsgpegIuVSs
BUTjWnRL1M4ypBO7E7a6TEDoV+fTNE1WoyeA2ipOVdqU85Em4Gdg/Ie1b8AX4xeYCI8wOyK0HuMu
na4WVIlVyIcOs2fVI2oyyjc5njJPnUNblw/9sprsoRp6dR15W6NXKA3W+TrFJ4q0wi/N4aNw+djF
TNIOiuoaW2R04kC8GhLgCt370ylavgD/PfSL19VVQhyRq9j4tEJyx4rMztEYsOr6tpMWrvQtH8yu
2qmra6T6mpPaI1oBQjuFgYG7OfMQgIC7hb0b0a1pLQU1w7PKDlePucf6Krf6bg/59cwmfPOF1Iud
zTlReIQkvUXTlkpQdF0VJol7OyM4mEcyDJA/4s/Zg+S//xeswMcdDyR1M2gNCj9rJJ2N90YhORHH
3KDOdXONufHicu0aVH0/bHGTmZVJmyhFWz8u+3as5Kjj8cPSoga3GauWN6DQVmoXb0NiUWOHWt17
Q7+L7EHnkBphMV/G9XKLvRuHDxa4wuMC+BFuT+DIO0l+XCmhSzx+Op4R0EHDsgp2xI/+RCxWYBm/
fCypnkInLeK5N2w5B8q36kpkjaW46iacHwkcK2sGJL8biKDa89wehURQjEeiAtXt6JQGs5D+RoYd
JQD4ZaD+noPcpivpC7RBtHU4M/N6uwJYSoEQg697GgHlANEQ/h8YdFEO4wS8C17/p+j1H/sxEjKl
Ngxw7zGXYS64SuyHusLyaqYf1JWx+s2Mg9U0RBM9T3ZOD9l9x11J6Ga+yAXCgLSZPTOVI9CnGQD9
qe03Ay1ZBJSpxA3YOFqeRQOCXJOsDRBxt34tjMzZTEZmciVrOy+2KbhF7qyUdf0aFCsA6srFwwco
HA6sXDEDeRitZlgABVfYkeeSaXsYSCqxo1WHzA9szJuhiMOGOzQtcquyioKecoAs9Rk6IQZ2oUTu
fkXvxDBVXIjDnIVSWjLcNLG37RI0EqodLpMrCjIH4SFdrn9GOw1UeSGxr/J0GlOrP0OeVSXnNwxk
fde/Fc4PeGo70DYdVJvf94GvyUJKOCKF2/F5u4xCbIFHgYFXJNjMnOs1M0Sq4dseYSxoQVXIFyu8
AUHhisi6A84qPOWeJ9KGSljuxYBRt5kolSGvDnKzMD48wVFjP5ROnAob++vUgydLeyawk29Ee1AJ
BdTMDfWupZYhRG0Yn3I8E/79G1fymqW9URJgZGOckT92Pvq34N6hjAX4vO7WPWU71g/0ibS32MAW
lFUVOWcc37lNKVviHlq55ebp8oJl4LLRbdVAUatS0Wj4vk98qPkGX2cO/8BqLajaqlmrLfB7vK4+
qajNiDSH74k3wG7L0XBZXHHVfEBrBrjXxAII6c/OkKWDG2/au70P1r0Dp8ebbxuqhPbaCAucbHtx
TwhE6rFbp1AB5c9Lqpm3CqeCt8mOz46wdGGY6URqIxhlIoexvL4CMgVdlkrrC0H1OTUmMbQeMcRg
sOShqMKOx05IEIlRHmsJ6vPkB+Lc5/uhDdaCeBpL/+4vK2dInSgs9BeJgRH0EipbqfOFU4OKDncp
oeKkecmNVh+dTH2ugrv0V3OvRUUjwPsNSGrdqZLfe3zeR+gGUXCP0291IzlgoxtNTRTDKjS9wqjJ
CQEUWWfW0MIu0xtGxDr0FH7nnQyNnkEqypdxVwWqoY6E6ejmLY9cRBSabbJrtTCZn3ySqaRYxMzS
LTM7mY2oPFQ6wXgB2u1S6Kzz/MBHtFX5XBv6I+OR4qTebgSLGIp9jgxjapO6cLxuVw8ZuSQ/ZW6b
qP2w74V1u1mo3lfu4v/STWnzW7gcHfrgOeASO5ZdQjvjkTVqpOPFHdnyw3R406i9Q4BOY9k823V2
wayHcgIhVgaoqtNA2agrLXTGl6KVjSLhzWUI7WfkcE9jpWs2a7BLBZr5mQitDUFnCM+FP+xxRnYj
L2JdGUUaPM/Lp/0CX/DWzRw98a/gkuJtbhcZdZzIP4k9QmVtG1vXgYUkuox5eA4K6uMChZu48oZ+
SlSeZlKNkYuu6Hwx/WcszECftmjpwLkQa1aIykFXXg3+ZeLtUgq/IH2hxvejacRCLJxhrhhO6sCA
rX+aNoJLOUO1e/MqZeOjB3T9jilxTvyDrQXAVEpq25DIux6SunTnTSN2Rv1A0w9++CTi4Z+UV/Gx
760+4HTVNAi45FrwXMWMNzLbO+Hjsuj6HdtA968OCdLZBaoXKTmum9O/7YYsKlMHaGT3FAikTPqf
IQJPLv0EsaR6Nj5VKGU6RYFt7OEjQaa8SAFkQuvTKvDnhwUOIW1vRVYl3yZ7sMJvCO996qHb9rLV
TnF6rQC1sENxZHDQCLpas2Lud8xiVp8NiK8kDJQ26cq6+EE3WRSP7H6+UVvP0IuBGYG+bne74o2F
xt0Gz5fg0ODsJ/XBbERIrrpMxc0lTnW/0Bk8LX1DZBeVNcaK+a4dPf1XBYwGcMMcqZzrh88ppwo8
g2gyAoKJPtBsqeYCShsr19nXcPRclVW4qRt6zDw61ERaIy/HsmajhnXoD9f31/jgPkqm539vYRFh
mZWO1I8cvEupy1b4oN4XojLRlbC9D06exKcZYH3JouKZ68VRBVHRMx9274loDlcF3vl16RWczZ59
sQV3ffkmN+50WlSQ9jkUBU7Qfma/iHKHFWlHvRNSfmD8Ji/N9r3YajXnGxGlrTOH6aRknteExMH9
Xvh/QTDrFTQhbGgh8C+l7T69Qpe6VOSK7v6lR1ebsIKFS9ky+fOYgHY1RzaBiE5vZ3Jch9ciiyKQ
+ip05tEOBKEFugyTsuR/fhG/Hg7xsWi+K17RlzvAbaCjfCzF1jpwXgjl4jkBJoQ/apm50XdDqMnj
iJEIb+esan/p1NiGK0In03XFikMw9/Zw5fh11sTmhvjXoFutGNTW15Rt26uCpJ6FvlxaYPH4jkFf
+ROzmBluw3SNPh4tkRmxqMTXlYdN/IGNV66q5PkGr8ltE0rkiBdg/SDWabMWStqS+I86RaMuEOez
hbtyVdE2E/J4bN1rbKho9qu3xYJ0I4FGIU0uuJDf/wJmf63lrHSoGq4GbGVRfi/A3G7HcaHuyulB
33y+I6/tvPfqrQl57QUjKhWUyVmxQaihqYJk4+lNY9swQAjcIL6+O7z6kFu9KDgQCEWP3QJZeOsL
Svr5VBy1POg2JbyTE1lVL1Iq5NCfaZJXWT88RyV2d4NyOF9gTmMAGIU8OSacEhzOSzhd8/u27zc6
BZBAd27IEBda1w8tMjBG/RNWvlWkQ+R061jEQM0izJglWPyYTPJOEagAKLcNMVg7bm3Rc2mKZrXl
JQMemAddjFfXQD5WhalbC2R7ig4qZ6FnYXnJijnrFlWxJBDUAWY9btj5SZo+y+Ed98p7DmhdBmOR
qf9G6o3vWfTwHBSHDAmNwjb2s6kGvrSDb8+iKu79ZbH5oKC7hLNovkJVLntgdJFZvEQvdxz9D5NI
4HFZhdtmhqoJdw7WAj/dnJ4v7gVrL+aATkcxMbuSOd+owFv150ImGZsMK+V5fIwsG+y0UefTkasm
v3NHILLK2o3assstDyDAE9CTYo4NOcxRX7hrvHI1Vhn3/depOIR22++AX1tRLk3MFS/kyiKZeZrx
NbYK7z1z8dkeckr2phpXO53Wwfgc+se2OxzBn7GFErCo4cw0oe9vzmPuP0SI+gU752W9HK8uaMvb
6LuEx0OVGUCHPTy/zwGnZEp99glWZPOsiw0hO3P0vMMPDD8bnWA7dW6yFWh8EeD/ryDzCsnMH2Oj
GzDozf636N0exYBlp+afWGUki6bBgdIMytdWDkqRYEXqhgDCLk30cOaOsHVlxpQOrPfRdAUHdh/V
d6h87du6bjr2azGNgsh34ZyBCT4Mp0loH/Vo70KwCsEM+bC/hkMhd7KnTOhics74z4/UCWWnNOzH
Bv6H0N+MLBwkkAJrBSGsbdoWqvW6d0UHAIhoEc9H12nAwCXkRmFgQJjkTCKzJj2tcWLECrmBGcpw
UuY6Zl/NchRJL7fo6sDwO7EyBMb9h6cLO3TrJYDSFmqWd6bqdWisV6ZDl4Xt5PhgykcorRFhtxT8
yByTQlCYzAMAAYKBetjY7V1c6E3xmigTl4ZMlswfmJEIuwAUUrT2mxjnip48PaiYMHw/Fiwp3z8Q
NmclKzufIjDkT/VTkcWJqLLV1oL46vWOeegs3rL1oAjzgLq101v8B0YDqypsiopBu5+un8cPsOv9
YYNtHCzwEa90mF0EuVCkBZFslnOcQk2Qto9acvLe3prRKzD7cXczVuEYS5wyiunrdPtD+cnMOPUu
ubvzAGIuaGacF334aUHgqZnd5utBn4W5RVvXPFpT0mu/sYf5E2DrfUV1sQAo9Paheqoba+Hjqouq
VCBiyrNByzEUfFqphv6Za4Z1ISXqXswZhGaClBFSdnK3TR6Gr+48x6WgUnJ2fJ5lgnG1hgJQR7gj
EjAWi3dKfn/fm7M4MS0slli/fL+yUDXlxKff5inUkdt1bClbdtIVuspUtUpi/V8gmMGQJ3UFJ6AD
NiUfKNEhC1Eebr6X+Y1Fy1Flt5z4+zW4EKmmjLTjTjfLGtfY2bF4U/rs9qaCsk8FjnANvt9HtWp1
N/txw3zzvg8ZxExC+x/g6COq2BEGkNgDoprqsW08W2ATdu21jajZrpUu9MvnCIZ5KwK2wWxK1Mor
pqN7v7wcEdPignvS/sQz2iGA+2BoH6IuEDljBu/65pKQDknM6xE/pT6qsCmG7OJ1RgdgYyQY4ZkG
cUOoaWTO8f6lZT1Rfvk8cTOYjoOykgeXkl9hFl/2xq5uKwDH3a5L7fmlL2PseIeBqw91+AufKfnE
tRqblhwH5LVCRrQa9R7Y0+cSPtBwRkD/soYFWbRqEpfKZEkV4MOuXuIb3cM7jcBy02Ol9SAZhVnv
Mu6xFSvOS4ejV3/2o/mikq76NTuCqju6c7k43psw3hG3zROog0bdztBBEXRSe5orPUKCeu5LXy+P
Y0nsaDsL64ehz6+qBQxuZgtt2Zu+TWoBKOuernannLVWZ4/Um9pDa2tfPrTg96fDRoTLxeZlnnCc
E+/SLA4C/o62PxGzZbzEnpgLNFxq5ETLnJPGMAtU1ULIFEwjOwFc5ZRjzLTHZ2HRwjVEtCKFaG3X
4fduFyINZ79c2A/YzQP4p4XyJATRA8/j3tXEEVBQrOa1GBUi0emTJKRIm9gN5aBiQBr6aWE4Lk2b
YipTtZAXcJLMLLz6lela82u++DsKCEPWR/jfnOZ5Ob7AZ0jmM98sC4NbiUwCoqs+AJeuHPFDhr8i
h/LIBWWBPoGP3tqdyhc/P7tZo3edMBjPhvAdnpfTqD/us+G9BfNbtxVkSwgCSdGLopi4kQMONham
kyiDRoeG9udyOY83eXsBB/+e9n1ytLBlp2I0TsAejnuHkz4GE+wNsyFYjMpu6n5SLhhNaMEp0UEN
pM7DBRVevVJueMypSbYnL3+rH4I5K7ZZ0NBNU4VXsfaodWvhcQfNLGH1lb3zwt+LJKuy3ntOQ9g7
5Q+aBjrzyU/a5QDPLB/cnj7XdIsHZ0WLfjQCLLX6KSxLwVWmlYtmRyI1U37kICgxgN5jg94Bz3CL
jAMoK69c3z1Fg42FEJGkwIEUbpAaKiN7toeEvuK4mURTv42lCWyHNMSk7kU7banKlC9S4p0Up8wK
sbqJpGYKJk1FRYUBJ49hhbPcRVAYYc4C4Qcmd+XC2TyZHQxsVJyOXfN+pn7RnKs5NSyqarVv0AmI
WYJZgl3TBZrGC7z3dzpUNLk8T61S73HkEzvgcbDG35ZFmzFITyepGp+BbnZPyO/SPCIhcas+Q2o8
+ceFjjxirkrfkerQYs3+v7bMhg/mA6KnaKHluP0OryzhHLckRzGNzgLzZK+bX3nAJdUeUP9zwsd6
TAno12KNCFIy5tSBgv943c8AhjT1cwxTTenqNC0hxYEY4h6j5rhARMzx972kJguPH2oumibukqP/
+T+QUklYcD4WOzDFp/aWpFhLe4T88NoFuoTjlifv+fu6jmacGQer+DPrjRmR8UThos5Irm/gQ8Nn
GHGen+k2gEUotpEFnLQ9Kc/m+kxN/IqkqxBuc+yZ0SMSvWK2QW0dRzS6oMunXuoy8gjHz+0H1juc
oJ0GoE8oSPhHdRehqmHsWIG8aNCYU+Cs0SSWqvooKKaJxRfmV40V0kN62FhAV2MECXpsbZr+iVTV
75toGQszUpunGsmhuhpwSeRZE1cmgBLXNSSjCOQM0Xjar1r0fMpLMLWVeIvtyn7SWYR+SDCCzeHo
dXua71ar9rPurQDcCoD0fabOyWb78Gur2FwXKg12PbwljRq2F/0DWreUG7i9TCkyGN24apHZ2FSC
AFCi0dxZ/JopKnK/2dtNGm8wIH52Amk7+fY+2vtvAjHNY6dUpZUN/KYvIOekTOtndvNtru/p31v1
aNVb/GIrzkmvooseq6nRjiQP/3+8HNGN54aY7+ST3t4T4Gdobs4vHaGwSEPmVcC6rKjHZCfYXHHN
6+74nOgh4Hdp+mrclhNzmTrKdk6dIM4PQJ9fXHNdpZhziOx9yigeunLHSkP2IznVZRee9Wk2v7x4
mdF6vZoc59OiGroKS/8VkhvjITzHUmbB0Z90sV5P5NoLMEAST62D3/FWTPr2p7OeAXhxC4lbPIlY
T/PJcJsxZ8m1SDlTAlufQ/jxT/FVUQKnoM/GR2Av7cAFTpsHhOOvHebAtMBEKEdgd3YyXeq7Cwnk
IdA/e9HA2FzWkKtpdkLKNUN4Jr3TrAvXagvFdgaej1nFgPfP73mBqBJBBCdGJeJHm5/RTnFgGso9
fhNRLqXzCRjSm8dRXvSLiLKY6kXhGHGrPZpqFDYBGdK7URtofgJrRqOhwzpmUvbhiwCMq5b4tdne
YZG0ICevzw0DvBmQwGx5Pe7s0+CTERnWdwLIgUjz4q7udBRH9wrp7fZ4DZc3CApi2e/ELzrezwT3
v/dxCzPrl2xQBXVwH6+UAH9L7tIrNvPH3W83bsabXf9DoOW9FuKoUjhdaSEdb5xEKdYaM9gh966p
NUUQqaH6fFAlswRiKmcs83M506XzytwCkdKLSGWmFfR0p9M+8LxudlX18zlEbCan6yRYcTVYqX90
IwBUSsBYj8/xri1tH4tOROkgmnBaMPWHnh6OKNZbSeyJHoDamqVt/de4kggHg087IAvG+gNelfM5
1tcDMxL6JrshZ9hz8PMH6hRbZcKa7XOwoyjNYUS7N4mvnJekEMfshaUQvSCGrQ7KB4BFl3FwcqyK
q6bPfClQDp3cH/lbsMrbXQ4Nk2xYcCARicrVYBzNA1kiXFyepN5OtrRyPyXXUKtGqbH+B6hPjkqO
BO726555XpS/0aNDwH+0+0uKZsB9WQzf7a6btbNWnps7NavVQp5dLMTNWW5A6dLhn+LtNEzaV9ix
oCsyvb1APMOIATyJJWRYh94IukV2OE5y+d/cGK4v0Z2uic3YphST2nJ+7ER0EoytEsCME49qYIL2
C+LcL0LhUR4uWFGU3DaaWe3laSvCNlvAHKuBk7EebQHjuW5Mf5QcLuZeADp5viSPyJ69Y+YOi6ra
Ck6N131rwTqPQr2Q5WrRjNJau617QvXNPksZ6tFeU2CR9n8JHE7coXG4yiVuRivpXucKyga/9lhB
mHaKKqAKTPYLr6UT+vwr5n5pTadhpQrdgyk7565j/J28RSDRt1zHOXZH1vDi2xGAmBgseJrle75y
Ov5OxE6z6bFauD2XHXKdyvHMyc7mZXB646nBpelSblpk9d0OJLIo8vWTHOJO+iqhMhzIs34Zpcsd
SuRR5xyHzM0rfk8kknvdXkzh0eijgX31xRW/Uu+gksYGjTG7Y05RRiBLu3Kez7oLFa3uNJ+N2G9C
oTcLVY/eVG4PTnD4BlTeu5X8kNiiMzCtGgaORuDQBY3VbrHjHjcZ9jRgZvLPVCe1h3/gLMtUnC4R
dT74u+2bLRWPuhRuhzFtp0zWo7Wu+WiM2/9PROYW3SLHQ5+VecyX/9oN9ZT7/VYYk4IpCwsluwzi
/CnVFahVmCq1xtGeT2GoRMOFQ8XkeoikA0EHNpt/Uzjl+5nTG5w9oRIXF9vzMVVVKExNCXLHeqRU
iA2qzbh6MlFhiUQwvgFZzch0nKXbZDmK2W4wEuOjfOz+4Yoca2kxZmH2JHXObCRTvP1bVAx2A3NN
PR1BfXouqYTd4vohbQaMGK0r/AmxwheaITVjCu4klmEGIiL40+rUNGBQipaozGEEbuRSNQ51POJz
cGxcomREariXFILzbHP+VAmttmcQCC2RTO78Ccto2TpPfnkv5a27vsiFAZWnrWFLptI7QuaK06Ai
+VF6SsPgNY0rMsk3j957DnuZlFmTvpzWwhnweFtX9yojAa8WjsY0o6A+Fordfw7Xiv6Y/xiom0rN
C4RvtzrviZjPj/cNJvHe0rb8s0pGmzJsVQtSL5SGmVjI0VwgspO8VQY+XwIllEY3RUckLJZ1aKrF
DNYLIWmSLcsBPZ1VSXUpuAhi2eSYwxcXDsOr9yEtAv3rw9EC6WfzwKksdcsfw6EN5SMZLwCuMv2d
gNEOoGpjb76LA3VdHoM1+YWssdmjdJgoqf1l/rnJ868IzeZBoQli6oqITwqnYVkvJaISYIrw3cn9
ptblfluy+rkvPOvMqzzmAibB/jfB13OL7XnPC3bodx3uT0Bgw7wpef4NQdlh6ZJZVX432Qg7hFaj
79rLYCZsuwrlytHgoZZ6RzlN1NxPiR0COq6JN+3BJYfmwLPdYemfEtAvhvpOhZz0oTVh8iSub4Qk
WzmguMrEwQM4LdAQekfydG0EMSTs6jg2B4wBQ8mUsJUriAN94ke8pTNKJTJg3DI1aYqPNGtm/mD1
q2oBHkJAoxXXqwADP3MN61JiKkr0AJl7oGMXEvW39TmCQ1+evxI4zd0+ETkS0yVYaojdzrHoVUSu
IOv0ZSGxHQzljqsQMEX30LNAihIV0RZ1sadGCMElsyk6ASdK7vyWbJQzx8L+KdHWpKnHHGGKuX95
NkSVPHSeZqZOR4VhIZiQWG4Ld7TUXpnijECgJDQLx7Mi3hFqHUL4r4CPhmVJpApIQlQlwDm8KxMN
0TsHnZNPkkVYdpss9EsJiJLSzkV74jaWoabttOkvAyHnSdjHDDlK9gEznSKhtYo2PrXT49X96D18
DL8brDlejOlqNNqJDv/ikxMmVQV/qEnXWYFwqaGVkb6gnczjlD0thWliG7toqjGmZkqdG+mGR0eq
WzOZudhiNvD49r9CXcLdXg4y/fWZS/eHV2pyI/vC9N/tkWLY/kbxiphFwaMaxzsPf02c4IEjiQps
Rx5dUUV00Mns4kX+QyJ0WAbmvjCEVfvKQA85Wrrv3i47PDDTfbOoWnaJ1LY9rcXM9zbjki8RNzaZ
rT+KCnWFzprIyx667bFX6w+kajp+vAdEe/luDvWLv1im1j0l2jpTOaXw4dQDNJeJSle6DerW4G/X
chRHwGrYjLGsve7pYGdINieLphS55Wf+oksDg07YSGxfW77EPY1n8IAAbQDA28nBJ46zoCGwdjuB
dRudHGw/mgqCDvBg9gYjtGnDa3RgjH/YCdu/xjQmjBXh/ICLdFFg1GqpNwobEqNOD2E9/LH+YgqR
ufv7oWnmlS+/AsfSd1wk0fJgMz12XdfE2Rr4GRGvXwGLX/iY6UPw/tv8GJB+3TaTOOzkxedliGQx
HBXUP1uxnRAFP8pIVgZE7cOVntCTEaWhVBQ29JMXECcIup9pfEgcViAcnyK76uJPAo7/0t4+n0lF
H8viBtcGoZl2MEBe1OX3ISQ7zfw0JONfG9Wfj96xnHfeeOGNakwRGQuWLtxfWHAKUfnf66WjvUoI
BYIJzfrD6GS/g83TLfZ7SIggZ/yeVgX6LrejO7jM+IwlW66ZrRS38zQ/ALaUP4a0d0L1Ukx6AgPh
6HiVYwSRgxf4gNkDnr1GmD3CeoWUZZx9pDhdTRvp4Vsrg42g5tkbZp98zx7D0ZQBTxdREEwtinzp
LksY4fZmOp7tiopgcwDeR2C7av/ZOdlkJCJJRypSwQ4fE1w5g1I/9Wc6ZEBRYbN2v5kF+G+b7SpV
+2dz4ThpIOT+Xv+B7Kcm/C3CE2osm3dXcEAkE1UjCxdIBKj2jBTzTU/j1axn2Ys1zv2T0WfSu4+5
fUh8CbnJUt6lOMo4byfjRA0041yB8weqtzRvi6kaKyvOGb6U4sox6KKjdf4q3I1KTle0v3NwtfjN
B+ckwciVjituxXdDBZJ/tQVv0tbYRelzdEqZ6cUcSHrOXoJQlZXO+Wrzdv3A6DSsOyZT+KxYrgN7
Z3AkA/yerP29xl/6Hv5BqDv92BMnyZH1SB4/nnRaymtqmiFt9qYbDmAxdByXF4uQ+3Ce7L7B6OIn
bHuPnq+bqwnb2ojJRQhmIPCfDaiU8av1YAfERnyFavDmUnxevS/ii+XLEAgaOEco+WCnWF6SHASD
hEnAiMV5HWijzUyWWj1eaoQJNh2fTpgkzIlOKnZ6Bqz7SfPpbP/t/FaZ9e+iPM7iTj+kXdcAxrVT
HteQjMmIr7J02MGGGlWYA/LZmvq8MKzfcaI0TP+pt7OezdJa3UfFhdNfKZRS7VQ7/HXkQsTDsjyA
ow2DyvywjSopSkio5FJXj1LGF4nW1wZKoy/uw/zDf98XMyLsT5qD1DIoSZh6E1CWc0cOGI5qp+z6
zDydTvrb3umncetCTNP7+A58S30DDek2XjDWqhtpFP8KZHf3Z29iRcQuJut2rQCJOuyRXN70LzoP
aYew5DOD25S2Nvjjv6t47nn+GfljAfY3hc2zCegn2Zu+OM2oz1fesPafihp/sWdFcysU3t/n4XNe
OAxml1C+jbmLAnMAaICHS/5rNE7Pr+pFcSIVCVLTSRY0ETIXNrIlfypf12Qh3izDXOARG8cvp+Yu
31rxHh9wOVsNv48hNEztZCe9QsnaWz+6kWeJU3WkN6mrDwujR2Cgv0AThILYoCxbVGKHxio//jVC
Q6CX01GfKvNeGG30089avDWP3IBBSgexYDTFrzmic7MP0IXdomUHFy5M+1udrReUrmEyNsylrwBZ
cHc2J4pwJkD3HcRNdm72w+gkaHg8jVd4hO0FpunLgi14lNMmZot2QNL46pA+soO+litCa1qdrTWH
N3jPlOOdWSjn5wINviyFXvahy/s+8sSgx8jmA5VRXnQBAoLR4ImvQDCaoSsYZkh2uZV1r6u1znpv
YMRB61YY3f0FBs4wHNwGt6zzA0vlRKKmE/YlnG5tbKYHUdz/d0Eqbn7gGxa7drbkyvmQYL6I4L9s
XOtrGz9WLrC4ckWOzGAQCxwvLp7kh2GBNyWuQWb4B+aXqcYtIayqqEUg4x34Lf+sGlMIRwO1g6Js
r4sV2YdZ8xcXOe0NEDfVMhyS9jiPEQJD6WLKuQ2Okx2R6FsA4Wf1lAcwtnT1xeDBXh6Fpmwyoltx
Sc1Ih/cTJxa+Yw88UySQdDVoK8oQ5VlDMnyWdapyQIxXXGJm4HGhiQvmPaxU7yVqIL9mD4+QS3Ze
cxNd4w/q1Fim/UAIKj75WLb0ls7xfpGpFI+f5p+hZj7qqbaJjf0LQIpy4VNvOvRdzTLoNtejMF1j
e0HHQX582+kHTB83kX9CFEy20kmibfUd+a2v6RopXGHk9DmzH0cnXm6NYOtG3c/kOY5gGCbEx2Bu
6SxgeJpy66oe67hNsA07OFUXqyw0fiVIQg8FZRZ9RN825zbHrV829Y3hRi5eqxhretiTKh0NEsuJ
rFwGTDRfD+9VoD3vGPQgrRyRCd9u+4p5SoZtzITAzE1TCJ48ujVwcky0f9vmAsLV8gkI3i4QK552
gKwf/2FopN4cCc24Fqu4R8EzqS3cEb2trofJJ/JgzB3c7cAkq128yWoxmQAK1W2Xy/wzFFdSd/Ni
95eDyl6qBsmbeh45Pk5tjd69oIMooAMPgiIv1nIgBU7VLrUdW92Not3uGN59py09Fm9F3VGcIcg4
VJeJu2EdYl1hJFK5KTud9EV9K4kMQgreoPlAy8AzPkf15veiabOnJSHyo7DFzVHmDA9iAsJeR+Cy
KZO5FD9BgjU3KfI7XH5OJyfnzngz/K8fo5Q6RM58FsdGdRT6CA5/EXW13RB/jhscCg2mlyfu5gXy
lUkAgQzvxHZByJeSSQOxCdz/Fx2FIAGCq3JOTtZgQrCAUfP3anIpB952efbdGoVqud5WvkkC/gMI
48g/AzLYe7vda8c2x5q1cJ2evzvbiC1ntU4tjxGWLj38gKqtcj3qXDLTW8PW9YPbZ/NkN7C6+N4p
ePg1X2PCnq9YiV5E45W0Tu3OXbmq2ljoI+OFPb0Yhsk5BI6RvwfcZ/65+hBFgxFTZWrR7BjhxRFo
hflkCuDurbslH8GwcqZe1w/cNM9XaBxgVBbgXT6OKCfoNRBm6G5bLo+GtOfrirJE2Y1jooan6IkR
hNsh5gSxSgOATsUVfSgCPlfnyFX5TLu1ZkPe1uUQEyoTilthlA9+sOylFsimmo3Bik+ISXwHApjr
BBed3VKN300ja/Ep7ncrOdTHIwpkHHq0bF3FKQ7NN0XomlJ0znbOF8aZ+BKrcRvzgGi+atKYMNrl
S6aEjG5vYTUNqBLHY27tb4Kj3DkL0xVanntn0iSYhcYBbNh1W8J5kw95QULxh60sKAOhnloLS2LP
9Slq6AibSFJllUNO2TWGjICy/I4VGjNo1k54YjbtkRe3kaUXtOoSfz2H/OIH2F99Ok9R+nBeLR25
nc3U/LGHFACcj1jGDS/o2V+hZe6eRGt8NvKhQM0q3ilVusgWFSZdkZydE0L4bFGOvcp8X542bGxD
RtsvJoVJqN1JHxh2bLLYFN0IHlJls1DtxCppWoZAoIf1bmByWiabKqCXbdcj3v7xpiJ/WddX02cS
fsgECZxkwNmAh7x+a/1SWXyqbTImCiOieBWkF+GNF3+rmVARKxO3Lc06/Jgxi0NB3KQgFivbsrIu
vpUCiWcxEQLD0SXfR+PtUIhQ6MHtQlJ0ydYdckUOip0iH9Ba+6fo9i16HYsJWdcgjrhefyKLs6FF
np7d/Dlpzie+Q/loFbjPElJluC0DJrcJ6E/Nde0Zdyxb43S9ARP7wpXLbrYMxOy0Ss+1S9W5GuIM
RN9K4GEi3vyjY/uXBy20n4TVUQ0LFlqnRIy60MQOVbUTYFxRTartb+PMP6HyashRDnuQFxuLf1+D
gs2LAQKcSsEyjogUurBYzjEpk4sCieNo8WwxGuF+RELRK31+cTk4U1X6v75syQBP3/Iisf9VS2X0
IIocq4f29i3s0FrEbGYzjefo/uxJMRGnC20WUuXt/YKsOjuf3c5uGVKIXEm5yc6KxHC48kGDVIHL
wBdQ9rOancXNqaKakgA5cYdjsD2EguqXmQKRIp5c7ICNUfjRp5JMTgWh6rCYY/nerZ5tC6YJgGOw
+1huRS+vZ3fHSbebmFR/5jB6MKFt5Iz9cDwz3Ff4yUkMDszDcEVfGGu3byUIK/GI9fVeeRFzKBEk
DMz4GGKNJnV4CrADfePFl/511lCG8vlJLb9rBkWNCiHG8//MMsOtwj5MHwxSp9xcmZg5zjDkSq1B
9O1Cqr38u5lt+RmikCWmfBZcMQjT0+C08PP9D1w5wo62It2q/3o1KczTOAlY8WjgWlTR9xzVfv5C
eK18ACfBW7Yg/gBgk9u5QuY2+fatRRFo364Aq2m7M+YIAl5Su5ussPjC7J3q/u5INPKAKOkeCBuG
F8IwYb/o6fJnm3Pfcl5UrPRggDf1Rb5/MySmpJdtBJ8t69ZUJvvrrzRRrkkM5gaRG7AdQXBtZ1rX
2alB2qowU4YZVpUM0X9SMTD4HPFK6Y8SL6y5KUHGhqDTqoQ4YXzs8GyJlFjAHu1gWvuMLrisCiso
EdUBec/AKCcZ7PAyTe3k12eByq0IT+sb2sDeciUhWAOXvrS+lee2+bl7+OP4toxpAkU0yRDaLZsg
UCAg6IzZM8LYih6QdzCT52ne8v5Qi+KwJyTvC2lZWOQ88nKncz9dxJuF7gw4dIw96rI6sMgSJsTd
hYBFFV+RLIwXqMzLb5qNWiva7M2YXasKA4fp3vgzEPBsdgPQcksn1i/fEhAjXpLfUyfJUCCdTv5B
9WMpMfVh3VMk1LzpvQgJA9cLo3zHutwvLGq7VpgJlaZgz2w9G4pziGDXOYxzeZzcLPUktoO6gUJQ
8XM5vmwwdcLlw5xE7G2SmxaBNgqcISrQKBric43aSR4FUgIDRfbuklI3Qb5vT7id2NPqCdNzpha4
Rd5IjP+LfnP2crocrFWLEqHL1mkpBmU4OvoO0ZwsAhaYWdgkD0fjlXI0gE8FdI7ZJlYos88K0BG7
kabUvE7ysCZdelkf2s4bzYjKIsr89grHO2OyCAF4TvvsOtdxd4ixGOzbYOWxTW4KLnN9ZXRRp/sx
oFN+N9CYeUKroMnWVvWcHlMwJfEz7+TnsYvyK/ujR1c/VqsYf5UuUH/e6JkC1oe2kRI3BVVYrRPH
0RK8VQlPmgOqFkb9kgFaveCFGHqH/PQNgK7MvDzO6Z/6qmaBOuugtOdegCcNDpQ5J6JvXf8bEPlB
C1z7XMMDWL1VVWWE7wP6sS8qoNoHSozRhgNe9Fq+4C7i5FZwLvaK1xzEu1LNZ1ZrcXIVGKdWfHYp
YUt7Q3J56D/hhS55mcSmsD7Z/uR0OGgOTdlKS2P+b5zP+db3EtoNngJAlSai+aRrml36A1uxaYxN
WxWR2TqFWp/k2oSZP2PasrTXTE26VF7CxuO6ThdsgkKn8smV7uwxYoEdtywxSEcgG5bclZpkdp39
I1cBTHHGynLo/DhntyZ92tK+in1IuZomYsspcR5cxK1TUbMGcXGsFsMvSrjRXHSkpuQjyplSNPQO
+l7tQ1vxS0+cSsWB1mmcJ9SP2m8CXRaFhbvcXwpQxBihH1BM1jCoyGhmVZJ21KI6gwrhQdc0gXto
JY8KfLqAs89+eaoZjs4SGsYKkgDORQC1GPI2hCqgj8mhDm5pQ2LR06FRblZ0Emj0cNj6IC84WOq8
+gh2x0rQ+dEVIfVHN2LMPFEX9KFgbQoT9O5S5Rf0CqbVDbF6Xm2vrVZruFFPQk1qOxx9L2fNOA+L
eFbKASy1QBB6d5iQxxAUHJvVHFwOmjuGCzoFfLMJJL5sWYsEtuuRMwErgUUk8LYMWDY/VWSI6u2V
AWUUOs1JStEpyMZlOtgi7QJMwc8L9X4kV0I7LfPTDAGQnrFh+0vjlJ6lWpwlh7moxH2kFx+aILPm
heeeAlTXcXCczPZrQHvhea0Qp6/zyFNO6JvGiNCUkK363nfc0+neowidLg2vaFO4nqsmxu9CfVHD
Hwh/fC/1cQ28jtgw3gz4/GQQPmpyFTu2dqqeBfb2NMOb8LPLyleIp9aSvwflO3BVP11ZJ2k71hfI
FjUSuiwq1K4+Rk66kUqmyeTML04x7aWLG6YLlvAC3E7yPsE8jrSRej2IPTIh62JLJ0DB+dy0y0p9
cm1vmReOny5HhMt5VWSiXDgJY9BQrNQHxfW420CMHOTipsboa2yWtAe+Vzlft2HEEaxAQRzsqU/p
05YmTdpnWu1wn+l1JUXNb1MJNl7dn05txDpLrFF5Psc00pYJfl2Ki60IfFrAbxCZEI7jolnZTQM/
oGKAQdA5V+kfDhuymyUgqasWYstbToGRzlTNiX+cqjDratI+wM4lvQoLjzKFUcBR/Mu2rxYAMKcx
IL3cpE2YtJfeAIZ2bDO6Ja8WAh4sPdmWqSSdAVPL2pkkfXL1qfSClCjL4vBgzNG7/Yb15hsaFcHE
z0xHk56W8XBK7agvwhThU8GXVfYG81Z0tLylewYJUqZT/7Ue2iRfQRied1iMS4nDgBIU6bEUNVxb
AKlxCEmk8X84/ZoB6VhBfMeEorRIRVrqZ6c+rQJtNsSPY77DcAbefu3bmLhO+WpUQaiTTkdaMegu
5eDdoq6DC3cPxH3zViW6BL1guHzweE1BpfavQk9p7mi3JLrZYjMkb0uUPqEfeHck4AWId+ANAJIi
zGzgQF4UPeuHHvx55fkzN6JnT82g3csUI67f2p3VzLFvQpsxNP25kRxD+ci+80TE2z2gCLERv1hs
T6RIDA7efMCRqdMy7DQHppayMEiEqPpYqstgnrE3nMYcJP3VUeMOV6aAPCzgQDUBkDyU2CTpKo0P
euep8PEUb+8xDhntNhg8U/o2RjG5bX4LE+EvecZyTyzqz4TXsqpnxdoNDLexoGFBTgCs9zY3mg/e
9ZsU46zEsBhzqylTEuMx5+JbXXlKft/cS0diQAzFO6XnYquOQIbYfEGyIp3/HDfjMzl9H18i2KeE
RTFEzOVfbSDy1prvxs39ifAZzuevL0NyoB9JT455SdjGxBR3YtQlJj3Vt1db/ykTyw8bUk/ilZbs
Hr0NIeemL28AN3DtpxrwmvZG245ygftI3ZxDtqY/5NB3Nk/Vy7E5Klx3LLlXbhx5EkFKZ+3h/fLY
ilX9zKc4VCktwUqaqmzlIu8tXO32BfrTtIarxTbl/1dyFBrF583DSZKBnLZHLGXV27BP7OjI0yBh
jdr6yqwzWOIWZ8qhF7zyk3PJ+qH3iWefSnyKPmBEuskuiED1T+pDREJCVLujTPfQJHJ0RL31oQtK
EGbmjtRxzv+k+hmIykIpQka2zuNzlxMXZ9g4+Lw5jg//qej1xHjPEi5NmVsdwHWlUcO67S85Ckde
DizQKxGn63W02LwrjxfDsF3s2UTM7yM9FlJKV5x0ist7vXAIxBPJ22RnGiQ1Gq3kwBfcZVttMvQG
zb3FSIOhdEhhR6vwW7GT9pOOBdZFZcdCzIeCoOb+kZIA/j3pLuY7rdvCtDDXkWCGaL7M5ZXPOvuY
5hkQUXIrSqX37PbB8l94iwrs+N60BGd1xmGzXIQN6/EXccTRMqGgoLye1YYu9f1MF1DnytGRHWa1
qXUfNLJzCJYpdbxabyLUICbpydtvTZRs6SR3AF3cSqCZ/WEOSGTAnSm2vVNMXfUxEl5k585mswsJ
q7XGVGdRSvsaW1qNuOAnuB/cbQ9LVXr3G+rJuPSgf79H6qVnBwvvTgQbCYJykqQaF25RJ8zh7P8K
IW1LSeh0ObqRXo3z52oNWWQR5i8sg/IlbB5Kp7gZ4bOClZD3wi7KF1gkxz4WKJIvEzWztrfd5vfy
XTkw6bqUVCnt8MNBpwWWmMuZX7tSTj0mWiwiltKUXdjcunkKRphBymdvsGawfSfLXxA+oziV4I+p
Ym8ZErz7ga00/oLG9iCZ+gZ++3hM1YIm6LeSgJAved1ao2w3kOCNoUFpAL/T61LoUcxBHsS1Lj3E
+LvB0gvvp7DvY1j0V/lVBf6e1q5bEAtiojlpwOPM3gxUqK6lpwakVDSGh/UWy6JUjXvvmonphOkR
bokeVTxpMS9qn/SBegxVVY1gRD9uxZ+iTrDguBkTexKkoNBtvMV4smHCfQPY9CwjQPlHcSBt2Dv+
Tr92Cdb0DLs20TNYjCJJdQ08XhQ2972LnwOctiGd9YAQNiGmLvZYvyv0f9MgdQg1ZzkH5JtX7jq1
y69CtV8nhVcfOrKLuh5EI+tnUXxTyaCH3qCTaTFTIHSMxvmitSsTrQIU1XSuQ3XfjRq/dmqjNszH
uLpTG8e+3kTg43+hjQk91dJHFJ7FFG2zZn+KgO0B/vabjxrGM57oRsMuTaiTdHkW/GR72dXXLVg6
4ZmjULNim2fWhPWVtShw4b/aBpLIZr447Z35W1trwxFX1EKJI5fqnroKfltWkR1AsQLqDHiT2+3j
xybFFtajuJ047tL30R5fIsXTveO6KZHieNmMoMNoJ/5+thrI+qbctAJ/oMRap4HRo5VBf3O1IXI+
em7q8rZMHHQrb83O9rXGoPf9CWI50MCSXlyJN2AnaCZ7+oKc6DH5NZky8+vq8ghsT4hypNB/3Lze
E8RlcOLTMEjziWzFE9gxlHNrfVqCcd10MJu+LtaEVw8pYjaVYexATT9D/XbI0GssKkFTfIs3OU4Q
C/+3mQnyFUj2spmSQowM0fnhOYfk28HuBcK9FAHKQL5HerZ5hbAnuwZMHtw5ka9qpHGG0tR9NlcV
ldDfwZOrXBC4vbK08bT7Z0H0kvWTbX53WO4sdz7LQPl0OqzT/lunspaZ6iSWwMqdQhYiJIchYtxv
zBmhFjuLUD64HBn4n/SktX/xZvEV+LfAdJgy5/P8oUBkBj9vgjXBfOVEuH4zvNovjteuGSo/4R9I
+yYAfmFmJsTNVIRPpOQLyRs4ZULl4PW0hzch9mhZPdFN8mXrErdhWfedtwwufCTs8bxMewH51lHn
4kL16TskXh5NWUjQ8rr90tmi8heSVVwkHpAkJjVSdsHczlAWI6MQPqyYUuK9uLICdVZhVisPxGwn
YmIj0TmBtCz1EDUVu7GpOX5QksVicUnKX/k9BlVu7jiK6qR+kEmRKG+qSKrZRRIdyMH4GJXSrXLJ
9GqMpWRstM0TnPaSxpbJrIFy2W0TqFfUjbeSZJ1M/lSTkFYpCu4St4e0lF9H6yoGfVHoGU3354b7
RiJiiZ2cvosYCys2+a4qbMFdgFSE2n7GMJSpNeXzZSWRQmvyHybrTqhGt10KQDMD+lzTdPeWMTNb
l9CTYhrwxasmxcZyys9naoeBrStwwx7fSK3nSHLDtSEus9vt6fSr4b0vaXHJYwTFC7Zs8b1/k0VO
DXdxpKKx6QPZKiaxYrklSVGwhpdmMl1ZoZt9lsHpJPaAis6UeCL4U2dJAnidT+JTf68+6p+Ya/Sk
mRX0H3Ns3H0Kl/3jXq3QWUPpr+lrfCy/btNm8VQikvVkbgCEKM0TkvjwWrE1jWxrF7iujESWXyfP
JvkqrE+g63s4zw0UhAyewm0WdOhIIA596CCHY4ARIjeDrZYJf5yd4MVKYhhfZgPgKSbbKKAOu5D0
EFfnO2Y7x+szohBa60YVkLpRZcI+r0NrhUKE806ZWyB17A0dMmkvM96X9xUbipo2CPbdzRoBV62U
eOcYFhVkMY4Jy3wehFAGTOAH+pnpFEZRdUSPQ3x+bHDKeMIw7/GkfT6mBTa8A8SGSRr84Ddxy1YJ
0cWFrpM9feyGLnQYc1QQEkzCwY1QQJS1Dy2jd//F/1Xf/ZLY9F3EDrXGkLAOrPAZHaQx6ff9Hnaj
wdGjlY7wqvJvlstE0EfGAjK0VzWg/qfEOR4c49RxWnjnaQgWU68TD59tXBdMvAmcsi9RRvcAJAR0
1fqO/0IU8lixwvbWaMGoq/A45UiaWuP6hNkqGtDF6UV8YGexymzqxbIK8DjmEBhQUde/EP4zYWeM
9qcvL5Kcnx72nMwM7caJDD9XJAZP6JJxwEtzvaklkh3anGDLSYWGnvKCl3cXyNa9X4NvAS1uj58P
vj/ffQpcLZOBXhP2EicElAT5Suhn0bGB22j1xcmauU8RKrYRfrd0GzdHs67D9+nvVsOwYLiWVMsO
I2mmTVrzN8V1nucqGlQ3u2NflOtsPwH2p3SibRYMF+Qhzt1DckmVqrAn7PKRxoIW0Y89S7j2V9hB
RuAGq6a07AHRgTMtCGTy3y3eZ9tIFfiHmhyvOlS69nENn++thO9rx661v2bTJsTck/DOAgrW1I3K
oXxbdspKYEdtImMRSWi5LAfyPSUJ+vu+KBcMsJFR0RpUyTCLjblly20zhV0C5XyMi9Cx8S0iM8uQ
hjDM4xAZtjmJWi4zUKu69rUHTTh54sAVjedBhOaAllYPgL27Pij2QKaKOoShgk4R1bSMO1Zsnra+
bZx5Rq2RJBxxTAcQzGUTOcXYNhpMgABXHRjtbY9a2yxosiJvAHHpNCv0X6wHDkJXM0tz/zlWeG1v
IGmxQbdrwGfs2aXw3zMysknKumD2I7s73VYtCHEwGhDqLIhEWJhmee5TJRBsek2CCNFPFHRThtNQ
1+m3dxhWOqfG/N7AxoaXBo9GP1UEwS0cHTBe5irt+ttAZ+PnZSewFSUlRIWgq8HtSW9jT8Nxcvvk
JU8E4FZvJ1S1jFYxzZyLuUpR8xsEx4kZVZ10kDH4gZJ/Z+yNimIUnawH8H/xEzlgyFOMAgPI/17u
MN5t074BY4Iie1VB2eIjAcl6juE73bn+W9bJq554hgEWX+T1bfRn3eOgbiFuEBs5xJhUxzle2cZs
8uvVaoK+gbJH0QGTH5aXCwvL4KZAjtMqqZZ7ng0xMa7gnKV/XGYaSDIC70OI/JDN1REVqwMLc7gT
/dmRcjYKoDL9oVmJN32CT9tZ7AZKAtOqD7iBTFU2Jxzjod3pBJAb4TynQFvHwIkTj8Fzvn+/NwsI
yBfjwXJrYOe+XTSOvKP6jmoqGV7EYCLp9D4thHph4Cv3d9LsUJtbVvG+tLkFr4XyAJsZ9IS1JUEv
XQNjMvnzIrgI0I2AL3dAGaj32YImtSLMm0z75AmHWFk1Tl3SDwQgC2045Rau4I/ruhQH7zje+wnE
i/mt9G9aFkzNe87El692PDL9R2+DteOvFFokDp5VsMeCeTYTFi9j+86YFssNUuVlnvEbC6fyWsXV
BcVQ7C+l1HfmO7TsIUn83RJZR4tUvf/hzLFer6KrEUuxCCfvohV9MTRCuFm8xbynlSoXI5Awwuqr
AxemS7iioddKGwnOR3mR5VuZt0Lh/5TjiaJ1/hKWHuZZnltuoGKkmXa0Oktrb37djJrrw6rJhG4I
w+raqpV7xARhsddW3XdrOztodwmONPDlJfPUvIarBMMv9B0fRi0gQkrO3Qn39NtIILztJZ5JJn3r
cZREmyMrpcVtDDJiO9+4+T9lExzvQFAMnAZtll7pcjVWRX7HNCTCn9lSilUxX3BEVdCSqodLdvjw
JYCiqYsFtMPx/xe4cJxPGILd00Nf6uGYWxZBzl669kOKaf0Qn0Q5/1yAEj4/kwVNEvDqETK5LVAv
E9zPgG1bWpHdOgkzy7ANRKIG2og4u6D437Ka1vFpSpXo4+FU9xmO1CdfGAGaEC3UPDWTAFThAIix
gcHUDe8WiDY0IALHkcBIaPBdh2qzqTnTu9Be24cCcFnRcItIQ0UFR57CSJ7TfJXUTtBgM7RgWTaY
8frdQyeuBj/2Mv0bLI3BXsYLiR1eQ5Nbz3MzExHXtjG5gL1+cG+CyJlhyprgWTwtj4Ixwgw4rGgw
8EJ/vN3d4agm57NpVRQHhnIte4/4hREuq1LkQO+lq7l91pj7F5kSmEAU3QFY5OQYpD1xgEQE9Y/6
RDWWOCnAbcDkVcxhnTKXzaE1/IYlsao55HoW8K3Dk6qm1GqqDjQ2QzHyC/qDQFxLqyEluHrZeiva
7nmpx2+ECFq/ykNeNzQggqXGxseOImOyluKF+OnhdRe3ZS6y9BjkdHW3qXQXX1Trz5Oe1GEADto6
Fb4Qi+rPukO4MDSBBpt5E+g+Y9icCHHQQkjVAvXa+QKXLSxh+zj62tWAGWCh1UbH1bATpgEJ+asA
Nioh39iSeUbbM/fwDWr/tP8luM2eRtvJErCaHSaTwGLn9P/tg1xmc5DeE+AVdIXy5gOOp5GTQTn2
86lmAUOM4PJubhqfYncxgzlhsKmRAfftRq0JheY05F/ysg3ty1MlPGDCJf8HgXLKljSXuiSE6DCR
/D8ezF5WXI0fwV1ODr9APyzwytgnRn1tI/UhYV2fAzGL0syZsU4OLLxXQ3J+AF2w2PWWEVIF1pSd
q4//tXuqTNpyqNNu0TTxX4+RWwhhmGtQpddDIlrXN/b+RMHuu3rtm4dnldVdJeMjX8I8Z9iSXzfO
PcNS7dVdyYtVPdOSDAH84tpIVCM3hwDbLisgWFSakRBK08stY8e32QvZHbLuOor7F1fdOkl/spDR
ygTBSBeggZBP82OPXIEuMKRSCHvRQyPvBkMLyOMg6nqYsfJuFhFbZSsjiv1VyWzpSfCCW5z3xSG/
h9XacZcjDjrb5SXz9ZwomC7Zl1PL3xxvAlFL9lfPV/zSXB9FWOeZpmKUWfDwteJnuRrjWshV70Ca
7SUxU6xsGO73xTu59iZlLo0uM4IkKWwKXbMFHcvjns6bOzXvVKA+KhvqnjkVloeHcIR07Ildvxro
730pVaGdkQnrWnx712OQmZWNltbQVn89Vw9MBWFtHLmmjnggP2IMg17Kqv8meV+P+S3A39qwuTfd
zo1jMuwY3S/wg7Rzv0J2Fyw+TQyP6MMPVHTqrLCIgNUhVP1YD5z15FFyRH8Kj6n8wGv6qarUeboC
Tuj3bWabA+dYjiB6kzy7LVyPW3RSs6gtqcriSGbxYiC1hAcBwluMSI9z5pj5DUOYZW18zTn/fvDI
mEfbZAdR06HUNfix01gpZ0GVncUOdCOo28mROY+P+P2t0qntKdtFYXwyapHzFEdH1GsVNSIi824o
l2uPtRNhUmLPfLLhz2zCZDjoan9qCssPkY93J3JPXv6qsx1YrWfIYSoSocFVDjZpDjC4gfs7udNh
E7L2RhFBeMKkM2QQbM6V8mnsceCc+MgTFoUketrDtCv5xUNYyuoTjzq0ahOG0hX9GvAaPHtUW0xa
tE7lj1RqvIeRBCm8ijCPgMX6P0tNQw4zrkJpDZY2y2Ek/XAdB625dwykWzkVwSoI4HTp+xbp+yXc
+G+kLnarjVLn6acUS34agfHoaj9ZcBsP5xpviHHQM4vtzsrqty9BvN/Hl64Tum6ua4PRCaWNWs/R
PeT61MjFf6O3a6XXMlsTyZFmzctnoBJ3zT0yD7HFaI6ANDn1n37WFpHZngIgpcmibsUt9ZCdIfar
BE2G8jZtJ4tzV9UkHuKYA7QYMytddROCLJAMcFSol1khstJJj1KgM6mj0pA8CXrNK5ADgOgi5Us7
mwtr57zImNyRK/S9PgpPyDe3cQ0lPNyKOkdF8bN6D280MPtRxc2+BaPyk/K9L3yhyWjfwi2ahQ4y
HcuVM8dv9+uPpiKY9pmUwECkBnwZBdNsPcGhoAZMwQg2FH4mnO/go0liervv+wh4MuVco6kqdGsB
5Jd55NskHvA/0ZFtLnaD+9wAs/9ZtlLbn47DCmz1tLueUo9PHlwq+cX3qmoiLQ7Jp8ltZA2LMPd0
3AQVda+swF7FXSxxgZ48TgqX8WsfibW5LnvouAAT5TFceB0fTwOph1mkCUrrW0GfZdgBSgwSwLyZ
14nKihmXLyb6B7bYQO0NLC4j77gzLWX8eurU6Ly1qhC8GPRXYmxLBeu7t4lSzN6wE8E9XtjwEjcq
8MtDbyv4ppfpiYO8HGoVVYhu2tjqWhE55wf2dMY4WAlHeIYuGlLSDv92HIdazv+CD6efc1fsIc12
4/vFC816QehfiQ4xMhLeDKNzONyY96SVEwAWexFtWepufwup0tPHOwKgDW9oe/FYpv9GVdDRgadv
4bVeIK1Umfkf/wWsDgveshZ/9H436x8XjVEVIufWguF16T0P245LHor5w/Oz7/GreOMjmi/5g77C
hhbH36cIeDaUG9Pb/ahs2vUYsBj6S/lvxLFUm0/OeG1xk0xocGP0LP8RwoMRdBZ9OFMDX35cftTg
PKcpRVyrpo0peCrrpJYESDVoQ5u/QMtN0lzrYiduoJ5BPC1884ooCnWGCY39sDEJwKMSIeIF9hWM
TdQLNvXYFUulK4JKmwGScBvbuRBbr5aEzgof7dOqUXBs6WXTKN/EfZkjxDy58Dvrxf4C2+h6cWv9
9jm2m1goQ/v5zlZf2KWnqWTgSh5Px5sRBgjDWiBkW7rwJFppwrh6rVvBGWfbpyr/YQkOXxMeCfCF
jpmylpz5UbQQiDX4ugN9gyEPLaGV/19tK0Jmne7graZyiNqjq6c8e5yIZpTJAoMj2I/NOeuZlg3+
lk8tH2Na7sf7WLoFOh1aohJOoC2COa5VQ6d+Kbc9QGLOtYVlPYyqJPGfz7TI0/QjZjx3GS2937e2
2potxlGY7ACKfIXz1R+8tuPox/itH07z7auGcO94znERzWhRlqDQb8G1tMpDLc4WtqgPpUTzO2Tt
gxttxdwYG3tSEKds7RplxsVyKnp4jssGT20aesPlqTiBmOknkue/Lwp9BY3ZyoPM6+G0S/YJuf1W
iKvZJwYKbfDwtXi5N6YP/d/TBjvNkgKTiZuQFnzbQwy7B3ex1Di9ok1WWAZblu73bAeEu66uWz+i
RX8DOEfUk9f17PRrsaLaeu+SiQX9KjU+7tjDG6uPHux3QBtwoNOQek7rNwemt3u0tzKMw/2tp7uh
2nd0NE57TmzTQDqoEN0wq7QRu2u6puGTr/HqNVykzwuW+1pSlOHkdaBiAcwTPy2vcRGVGywwXVZs
VBJQ/IC2CI+WgGettLPbbnb9Ki7BRxnnDCABc1+IlxQlEmyhoZgN9j/rEfX6tXBUGTpbvzLUMnDZ
QmRGiuFSFSClSeDYd1Cx86bAvcULn/mozhi+jvMgkeoRw0FT9GoDNGDJw61/2A8v1KzRE2Fma13k
OE+NK2RVo8e+Mtz7Y7vSS+HoagYnW4uIuu3Q5db50wc2WD72MX+bZf9+63PIvWGxdFOejJ5Ukhnb
T0Hp0FawE5lfMPauaOjDiUaqATxsZx9OTsz9Bn/iq6nfxm3yiACZGRMejSOefTZd1DLFtuBizHrh
S+ZIkC8u0vjfTKxmCeX5HvHSNuWQsWhy+oPJrF8ZTKCKhcBPa8Ckc7fIYvDsJ14pPVzQ/7DgYkF8
U8HGOIgecwrtf5WcXmmdzmxlBAxJtPnDOnAhVphgm7f7OVVXvAZ8bebptLmtB4UhH0HiOqAkw1KN
9KNwZgKJF2gvlzXzmMTl2lCqxZWCgqsjTqjgbRKGwfR/n97jZwwRfVT25User6HeDam6KbR4osoI
iDC+C4Ay7PfKjRE0CQB0bd2n2SeJyrHYwFUWwBtQHs0UWgjqZM2kp68fOWXctxPeJqGOKhdwC43F
iV+SGFM8jJCGWGVzmCwUM0WPIFkw5L9zoq2f68cIYPg056bvhEs1V+Ftjtp+RZj9eQL1UKIcTOw5
Qy4665KJ1htu/MwKpd451jjc9vyTGisLETPZnWaRCuD1Gjvb9fFdhrZFMKDugkSOu0BXqQLAxPPW
eveltEDMEV4fK9slnzNJ/aQQfz4F+ifsvME/QjiXqFHhigYwYMO0w+eZrJMfYO0e+uNGHLDuluXo
HLARLnTvtEK0TJvFRtuwsiHMTiyQ8k/RPMennuSP1TSnSXv0cMRdvXEcibutcINGk1M7pf806aEp
5edyHoX516ozv6vd8jTBKGI7pRYV1q94gizZY8K/inqMiOucAZgA3lQyFEwg31AGHpuoYGFe5CLQ
NrCbldPHiihcKm/NVcoy0q5dihFL2fa7eo42n7LKBCYVw8IYrYtykOHCiFkf9NsVwFC3qeRhnaCd
THOvavDd9EFIcGyy5DNEhVRghyLmXPT0yNl52cO72tPLjHssB31nmx9xRSh9p5cVCb/1+f4WptuM
Dmn413XrNTmVb9pYyx+93++Y+AYasWbhPuIX7SJwREyuaJJAKL5Fe3vw998EqHF6BrelxCSjEQ+A
WaqkBiN0RufF/pZc6JA832bU8aEJHdKr8dD2LHa7qAVNWF5kLuYJZ/o6ge1W+y9wLEUDWRQtSacy
TRLlNB36D/4g527i1asZW1IecIL0Wv/3POmG/4sNgDtUMcnmZYPdVPsN4jacxeHFjPE/F6JfF6LZ
gBV8AUB/eJukWuJRw4+ClN+ELZsMBAeRJt2S4P5BmngLufsSUrIjlg5wdzlUtQ0T6BHTRVX9qkGa
pRxGOhDalAM4RhrR0HbNwaCyBJ6IpHTzoDUWsUZMmERKZGcIQM3oosjjgA21M2dKFfhNdQoFq0pJ
X2NGJRkcIYpUT76pITFOZmd3bgS8oGn9PVoJS0nRLm2NgPZidHwn7sm1DsBiRbJrrrK/3eWySSvU
Kws4LAUOt8lxdRqztgmuILDwmc8oItOUXWF9bl/YxvuJTFNdkUY69ebF9UK7k/A9JSBtl3zULqKI
swkpOI9mY3ByYVD9DsD0RLaTPaHk3wR1fkmariKbcLhznXeHApxX8xn+PJG4FWi+3dFjdBV/LdHa
5Q4KGKk8sJtTCvSC+qmH5NSpIEuYIuTjN03hDAr+mJDyy5pPvaYSFbIK02t1XmoxuXP1cO/+tLqo
dC4l/ZGtyTlQROfCWYkbDik64hRaWwK2VV7ndVrNR55WMXhE7JuWTRKfEXHx6MFd8+wJDRqKXrpV
iVIL8Qc+rOyOGamtlXIa1U6Y6tJAOcv5JzcXHEQMomn4OzuCEuHJGsg52GIOCWomvcPmQk8A5YYw
I/u0ICM93NV4UCLZRY9bJpwzskc+n5TXRpa3Dt+khKreTbivwlVMUwhyzvoeU4aw7fKuT+72zjGm
Om/MHl1O/xULyefCXgTRaJcr9ZGxCVbhMrez+ScAMjRjeJEKkysjB8NKE6MkwQddX5Udeus/QxhU
iwImudyz+XrmoFe7ud9Hq5dMhM/wglWWy1ncoUTJUkgQLQJPTyFZeS20v8zeQrG6+OJTkyHC4quL
u/KzaxctRaDbS5U6KFxDciONTRoFVqLe4ZMbNAl7o9gHcrxQ8aS3LEYIYpGzjsMUQuuwOvmGDdMI
3aboUMnVAJu9Mtr33rNuBFUGRlvtkmPTsHyDZezR5ZZyXSEOfBRKr0FloNqdAV2cwqaNRc1GdB9w
GHgVIEnG1GWz7C2h9dr9l+GA6UHQhmYsfY6UlE1pI4mWgisLIAIQ2kDYfj1sq3s06l3KQff1FvbS
h2naepz2RwRsLngbF95eIhlbUQFMI4VeDuAOIzxaDcFylwf+eebtRYmGajZUFe9rqlG/46GNVNXe
2PCKhU5SqBXfX84gVVzZLq8BIBRmr7+KYF3lIFtBa19GJ2ZvHescYwnfabeC39CsmA8HfBOJdl9z
5eSkk1ZUymSRN6w/noJf2SYdNjZNAoYomTp+8ycPoct7wiRpvx+cy4Z17QK9nQUbdd9LKIckPUv6
sTl9gL59AJgm0KF/QRezRHubl02Ut1KaXXod6kaizpi+2T6brS+ODywbnzNC8qPCNAOvp+uJW15q
1mt9/j2HnPZTtXVl5fSDlU4y/fjjCPhjeZRWs4Tg0cLCyjJr0lWTNLMRbHNUv7ZtXYd60jOdqiFl
AXHyxpxb2BRzHZ+3BUpwvFUzVoC9uYOATlyr0aDGEuE5bDQ+vTeoRjvg809u1nJM6K2XiCbk4SC/
FO69hMcBx2VcxYeaUMJEJFoTRvFfMOvSKF6oWQZNPuUL5h20xcxgR+TUWBtVabE1Vns2CGIDjMVc
7230TeZOmwCOr4RFYIxcx+9HcUVkdRbECH3bmVcWZtVnzLnWJyvVtjHPNXabyg4rRrZ/cf8J1Nee
hwFXEv7Z2pDX2LuOhq9T4jWyPgujZroH99SzLLyJuaVGYgf3RboYDLwv1OiAAsyQN84dwVXqrRmG
IGRMgBwWXX5THjix2jSD36XUstzL3CeBrfTbTF3rJ6p6CyKWuNWm4cztXJ81zwEBt+sDGet+9ZLq
GQEVG+5EEgwS0f/v4RLDZonqGFvGpF+1aHAp3yGomvQiWfb97pepcpwdxWqR3K5oufgE1ezzKx+w
gDZS7qtIkSYPmZrsae131cHjV1ke+c5LXKKiSuQMsIzfs5lXJbyJCmltaQZq/ERHbrtRS8thuQPk
ivWM4sl5HbZg386by5Xt/mWKUn0jYd5G1yK/50QA77cQTtmnhHXCthjU2gatQvLchcPCa+wJEhA5
agfNqyzoKTdgKksnzdUW02G+FrN+ndS2OAg4nlV9EBSP3PSfry5WS+MsNblrKNtWAne1cP4Vpyrk
RvomnyDFabopnbX4kQ2GJtxvD/yYKk7gIJ3Ppv2SeXq1NGoqbiqUmRbYDa0gcCIGmBmCqDTmoXLj
F9hOdC+STsedIdPZ5Uduh/HWyQJceDSgiYY3ACLJie/fy0RKORBgodvNDNNJEje+aXMZU7IXsgYX
kph9FLbYg9ih0RXfsJo1gvCzn+Zi4xjp6ZKr7waLQdeJuYUehEtYkAESX8RCufixB0k355F3Y9SB
KzUFrVvapoPF/T7XPJkYyOKf/1qHqtFouU+9NeF7Leequ8MtQi6GTLttOWuHsSJgd8PvvbjhKyJB
gvp4jimcB4Y//CAWRqvgf4de7tx3jvWHvKuuE4Z8X13s+a0JX1BgoalysRb8X8sS9OVhDK09N7TX
5akT0s9adZnE/EMihKkeaGg3OUdDmp0zJ9UMRmaPeTW/hWdgwLN8dPFrG7EZK6t33MfEdCjaVW9B
5Y3i0UkNKgfpU85xgREQzzPcYIqxpCB293DIcSZJVoHg/DJB+sFW+teJqZoMSidrnSbCyia1BxjA
6l1t1cegqOSNP8H3zI/sstufHBOPAjiJqTPEK4frzlfvl6TqW4XaHmuDSZNGrJtitUoZFWvgpJLF
iLKRozT2S1DC4OlLx4p+RoflRK6frdj7EtkyhkPs/vXOxIa2/7sdGSagaOMsCYmCBIVIir9ZtuOj
qhD/MeknUVn1CDJGff7LFbcGbmYNaSnk56wCSBSNmJi5wgc3YppDGvGQRRleDw5rBz6VPWh8Xa2w
GndLyU1D1z7fyJCVngUGFo7RgCDy6lPVe5bFHoS/uHOw+ueGlOoIszOnPIp5LX+dmJUqqcoHbCew
/yyqbQOn96HsVKLsbc5H/ARdJv/hOhKSrcIpiScMwkB8cVzfw6VkfWShvlIv9QvAVwWEBCtkeFi+
APRdoYL4VMDtMZogbKbhHsGeAeNZodE5hNMJ6dATNBVYNV6bh53MSrBwVaIS+TXKZIriZ9ovLjHY
fQjcIObtrJMowYzCUNV3Qu06OkXYXlc5WRHr3LPFucHWu5EMp+iq6zQzQOGtBhzd4aMO4eD88S+1
EbWQB6mfQQhz0vDSfx7sRnnTlJD7lInO+NgoEx8HLi9seN4UuDtoRB2c95Guk45tEc1nPiycYj7C
enHgjUWFOQrNl/MSPUaZHia8kSoGH/ZBW2bRuEC/oKwtZBRxf3wW5P8CfA5qa1wJ35mDyyzbhmfJ
oPpn/XZ2XwcGwROYNeyXIVF5JpZJDu62F8QmGDSjqDIuWGr8cF4+qmHSNmICCz6zgAgGobauuyJc
enQznmFtYISXzQTYL116E6zCIZnl7MpGUcneognBuA6CoxDOuTHA+Eg/dHCPLejtldyrKNQAQtVN
/kvbEec8mReLuGsFKwWKJa0/pWKQzEd3ktzjDgsgXo6UlU7PYnvKxgjmiVKqMgkHo5zcvx9kS3Rn
RzyCCd8fRX0EX0IO7J5mjWlw4l/G7QT1xq03lF6yNPq7S5mJrfxYZziLNUlTQlviTP0vEcRZ5Umu
iT6V34uUdYKmuqvet7fl+7PCqUyoelAjGEPM8W6bT+QlenJyIW2VMrYzwHT3pYgcD4+ARk9d5lg8
d3oTHRyMaJxlleIFm/pxz9Aqk5Lv+GzBYXd+sKsfelu1cnBfbOsv5M/+wXXXIfZyTl12G9RCbtS3
L6+VbF/8M1bXb3Z04KddfBONIuqlMs8KqaXpLdQ/Fv6p/XTt3sDyi+Hw/klSApzRhlPTiQu0ae6j
Xg2oE4LGVB11r3+20euRgz9GQ09fB66jXbBdHgJWmdKBg1KDRsozOlEnL7kPBIV1fx7fHyOIFlVu
Sq+0VTZfNKSPY8rEW6zwhwHmt3Hj5IsJ5Nu2xDUyj8B8bSQx6ZLHILEOH4VODxUeWk2wLJwkxsEp
1EN3or5UAQKNi6GbuteMa0AluegHqrQW09Ttsz+pIpl18rBi/CcD0WEDKKRGpeYnzYaXQVJ2T7Wd
HEoCjwHWDHpiPCPUSOAXzFN6JSh0012ilsejXD8LYnlawndChL11hk2zeVbvY8DrZfVUCcklmt8V
ef2EbggUurTO/T7Nq15UHWdsQDERNaPpdeRwoSBjkWgvF2CPgaTxp8ck8UaQPC4d4OJVP+bcLQ8o
VdLM98xCOlKVN8ZcjUXQOA0/d/ptIDITQ1Wp5ntCGkLhL5mqH8ZdTHTStSC/K2VrS4jX6w+q/KRq
U4CozQJdv7hy8bcrdLm2KSH0sc1vD7m73bLd1NKS28xEQfdzQ0dwA98HjDiN30NNhm7foI9Ihr0c
3OJHhRtH0Ce3gcGgbyWD0pobKZek5J0d+spu50Ey5DaQNSJaYp4mFxEuwiDtwad7fM/ssmmloDjl
X6kZF3FrjbtiRR84K4Adj4Hz1DofDNQonvEUlJQ+CUPk3BuvaCult8mZHlL1Q8/VI+wMTUSbkXUC
LViUoRXoMDGfR0KgAd137OxzpgH6cSYjwZqA8UvpZIvitXbcOhRRmeZCU4jkGsDZbZ96IPIY9Da/
6QWGlbY9hUVK+EQM4PK/1mlZPKVU3Usf+SzibLiD6DceWvL5dqhvPEzWKcQw/F2SHvJEDwUg6yVB
PwFnXIiEyZhvNOwsEv61kkgKotPtGqUmhs5PrFEfifFI9UW8rxfEPZtlZvouya2+neDbUSQcKdOF
tFJQAOTFj6PSf1mNmmLXUqATGqGz5+asAdm3Sygep304vN3JardKVWm0cGtEjdcXmnhdK6vQ+9ps
P9ibZRPL1Mw7A2bPyVnKQPahtmeRELabmj4AR5NBwFuhS8R6HbZ1AES54SiohThhG3KG6whWXYNE
7cSv2BrChieOLI6H10RdkiKxAJ6D5v56Pd7MveCm4j321lKFmWt/pmNuMbdRqjXN9RjO15VX+Rtb
cjy4p1b4qGnm+WNDZfe2+5RmWWS82uhK4g/EqpmnQhBoGCC59xdfbWryctn4qnDnH4oT2hylAB44
rIfKbk+Ihh5T/sN57BmLrZSyUj90GzLJtNGDYd62W0P5rtJLCfJ+WeaduyJw5q6URg9ytiwXnGbs
FcwVuSYdOixp2hNg/AlH9UnGMZh28Hd4w7V/BH/ZQjpYkJNfSKzEddqkBvR63evRxwCtFaFvJ/R9
T/H5Wir9Bf33vThAtX/BFnYf66yQB9NswAq+M2OYopCx9qQNieZwlThZZpyFQVy3a+/Cb6J5Yec7
hvrdp6V7kCBwXc+nxmJT3jOorsXkHKhzfX8bSRWxSUYsl4/dAD1EMpzvdvRKBPIHAPafW0u/dX7L
dvMwzd/+4VCGB0yIpY+NFaYKtexLt9ZFp1KUx9y/uode3mr+xqjZVIshDSQvC5rEjJEvygHOUa8D
u3Ys0Biq36DsKV5KDWWI1sR2I4wAVRd+GZdsytlpw12SsIt4olWbY0Gtg7OwdBQJA5iDg5W8QzBE
A7GuoLPDkzHP8ZJbOALApnkO9O5PCkZ0cN7RBJPE6QBVvlI+TGJXKLCdprxnbsoJEH77Q4QNBVxt
viyyMK3dCMI7pEUJ7Vn4pk9tSnzBhjPhpTx3baP9iLnvAk5RPnujEmfPce4XnmL+CkSLGtYX8ffG
Ad3CtEoS+vf3yCHXQBv+Rxv2gkx8GjeaRphiuciTXYSxReYMQHsbHGQNmWn3drzFS9oPybcqrr/k
6t8rZWYRkeAKBpx+nrXphT+/Tv7LNbFOEEsIYOwQ7uFmzP6Zcoa7qbZ9RPR3K4aDHKuuQ0qjYKvC
AUbfIjxGYHGcgo1Zvr+hIASHwP3nC6Kwnkz6VKbIzWiUUMctYDMKRNE4lPkBcQ279qlg7jszbvWP
2euUgu82Rn38oA7CozW4Z4i3vzBE1+cX9b6/wPfT/f664Z9dsUFvHTxoxxl4y66/waT9Imoq9HRw
qSEjR6PSfH706w0Themk+SGfJksASxicgAIQc/cE6zIbCX8VJ0T1ilrjNCDYE2+E6dwiGQlKHcWn
loXCZ9mc/itW4MxM5pPm1XK08ATk1C9m4FqQvDyeC0x8X0jF4JDfdGfZ4eroq6rjTpchh16DM6uU
JTxihKpX6tNKoMOPbAVxW/AmrsE7mJL3+xYNO0vJHTLmRPdzdtGBvImFdE9iROXq97QOoYiDTCju
C57l3yww0uBf4VdjiCMAv9rLbSkmPBCuvZBODQboU2IZa3Wk0wjv/I4ffmewm9OMB2NXZCbXZPJD
Xm7FFxHbJTF97+dPXaDdaRnGxjF/jc+AjrwTVh5HkHvMirEnXIlzwLcJNyj/0ivc3U2jVGLKi/H5
VrupqIdqAp/K4CFRFyMnveT2xhjskFVKg/bb7RYthwZcfpVKb5pG8rjSeHNMoSjHNc7LLcS7qIzX
DEeMJ57afvqLCLIDy1NB8rxNR0W36wlYbN+VpvsLp+gGZikMZHU7FSG1rTF4QyOQi7qezppW6jww
+1mb1rtOZCf19iX0fCC8L5ALvA7FNXW8WALknwlYCpDb6djxtEvgzLF9kmaN7PBufF7FTwFz1V/M
pAu0v5v7eMOJbTJCFdtEuCWHUUn/LV378ajy+rFvbM79h7dJtJQEEfaDsFlATUgY0tG1Dus2AfJ7
qFVQindiIG7yWKCTQeSZ698c1yU49T4gU5/qjB+7FRlRqePTxhC8shbc9X0zq4XRnWjpLqn49mQh
rH3I+cpF1EZdVsq43x/sRljWGoyzeIBo3CwDmOXEJlYtwSvxtkcY7UCgMOwdLYdvnISFrtU+f0zr
CqBVJKalI1XnTRQxwYyQbsAfPggkR8kmLqB3ZYvnsY8HSotR/ftLM+ycuPaBzRdkxXhBMHT7zETI
yEB5MsqMvxcpYMnLlXfvyZEYlYlRCcitVhJOrqug1rSj5uYGfz1WBSFsGhM+u+HTS7Z3eqETzJ8T
E8zW6mUiOCrQWU3Rh6i+JB4woqKndVBX3kcB9weYs6N0mXJ8MgnReNHoFiwnXNBVsxvwgBA36lGy
c8v+V9vIJWDdXljeyf5tDY5qJn2mSGtGt3Kxr91zPpr7bshzKWgyBdguY5W929grID/kqdPARnkY
PR4tlC1AtdOAM2u39nil9IZ5pGzVenvlESfEi8nbfmqhDfH9x32/IWVHL9FEKTD7PCVB9bPdcchA
R8cjtIiyoYW4gb3siobkTgKvu+gHBnAXdqxnn/JLX6zcEe+B5bT4GjN2CLMrVJ734pKVefRu0ap1
+o7+hpuzk8IORHwGMWesko1zDJzY0nX/Tf4fCrSLevmNqmM5dZesGkHI5IOcdNy+W1ECdZjBlVw3
LDN9iXozEXQvM9RjSXqDYAywUemlIvMc03f8ElytzqxWCZYyjevwzybtvqoQtYB/DpNqiJSjBBor
QjpjH6mqV7v06//DfuoLnYZQkvuZqsMV3uFQv/o+/I891bYncxN4ccpe6aQmALrNlibMd+dlC55w
onBDpZ9UQAKmlvZ3gy9RKZDD2/xXTc0aNG2eumiOwche5jojk9g8fzTMKg4bUhi2o3ih2xplxwr5
Y5arAUdyhhPT1FOZrx5w7lY/8ABkuevM660/OG8MSGqCeQAW1/o+elRyoPsVveys55oJ+7bfirOY
Z/apLkKpR4m4assbEl43MiFVkQQOgd8g9vQkqdY0fdK2sX0+xApPjrIUiDqjTddCCv+mZFp81GSN
iGauBD5tcqI4Whi7/3r1bS6xW5LfkzHB/KH3UDqHWIlgeFX5gB30Pd1NgOkMbCHHRZ5Hoz8SYJM/
p5yN5s05H3MmGnKi91QYqQy/ndkL1clo7yK7KjBouQ3ZcdDPpN5b/x/x8X6ehGSVUTJ16Irv9WYO
PagHvJZxZ3mCQYB5azF1oxXxPhwEFXnB4GoHbgEp8wj4kf3P33oCyeEepIQMvjAXFR4AS2HE0kZz
3glgQa509wO8Ix3jy3uho5pdlyGUvXs/icyOZYC8qPyOb24hntw35+Q3CRYG+ADpxDQw8gHgxTJq
9vJ8W3AmJeG4SLJROZE14IZW+6kQC6+/xwaTxmBijdll/mI6p7ASAMTQGcnRZRAlICodeUXApRp2
sTpy546hGUtAAc4t1Y9Zj0NyzlVxf8GAKcdQaWDSPhuZKBRyDEf/SkphAY/S5ToPg/TEfZ8MEKth
0lkEQpjD3DgwMSFtwcto8L7vxfZRXYParz3js8Skpx9bLNzmizMeuCGdDQOPN8Ro9Rc3YUrewbDa
qu902HkU2tL7uwqw0k/oJSu29WIJIMkpLBYBVALFJWJk/1n1elpJudUbyDYgHJqkkLFhqOgs5dyX
r8CRDEfxHP3UVsqbI98QkuKoO1KeptFoVFbfE3DLVi9Rp5+lxl4Ysb6mhTcMHxu/JZy4O66MGEZT
rYVmfLWmkr4NoPkQTqSQOi6DVQEQAa7hX6rbeLz6TE+vNpMADBKgoSxG/lZQlAs+OAhNrvs+ts9A
N6uqSROfJB+0yYwBymVyCT4plEwasJ1LDgj/ulzZ1AsWRc1B6IQGXtUwxYrH7IgDSNIn4G390gCW
DfBTa5BHU/dHJ+TKs1k5V9dq+xnuu1eFnnOocATWISaTGX19SMP3amHs0Jw4SyP6n8SOz5lEACML
TS3VHE8GmOhPgmhu8hkwr8r4fmm+OS5zziosTq2IRSCGWCx0OuQVnlMtxuIbreBq17/A1H22WUCy
x2/kn+iSg8e7nW/t+XZ3mk1D1RU32YzxomF2x4U2xihJTSUSo/CbVzVdg8nnqWNnupBuI7adUPE4
e3lkajeX8i6LLAdu95OPm9LbeNY93ji/efKmwqsUtOYG7HUVKY/NPhVWHc4OO+TMUxw0vrzHMH6y
QQ12Hmkq6q9WskRSxTS06og/KGMZeLN1XxSaH0yQgcs5Epe9EY3K6/68EKN1gN61dEX4NDCobNMU
zQ2C4TqKVuVFviUua7rWrGxSBS5s2/6fxsaIKDmj/UvPMT4tppJ9y3bdJbcTAR2R+hFplzj4hWDA
77S+8AtOmI3SvRCqKep2pFODlvHACMYAIh7igkEzSfxzr2Yq7u/3psAgWXstsK6Pxfe1gAqHkD9u
8iH2fwS1EEumOc3nM4GvnA03iVXSxdyL1wzQTMTWLSO4zf5EzxXcOBuSA2WFIzEvNonlHFezOsAe
3OnBP2jq3UWklZ/cNIAYtKPvxkEElSv1u6KsB9x/wC9Ekvn83zG2f3ZeL3+du0EBwVI4r426OV2l
kpLdXPTsfoSyfbVPrcYuzND+w3OecMGrQySzjVkBaFeV2vXD9FqNLtQ3rRQRUq+zDSsi1ua2Ag7r
qqH4ZazuOHLtrMAfZ8N0DY7+6qQybKH54Q51qM/Eb1SR/EP11KZAoGm+Wg+EtYZ1AH2SeTcw7a5z
bXLuWReSkMnycug4Rk8WFlo0D8ZXlrQmn/5HzMb8VqaV6TX0Ij+98mzXhtuVWEaT3Oq23N6jqxDO
maQaeV2Uv55jjw4eSSD11lkijwwug6l7ELuIDaDViyJfry1U9BZNPTMewykYfIAf4MSpvLG+u/gu
6d65oP2Z9PgU5lXZVLEb1q1mIdz/Uzsb8HQyn0bVoK0/x9YeSeIcH5gn40yJiIJqaqQoHjez/oLw
7/ShP7brFjKj0rH0kxuDdB68q7dL6nI1gW9wswoqqCDY1Esba3nz3PfwT/njQOBIaDviijBN3M8L
dmZNuxD1HXJ5kJQOgtULuXPgeKCzCysaT1/OAPwK4QWjik9vPUosaTyjATu6pdMqhJzIb+fi3/Uv
qc9D4abkIO3NU/qs8Hc7dzrV8Za9+CNY0aVLIToYOlK1uqtQatNlOGzb1cjbnol1154BrVXGNMQp
h64XCVJQNF1DYYWLY3ydsYxPj4q2ZGtnwFbXCCs2Rf1MF4Lrz3np6I8ooLToTQkLKSldFMbZAk4a
nAZ5WBvZ7QfQW6GmYcpEQuitFOVUvuGI4OVqnQvL85nn9Z0U662l+Ib2iBgKKTVkycb8Pf0ftorM
31VHRKwsnXpy/QKDYdEx69t8yblYjpWRopJMJi/vUb9xGO+cKu8t810/IRGOwqJrHPOj/zsU+o/4
oQzIQsuBwOVe8/IRBykbXVqV8JGgIeH44VIqRu7VtenDOk+9LUgdABOAN06YnTvSSkBwuI3HXo0s
HSo4LkMBQC21SrwdglV2UR/yfUHqJH1qdPnXXFuilEm/XHQJg4e/PqEg5bp1rioGPBLKnd2VZhJP
l99uu7EZmDWZikObGwJtjJsMvnoyFdMUSWx9zRix9D80D0LAGzYru/jDfRRL19849yitWI7u+dkl
pbECSSLq9geWaiWZ4nZrq/3HHDsntHfQzjgm7l3f6ZSJNltwnurL2xDKKrALgMuVyPystBJB5JJC
Bn0jdMza6L8VU/XVKpPFFWuLIu1HPeD3YpgTXqw5YyWxPrCCiGH7h4trETH/rbuYG20UdBIJ5gSF
4G1Mt0dytlJd+YErlk4J2E7X8wloBi1bD7xq/T+ZOQyObnmbfiNUUXQ6v6j0NXaXGklcX646Uiaz
MsvhEmKf/Gz+fwQXgI/fmZB/ALGj2q0C2AAoTdoeqq8cls4ABRXqTvmVla4ee0hnwzNI2Ldhcijl
pBjmCbUTWMZNRAPB+AridglS7yurZwbr/Iw+A2iFMAzSCLbpYd7onnslpikP76+LnMVG+rWj4iaH
FOMIB4gU3Cw/ShNLZoQ6mIgFh6qjd3JmfVzHA9UI+/13kZbEqQ5mMAgbXI1Q/pD7FuE0RiIKJe5v
AKztnkeA1exDx4HKxtHLiBn8VIRxPkANsuX8+80Vu/59GjQ0k+L3inMDsDsbt6ynVNmfx8+1CBtA
odPggEVt+dtQUQ5OgeTyZRoZjOlMFR/pYMmr3BlOsbWd5YgMEK4xOKpTeo7lidQ9VC3mpimxSWjD
a+e3yFxyjkQ28RaNBSmDgWQxFm8obd+iSvAulrFnHgt4V2iRceBLWUYl4zOYvN8pG8DO3NaBtFyQ
DBNZ35q22OJD5DXxLjdVG79hiDEabKNArI1SxVvI+klVd9DP+C/pQNs1JEmSuwP4BLoXaoFmSDs9
EU4i7HGgj3UIhsUAhqES6rkytV2Q4f+tZ1Ug5LSooriRBVCYhOlIAx4V+GtI9VbPy0J0kclMSv44
SUhzV2ZTqAQAJFXb+K0Ke9s0SD2wbtGhHVrG6sPV05qhxkqp458l33vXM1kEu+EBLArCrg2/+cYp
ZtinOxJEkolUeDtwkVak3apuC3FXGiRo39eTFICcxqVNEAPiodHbnsEopmkYKmEnwO6dB4gzDGrg
Ll17213o/Irdlkq68Ha5ZT9MjJeWOoBJ7sLjtI4vmuOnu5vnMzWkv0TSCxQg2NUB5vSARE9PigsN
eX+XKkLTKBorb/ZZkEDSwIfuui5KklrmFxceEmmN/koRgXmXQ4D9keC5pTtgZ88zGTyEuWyUvitH
giLYGZYl9kRo4cdLPKt7dRR82WqxOSAOFziMK+lcDSdJRcYS2/bGPbigXrdVr26erAldobSEmP4C
g7wwx91PKbz1C2+SqqTDgedbA+O4PW/93KhND8JrlCFswCYpANYjscHj8T3DNoo8vGLgDzwgW6yg
UkPM3AmTMEe8nBxJ3Hu59oS1THmRx+ZGOu0XFQttm81ds2EuFiV/TzNiiP/WcJzP056EuSopMKWG
vMSUOguMYEDVh+kwNghvmEh8qc69XYuyCchzzRkE7S/sarb3kIRreGf2292itAe+KPNoP48x/SEi
KQncINC52f6UBmZbPcN6d6Hou5ZAuaESmYIiL2du8XogVU1uee8/NcL1XYY8q1tb4QN0DZ7AA3/P
STc0e0CVNvDZsJR9TU2aYgJahv+xepm0a8vliJ6xUd4SY/OzIbzSKARBnIEw9sldf3tqgYgqoyWH
BQ31WXih1IYoh8SNpJ2qpx2+HLNsz1L0ZMZjHUgqLv2qzFH8KDSaw8yjm/E8ZCEoCMxMyBhR5YOg
AjWggArUl2jy+CnxUwzYk295N6t3z7T8nT9qpkQvcRSQzsHk8fu56xLmgrDhWAnLl/cjmW4iKq9o
acKElsOoXBOnXzjseLzsFn6EyWjDegN9M/uCvtptiHtpkZ/0nZpbOrC0fJYCakLlT4gLQ5SvezBa
k9I7vgQlDX4GxhR5lua1um2p3BAw3ZVgY5u9g/vGL427OvaulCDOXoq98KIEY4DWSSySmKUNkRZq
bDaruN1zteDgA74V3LgtwV5XlQFEPh9klajVZvgzmdQZldMeFYGR2fUK6u3F7lwrY040F8AltG9H
ctXCa123uyuloUJuNbK9ov29+1FsEBX9QeYcgUUPFhcE6lj305qjNZuTrtJqCMbMv5HF+07Gg8aq
gKD6iCxUUAx587d38Wb5qSz54owBIG8JW4g0mHyBfNdGdwpM9kBom3lY12V+uVaITQwwVHffE2s5
z5KORIXURWiJyRuoOF6+kgRZHYGmrtblbalBgs8tER9Ls2gy5VEtKuB0s6kQx9vcgoJFhCzQBtrh
Te4e/0cYsqYGgWL2GmETm2HcY+rgNoWwSGZa33G69cQ0+CiZpcZoHa88RqE7fjoSULbDymbUAKcH
e8a0vWrkq9bu6QHDrd3IgnL/BB66cmNHWXHe+65frE5doZoKYJ5hjXF9xv/2NgSHHalQoLMjeXSS
pHVsoMyunYxZedtSEIVOUihhGy97tuZSmAyqqiiPA89l4Izt3brFlfeQGQz5AWYaUK1kM9XaCdMy
chA6cTSgDrQaHFAZsrQMfQZfqRGr3fife1pOoZvOGyinB3XsWnGf6B+8+0TDCGgkXJhFYz0U3J0/
2SC1SrufNmD2hhLZ5d0LbVamJsneo8BD2hhuDthEbepDlEtOl4VyxOBBY5huHkHgsElkNa7L7SSF
LYa5LxFGZwI0lI2q7n8zdi2xjQQ952u0r7pqanRioajQi0egLWsO0NqMOhOULkSTyw4XQAECqx/9
tk+Vvvxv5g57Kg9M732OaFoaM2OJHlXZ6b53DqNBsL/NQszSfgjVYFiOLskLoVilctMm+odkZ8ph
0D+y2mFWKJS7TCG4R50noCcRRV7CiytkAKoxk2gA3JV1OyCS5Ju5mTqxKwJz+owb+BqB0mF9Z6Dy
MOoVQIn368Te8IyJ98sP1ctb7lpLKwIwGvrPNOIrDjVXpR5J1FUhdoQVtKi58p25oKjwvG0S54eW
J841KGnzIPOrzsrGP+6Y2F6h57syQYsqZ9GrH2VLT9haxU+uXvHN2ra9bIE5Rhh31X44V7VOOcef
Uz43XSTPh9W372t/g/YBhIimB1zOS8gzCZxyh68J3/BItfg6namz7g5AV18lWQbjxqSFpMwIzGbj
guz6qKHwZzZYLrcgnmuzu+orOknDqSbuhZWEkN2IDX6mwhV5FNbfT2RfGbirJGSVbT3YluUFZoLx
e4tgWCw5/ePx6IDrFYS5wogjkjG4ClhFfVXoLZYRhuAb1Gp4w4Lc3SqWlbUWUtAvmLw+Vg0Ukr2J
QtVVmOa/jtnU5+cuaP9C60RlcfGeHbqymMuOgJHJe82PITYP3CnhLN7HJF47iGCgG3vU60h7a0EZ
pqwBISvhkybnpQ1euNf/loMUcxXcGq+TSEHIzCVbTZ+gb+Dc17CWEvV986uhdf0Ps3z1M0X2kjkY
lbdRNUVKBswNYM2tGvQi+/W4N/Pb+w60eTpvBzDWDyqKdK9kdhr9+ksA4+XChcSHR5t2tQnfYiZb
mPIH/LqXcFEqpH9Ltc+YsgWaAI1VY04qapQd9MRH7BhLFVoeKFFFrJL3QtJ+4sVg+rLU7Magmes7
lH+gqm41vJ3kWhoetlA9VA4AczN2Lyg6Y2hq0TiYsJfAQLQqxIPGy/++DGPEzA2Zm3m3XJcXt++O
kX5LOqJ9ue368uUhtsPI6nH3sCbextJqfSGIijwk802hdQOq4fqx8lwKOLRFfnXe2B/3o6ugetMo
i8cHDs2up+2Zhi4M36reHl1UYQjRFD7J07K6Qy3SMDjF8T/0BPNySucMWOY+Yi7t97n4vEr9KtjT
YMlvXFddVxSxo2jn0lIvthPK7+I+GFcGzH6+hh0yzRArRjgF4ukP/erWw2vs5PbLJ03KNor8AJqA
wwMeC8ER8/twlzLyt0bjosa5u+OzdsaMA5+0iowQ/FK522KLYqO5qjAuYvLw85Uw5F6i7nLSpTTu
6D/2kyro8uVjhje3abFr/83Ysq1+8ISWAivKGjeQ8jHqppKmnNC7i521YSNAH3GcymfdIy+Ng9qu
eP1Xbe28Y/buRqPxjKPw32VaRzbjaiSpBfVs+UIR+0RoD+E04vuXCENLRxzvmzN3m1mxkg3moWk3
1ht/6P8OqX8QkQyQAb3t3BwE7JZH9blSUd/z0WWvOuvezj8rIkZNkoZpHi+4Em6kscaWZKtK34mP
PChgtA1SCTy0Czr0of/R55W1PmaAtoFynQL3pRZ6dgdTJ95bxkjN4GyfCviy1Nqs/9ucOhvlFjth
pnEk5WbazwMR3yAk8brJjfKw8Y+VkfoBxuX0Myv6u1/gOkkUYdriDVo3fcghrpKRkreYkQoa6VMy
yQs4Q+U6kk9B3D2m0qHv/5/Kl9OKFaN9H+9/XMy2ndBNcckHSgAvC2JTxFa03bvvi/oXK5AH0Dau
NPdLNNQslIUT0Y8Awc8DSagCHtgxYUhOtNdv9FN3qJDk2d5+QHvg2inJv/dzZ0/wMCF6xtEXeklF
IVIMOKADXE5m0/cin39crECOa65VaR6YXC79k8h4GL1v8HFXwBIeTyJFkeUC4m/bvWHCizk90Ibp
DMOl1JL2dhyv9AuHPpdIHgVOQoYcncyGjfpVmNQORDnpgZ/KRY0dGRNzSHzOTjqzcE+PxkaLSQVA
arA8tExbQM45+DVu88i+MDKZvoYoqH3KkmsjZ2GM6FLxt5tBNjLSY/dLa6W8wb1nl9L4RuI+Ghkg
epopzfBqHdBD8vIW5casPWrBaWzcAvSF3VqbCBWiktDJSA4UeUAvdFlIplMsaHpZAyKD7+DKp0nT
tFkTnO8xxmShMZ4MGNXqgx0xGXgccwzqltWidohIlgMpBvV3xUGjcE1hnGl+W/qsCKQ5JVMnf6Oz
4XknivRL/SkDTbhYQpZyDwmlyjrFBCXaFuxNK05YVwLOQNU6epj7LvWD7DcQi1n7YHyZDDVKMJlk
wLMZXsQRoS/M8UwnWJsAR+aLZvrYF+o9kjCirV0zir/q3uMZ+rwkCXn9ZJUTCnusjVcSUwEuRryf
1RTYb19ap5ixlGUFCQ52A9K8LbmO9VfxqF7L0xF+CNo8YyEq6l7y5WvI7ui3MkIzEOo6mNWY3V4J
eH4RcG5/JeMmroviTmAX5HNLZxtb23dtcBD0PpzPDdbLt5f2ZucAZ1I9r2MYcoYoE6Pi7rBcQGib
PV+gQTyx6guF3JSZq0jeyNasUwRnCAB3e3p3eUSiHgauC0GOVJPviORTow0YgAxcep40dLlkJtQA
NiJ5qPMHIgkIgwGxGa5hR2xhU1/+jCLC1DUYZKRdMaixR93Jhtp6cl6w/wiTNf9q1GTWJIf0Be/7
SZEjE14HyFHx4BRYjD4j4mlWgXSEY0G9Gbd++NdkCPgc6GpWfcPhbWFcttPwY8XXqezdJGCvBV9S
X3lEm53nEXe8iTofZI0xq1EvOyGDMkTQR8nDPCoIGJsympWZr3keNojaIFgN7nWUndWDH3yYNXCu
Qxc+W3Gm4J288JRxwRyxtozPt5rvL46VwQgXuB5uNkCwdETy5HXKVerWZq6cieddeDq78cK00kiu
tZXujX1R9zdYF8aeg69708wIBAyV44ASZOkVnNNOi7fD6LKW7AmD4iew/0FSIfGi9NViTZjaDTe+
KsuOBLNNUmawv/z7QMUNGChnXWPeGO0hbc5Ol6dEwXWHVcgDuhFaCFS+BykAcxvcU54K17Mfo4IA
GUGaZnL4HrDKOITYwKQtv5GvbekZr8LbqMDgeZCO647t2EPEd5rEt552/4PeEUj08z7rSa/gDcb5
69yZd3TdSDcVb8LZ89FCoTLh5EYk2S7lAZ5999hXtovfJW9Rm/0eFTFNfw6ouyTY86eaYUXHfj+2
G6MAaWfBtLKpO1M1uUB2YZHBrm1QJd+YrdxlKSuqS+g50yRrGmQEqjwZDvLb4DjAss6ypNYj/V/n
Hmju5Aa5ctc1EtDxHHYPZyXyvID6ryLL+r7FprB98NJJP2p34Ff+rYtKxrNR25I48cwRUhAOjheq
LhS0txxyS52Sg9txzfEa2vb/49t4szaNZjmaldCr76Eb+ADi03ir8iG8dSlEp81CEc2KC7HsictJ
Fh5SzUsk+S91NWndzk8scYbr5o9Q3qcF9O6xVACfRoeOLfUl+La441Djng8P12cc/YhP6RYiRIEZ
FpurT8PURBTGG8yffOTz6PwrQovGvTmssSHg3Tzz2kcX0GLiUdWknY7PqKQJ2ME2T3qWWOMeaaUW
6p3hdIgurbTYgKM88YAuj0ExqnciAKuG0/y3hlbE0y1ga1r/5RtpRDTWk2EXGw3+qm3DLQXKoi5w
hv7dBvdzEJ0NxYLu03cleHKr9E8d+MK6gFTPfVFhYVVPQngPzEKSuX0MjP76q2bOrVCMY80qbs8U
s8nymT/aUPhAGCDmdY3xft/dtbPmEZrlo9u9KFOwT7z/YOZ+dO22E34oB1k4DEAaz1iM5MHBtOHL
ZrT/4deU5oKzTBJFTSb1xf9ApcSyhAhPgKSe4GO0vV6bUlo3u+d66cxoxUVMnoNXvqEkalwmrgiW
jj4xBAXF9yHq26NLuET1g/KT7sKm++UbaeDgXjVG7EILzLsTlZc9k/4uzozx44C2ODAHVxvA7l3L
SR32uuBW8kh1zwCEibEl92UOaFbDr71QarhKIqtni6grT2VPwjPtQz2YA1HgMrsjQKx52+Ddc3XY
MmHlhtrrqfqBpGBgdIjIa4hhqFQqm/dRdWGafMdEZjpk51nAo4642CtC21UHNiF1GhmXCy/mObBk
yCmIk+wdPYh/UsxrMKRKYT3Wv3KQtnTYVibPj1xqdZUty64FEU54Mt3x5u2WeD61DCcIjYJHxrDa
TH00QFQ1MSsQiGl0BB2V7ktCi6vmAX7IyNYnGrS6kIwvbVF7vPw0ZnDWuIFTy84YnBqUUMBaClnB
mAmeWBeI6owkq3Hn6RdCeMlTRBtgGJxrJMTj7NvP7zSc3WHpN3Ahh+aME5S7qcSLDYoZ46pWuk1P
HSBWccxJqzgmHFeQZ1edAjWC+taSyP01OVPQc41UytDTU+x05x7hmPRLYSCIaJIeNcbGo4m5o8vz
vZHlqvAdSUbKyJqSWkMYr6mgEODJhVWzHIUJcq5PdgMEkBzEWV8ZLklM2GfBYbNnYxf/tm/80qOA
aweTlH4nKUjNf7JZ0Ze0ZVaubtCtUkA72Uj9+W/gyGiQgD7xF6u1e1/t9rWTw7sqWgA7lLb23+jh
QY4HcKEq2IWNTJE+M+VceN8senawDNwWyjW+ESJFf20gX6XYVCqiMGgSWbXmUS7lrZYz6qDtz6xC
SJ+IZqvMUg4WqR++3Oulzi1/qqm8w75UiLqRZhBJfbe8PyweGjfRd5EJCcRsmWJKaptGxOAd6Ihj
3Oo9jKCtFC4j2Fcvk3ONR4hH2lhkAlQRjgZGqyubzKtwaLywdPryHppRmvCsSUHNE+hkQrUE48bQ
kryCVZuL5L70jLZ9G06km7I4kN6XQVqmnZsRqLYJ+aZoLPQSvBybmtwHKHshcgqt397nO+XaHJ8d
G4BRIJzEG5ZwLWVViUtWkIsJMbJ7cua1hptlmrZIQrt7wJ8A3DbhSZfsEGb8X4aHV8mW/D2kbHp1
FkMWKFx2c1SjamI+jplIOLIYOvde2r6KmdHObKbbnHXHDa/D5BVvUmys100xRiYfaLbxh7BnR+iN
QMo3eSEW6H6ROpz3/hb5rmbI9cNoTrcNffN424BEi0QCi0uL8uxKh/olOiaWksGFh1HgesXt+gkT
w+v0FXfWRo3g6t4uu+1cJLXwK5NKVQwPBNthFWSjyeFHJ0gXZJ3DfqnpzH63aKnZ3emqtTKd23RO
Klns535w7qPOa1rsEqiQQTldO4ca5zVh/zXXeRN3W5MeoVFbNc2eLqCXqfhllPXQnd5VOHcVwk3q
OlIG+SMLU1MqsY+7UpzLn/emggFY1elz8/6iGJkTzzG5iX7fkrpNhNu2MDsO0xNghcJYVMWaGxBB
nfo22wh0sdDs1dAgErjia0HVZDe6/V+h9V3rzUOueaV7myNxIn4AHzlRbNjzSNL/lUKgmCLsdloq
YQ8a5J1nyiA5oEroTi+BezrzICfUq1oTdFeOUHCfIFZ6j9/N9b8tqtpWRbL1tiu7V7Rk4iilvwAh
qTJl0LykcWgXL/67pE8bOvhxaWa+24q6eZnbzg1dXHD0DFb68v4XI4HjZQ3i7ILbPW1eikbZo3g0
uKJDe6Vvy9OFBICuZBU85v6/PSwJ5MdLobVV9YX1vfx9qWgzbgQPoWtjbJmHMr/OYRCo0sXzPTfl
TxWELqNUYmF6h1M8qTO2PwxnQBzPG882uOnrtOv4e4oZvLnoqkrIhIEgtFQ1TdUoGRokeqO3pwDp
hYkS+xP3fjSqkfkW/eFsFZu6up+ESdsN8hkb6Q8xH8NXSMCyJei69tdoG/rM+YmY0pGIzuvZ3IQ8
mkbpdITGeyrVnH1h/J8pQV/8RzyRAR163jaU9lU9ifbVNxbqubczmYaX6WJ10RLwy0hwAWB6dXma
s/ahShsOd+l2ZlqOfkKszebc8YMrrvZmnHfR5+SsIwTDNIqRT7ioDekUg1eYzKCCsYVy/ul/6bgM
QVdvBrdNKKdmXrPfzH6VFyCiYCyTUYnm/qzLLyYz3AEh0LKccaOGb/dQjCzZlP0y7fsaDEVD3Zmf
IZxtBSTuqor3U27PiM+Bg3W1CeQChGOdqyxckaHMJfCx0Ucl7IRG5Ecv1eDSgmL0nIti+d1qYgH/
wBYN3o9QocPVms8w9S/be5QicL6xjE6j/TzQOFvq3ZBuTGH29vakNik74r28EAD8B1vaRi6VWBH7
IyEuutGtehihDFj4iTa1bX3pGOu/EwhCptiVGK/z7n6YwiCHiyqKloKhJ1Nxf5kXC6wxnVAJvEDu
AB15oO6VrZgIJYRwxc2pjpP4qfndyRZG6n/DjFqu+MhVwRBR9+B0uYm9Nzo4GW4MPb7+zK5C5abw
FS3rj4GQNK/zDwSuhH74pO3pp+pOIGHve8NaOaNuhIWU8l0WIDEOxuRYYHDznKNlK3/PvhTkXdGj
w54PSTpdd5w2tjB9ABby5cf2z+rS18V6anHtKQQlgmBXNpVKAKs43Ywo1YcYIBP6uRA1aXEUI3Dp
3SPV/nVi1pCkD7DysTBzTS+73gaKTmO+e9/4WUcJ6Qrqq3DCKiy6uhsUNTi2ToBZYqkEZOTxEID5
Cd0SPspL5OoyDf3m8YG4hBI52R/sfzy8bz3MtviAitNFeLvVs0InHuCWY+sPwmQoD1QiA73by+er
fW3uZT1q+XH9CGEpGnu7lM/LiREPC5UAi9CL2TMhQpqaK56e+ZG0MF1dkqX4m73RMpRAKBtCe2XJ
FZE+xhcQzfCwDYmqBAfFEbnIVb3xb7znWHly2zCCphpB4DDWYX0ykVaMwJ0Zpd7LV3He0Hvjwe1F
8W9xVevWsUR5lCVeTdBB7jRdAstujv0fTuASkgtK4xkgvgv8uPY8PKG30NMgWuXw1LoFBMK/d4fv
NROhE6kIUGt/vlBZm/+Px+8zeW+Nws4zNpygQoCyYr6Ft8wGOihSQ0XbDJ9pSWH8uiFcJYYWPZiE
IKl3TkRGa5wYhPJkfWe6pU63zQQkTiO2Hjx7DuEer4pkj3WO+CKWncb5vYH+sAX5IhKDco7UaUDb
IGVRp8TXJtKF2MV5KqdypIQxoP15jy6XhFvjDe7tmSnZM21xl9eECYPm21v0fEfAeEb7Bd4KRpCY
OyQ2h2N1Kozf1CVk6ZRv07LEEzeR4bzo2sV+jfae9ZYYxfWQqHHAg8BL7Qbtmc3QyChQComO9OVN
eO09RZ0qPlzPLcwzhSu4+wocl1JfAb/fGAv8vNDUcHmwt3JCBQXqXdZIy7U9/VMQAG+k0GES0C3k
oscp1qQMToJwxHJ7M+lCSdg+4KqA0DZHFHnuo7b7/wQDiCgUS+cgS+N7JsZ092+ctBQ5e6yuniCO
UEAscgM/o1aBa9dPEATrf4QYoXT4RtOeS+cYrWWJNjb+2FO7n1bLb+aN4tXarnHp7d94rqrqflQO
mFv70lAmaADWf/1hrNSlZ5nCI34KhmRMr9SELs9BEOCrfLzq+Jtm+ubngi1DOWgWQcsNVRJEJ3QA
l49Da6uLTSzZ/Aa1ptqqNO7JSlr1RvjFpX4LAKA2CKT/fiuEhmxVXydXrJBiQq6BCJhYbdeE7UtP
zRL479ephxKSlD6YaSAZlp1QYPTm3mTOHUOJYVNFnvXMXGoGzE9uH3PbYHAPhqrbtTJdsg/QfZxH
sdZVg/oTxq1dH+MknloyCfXsCFTarEywVLx5pqPvxD4Z/BpcS9fdpAAXzmdDP1yjN19BzJMlaTNM
Jp6Uwf9wYzpMbUV/xIfkpevHyb46ceMc63lovtuyllYNYBuNElrnTbxxRyBKcg0ww/RDDisDKCJC
WiKzWOhinMO6SQz5OzDcs8PO8oFnQi9EYEW310tIypZJ5MDhCgq3KoESxUERhUZYHUUEY01ImP4x
3C43Lki1A3mDVjRvgkFy4/rGF0X72PXsk7WWBiDDW7GP3T8MfSX6azLqzJdpOgBxBC7kAHpHUftr
eDPAz0/NillJ8dA/pXyP9gfNMw2zSAxgqgPMVRiK4Q+81uihdgl4BTmH/QZbV5/ALiSK2IXhnrMR
LHOQ5qcX+p3ixWJVcIc1EzJEPAJBeHJr3wLE2a/ddO3IRGVnbY356NaKDTRdKIl+KCQV90zNFlGs
qpQD/2xhsLEmo/YhOqj0xUKag5A8gDy9eGCtO4TCoxLa30zaoFN1xfxf4BOvUNWvj/8/qmt/+Odf
5ZM70AoJjCaTJRRlIOXIh+hqmpZRX5lns6JNiq0+TE1B6VYT8jpv9ZkXAYy+HOkd+NqE2VH+E6Qw
cYwfCFjEEBIIU68w9ygotVJdZzro/yTjjYclBKSU3f/oJRbVeLru9UIEppScbsX7accFvnjxtlaH
tjoersb3+R+XQYp7ESlddopA6xBPMQmDarbO2nbAgsuIrBFvjHa7H1tkF4wQKjvPR5Sc7oGT/gKb
ui/M1KpBdojw4ppqKotREhOgTnL8bEnWoAOIZNoaR7a4hr2yTbdPcOJESOMOvvgwxpfhigGZf0Gr
UXz9GdU/d+4TmhYsvuajLhoyEDCrdfJpyoN1wLTV+/RQ7B6jpZZpZWlpI1YDos3on16fT20Ao9kF
Bp5ZjpaDetmW1SFT0b2qUjB0e7EzCLLTZQ5LdNE0sykBi+8AnIuaXjfFMX/cxArhepRjRrsSS4r6
WelriX4tR2AwZ/o+vFyqT2yZV/nekOvU0RDsukFiWJXr0L3EyXHA3LgJIBtA7CWR1lQ8ayucPw90
1uQArJvN4wUtuGo+fvOalW+aZ/rfDVTa11sbC3UZppFYBmSQul0sPQLkrFBc9nmvhhyOdNJoaDd0
bg2zaJ+6+HHMXjoaHziL+MwAdeP1syJ4BJbvU7VkQ3Ct4Xu+x/nDCeFGUIYsSRQEVfbNf5SFw0ZA
vQ0P8sFVJVFEwtsQnROxu3w9wA4lhBVZJMPM5HxXoUTAHY/2N4dnS4+jPOLa32i9m6Zzl+0s7nqk
HmttTJ2g5I8g2XbM0BeZdCWXAoJFMClVn4FJHMneU96lsYgsMYXVeVH63oz0jV9rxIHzi6lR2hIX
VguHL2qczCqlYr199aZG0A/HyM+15F6Je9bnBpNZEHocuCH0pLoBgs1rGCcJX2Vx8zxM1DQa4wIu
Dbiw71WyCAzp3btj7c3DAaDyz7DuNVaxzWg+s73gkgDUqK2QcOhgmm5tBRjSxfvFtmZYUKGvY+UR
AY1nn2iyPB5XBEVhfDhV411AohQ/zY9pietUlLLOWDLLRdriIlu6pZcOxal3dQgeO0KHJtQmsWcA
9PbynO/XfyXcgLy561+0lKLhH9CU4rTMyNRRJIfwba4AqLk2hpomDcKiFHFbaPPlgAx3CZ024LKa
y/p5A17OCqNbclp6vevVP6z71N8HH8vQdfFQkw51omD9d08HzsKxEKCFlQ0eMtfLY5D1CX9Kxxlp
eIZeP8BZ3yobQIq8UjjAddrchMJBs4Roe56NiazKYob/wTJ11GpIMeyx0C0+qmAgFVmPpKVa0FQ8
IOeW8yKtZLBkeWE1C/NM1IGCOC5GRV+UKjJkRd7VpO7Yn1i34Opn1KCh9pQr8cFy+TaN2ROJUsLA
xAbfKk6ECpfNa+9paEQjYZgao8gR3xv4zVG/ygSF9/rdCIpmc9RVAcp5pxj1DQQl9uiq1slRPG+I
ovjgiGPmrIH1ZeNDKgXAAx5pYtCQz0OPHrW8BLVZSo1HJCpL5Vnj+TnKc2dek1A1huGFEmLqghla
ACtaSk2tXMiWP2cvw/T76S0w3IeUAT1DdtUS26/ELPrK4/2D6enzan7r718FGFLK/6SAniWtuoQX
LqR+91VOAFV5/PdrtEtjCQD0QgXHoxy6mKZFNCnNL4wW9n9QltwTBsa7iq4KmQ6Qio5Ttd5q0b2H
+EHYelgNG0oAkb8QxOzwciXraeMd715FfwEvW5gZC4oZ3npUfuqtedrEce1QRUIRncVESiTyD2K0
ZEdJWs/OyYknprXsnAPgyjLYLhNbJrcc7g0RstAYCVvXQpEOTCi+x+GqBG+4MEdhCKwd5utVczCF
immcxLLrbbc7Sn1p7JTrVZKv1ITB8o8TJCbSxfLtCtaZCJ7+IsGs4IJRmyH1TivB3hSPfM6MJALm
Lh/0pTPpzHeUHbjwrkXG2OblEeIt7n1VJHhpy1esTiFwtW3CTcC7E+o0e2P+XJnhww4DZ8IrpsJo
JXB0gZQjq85eWBJZuu2SAZdavdf/HSeCWJQgNUbd1kpSToyGsj9a7Yj+cR7CbrRvRy8lu62FzNTe
F61hR36BFH8VfT1lnp6xPGXALwxqhrhftEGPdakrS1Rkty7oSDKEoqFSKmNGlzzk6dAWj4n6g9W3
DnNwuJLa9bqH2L3qnZuyK1LF7XuEcA2E3rG6hYaJsMFrqtnnmTMTYGUZ6wyczbHNpg+waOQzpM3V
fuSVqVkS1hT9ZvSkT/r/LdANITBKQM+kaXvRuLNISq9mWNvECPyZ7WhkAnQpvjyL36C2s0rgh7or
7sOjvm7YaIo0mzm2FWT6LNxG0eGDPxVFSyRaDoqfxYjc5Ph5adCpBBGYe/iKSYyM/bxEg01OHnbl
Pucs+i7fnU0sGOzeBijv/JXb5Iizv1Q1DqtokFzckVqCu4lKxChR+RCxMIm/qFnO1retzhRQTzVK
dKLAqoJddVWr/SoZMkESMwb7RQVLpCGS/lxrF+Jc4YT7gkQZifis6LoccYvgOfNxJ/4HKk5yzuSn
IbPwCDv3QNo+UywGA/qg5phZTFEpE6GGsr9ntSGLEKOLHhs0h7BvJ94ZpU0dGXue035BG/JqT2sf
z0E5Z2DGb2QkroIucSF4w60yjh8d9TmB/w8odFvnugHUJGZldHgGZiQeeRRgYxfc/GTeePDmz24Q
G62FBVy6ioqZOrtS2UIPlTBUkukBUQM0OZhIupZznJUVUsaInP8qmJ37dME4IMAalkRv+ZXKqnlo
trXTykyblyqAqGw6tOXwJKOqp/ZzPafgukDSZhU97/rG3IOL4NWoB895j5SHOU+lKyhWOzn6aYyo
ZfNSl+QRaQeS+hH1wpxzTtJ3tXCov383sidDyGuwCTTUB3eJRPdjH+HbhIJznLAkQZTrzy24qU7Z
Uc3uxnqB4CZ8DkaaZoRyvvRlJr6P1MOUvm0n/65Geog4WFKzZASe+6OH9WpuIZuYLk+pu/XshR4d
6rMxRUNoUUG4PG2dtGutQRAzNWeu9U8XgPuBU4Gf/AGJBFaWJ5+iamQGBvked99fFaTomiHKYJxH
IwsaiRJcyd27W6da3IuLuzhAeS7R/9oltC1eGMUXOjAH906T5M978VG5DhWOuwIncBaAVnHv3U3W
smU08zzjRK3VrXxB4Sf/WUdlj6QzCCOr0r76Zrv74LLC2LGGXVmk7SqS3lpJJns36CqUsyM8rntp
8TSRISbsNPDkGxpha2EyFvo5fZufS7XL6fGd+i3BSG2S1ubE1ekKIIVszlphl3n1+bSUGdXw88Mx
FYN43GSTzTuznLE8VfH7JSUgF5ja6WHhKTUwTtBTCZ/JPmc3IDzF6cK9GMbQXNOvaBEdEQEwPTWr
3zfM/FOZEnBaZhjIgvE5q9VCWkuQ+Q1td0MWfSuwhv1LeE1YTwYoSNNW4bYcabNY6jYKxC5fkvzL
N6XMAKYBwRxxXFH9UtAhgOoLMA1xCvq/RHmTej30clSvoCiXgVNWm1KzyIEKa5l0R1I3w7cfvy29
hRaXykJKonqkhfDMWEgkQ7RPyFBwkgw86JWLW/vVx7+E4O2Q3ZBhKFc3eOthPAcdd0JTX56hIfag
UskA+W80dJstb9iqCK5EjCc4AerA+QBkwUO4t2cVRIaeUDuZAIQJk2c/WcSv19up2HgOxtu9u4x2
XXjCxhseDWGEz0tQhsNzF/oZgfoHeGYpg2+ZzD3mCsVYieIFmzTIBbEylfYzSXhfrb7pL6+WosC5
4dKHI75zHYD1fDPCUQFQ7pfF9+wc75tXFrlmat5lOPGKXnGja0Ic3CqvMmLZtkTPmAfVk9FCFVB7
Uaa5H/n+UgMSlBPJotYCd5mL/8Iug09suIK7lnp4n391hv8VT9zm86IrIugw1viQc2YIXa7Uv6VV
va12JJplfhhJ0tPOzbsuLERjjzkO301FN130zdg6mVSOX9BGVIByc7pEUB4pw9SzsLPcWadykng/
pi74xD9BLxJHG1lVMaXZWtQ8t/4M0JV8fCHLvTPqVVXQRDpuxLDcUEB5du7gL7nEIqg1q0yUP+Hz
8lYdl6zyNub5eUvHP0Aixtpd1lkyelFXpvA7Ia75n/ef9gWQUo99KCRAYMV6x1lM9H5xmVzhKW+2
ze+ioC1Vmxq2hOMCEhSh7VjTuZfs/Obclm1ZqpuTBWyy13d7Mv+FtbwRB8PCWuoZop0HYnfJxgr7
fZigP99/m3wfTevJG13l0wj3n6E6niLzFCnFPkBwoGXzl/Pz3+bobg2D3cjI/UzlVkB4mByv6wEe
9n25ZpYDe1elXeXb1jkFluZC04V6vR2wS3L1dGabTYzZTqw7Y7ZHWp04FscZczGPM8aSqLwmYJb0
oJg/9S994QD4Wf25ws2lj+sQWzKEayXVZTxXvk7RNYpMR8UeeKkthSHcyq78wXc2HpoR/6UQNOly
q/nAKcQpCd/wvLwC7ICqS1Iz0fS0Vp2mJmuPEkcfBwXNSbCsfq3FDBcz5FVSz+lCOrmnMvYxp4rq
itpKtQfxyKmPJB2bhXJ7JQGI211R+o472znd7t87OgQMbOMaJwdHpmAX3Y2NRDG6MX79WpEIlAGV
u5Srb+8EoLUZi22QglQ3ZD1B6+DJRRsY3kqLsTxEFERINqKNe7gdBREn9mWjK90AoXRZJkPNBgtD
bwf/NHlPOaWISaXDPR9TmqQ34rXNreeCMP2R21TQHzlq1B4cmN/V+GKWJ2aWpmExbxUTwqhW7xme
70kGj1dzzRv545OYeA/0lQWOviRQdOddcjoIHYRG8ES6vnSZU1Tg3fqm35J2+S77cTfOx0I4RVi5
/B94udnEnsfD9VC4mJTny4nPC1h+cfW6a3mnGjuinQ3frADqA/rN2UDd3dv7+JD31xDikvtpLgem
C0+OY0RupRkuQIrr/eVGMlLU4kSVe6Z2jl3D70c/fJBUkitGUHO678/1UZYhYPXKsb8/1tPKc17C
glQcwavW9C99rTk6SGJcYrJB+bkn6QxRvYxMvR7tho0VPZVTOgy7H0rG+QkUI0/WUNMkts0lL19L
IaPwhMEGEXNK2TRB/0edjoFAEy/cxpSYeYbaROvWUFqixwun8mZLjE8paGekur4HG6Hmb/TXlPkA
aLPo+hDSNOKP4UMG0R5dZPEvDENIb7Wbk+3s5BvTSr2c7Tf3e+rVSxe8aHWxN/A/v2O8hXyOLwAu
N5xoc7a5zIsy+UNb0lfGe54DBknIVxJKIymqmtiSP0+7LjpIsZUfOT3FbLZ8XhvOedNwKMjpfnc3
pfIQBlOa2Oo3RgpqT1m0+dnaB+ra/8wZMrwodyh9JU1VuTfq9386cyCd/bMafGy+qu10cl+2yHkM
K/kzKU8V2f8CBDvzNkJy2Yia3GhAupsdwXOw9XhwJZ5no4nqLIs5kOf64hFkPPJ27MSenGW5kqnk
IxtamOo1274nRkt77clX6PPnWu5zg9Ejs6AnMS3fbPRN4vcJiS1OhQo/Sq2vC2cx/YVv6I4ZLE+A
713LHzH2Q9mo0He5ODFzNWiCSUIxFz+ts06JJdxG3VjA/OmPGZbGVYTmIMoUdq8QRo1fVo5thGzn
8gbeBFv5gwSkXqaH856HNj3Jvqty4DrEb3edwVW8MIsuivdH/THEPxnUCiWXj0pCk0BbhSqQ05cq
e497SZtlurbUwK46cmydDHrbfZozHDUZH/hqL8siML/O3fLnqh/jTz1Mj+yEotHVxbiJYG4HAJyR
ZSHKDlai1+th15aghzghHGFHde6WwjHC3zB9LsNkfuROVqlpYnL3iAaHyrxl+JaX64+q2m72HZCL
Anryu3ONnZKlHUb1fVdrRwGn28SpZP9mpBqS8ota00CzskiUaebdNVlzdol/ZSvPwaVRfKrtYXPP
MFRokhjffdPgTJWMrtzQb72GxvT/Gaga4xrtxN368cNY6iIpwIRCS0Jv/tkkp1S48XQESVpmLeHA
y4v9ZepQm1zMAKYH+Bjy8ly5wmkRxbEmma+861ircq1lM5BCgz5MDiXKeEDb27oUEE7QX6PvgHNA
liYNIKukjA0D7ETPp3KSHfjyokiM+HRo/hjYldndc10bQUGGAWeQtpJQSoZ9t0uYlVQjbF5tIwgB
JZEp02mJmQDQubiI/Jlb1yJRCw019TP7seqNu6CSiq7k6Mhfh0uhCkz6e8TFiScCoVG3BGDIlzY7
ORHLYFk4D+10Y77Ddf20TzUN+nff+rOZd45Ta2zXthfR+GJE3rd+rgp1eHmKqnjR5oI5x39Ze5V5
SLoWTkQa0E0K6q9u/j9SnSvFxBKqfnx+DukD2kiyebe/l3cIxGJVu1E5+8XWdTkQNOHIwUHUxwa3
IRQHIJ+CLyji5//9a/8eXn1OZ377Y4GLpAph6k5AVTpoWwDVX+rYlKuYh6q+wX9xAuJ1FVdPmkVg
u4kzic/n92kyN1sCQS3F8AZzklhaYByTYjCEsJNBYvJ8+vtiJ7DGld0S6awR6PhLhNdLZTzgCohk
7xeynLveKtmIWqU9+cS6IS/8+yvT1/DIHhBJ39e2f2ZFl2RqV4GA4GwUlu3nbsqgTZ7Eobg/bX3a
AK3PiZi8uMtTnWeHUeSYREggkOERXSZRbrSpYcWKpbBAFrjwjjYsI/BvTZ1d6InmiBZKaFr6EeXh
dv6NxT02vMVhGyKwsTb7NKCnNHxISaz992y5AYcWUTiiNx4+1lDPld41oBquRdftM44Kfsx0xqUq
HN55PiCbK1JCC0MECnvmUeN7ViM3yzM8bKFW4fT51wxJQK4QyZ41dehVNSTjcWzxXWBvVXoo1Ryq
7un26ZCjwp9LaM7FcYy3X8iEwEk304ASMVDBkLvL0D3qoxbgWizKMW5AvM4GOe0q//ImqUtBFpYj
wXcrb0UjG9DFMIEFpag6PFYkYmTHWNI5wdXPmjRlrucxZH3E2XV6VuXKQ+UCfvrYbTOxmIgRF2Ef
avGZPfCHASULCInZkLFExTVEg8QIpMwajFdjrTDIoQu8Ttvi/GrILENFokEHWDIYxgErMOemQWDq
aZjjLkFSm7NCk26xjAqMdC6Kr+eipFX18y/uTcAXUvyypK8emjbaNlSXXEofRj3u/NEnrFGOjmCl
iSijtK9XF0QmwfPZfAWIThPKVGkVFYC39Vuf6/RGztfqv3lXaMnrK6Ji3xOh7M66op8feqC5Vsta
qx6UO6o3iizsixu760qeemPtGtKB6jyXMKQRWT7hXEeXYJvC3IDm9JDCbgTkv2GqGnvjhIrs9zNt
VN9FLxRmxFrMLZ3bLQzh/NXSB4RmDxzZddkX6/sYaEMbGq8eLRlqMq5+hViz/e6VEHZ8InOPdWYS
3psL94II7HhQxumlX/TlT1/RoUcqbzGb3R/pI3566lEcBN2h+qAKq3R3EulMJkQ5FThuHL+z1qlf
A+Y4cuQpv4yKpgwMA1DwbVzz3jkVy0QVhgnfMEMbCnhle3r8ac3cDJMmgNtSKCMWmPJkIjRUdYny
BnAweocMdgGgQbnMB8Oogx2O1IYAgUyqfueXHx10dfy3IfZpki0eYF200ERCncVYzXbVVjCCF1eB
oVRr8soMtpXK/ITwsOtIOsgV3b2775wy86M4tXwoxQAo6QI8G+jDkeCm2sjrQTqarqRHLP2T7lqn
Ntaufqovo12HOhXiVtekaCABQ7OC+4MCI0nBHVDjUu1UpmBzEWfG+1rPnYr2WYTKxPgB8ouOP/rm
Lh8KIOW1sMyxKIXZtty21jvjx1pGY840+jL8zCg25VEN1HkLKl5hEFgnmRwKMe/QiqAxr5gIYtAO
l+CZGJp/4ioMSok3CgBEEHfuyEz5L2HpmWd9/4owu9jLIwEkSa6OoZl9hP6DqGXDduMn3ThDzPAs
Eif05PIFgKjsV3BYwEgwCnXtq0GcazfAOtHL3QE0/dMpKpGE9bE9QshBL8TkVRBRFi5UsSvB5iLE
XwPVegv7PnJnUXLN1DDdHPgX5JcNSn2fPDMEjlxSszzZIRX/SZ7KlSixJMZ5/GD9BuuxzY2hEPHM
fvA5YcogGVvFQO4cf3xOSgGEYACBkeKtz58P/QL5Bs/M2CTt7wdtomGQIJcHqPGaWMjdQ9uyG6u6
Gg7aVt1C7EgPn+ZQaZdbUQKx4jsbl5PLxCFihgBwaQc4We1Asnl5f5JN5qcapeUa//aA4rpFvgIP
vyzQSk7Hw5/TnFX3LWAIEm9CLuO4vu28m5r9R4h7+Lb7VUu66HlSbnIWiovmLWNYsBRn0vSj/7Ci
sone6rBRz4tYjtv4zcVicqj+6XfuyeMOEH476yywsb6zk5Hj9ZiW4aQiERgT2yWrK3saHRmo3tA0
nGF/tvl4mEwUYCqAghhWrN+nkeS+HcY+eg5ACvDGdCO4vlrHtJ8iw1b36sz4wPFoE/ABe4ZdP7kL
cKTRDdM549NZEysAL0IxwWfUuP3uQEQVeQ0mU7GaZGliBqWmNSafQ5Qj+I/KdCy+XDReFtnKMtwS
tv5LSKZ8GuokQtmjaMP8UA/HPzQ235BTel0dgpx4dMusEpyboCQRwsX8YyuKcYUVXeJlbm+xd6om
m9rFF6hxsyJIJshlgTTcj8a/kbN69sjLJ4V7Tb5TA+kFHKRWpnARp1yoEXLIWrSxLyfAH0DIw6Hw
y30V+/35uHf/sTYE6Jna3Hh8Ayb6D6IgjA/Tji9pi7X1yHjvf1Vch3acAdmrpzEHrN3Nqksl/uCL
tbIxMji5dFfWQy8M2wyupd+MHub4eFGWGMUwJiXrIt0cDoTgJsssi8Jv4Lscu0TrnaZxYi+G0oMV
k/1aquIMnaPOxpqqByzURx1ODUWX0wHXOh0cLJtk64APT6wu+vJyDXspOC0uDiNhQhQq7lvlBVBC
iDAw/vSnc9o1XH8hVIeM3G43t9445VhqmJeY+7o9HjERHuWTrs6wk49itKInaaFHkTLrEXNfM0w1
Xbcs2DC7Ksf7N7aiDMXsNRIOJIEX8C0/OxwzIFSh1AaBCxbz9Lm+f2zydQZZF0Ucu0PXz1TpDZ2f
sELimBRyFNWCrGJo7GIG+EXOTk505U00xfoIeQzetWTbbHOn75Xo0j40xp6z+572D9WsoFEr1uRr
/H48OYcjHw/DW2S9nOZLmZGmt4Rhm3Pf20jbWCqw7B9wvfMsxkUg8GQT2VKbekTskTQUnZOr6lCz
vdtOImRLRce89i73lE912gaKGJHxoL+SbbK89Yt6yO7ZJoBB3Wgt+uw+qe2XbwcLkC9TTgRZVf1Z
2BxsXBVd5TmWRuOYFlBQ99nI1P+VLlnTDSo3UgMItd/gEbUMdhSuct2I0utihx0cu/BlSlugmDqO
GOApEO2Vlo4mXAX1Bedl4o+0oivFqyc+rLtI++dkNV9s92aYaqsPvFDgnKOb73Juj5jwjBavud5w
e1/Yb03hgKQfKQfZEuRuahzW2ukXtEPVMndT4o/2wE+PXydrPxsWg1thzaFofibi3P2KjstWPIc+
XuvQcUy7Bn+dUK5R9CnT92TtrgCJ1ElWtfNLFL/M7KJ6/CN3qzcEZj4pMdUUHP9B6kjmbGa4gskj
yxWeKsGxEA+179Uc2285Z4hXvxKcvGmeYRHZ33NdknRyVJn+Dw4Gbb3pNlfnfuQGlYHMdXnEiIjv
AU9XnsJEEMmxrG3aGu0IgLlO6qN7oopdSV+34GFwIFY16okwZ4AXShde3pUJe6otMM/ri4g4vrhS
HLNQ94CvHYvF7MxCy8AoBFcBdw+aa/3C5AXGqTMmRqGOYANOb6VQ4rplUQRFDchjJohWN20b5J43
6heCvrQegvTNFX6sg00zmE3kWNwTAYcYzBmaBy3v+D0P9iDMGLQil6hqvFwvP5h8DYDY/55ynQE6
xrzO+Xhmg6AxYpws30jn4KTuW/+UX6DxUZzV4dH7crdZ0Qn3C+QBvqaHTqOL8HoQbsqrRtllpk+I
N9EHfC2IiKTulEz3+ct8L1HebJBdgow52LulD+x1t955tHuBRbD67piY5uNxja48sEkIxo1Q72hF
+3MGnshAdBhEo9JcSsLYkpOSYV+MH0IxtDh7xTCFHHJrVb1DEgkXXFd3UqAdF11ieKwuzsbatWtC
6pJWf/E3zm8Eb7YvODcqghjelbQRW56Dc5hWwdxkOCNrs7ECsaZHvg50ddWYUxoWngAwpxS8KHDT
H6qThgjYbhIU5yINdGMkaaCSOT3E618fytkQK4uv64shzGh9CK3nCwvntwXAIkQb6n5HTcoXaoAL
8GESG7H83wz58O0BlmtwwKbFZ3DqV21jlAXH+a7v5npmpz0ntWvy/NrmtCB3c+hl/lCukTP2Om1J
Mb5HQUcyYFpOK4ge6PTojwOtj8QrWQ3tE3Zoa1EdnOiV6NyN4ekHbnx0shVHK8QMcgE9hOzSKf14
FbwCwxTACwSBtceIMqot/VokaUAhc1a3XZ5LaJNDlfUdj/HEVXX1Lf4r+TEhZ4dQCfwusabvD347
fRW05RxWAThmyV+TA7G2ownX9fjcl5vFqu5kPOQMqvTL4HMFYcRE2+hxOmBNL0KO2q9Nvo5bci9v
Nwk+pSZwdy3mPVUmv3WpfyA+K8/byPRl1ceadjsPB/UmL4PbbxCJhkQaVxAaZ2ahkFXMZTHLiMjC
CRycT4YY8u5K81iNwU3dMnBylaYU0CNg0+ipfQerf3cKgZFkC6Lu/0SQoWsUM2djkkyS55173/nm
k49W642PyCnAulvqMmpTvylC+Pb5cwg0EOuJmOTVMWv87VCR/TUaxEZ80m/uGxqK9Q1HHrwqdLP3
Cf4XSR/KWsORl2+zWO+BTe9SLEFCGQ7fgzbBSwWrMkz8BzbQZOfR6sUbXAiDvdOBmVrF0LyJ6tpe
nZTFPdANYHIQqx0FaFXO3jn4YdXzdUIV0x3ntMhthPlk6e13XfhJLSi7PGMiHZQ3ZyxzFX/unfPf
6WUmGuX4mTfrqc/aKregJlFWfcIW7C1T0F0Cj34bLVG3MMgLxvfbBtwoKq8fczmeW30Xf4ZCupPB
GwRUhsktH75XqAzjAzAmv+eEpCN1gcyhmqI2YsGvs82D9N7qDU9pvaJ+KfGP7fCL/W+dNhnsjvMW
BaPwMaMgbsXhfxqIx2XxIZX80ycvZ2Vtru4pcVthhR0CvS4ioeSXUyV3RuqL53e8bTCJn81wztxn
fBPHrdSIOrbLokxyV2RktTbTKF1BSosij50r7Y4PzkLaGr7eT212x8QsLqWzwlU6kiyFkoh3SpmY
dIRBm4WbOKxg/fDDo8PCQme4MhDa8PSymeVuAuxIubQlH9P6NKttSpgXDcnKABIqJGdetJ8XEr3a
liv9Q+sCZ1mzUvLOD8HgxMxpr8B6lYCQd5sEaj3sXweCetgKvoBPdCxbe4+1vFpqcTlpHj0Ez+0c
faQK1ix/rNZoq5FTYLega+EIaJOWKW6kshY0elbUMG4ASrvuHsGgAWCUuDTNrgdJ0kS/chUQ4y8c
A6dIa7i6fHQhp4Beu8c+HZaX6i7lsjLdD4KKrdntzMTdrpYwd+dOaaIrs9b2Frs2BveEFncU8slG
lIZuUOTkPLu5WXY4/UaiiMfholBvtkxaeTC+iBVfuoFRfvdX7q9p84g81iEIUeUCC5TqB0oQmXnw
x20aEigfde999KzQPEf2lcO9omxVwCIRDz5BClZEC+ZHYYJ1JsMDF34Qdy/9uzgQ9Jp+MIGeSfV0
CnN/SWNHrjF1pRZ0ilL+1z/od7Pi+W5SdHzMhLAfKYTHwFOcuAXfwIoUcV19DXqrXNDf5I0rHhEV
WAwHYlL6x/Ktb65MRVft7p2I2QQI4NpxAbAKL2y6gTew3bt3VcPR8B4yN5XEbr3JYqwPYa28jVX0
acJHSF3DIDqAglPuBYxA2p4lBmjR4byF2OEYerOqodat1c2IrN6NvgbNFKPViV5JpDTUXLSL/h+w
NR+R9k8Y4EFqD/Sno7ojuCqHqYY/hos5V3RWtIuF78mEDJ/Ii7MG/z7oUuFDb50nhp777WF4LKBL
ed2+XSIt6OP05MHIUylHrhdcmlLwWMfD2WrL2ZWdy+a63igON2QmpNLESBu/IMgurG3xQsbKWvCM
drYNIfwSuDUnALits6VG/BHvzMsPzKpTI4dv7o3Wm7HhwligvSNejZ0fDsXBSEGHAx7Ce2oWutjd
7Zdrm1FmqDsOHQ1+LsjpU8mVd6jowszOz5SXN+CgGMS/PkdYwgfofU0sR8CZ+6OA2CZ76t45TFbb
KgBDXImlooOGw2M4zMXdK3pA0qwOENgV9YGGEqwHMuFTmCDXyWRUlWlGFXp76qfw7AV/d3UgDf3D
RT1GttXfhBZcgNU21EqQ91RxWby4wPXkElU00mxMC3oabBbPSaLacSDgojZ+a/nb/oMZR0wVsjRA
4iT4y5b0VFte9kI5fsMvHPIybcC9IooT7kUGWrpwJ2NxLfF/IaFPmSBrWdYniyBEah9KmfVcBfPk
N5imvjwsytf0b+EtGAUTvL/QGh4EmW4n57T7sqTcQx/1AKe/rLrpGMHn1Vrbj4cegT176Xx5Aalb
GGGGLaAP/kRXNuTWkAmL1PgZGQF9EtH2bSlrnSiPJnSM50dwiHeEJoW8LGhLBIiVE3oobauPeaoD
AMpT41B1AsqhwZtnKHlkYNQKJ9XYoykPYGQNT3l0nomyodMJ/vjN1GOA/I1oXDWCjj7YMXZfj3g9
a2aAJuwFs2FPXrIJ45lOiEecfYkEtJ/IMM5zDh/wQ2SaoCBQZiXnuyK9Nrcrs5TBR91vkrNVtjy7
goylVj3kikTJDWT8E5mQYEFDipqETagIlfu/YJz77n6AqTxpYWtrwauguSHj0jZpRi4oe1C4gctN
besPimXuZD6XsxYxs0j7184n+1PZRU78QzNGZFfnCDQpG3bFX47ixqmzrzjTl14vJSNHIATSsHGP
ojX3k0u/LjSz23UAGD94WkSm4+TEf6aHGjnFIq0DKb10IWtaQPT2rs8PnicvfD3jLjfNKhQGD79A
J/laZLhak2lekzjNX7P3Fg/bxG86vtKCKGcoun6pSUk2bvlwazN7lUwB+0O+u2b7j/ACts/BN7aw
3qu94QyJvDkLwx7NknAXeRT8oOLePXoG1qqAYWU12PA+SDRbbxzQmT2ZFqM+Znq0ZXF6z6Iw0fxi
w6S7Q2rUrCbjHj8bUeeIxjGZOH3gcOFDZQ7k9mtTgCunVXJ4y5cbCcLgeVlJNr1EhjkO4BcWrlbj
9gHu4gs/Z5lwAWoc420OYBWColHVLiQsFi9Myk9T+1gX3U9coyfAuypx2UusxWfRrzJZb+amNu4v
p5diy6XTulWWmt1t4GCkfww4wxc4vL5ChdPW+JQhqMd5wEQ6uDHcIaYCWUaDdQYcSNgst054/8Rt
oi89UYHl/FrnAcJqTPeLxPqaafMpvwfLfV9cLTDWl+WCV7cp8ZWm4HLP2kCOrAQ0u6cUOhk+EHap
tan1bdvxUdQY6H2Z7Z8Ayb5tmcvyM3OwTsIbmpD4MEXBY/Wz9w5ALw9MzTUlQ56nY9INQEB6YsgV
rzPa1GbkmlXa6qHxxZz1rV61Bil8fKBQdsDtNMSYn+zF3sIhPXy1bQM1DXt3QHmHJ1ky6uyFxBbe
VUxViRbI4Vklnde5bJ5m2jPb2jTP7gsH+aMfa1XXfvZNeWDNQFX6k4hSV9lYYBUp695pYjGiPNvs
DAmgwmVWjbkUoP3PYh6s3FbBK1vI10Rhk9b3vybVO2T3Ydzmu2pc1WxBub38dr58Rd/20VsRo0S9
S82+Ci+uldqKaDi7g592KJSShB1im3JoFR6ZXwL38RsRkbliYBb9HnWxeNdHTvqkkoqL87lDDwLv
WqCmotsqCa2AZ7Yh4vLVLzkNN9eoOcZ8JMkfwg4cZwIizhQFqoeNjNXShEmi5MRK1133cDnYtFzk
TzHrgXFJ7kVv/K1C9t/6RC2X6YG0wRsQT+NjxKWIl/296Ryf1/dUw7jRdam9ycLE4/zgJuIgsvlv
XJfdidXW6w63TR5dtjfEzj6Ba0M8Z8t0gx1GKV060MbxBcgDArwbqwkYN4ii/95H5csdv4FffEg7
8H8DrQ8uuUhABDJa8EcLODGCt87WDKNqhMcXkdJSp/yQn6MLqLyZQvgOhCy7KINgzCHnZJquHyBt
7Wq6UAOYQ21nfbYyRjXEUY/E5Xqvku+bw7DzZBiVTiXOnlDAkZAv72cwVrmP9vPtZ66iCKF6yyR+
1QmugCPvIPsTG0qBREy0oVyeEr/llWo6oP/ltU6q5bl4dPYWOGisvNYFc2ZieZCizBgSdRaYr0fg
OFFBweEUux5BZThOS2ZKmLfEhbW/alRAxd4dyJmGnmb8IXNKKvEeUVhXsF5W3tDXMh1MwDddRiL8
Z4bmETw8b048CChSxd7H6P1/uXHXvP/hfj5w1X/tjt7dsSciFcqUWFSa3tC+fkx5A6FZTvphjvxn
sjA9YmUN6I+YyeS3y9Ut8JM5xrvhxQytf1uFWwfY5OAwCXhiVi0PDxg2vlDqpYRhtciIRxnFHYUH
QmDk0yKiXkgShaMUVuH/dbpeivv2setS92Fg7zJm7z6yES+rbMtsGJxdr3XaMryazesQfWUjlaK+
BPqimqWHtkeziz15ZVfx4vnnY/eoUdJttksli9+lRfZkN7MecWbCvgCIJJm+szNmBa2qnqvB5LJm
CMoKQOabZzuyXm3yjJt2OGhIhThKCj3nnJPyCTAVtGtDvxRkFPNocLvzWbQGy81reOwk0tr2dndN
M45TYg32woW+I8wdlVc1fiPVd2wdCFXetwEPnnnlMyeDYxWiztu+AZLrzgv7OERx/J8odfaS5Npr
NhVNLQapB4Alfbnk9JvijplSalgyrrk8a8Eu6nWCpQeqEaV1Jc/zsbWi9cvCfAE3ILdwhAt6EQGu
+3eytDdxs41LiwUCz/GOpkvzAWkm/fOj5DSMP/Y+amiSBZJUR2d/pCcJ3L2RoAOXom2yC8ecOnPd
xTAIMJ3eoSsnN7Qo395pGUruKmUNCRMbaquHqL3yfR5rsa+032aNsttPhph5wrI0MopOhQt26xSm
3TZrCDho50LX8mK2cbOpLxTLRYC2bwB7LLZhlvVt/jN/EfL1jl2XG3wMlj9CkDbednGKRVp59fYy
3YGKCzJxWBjCN/cftbJyX1KbamTWp98i6VxnLDNBnLKh3eKoYPWulaVFQE1/epYSsKie+MwgFi6e
cjfAi+LJmuQ7xAPXKhqtKAEB5FHSudWp8ilaBRvz55S/qpuqL0kwpSCOk1Fc9uQCqYlb+afLSkey
PH8gsDoOgzJ3Q485H8jbMO1DseCu7qf7DPUg/gvvBIfEtu76gEbB6vWcLf8BTqt4qckw+bB6XhWe
/Rf7FArFxt5Y42ZFvFBSXj0zLqK2oWgdzvk9QEfW+aef9JDWoa9Hz6EnWbXhijgrt3PHp0oWmBc5
PfciiISZ4G3mVg8O31GnST3rU7NLNqXcoPfugahpt3rEzlPn9AAoNE0PNta5wXgZrVzA0KJoo1bp
6Dq6JNrFpQvNVadvEziMh1usjzEWKrNIUkUEfAR79SqNcHQHUdSASdqezS7xNEintUs6PGiu3C/+
R9vGwPjUtLqFBDz+9O1CIq8XgwpZttQo9HehMO3AjdELotbvYcmZyq/5uf6h+1VpKWVFoanK7V16
xmEO/rop5QD59EvMEsks2sloI5BgjEIvKKmtVZ3X97No8V03x/JG4HyzITvlKhiV6IBDkxmbpKMI
ueHYpT65qtuENcdkts/+HdNE5WG/R+nMkz7EUQljoShJfcxBMUc6CPiVEDImekTBuaUZGyWgeZKJ
7+aYv8OF8+IeNmyyYZ7u0igqQ//uB99TXrI0b6m2B5vS6DE6o3drAoBUfT8eqB77X67WOtPGXwiJ
7qIRTAWjrk5JNyDxtZT8xAUMFC/HGiFPhQZrUs11pF65klbXShL4mD+SROCe2Pmw7AjNhYYBR93O
bi4CG/raDYzif/THmqkg7oGlflhD/hHLZHs8DI3gPud/SWXmTuFvYbu5rxOTwKXpyWRWD1ZYYr7z
15Cla6Ijj2k/72gtnlujdwXi1rhAmhNmOxh8iBVubBwJYZG1Gq/EPh6Xy5s+ovl3MsBPzJlanM0R
pR6LE6Dd0m6ik1ibUbCCpZNZwjtPqMJ5hlx4N6cw8SIhS7s9YhVBXeZ5lnJI/x2hlZVf4tlhmnuj
7rWOW4LvIzXuEa3egUdZJpFVE6YLvw7JCSIoIjkjrJ9YeLzLh1Oj32WG7KOg+SSbb1QNjakYtNy7
ewuEJ7tV/q/HcoH1vHnSClrkD2vvxWVSgvUNIyVWp/04d7YKfXzJgT2NilNhJDXy4Km6OYm5pczo
ZEvPrtoQk8oc+xwe/6Vh+KU1YmWRQUrdMAt2LAwGza/IwydMJvbXpXnMW8uwSh8ghbohq/Dj6iCf
fJJXl/KuCoeyPwlQHPN/eTcrzgikTjjBI6rC6eM6vHZ04ruXV5znJ1rqD10MQs59zbbftHd8juMG
to8IQ9j9y4SUuHMhXm2jQJifArj+4dMrilcZnbcTWJdm3za6irEJEV4BEnovInccYTYpPL41qBjk
o9r4krhXUxnwnQh7K+CtjuIzxE7lt6NxDIh+1QoG2E5TWzC5GSiOObnk/IwZtS4bPv5IjKBd1EjG
+dQhEVegKtO9Es7zLVQqy6qUeKyCSLXiVZdADyfA6UqhL1Udp/j7ZikO3Y2cZExLwMyp+igBXV4m
L6PE+MkrNKxdhSd2J85es8S2u7y8Iu1IClCu6BzSO73WaFS3wXXQbHaGRxVJWhS2dfM+GdV9Djpo
tM8EYHxbY+5gopL9ZmtraID0mEz6dvAqb3C5hiPuwRXI6DtXHbfeN1olkIcheFLOiq+Qilho6xQZ
NNZX582tx7tEEJXCwluZo6GAKufFcVAJx+d//69GdAHFksTmdcOAWkb/4Do/GszboRP/UGcn0Yy5
ReQBdWesxPgDG/MMf3lGE8XkDgZjBZAEdE0SbZEcMzJzWdd3EGb/hFyu1lEifTPT+Uq+dl1FRr3r
8h6MMKjJMk3GdeLdW/8Ka4gBIZEGtaIYAnZczq/GmK7JovnPbiwXxNuNCni837ydmF46zOQRhvyh
fY0jnZyGdBd6Jya/bHCgCDcd3g06rgWPCYvWnlTMsYTjnzQOhEWhh9bw35iykJ3cZkzT1BpDYf2r
CjRFqQhHAhpPPsPiUUmfCO4/JMXnZFuzdP1UX7PZWc0zjHkU5bfaPEpT6grgiK0eBAP6EICMQeVD
BT507uU9H1+ECnInH86JOxLJhtetyplbdguI0csX+fxCr3LSYKNWOYEJ9UirSapwVkW1/cjCWKnG
hoAjMRnZROG0DoHNyIQqminGxkaGFzsNt2SGuEhdKfF5vgLlGOCMfehU+8MafHuPwl+LLzfTgy97
LEZqKTrrX4xnUOT0PA2ccBmc0egOKkZE+bEJv78oEyru/lSr/NF2WDv2dZJSnzDPSmRtIeupKtL7
L0fy+zWhQL+m4+NTly/tdRwS3oUUc+nF0AwUTP4oS0ABd6ocgN3eL6JP3TQlAbq74BPnfsYY8nrn
48nhEWcf1u7qMWQMrq8q5LecKOmlX9D3Ci6RcOKC9+DEpJIrjF9nIl+M1z3J6/kWJRZpwxv++2IR
abk9P9JseIstPEhrnn4etOOBOS41Kft3Ogo9XOR/UZpfE78UgTzhtfnR9FLU3z5jJFoA39rPm5IU
EZqmsUQIugdXO+YuFbsw8YqBTIjevUPmMhWScemFVfppucwHCkl+hBK+GOkluER6llNkMX2ZSFEU
xNaBqxEiWeCpBIhRSGTg5mf9eH8U5O/3A7EucVs+K/KPa1guDp5QNyCAyOIsPWla5TGJzF18zEa2
ThrX2acSwq0cMFa6mODNjxlVInp2Bpkc78P0FH4xiFYGVRaciFOjo4uJqI6FWEUepdFItGOno11M
6/mFzyyv0gikHv6o0UzTITCIGU9x0IsP7nLzE+Bu9MI5YZpnYFC7w1bMJp3ZsESud9yDgLQAl3+Q
vwzwJsXOm9ml/pGYSInif+wzIcWVMPt2RHRPuDnEcVm4nPHp/ZjGfQ2MmcXtiGnOS0j2LIGYbIAR
bHLWQuJKG7hgs05ABhtZmcHCKfRdO80uMk9G589OxEoupbgOdw3etDHnVXMGMVrzdaTXKg/QsVOV
uEVLcgYwzK3fEfKo+QirCW++cOeOUPi7Q4bhgtE7DUCQ1hXEjeTHdVrhn7JhKTSZE3nZKr9jy9rs
CGHSv+dd9OY3qNi6pcu21iExFI3RxwFdZfD4odGK+5EDRCCyOIE7/nGXoK98BAWkKLLzGf1ZWl4x
fjRx80B8Poj7XIZmmCkb+obKLrwX0hdl0W41trBtvgGPL3EaigBBAYM6bNyKwqy8A67mtbtn6qjM
s2pMQlRTm9N2KzMN2hCxt46sCzK5wR+nARm/4Dwg7fDN9PFTzEHG0ROX99g5Ik1L9La6EEUAqTyN
xdK0BIQrofJOXo0lkeeNLFSpYARFcm6/9qDP2DkFesZI9aal/c7ZzhG8pVkknNi+DUneY8d1vH/0
499S3KITGpjbwWFwGM9AvJZw7r4BzuGhJdxSzks3+DQTS/8HuLQqQdB/3Ox3RR1PgWpy4neiLw26
S37f1aJqDQaonLAEdrq8KoIouQmSocx3krZ8+G/aWdoxaCtd7Nby74dc/t5mc4oyFvDBOiXMJJ7r
mraXFrTBpHxchr9f6THcl/Mnf4lXybWSzJDenQRwLtMGFCmSXX8dAu6nqC0tnhfYqJFnev9Tgty7
/Kc08mp1LekktkMOh0Zh5KVxIn1UdsCCbw3ljlS0BApa41zglkrDJwOR0zzGsW8otRM6+nEzMC9n
2GGPFM7h/mVIPFqkak17cq8VHTb9LCv16Aa+ElS9FBWDlnFZ2RlcslfaMXWkzffjO8V/ijTK0ysl
LNO7ZJ+a7AUcXQY0FWIc1DGIJM+KpK1NkAOIIvAMRZAG9Dko8TbTvGhIWisGIb5VH1cU+lwA3Bv0
uMGCw7MYe40fif2rpeqep0NOhYZvQH8H5tPJkOeYyCZncTTZHWLyyeRoyGkimzy2zPpwZfhhuSkl
es2LDvuFKEngUnusTIX6UTt2Uds2/DQPlBad9eyBO3MhXCXfUbfWcoP8FaQyXP1MyomgqXSeS7sF
S5dKV9Lkfgz+D6F+qVKMhiB3DbMDhGk00dLSTt0l4nym5z/2qEddDTjT8eUVZbPKI/o0G7eT5tki
ndhxXi5OTwfTmsEENpXwFXi7MIUlP+8CtSqrKeE68YY8CSic/5zhgHHk/hTLE1Ce4luhnwr9rjJg
PSJwy64f3X8dxEjEYhpICngG+irWhRvGQnQILhpnicTK9/3e487GOxCAHTnD46tE2dLcNESGLhbt
uROodxkerOn77BU35TQEIgQpczBa4yKGaVxklpm6qR+D7gNs/msd32vYXeg1C9HGC/CUpKDFHd/A
0W7EZImT7JSZnSq2j1/i7D2RyfbUL/NBR1Uy2fWP3SMcNqHTCwizLCCdhQtsF4TokEQ1gDh2YEGQ
QgHp5ewxTRlMe9YWgSPqw9lQObGiZUFQEC6wYkDdY24YepxG9Qnl2KnEy/65BttFVLrB3c9eBc8d
jVgf1UWOsb2t+S0vf4pn8XgFLBBNtcA6zIeOD234vJpxASMDQo+28lWU6i0E1TaDhqAt6hutFQ13
2qvvgf/4xH8n9x8ld1YibHU3dxPxrkV9tAgRGQKZYAIVT/82IyGuZ9bL2KJs5etZNMy3xhXblBAj
RKy24H6t8Zcf1AbkeGr5qVClMMgwoFIwVr/KMuvBSN6x3cG3UlY04fuOSBRuyCLirnrv4hQNsogx
9bXK9p/aZKtsCz9/wkxOWe1qVuimuMdU+WzOY7E/3rk3z29DGx9Tg6PYc64VssnsoumfzgWasLVD
kZwZqiLOt/AScw7SN7wbKQCsrdQkJJMZmzKjujJyBSIWcgW2QlDaDgJRbR2GwVrttBPyImGAwynh
ksRMDogkIt/gku0SGMDt1AN2rWFhOmcWpHlcWiwOs4TWn/+El1UFqSYnF8yidU0Lc8gOR+Hv1XCj
O8y6r/+yKPsXdu0C86ClXL1A2OHg9sC/xIcUOU7FUj9vi4qUgJqNzaWvK6P8VFG9Cjm66ia4MZ3I
wCJtT8ACMcy0CoFinFxTi3Az7O+J5ncta6t2ZOOVUH9NX1niYCwER68+PDKBHFjLcT6gvyFOt8qH
i26egOWr82K9+uuknFUwKAqJ51OFIHrs+7gEUd4ZijYA6EaCfd4/Oa9IXAuuA89l2MeHnqevGapg
mZSaHz/ZPVbqRM8Wc11pHdVB7b7nHFP+9ljYjK3kxxkX9i15HbOB9DOuJ2EMJMjtoZz8Sxi3VpZ+
oq6UCZBUd45iJBnIt0QrQHjWs5ySIBIyE9B73x4cJrNXXfkBe/q1XT5pPWxLNHM5X6NTbjMmCLs0
wUeW4X6BXNmJhh7RUmsqOZqEQ0u/XebInHfKg63HEZHFQNsO1DRkpFsXxozQJKJzDIqufF4EyedU
m224e3StrZ9OxyUW+y582eWORYUaf8HG5+rC4MHE9yUf587YJr6KRDe6DtUuI8a/W67FVhvEEwQ6
qhno0yBkfHVCPuh8yDE7UJSgPXBxqxeNygGlqLM/6FdTOUO8m7QCbw+OPSUDYuF7us15iwt38szE
4gdOBoJub76QGxDAGRMzqvG1boQ0w/wxQsErP5oPO0KvL93RSMFIVuvIJIXxW4C6SO8N46MvWhSv
83V7WAUXSiSWdCKwTkzfqkFQ9toVFe/8QKmThypWm1pi+Lyz8yM04nirTl0ER7ZvNGbxOGRrZG3L
QgRxtVIpDtSiaaX/uSwDOolo9D5hq3wT192NW0QFavT6v+egFA27Cpg6C5aM3/7/YLvKtLlaagDO
Z8L3pgU0OtgEMsW5CBmvq9GrWjbIXO5E8zY2VWsEvM1Xyvq179qlukXqcfFMy6kL7xmK57oYNZyK
JmeE9qDS3fT39icZsr/wXSoIeX2+ug5DDYVKOIBMhIpoD0S6RrIquaFb8wgoi/QwPDAkK89+4ajA
mTIuUsLRsBnWdBws2WaX0n/oM29dDjqmW+niFU08txbZMCN2QyPrI/EL0IRo8cizqLaM7w9+FKfW
A/X3YPs1SkXngzJRkXZGsCOa3H/8J0uhqFe/H2blrqjlJ8X6pZ+tnG4wwPRj/+roiFnSKj/pAWjE
icpUpixWlw1VQVdACfQ+3jnUwlKKg8ELnbx5k34mU2j68I7yOzGdJe/3P2P//gqI3pqP7xmLRkv4
JuF5uYNtZfKFmF08Cr9sNfx32sGk/2isU/GI+eEFv7GFuQZ/iip4dfYBXOiuENLNHqQlCS+LMFLp
wpxsRziByMaz8GFRn6hXAJ9iwpH/qXdvqpvTWkbPR2tKfe8gbYX4X+LTwA614iIC6IOrzQ/Uhjkx
QDJow2TE1icV4Du4Iye9QeVBEiWJMXwiN6zXHWqiC5uxnauJSwMMR5IYHrgG5SdHAsE9vB/Ocqgt
0bl/U8v7OKDdZRIJ3lpjMCVCGZbOzRzO+IfI8JDCrclsAHQtXPpJJKamoO0vFgzBorjw0Py8ZXtK
N3eM7lI+KwTREFhR51p7QYhxpn5RP5QKRz5UkExXMXwtc0/fCmQ5zWaLZBRJ4v6844A4xPgLMV/w
0nYjAh48dkOQaI/6E1NZqBf/V2md8ODfiYr4nBVypVZhVVqTDuyoBlTD7WK5mTZrv4i8fshNmcWj
4mo4RP2KjA7/NSXeKlTggn+S8ZRSeuffP45YKQSKYWuWmO7c2Y0cIXLNdOPtAxoeqcQn7+aT3Jev
IQZ6TtSJYLsYwDdAdSA+VL7I/WXEyD8BHTbGZWFrLSu3xLikuZuuqjUglW4jSFveGBgaAmwA/fYt
bzfKT5LfMJwDe+LVVghIYfaA9u+LJ9dggCmAo4m1rrIVaMEGrhrLSY8MGpuJ38tjkBrZWe9kO1E5
1lj4do5hmx82D9gckK7z3++oZCTJvbEDPiGW+AD6ZVcQyeqJS9igQ2DsFpBt6/9DqQupTC2XA3JY
eomqM3ynnTUZSiivRhEb64nffsuAthd5gt4crs90dJpaD0CiLEU6qOIJcH1TssNufhGRdkcZvuQ5
a6umWo7Poq3fS1hRXDDbmKP3wC+gPmX5/AuTQKb4MJwBr5iS5qowL4Ja8nuwhZ4DK7ahNohCCqZf
JpfrDHrIMJrsdsNmfiJTUdT+xjXxZhj7SaOv6D1bsSqZvd24ierMwL+T4ih9kKp7V+TezOQOCSfF
89kdpw3HZ6pWfOTSujEKBC5rfkuLv+e87YAdmJMGkBlLLGv/m7ibNvcHy0tZxS2Cj08kXMlrOg09
TgJLNfB0FytbPWdZFIvlf/vGqS3LNzVkVfSWL6DF6WrVCy6nrWo6hWQDtQ7oEC/+RR2+596qkonv
PiVTLpa2UYX51dbCqcl7MdWhaJ2FU8DzBQL+pRaxlBtD8Xeg6rTh/NhyYLhvUyTMgzHKPSUeai/K
TRT+gSaUGfpqUPUUpug5CtlBKv1uEdj80Dft5fM8R1Q9jKrcwMD8wH398mrOHeJPaxoTK5mgG3/v
pk2rKCBIz36twmtHlgikcw588y7GCCEK/nNe/0npK/o8HjT4CfT52ITNJPxOktZ1aNzoBFDl8HEA
MsnnSnrPmpNEN4+wsCvvYwIwSG1LpgN+DHSb6BUXibIQz4dK8JStvS2UDbz+tUS8BrDuwOVPRLz2
3TYyumSpQu5yu+8hhkuVAulQMNKF5p8rTEsH5b7Wtx0J+NZjgQA2gBYeJI37z//DUry1JRiDTb3q
2bl19TsWKxQsMnqd1lU068e9PD3q4d0FxSsIhJq+M6bqNRSpH7iwsJv+c9k668HrDiV9YqGkvIWG
pFTDYFmbWrQ7Q7nmyiWaRX+OYOMbzeZLXvT7V8J5+CfdoU1k8fRTWV4MyM3eq+v1ztsMDDpc+Ykn
xopS+UBtcF19ijCRIbOQjG8QuqsPdQZq2Q85twLuUqOAhwDPpYVldKfrAqxo88yE4F6Vq4YsA632
s01mR0DBIFnrxO0/Di+Vq9eyk00eBHQCR3K4ioJIvwP1LxUPzyCrXF64aipjQ9akTnTqAFSHS1hw
f9D+MjvCfZfWkGIgw6d5LESqDHg6VtkjO6Yqe+8S8tscoJ1Xos7h2rlhEpFbMNlTiwOnTH/LL610
h2MBpQo41zONKeDDCOMVgGvGG59qW7rxGx3pz5hx6mB/cXqR53pqoQk4KSPIF7DurO/boz7FKHDL
LIDkCROD+O+oD+s4LYt1jbVXDvU/LnzXSKEfEKVEKXi4csafkasNXL4t2WMTpGHHAcq4ebjEkI6j
57ViAv+my9tJ5VTFZT7TPeW4F0+rX1DynjvEs+07ZtAXsxTNKFQgzc2BaV9lM6nD5ay2pqkxwCvY
V+jxoBRH/30YO180ZcTj9d0qfDB4VOx3cqTxzE2kjo7Wcq8/I3MaKpvvr0o+j2D71dxjnhSam9sJ
eJJDinybqGgafZsUMT6XW00YuQgTiWUlRekdVIDagQy0RhoC0CrtHPHSF9PLNyJhGT7lq1k3DP2q
BhWNivzkfiz2PKRClBd8BCHiGL0kb9mmDZIFjQOXP5ao4fT9MIYrJfWAAqqwo7/KSagUifNQdtYV
4o1sVjzr+6j2O2pKy//AYIEJJEQDh6C1w1gb7YICAAFOyyd1tGbq/ey8M1WJ/UfFeI9HiPq22K8F
pD58h8uLxmZCKO7TNHSzOByJtG8a1278wqLAQ/42JerSDYpMA5wU5WyiuG047wd730Bs26YdJ35r
iaRgnaIrHpmObWQ3AjfFVR+F5IvrLO/cysIXfiyb1q9ejHu5t6KZfeTqdPXxBVpb6igxkwgOADyw
Pc+O+VCBakwVhiuiafuGvGkMXOREbLFRSfEV12z96m9TONj03JUsC/xwXNXqvHnfGTsYAxWQbysW
WapxD4JkP7i0x5el1y14gBIfWjghHiB1/aIoFq2VYcISEmjlNRxwMUBM6WSWZuCYjuezq3YEgtQJ
q6tpDc8nv6LemXcZj7lxj/FMzbELddLqyMYFU8ADeFO/QLQUFrjPjZpCedFBegUWb3m0KD9LM0Op
P4EWitd52skNWOKJkalXiSHFIv5EoTPKU/fx8dg+mNoDtAE/SjxQpIrVGDAtYntgJhhJ5Ksoi7AR
E098Oj4KcwNK1CAuVMmgoqtYbDiP39avdtPM4XI06ONHbmsi9/q3cu1NCAZRvDYh1vKxoKDtFgKs
ngnTANl8lwcqUbRcKWuvV05Ij34V52iqIPLf7+PAg8qSAo/Wdzff2sY+1VF1MoEeldl02yLAFu0Z
fw0XEsX2gzyWfwoA6SWc8ifxXDLAfzOjzf47f5C5vQWorAlsSi7uzVfWyWQ/xd2sUZZlBDVJUaEp
pZVkq/9sps0gdzbtHYBdCas+7xABIbQPqUEZoWq3EnnEKV4tGDXwTce9UEzFYTi8XiV9zV9pwZmr
YM3I4bltxEJCjs9Th9moLLtAw3OmCB46mIwV1F9JL7jlX0+E9zb6f8pB07uy7bAr4SBmytWmf8QL
IENLtfSDI8xrcjLN0/vpdLNsASgh2NC5DDXp7nRaJqxKpK5pjYHTJV17O7JBp9oTwVXA9IF/VCfX
+nhdfXSyqJT/dnlf1ZiCWbvwRnWAxfnDe5GCIyCwDN/DBoFn3HHVCIE8uSpn/2mGpj7gnSAzyFPn
pIOj0g3mYi17CZ7nDRzi0NSogewPTcBUdRbC+of4ONdJgZHcaD4XBmLiXiqZ5W+t79NWG1v7Iv2U
ar9nT20MyAdcrNyUCxcFJW6UtzsARjnm5moIdyuCv3gO7W6Eviwas/NvJWhEBdtCWZNuR4dp58Ms
g3yjFuJ0kCwatGhANbp5CFzw6ZPbf3D1ZoAA2he9mpIFRyL7H0jtgcUEpGgyunaW3lbMMFoAMb4I
w6joBt9peEk6kUt+2GMP6D7uGkr/kR+va9dJkmPQ4zkzHY74A7ohv0spc9mUUvph3huYaN15RAw2
PaKwP76zVBINUoRs6p2wmVBTmHZ5mNJv+t33RE8T+FI0ZuNy0lj1zTCFlFOV+y5Mh17qLZGpvkMd
g1A+p3GRrR7xikXYiJUSRic/JMoi706KO4bbj8LY+cq8AaeIytxU9OtzxmFZO5pwu5lt/ymB60o6
xaSGDgCUCOyymzCBw1hSbJ7eBd0HSdXMi93evhMUbC9ppQBJtKO/BLDzahYLIzrX5kVNFAzb8ysb
oyqelM698PpNXf2mHcVKVNPiN2RcbzbchD3KmAqjB34zsalCltpj059r8UgzMPaJLwh93ZUJ8R1h
kVWfEN8w7LxeO08A9DzY5twEVnraA+m3iglZnUyAUrc1AYZWZk1NHX/FTFfYIUWht52xTGu40Lt7
Z4JMTZFtWG7MYh3dvPbzr3BSUfNJd5a8oHTzhoh9oDDbXlunyJo2cym1pmmXz+tehknc/4/hSkPf
Jh6r7rCJGxpnHvjRWid6Wp+A63TM0GoY1g4nHh0MM2+pADTz0wzbZuS6nE8rpRcUby2Ww+l94WhC
HW4N4BfvvYW8kHRcnDdx5+tU8VkWOvOyDA7jVuI4SGDUKS/VpzuoyOJiedZlFhFOD90i5/D3WmJO
pmb/zwZyvnFQz5yg3PjFQtisNjp9ginon7CHztUDE+Ywk6A9eV//oq7OMb6tKwRUgvXgFHINITro
cAbJh+nXLDv0VPOJc0j+xfRmD7iL7K3VnYnC2JMztdgwMPwKA6gVZdGceLxjW98gHVrog1I9CfYv
VSb+xbMnxMOV4HQPezDLMBxKvE+RMjOaXLn9/eIiv5zCIzAZrMcOz3KIEs8DVDzvbylX9sQIpQij
QEydI6l3WTgjZG7+Sp3Ep75JwVsR7ZFAVU6Priw6vQnt7t4OXPtXSXzkx4R2Ka+qxOb4I0KSSjNP
2pjCb1/e9N/R4C1HZBqNcewIF+HQVRk2y/OiJ9lrCIVoBOTjGlZcOst89QroabnlSrTLRR4C3OGo
rEXOm+T4yn9OfHUk80xZUnS4/D1W9+ubGKmF/dasoFLnqyR72PA55izaNLs7hIG1wlXeqgP2eniJ
leD7x4GlAfXVcV/dKlUFdV18rheormK+qmsNsyNDWuSQ/Rp3N+x/Xs3E7YluSkmySl1HqHtU4Ah5
90OMZb98hECFcNlZDWIlhhyjwRG0JZ91Ys9X/Ki1yo26Fw1LqxAHKfChK1QllsQ5SzQtHum4DaW6
68HkQH4va9FkUiNRbgpUv1Beo3Q0NWUyTueExEskF77vP36sYD/E/k+Q2MYJ0tVZWk7yhKn2g6If
ZwKJMX/GLwk09p2JOWDKp7dZDUsINjiAS3I77Iw/sxJssb3eS2feA44aX3lQW8EvtTinRhk0Obhw
vCkr9QA6d8jd0ftgQ6Wb9rbhXLevjacctQRyoc4dk22xg8c9LyFtEYi0qpA6mT050yoKXD9Izgfm
P9J/ML/xaXAwm2mmftkvPMmIcg/VCaiTi8sX69iopQD9gTKghfUMLrLJPz3x4D5zKzKpbn6bzeTm
tU1mWmoeWxI72igg4YNdAGK+5RUbqnRX/Bbdl4wArMGJqwP5vwwMh0aNhKe6grLdZIKY/CSOquJ8
K0Mx1erSaM2CXdmFb65kOOwJLqQFrrnGcurE9W7FRl7/5Lmp/v800BcwlcyqusLWe1lY3XUlV6PB
Bx5DbWBHJxBIYGw5YIkWsUnfOkNseYeoMSenMtC2TVAouDMmr0siZVviIp3QJb7wRpy0RWo5b5wz
JWz56YzVGLbBmVAgrrtrZvoviqfS00plyZOdi3+36BkI4E230m5mfRGqTYXWmkxtBa8vnJnW81aS
p2w+u9FfUWfH2BSEMgta7iEPndxs11DunMEvBhP9c+b9MxCzukY+9+zoobQmt/UhguYcGNC1e5Wp
7M5DX0YWL4iS5wNvnU0oYPIWsQlZfLaufMcTyLvX6xZ1fbzWpz0E/ov9klztVcUgbg+Njo9/vVTO
pc/G03exO5qkiVHhglTvkTxevpme7z6rSstcbvUNXI6es1D1tiAJiDQa6vhFD/YyQ2UtfPvaWfnW
8LkqBaB9fherKFMfqBuSYVHxeBul/Kx2VAzZUAFj6cbM7PEIRaFUCqP4OaNXyrg63fc9yO99UZFM
jtI5t0lhN9DnK9T0HyfVCGKOgI+GkPeEfJAJ7jFEXW2jplAFlur33V0VKm6CYggywTjQhvkcLdf5
g0pd6Y8AdKaFA7hGnFgRvZpvMxo06X+98c4LrM4DkHxtMwHwjeMFa4fNedTWjtwYd2Qh0shzXdNY
+dAY8yxEGx2prTtF6sDqcgBBgu7CSKgOHpjKxYHTpMo+SzO2Q7a8ASdLZCjuR8sUN/sLGFY5DkxS
xfZWYxFqDOgxj2tCeMF5yuRpGePWHy1WeMe1mOjrhKf/s6k4s9EZ1esrXr63X+Dac1R2/8TNyON9
PzdMwjnce6yrr2CLkJ8xiaEIKaD+evYsXihfse72loXhGTKoWyZUMs+mLAORJjj2EHTbXU0r9uD+
/3VlOFvvArYub9XId/X9z0/FTjFt+Jn63x/FZttNbVZRvpcZxDlU7MABvcBxeJAn4Zcc2ClX7p9k
eJ1VWrLR8dgA29zIu+7QPHfrV5BV5B28r8lPcAinNw8CgcSG3ORZ7HxtX6PiCQedW25KJGT6z7ek
MTmyg0gof9S6+/r95sBBt2O1h4Ywbh/3/TLcde9IODWJ1xdG/7CwYHcNKCSd8zXLk0sF2IsebbKg
RvhGiPVHjjAyF6Ev4qkmMJkUOOLO4CCQ+CL6568BZ0fo3BbqwZjU+A5EqX+nlYFOLYLuPm+eUz56
fUKWzO3kjMK5Au1c5w54SJeApX6RtyywaygYj5cJdiZO/HohLBBP3gG9vMM4kbwGg/h0xPThZzaX
+UgTJVwQ7uYI8cP2aS+HRISKyu5TMUgpfDHLhmSlew6USXXJhFj89cEJ/OXL+nTVZgu4PsgczYZx
M0lW3sJMlTvYni5sqDXzIbbz4wZ/A9+fm0d186HmauGegpbfEhnb43vC9KexYu64Q+qHsfxLrJWy
NU9cxSPMghhv584F9qbacsEEO5zlPaQZZAxcZOO3ChQQ1SHFVFPQwB4E7O6w0QknFheiA3R/ztzn
/2pAh7xgiQfDsDe9h7yfxGrya5Qr3V+VwHk6r0TUPpWEcOtLsdE/AMSbdClmXJ8eJbLgKy7nFMkR
exGz2Jn0hKn/YbpBbkThFhIyy+AlpKzQciU/pccsEWTTPjxl9NJ//9/qxnVJ12HUz6vSic1qRz1h
+nmWLTRyvGVEMi1grzwiuQCr3+Ort7wkS7LwJ31Tl837oTPOq48bZjHochmW3lhDjIFbwaqgomup
pKm+j2f9SWdFRkO91mXXFj86xNY7+k71T1BrtRHII2jbDRp+PQN+/TgukvIJLn1Lfg7cE8K2hKe5
QL7hoVqfrie9UrriXM0pgFNtQnuonsquSKw4gkGVGOWoZ7GalORZ1+/3rTFd58Nhq09FzNbJsmp/
MqbvggDu3WhJBXHWthqf5lby+zrgSOujNhoh9mpvJTgRb2zkUuPvLI99aQtk/0wZaPmKw2qkFjx6
lumEkS0IY8OgyeUcJj2Z+z+FgzPWDAmll8pe6O6syDtkvy6pK8vh15m/DN+6DMMVp3t0+e4SMXEy
PFOttrRVo4E5cW1Zf/iBlPg4AjGwLVepFrpfRVtDxebSAYRoAtEFx58Iu6BjWNCQC1pbcOzxVIr4
admZLudQWnYmXQYL3w5SxFQ+45aiHFOZG+tv1y1acJiEEcOcAQiGZoKFBi+8a6unNCcdhXSj3tAZ
hhlRgadIjhNNolYeMzdB8DhILPamyARXpiaTkI0hcteIaYi73rKRub61zIFo23/DrdZh0LDOYN44
qepSz7WCaegIyvFWtdj95Zw0kCfdVoYlZe9Vi9ZmrFc/sIQ+Nv4rWuczo2O/JcrtTN1K6uYJrqqJ
y1nHovTPGefdQISAxdmoHKLhQPqj3aQ9E0rLfPdQAe2gfmZbj2RjE/u0HzvfXcLhfA1qx04DY0oe
GU9pkCi+lLr314Rgl8mxeJkpJlVT1HJaC+ZxIiHubakIezwKzFAwaA2BdZ/h3SlJdIuYHXN4m5Nf
e7+5A29EnCemJebW4EE2dKjHqvw+u7t3k8e+51AymAmcwcYwb4auCwL9aazgUGVPZKxIeG6KClCR
KgJKkWrqcaLf7R5BhRgAuydJMR6ZmK4fY8OdpQZkyOlRK601mrJjFiQr7CkcRbD6WRK0KYsm2YdG
xfUhjjDuc+FAz3lCXPJc5ckb8h1I6OXUO/fMs2ofcUNht27As+Itm3WcL0pjuBhQWHizRHbWFV3n
SFBpX4dfp+IyBt/ypb3RNH1XuO5nqQ19qHdoR61rcJ88dGyZVPtNKmK6/8owrqeKLHRQlAeI3Xgz
A29Ua9JqlbxpT4nGfh2eV/xvjiJfve9jc2QwDHZQE/NLb2b7hzJTL6XqX+aybV84cw9YHjCyPBwo
Wb9HhQvRZEeQy/VRS0bk0ee8l06xf/uyS54Wgs40g3dbnFQOi5UXIcQ0oLqFuG8SQLCjAdVt8X1Q
WUDU/ct8OSMc06nzBkWwMFwKe/m0jKETiP5Y5C3rVFaibumqOmgTNkVaUBxbPdRxSG///ctdruSc
ltgOgFEqJ/FcSiLmUu+pE99NyP47vpPImmKaUVx1a20wNkHGTeyr+XzKrjkeRfFtAvzFuacfn7dJ
2/Z5YuVfTEkds/76uL/JdJhTr11+ODgSp07thtCFWlrQDxI5tAw/PfSyl//1umHyCa7gnemcRkrv
I0POhHtQ2BTStq9ZPAuF7cBdm+3UZzGVzkQhsCavRHEs+z1Gd7d+zVbmmqhks7lArM6ZmFNw37o4
bnz5SQotaue1Pvgcbfm73rJ9jcZ8llmFmLJVHwg8DQOttvS53bndxQSEDAdB9Y5lPxxOB8gsNabl
cpLDaluBt1OKVXdI5diKHXHSFgPMLSJ+1TC9okSj7MKbCWHy7OKclqHqCGhK8YvB+GImzqeObObM
JQSBnkCpDqlOU0nFcxgaoW6u7nBaazhSvdXTYmKQIie8akUbBaY0LF8qCzn7JMqWl5lfk2LcCUnY
TGPs1HXrdpcYSX8mA1UbpGIdsAuAyIFVo07qDUnFC55eP5es+02izU2DF17aOazKtvb6ehxHrnc8
NOHogH2DCuRCz0K2KhM51ib54B5dpeoG0pwhfLcjLanqXHxd+ap0yVOPthKjDsNP4BT2QLlUXVri
iJyb4aaCYf0d9MKJKQ0sst/UmztqtI90renpNwO0ucD7Xak8gLigb/qVsHzYEVsm8BJmoP54eQZV
sKuws3bpSfmZXuXoyaB5BOebm0m5aXS/glcQptCY/k1IvZXbgeYZSmUES4KbN0K05tOkukpudUAQ
C/uqabkKPIDYe3/SyQA1xszP83NmgUwLwNkirNSTMLXcoEZ4ufTJeNQPl4YcpBO7it0RNrw5PGRS
l8SyRaO7YZ1mnwhMgO5qmhQt+HaR10XB4vq9/8JZilIkfxb5DewdQAvx6PZfs5wVuovFdnA6rlrB
6K0vEk9cFOO9HMdUBfiuH+Q9Bi6wtd1ZnuSP3IyLRxZ62A28l9XGa10M1uW0F7oRzbod6YGZ/30J
rVV8UXPfVZuK2ebZkmxRAcCo52LBFHQNttcT5UCNFJyBZU72ai947gl8i8NnJbK9wGT2BzlY4VSo
0ewhzFdNSpMV2z7vHMdYV1DX8ceTjq+D3R4583jNYiu0ZZcwmD7nPZ0FI5/KC4IBH0AwZswE9gYW
/lJqMetWvVaEGBf7evy44wWqzUtp5vLbCC3EiY7MXp5fYPBxIZop4+EEbda5Xj19cy+3Q0L/MMDb
8EfsfKWcXFZo9g4CAdBqGYMq9Bnc1pRoCR5Q8n8S+OlvFCq1eqpGpFxEmJiuRGJKjekca6aCDYxT
Jrn36FaHXPRT3CIHYiYKrRwvITLS704kPmxH2dEgfMGBNjI7Xe+8WOOWazYH1CoNIxnCpJDMHiTI
NgTAp2Zt6f1xPizQOAiRV9Rmkdd5ow5bz8Gf0nU7DSRi8RvlXm6tPvNIDY8a0muFf3X5VirApR97
e9pQ2D1rimMj8wzPMv9R58DVo6nsVgyQD4l3MLeWRGaPcbs9oo0SElrNd524whctk4ClFQslT7Qi
my6jBwTLasyHG1CCMdbb94APSaMQ0KZZ5sAzUuSxf6II3pgXFHdK6amVorVfciKQ9Jajh8oSzH/B
5ZPpmU9nBRiuLijlQH00cdQhEpWjoZ/kxpNN3m7I+aVDRgrHsqOCXJJFyx+1Ste1JDWT1fpbYbfT
OiIdqyV+IX9AwWCF9AIOHTIGkN9HlwYkC560IkZ2OemRsAscBL4XRd6wCb9it1E5urvbg9PWCdX2
7o0QC7uN8diYOgR3bkCcF6S+bLcIj0FrHy7C9Pf/Ie2NlmYSK5FGO8stw5J/FqI2YMcjRIvdBzYa
8BnO09tcCei2CVnJh55LPYBI7+QdxjmVcsMGn+Hu8hb/kXz6FUdT9NCbXzk5CuAm3P4M6B7CQMP7
mJYHlA6uA9BOqSj0RSbGr1b/NLDx0IFCNnqnOiZ/RT9BfJRvptWCbfGX6BjjLZn0xsz0IOpXZOVA
bVMU8vmjca08LpERYUZidKBFphCyZ5cklo03u4rVl8A8jCR3JW2MXqYv+gK7oUvz7Ae9AjF3fzkt
mU2QuUtwgU8QdttvWSubdabPWKp1hu4Rhf8BjrQXCVDzMMfOyVC35tyz0YAoAVuQRc7P/9RWtW0C
esBm3Djp1LHVRQXSSuyTPm9AlhaBhIjBM9xNWH7ZwUa0Z2e8tCvp5Ts6tVNOzL4GPtI38IoWf8Rd
+OtOBqB7uhMotbkkNDOwKvsB2SPwzHva/1WKD4HZC677YHw1cBXjM3TFolP6LdS9bOVlbrkAA8MD
NdQK/XS83Xs1dfvLVh0oJPJ6W+CYsKywYSBZcjpjbGyGDPbktOusvc8EJuKCKyREzuPWqW7s+Nmx
MzMYcf24BySTfal9lvqMxYPRuwvEL8BL6Wp3cg24GSYH5sbSQ7gFBvtTVzpnpMXHl9wdSp3zcwNm
UmVxoH/xmSYdCbEMQAotl9nZBKOpGhI82KXHE7npcYkhuUxnN6Xifjs1/6WryanIkGx0gdwFmRBD
sJWjL8sAAT46r1hshMg25jIhHaC9XbH3vSqdCc4PwiEm8JTWMq5lB/gUIb5524kcbqZ4xOPP/xGi
+nT4Wb+ou0P1MzwEUhclDjIzZGwwdORrNUpDVtYd8Yd5+58MHNLvIX8eAT/g9Zdmv6q7qmniP7sL
Nl9+LlhAN714fGiTeu3o1pEE3HCSE22FGJvoADSs+J96fDcyhtFU3iFm0KC9fxo3Nsk8VSkRGPBB
ojIdF/PcDUulyV/Uea+wJOfs0lgpNXCXJR4LX9J1GyAOosWLFyNW/84NRTPWz90OE/D4g/k0BoR4
LO4x+aNdxENGoNHuwv0R3OR3OufAgCBoZNrx1gCjdFjGpbf/htwnQBSGr+UM5jtbN+sCviYjA+Ey
ZMJWaf+gNGJJHwi703v6nMpM+iKU2X/cRF0k4rFHoDUwWMTTmztN2U8LMia1ntDby/vKWSrWcrd2
dPDHR2enRVAJ3agngjJeP4ChV73K0AJFf6KAMLvudsaXaFvw4gd95q+wejqiEAcWyAaOykxJI170
AuVafRQNEQK83OB/HSCHdNNr57hmovC0hF6t05se4+o8NoUErqKH/oXgyeV8nU+V4z8P6hFT+pbT
BqL/jt3KtvsdzEOzwpBocIdJmiPNAdB8CByQhRqfjKDAIyhEp6BzaM4yTpSv851S63KEkTtQ22JG
jBM0VgF1BkuBDZuPC9CHG7FbXSiUvhHp2OHSqkMGb4AI/IV+BO5Fv4tDWtep6Su2tzWuCVThV+Ju
wtxaAaHqad2aHc5EpzKaTl39FqRBFtiM8fg+tJJEtQu+9xtjeUp77b9QsGIDJqaP8sOES/PUvUgD
PAOPuQckubWVeUxmiV1x55S7kkJvwe3GObKprn+knNhqCO3AEzx5pSMvYLmF8wSUxUBzqQHQn657
tHYa3ViSqLY8bbUeJZto1yNvyWJwsMo4l1pf7qlzDD36M8FNMALjinIMC9P86eHLFVj/NhY2Z+OI
pNdPJShr4AvB53N9+TlXXsAcy+jKLHBVS4am7gRfy9xWj08KqMCXpAuU6/qGzHfTo24xcHV7ZvN7
eRRuJLDrIbVo+iOrMCB+aT/YH/0zXhRZtG30RNdneFiCzVQ5Kr1HbWkATUFAiwhUsxTcWcoJ4aTG
vL+9pZxcVdWET4W5uZNw42QuQaVOkVn1/t5LWO2WkCBXx5OQNjmm/E3vXRdPNOO+86m+Xodth1sc
AnD9HuBy8wCXNKPZ230lmLswWZxwdXSY2pdxMicVjJZEux9A3qjzl11orF9ft83MAgEUuiFZR912
DYhsOX95170tzKJHFi0XuVtjpngNif2WFkfkGSYGtNFis3V/d0Ze+icM2dQ3+fyf8vOc+nzUlDtf
AKWRrpeoG6bvgPqWVi+ZyYJRHirR0ktUBSbZK21Q+Lan+g9vb4h3JO18GUUxZmvJCqxUKDR96vhd
jl8gRZo236WH1M5McOCPwrfFyt4yb5/wXPXTkA/ftjTBHK6eZjocV4Ncn9iBDlVOGlRt7E4pW7dK
/OgpiCgLSOINEGrG20isHsVzPHAuDmLln8anH+ugD+ShoyKl4UUkfGh2E88SlXKL0UfUGPM67C6J
ErawyJWi/PVWhFWYRjQSX5twPZWgVrnuWBK+ROEi6b0Fm0P9D/+GFNP3N2sMJ5thupgy+QKXJAYP
DLPD4ynbwDyXDMkDKAh1Uwa58InQBlomYdnRcJaBwGUcBQ0pRiB8aMRqJa0aieDHN3mqovFeNE7h
2ocDYccLHvfQ4cVADKBKqmUKJS5YSMeIG0zc+3zMOVPqVLEhQ8qSLagYUlAfv8VuGoSQYdGlNXX4
HYC3e+e+8Hc9Pmlrt/WCtujyTOol6HjMoW8AAmfjqusUbto32PKTxtR8PJHCT/NMGdP8KfATVgUB
FwgEgOssGUIqTEVT2u8mK8T9bmumIAM777FheOGBeeFounNhAg2dpc8FDC9JO55OgHHkRelbkq0W
+RqscUWtzFSSW6XSbe1Mp8eN731Qmm/7rOThNNTxGjsLo+Ri8tzvS4AaT+bevYt9MZwjRSMTV8B1
c1a8b8plf4otv33g4c8fQAO2+WbJn/8bQhFizOLFjpM8FX324k7AQk220lZ8EW+fMZ9c3tGIugq5
aZ5EztH4Ek9j/QojSZElgOU8AX2UUII/vxR/Al26vJUDQoETe7D8gxBdsnAcpjeejDrm3W9ooPdS
noHQjrpo9tYxN7/Te6iaYyilmpeYgVB0z8JYClIJgubLqX+PtKeu94AppH5xPUbH/KKHnMxbdrb9
K3Gd2vBkWJ5yIhjJCOWUU3ncCJd6aVBBXVb2IeAN1H6eVOY4qA0suw/VBHQ42dt+gWAhug2g12ti
a/bkZiM7fRL1LU1BxKktylsHX4/G2EegeR7RWFww2hfwTmIM2dXxQ8UbpHWxC0bUfRg2+1TblaWu
xKtQ0BoIkV+TvjRePhgCYRHmrzp22L/WxH6cV8t7cbKwPVD3/utdO1lWpntjFrJNVGND6T03SnmG
8C879G/oexfslL4qQcr8Fcy+qzq4D1oRp+t9Xj8N856CByTvE3/HP8gASbNeVpUgb75n4/gpwdlY
BWRu+ftOzEkmCNbCp09K/8TEcfw1+FB8sxbOZ3c5ue2yqNAbecSP1ggHhtqhnBhJtBETx1ePDRO0
F7Owuz3A5j1OuLPqbIZ2rJMC9sbZ6ngRnvIu4r0mIbPxPRM49WBr6foWOwVtEi/V4IP+YLpoIgqv
GuQJu9ukfWx7vIP58Np0cEc1yyR2Bafv+IEa9EF3+zOddPLTCE11RmD3TRngflnSTyUng0lWQnXE
bcCnVAzqE/S1gkCFKn3LXuRlW6C3Qb1gSiY2gUVWQDwhhmXQY83pqXIBpbybzTLaWAb2wMCPPWDU
fMygIMi1Tfw2aJYxUbmeCMsiE0LV/vQ560C1exeO89IXvma0mZTsgRiiD/3vN2Z/Ft2i4JFz8eLp
gT69yBCjerbbbshTl1Fr6Qk20zUSTV+NmSc93D4/j36UGTETBM71mifg3Ta4H8UBimmWI0IjIQHM
p4CJqO7b+AgvwDh2A+tEG7Sjy1tHPAN+rNnaS35m+2g84Ga3d3qHpj48ozwZq26UbJtadB4XIo+8
72rP6onNmQJ6SdDN5+cx90qW7lGe6aFhNOz70QrF6QwdfXQeKDnioBBLAzx7X0blUxCWea+1W6hB
1KljOAwZ8DXTS+TnBrRG3+75ReZxPgs9y0VZlGJywFeI6xRKO6cD1NLHdbK43CTxf0XP0yOEhV2m
WsWZrBV3r5t3EptwV3jyC8od0wWlyXAX2ZZBecvVepksRa+7DdVZN3dcEihMHmYyv8vGqsCEKSNO
zLhmAHdu2PxnsOYCenIHKbzGFggE6hvHRyyJ9ctil0V0me4NaGF7bN93mWstH9NDkYZwQyHgW8bm
N/+lpUob4ImyPacYUZZCfe6GIp38Hf6H8PZVaXYmuU32UKeu0y4S8SvhTrBIUnbbcOguIYq6wAI5
HGCqoLioyX3b0PUNsjN1UMU+8M/WCvGTXwV9pa5SQwrQm31vskbv+kjJ87knb6wQ5BoFeo0PJcdE
WGX8wYypFoQy0dIhqnNotDWy1FNMbm4NLgdhdwl8yB7of4R8tARjN4qN+us6L/IE+fSnhLloSWzI
4FrjSg/OHiTO0+p72hVWoM4iV2S8+EzGumIiDyTIvbea+CgcPfv5bxlIeMhWQMLCoIUD7x49j9kj
uVQu/ALW86KAhRQQQFnZdlkYiuNzTATshPbGA0Kh3EN1G0bUEh1yvFWJwAb4s44BlEh+h4FnANaG
dgEa9ZvthD/wBVbfZ431AwF4vJyFcG6VXtULTvynAe1gsrpoOXNrJxG+9qy0EjLmao0F531WhM6E
gJjawlKGbT5IgGrqGjY3u4cud67GADSCMsy7gNg1ghiViIX851DAqk5TcFHXpYNeMVpKLHEWZUtf
xqj0wngv9N5O4yYcLJk6WgADpORbOnMGTDTT6WLkrsPmeQ3xlrVMUgLaJNBqzIT1GlhieuLZMdTa
Q9KgeffltemdLuxtxBtHER7nvc0JJ+0edJDBp0UpruaUfhPtFVn2abpThfNtVP4Oct2aBbjaXgGr
ac6j1myXWNvAYpYdfH/cd7VVBQlsFJWkdJybFtPQKDWMMa6fXKnJhxspRv4HyziaIOUAhlg8LoMe
3B0yveV1T6Q5MT74OEToJKHaAP6rwTjSCb/d+Rs5omYdRY+F93DYdZNwEpr6XRKpF9tBom38oO5P
ucPNZGYSK2/uNhZ4efYMadSKgpQ0EILTkokcPTkLP+TyllFW31Y5cxYfuHAlWyMs9kKeKgblDR01
KIxE6T3UDB0nibe1O102y8MlC/J40gZxIGjMSR4gxzT7K6H7AN5Cz8/sQrTWAF0u300hr/0PbBD/
7UCSqvFLMdzjVk346z8SsO1C5GrWDOVTNml6d0BAk6mTYskHAukeWixDcXIk8EggL7wEnGGZfPlI
1tvVakYd73Dj01oQ1xP5DmLBPVcUjbRS+MR9wZO9/1gieNd33NXwvVoqgdpsVPPXVxQ4kLRRtORs
H+LXwxoPYD5hJ8vCFme6tDe+tP6aQGzg+55YkEMtTI6wOhPLgJVuDHdmIuaqkKDeSWrr1MROuGJC
m1BgX3HfPdoU8Ho/p5M+jlzIrjYapPk8CHI3Gy8b441VR2nYTPR5rgVCLIdlLQJimHLIaduoQniO
B7OxHFeDAVjHUgFxkWLGTjLMRx6ls7/toV0RkyG01G1afyaUyqbC3poTX9y5KnZFF0wpwX0nuSAK
15dPz+mM+e9k/9pT7bY5ELRe9QS0B/dxxpyWVnyftpqV+GcZ2p258/LLfL79HPb+6EJpIFA+L37d
6+ohhtnarGTEgH1HdWLvrurd9oi4HxebH+q7/yDN4oBKiWAvITfPLwBdFh7/zJepm+ppR/EghZgr
oWdEYqZTxQ2WSksbgehSRgPOUNnqdG2/hRM+USlThrLaK/0RgGCu9rwm+R8terkpFyfJ+9+0whV+
Z7bhmxnEgBmZ3E4qbBlZxAWa5mxYQet9svR38ji//lBfF9EiPymJy5mVV/O4kLjDKXqY6FTV8ynh
Ql+AJvadt3ITTS6TH6pUvmx1cnrcH1wD3tFndfX60bxoU2t9oTeJz25P2g/1TsOPfhWNe2Ix7H42
V8PbZbv16oLgGBacEADRtz/Xv3YVOb1FEXXJ7SB+KLOuJvU+i6LkrHmlTcWSBixGgOoHWynUEx7j
p5gMh/SWSLgTbfuUNlhHonQAlESTXMpnQausHt5Jru6uFdZkjXwvMOC5MqKPjeaJYibMXYAfT2Gk
q/A79J1czouWPyDrJP+HVC9gVL3U5g/D3OdUDZZGphBp6ni7IjXS2zwKD+HhCz1Uox+8kKmk7BY2
mc0gWSPUDGIvWc4u6oOYRarEGxmleERKLhtcyuIf1HOegOlu/NxF3QBPoAcU/P4Uz/WJc3J67Z1+
cps1SNo6Re2vvZE6YijKvMOx01kYO3uKSYJ8FnP6KDj6g0R9foSyVWBuZ5e/MRvXdLOda3tA1q6T
z4pVhZ/7Ctgn0GzUeeWDPYyQtmYFLqUQXjxqcJ/600Iw9Hk5BTkr7q5ufAdCHmNhK0pK/CJy5qZX
xkXG1425aO7iWnaK+lTJORZDJvfa6byFL3/C0JcbxtKHepdXAGHBPseFyEyFOGCtn92Cd7hPeqvS
srzav2eQsT09+hS3vdNO77Us761yuDB2n4iJXsVcBF0FCxLUrhWrSOWtScwHUvzVWznDRb+87Auw
U2KaXShNPXZVxA0CIHf0uvTxgUPEcEURFHT9lom0ieaoCTUwlzUTwn5ajW/9tDBO+ORdFm5KxftH
hTBcesN3bGvu45m7MYqO7LPiBT3bwj/6AK2HESjjHvrVMZTh1p6yeMneoTBkZ/VBqVnuFDlOhhAR
X+2njDMQTw0lkdFyvOLsjOoA4iRg03hExqkpU3+WyLbIt+PvcyyMw1vysitRdZXp/iFO5XfIQ/F1
RDs3c0ghOx1N/oN5YrBhc3aWe0R+ylTS0U9ml+ynHhcfR3372dCEOIQXHNJhn1l2ELugO+orH9Ll
ePpjl+h7BUb4KprklCxL/+MeaX95+aNP0dnzSevBZ8eJuH1uQIpjHrSjqToGMcwDJ3ktnb4zTxX3
9DQU2jUEw7bR/UGgMF3cxu+XVh3FP2AxCvIKrxW5XsaOk8RKaM3p6iuL/blgv/255RRkRrKm2y6R
yXv96kIkcSvXN1TUBd7G8sWPNZd/m/oxB0sHUpCKSv5Ith1DeJK67M1OeAkoHn59DHyo0cnuO/Rc
Lz/qbJpU/t6W9Ixw8dB47H7/gN1auknk0Us9ikCcycnla1Z70VsyrGes75i0oZUf5muh2e9m6SWq
g5W17r+rKGxO7etOr2JrXdItMJmlEsPpHR2rEg3C7OhNWHgjM4bzzC2r6HzVrc73Mt/FF8Br71Fe
S4zWVJwult7jO+eWN5z0R9CUzuSPPnl6QedHIcKPehDaNamN5jlpowdeZSv47e6qjGenm0Xn+B7E
/QlAhERl6T1/FYgN6uhuUoGxCi5rEboDDk5CfGH+FdGbh1xoMizQyNkJc1P31ZW/tIAbH5JTV8sF
RqPmBOQJa/5v4m+2xCOT6pTmz1d9kh3FTtv9ySdizhZ5CbnY4tSrPvSFQuyurf7iHY+MMWb/tJAH
YZ+Sp5cGQzDvrYxyXWCxnI5EL4oAS03B3YZLk1bM2rwLQueqgwb7pvFmxSyEyGtn8wzEC+WtEfrk
9EAnWWCF8qCWrn8KGUgdfMx9a7lyqSFE3XFzk4WRhU3z4YtTDFeLmlkEZrP2xX+xlYZrmsTn8mlP
cNOgdEdsOLUGaTgSBi7V5d3568xzl0zQ0iR4twb+59j3kUWJOM6jEevAzFOjRmbFI7MD7PEAJq4n
ky0VfkOjE9/9uDSS9n9xty+/efLmqxG6pZz78vitUMOIfI9HuhCtMSR5qbMtrC0koSKWQerK2Opb
cYL3y+vKpGFD7wdty3/7rC+5PtKHa4jm4iy2R7M5auzHAG8f5ufurgZlJvNfbfhDrPpo+DngsOM+
xxQdSnAy4eQS1IL6BcPmC6Ex4TZN+skK3QWtmjoeXlddV46kiNcWlry89C7K/JUINzTrGIjJTXFQ
4dYszUbwIFSK7RSSBtfYWv6bUqZlxQOtI5lc5SSCJfT6iCMHapJoR77pUYZV0eTd+GnoFqKcfaMN
xsuWUDAyWXBdEOww1lCONRsDgv41kjk6B6Bmx1y19RLCNS7aVra/pUVgOeirvgC54YGeOwcur573
0BS+leZJJW48kp3/F1ujNKjOQI4+PB0N3w4OfKHOqoaPtBqbfx8XTBxjR9wH0imX5B29vXqKAISc
LnIghe6lyblVYt2SBcOZMTYfnil2Ar1Usa0XczoSwjGXxvmgspvwjqb3ge5a2Wfp6Z7e0DDMctgF
EhBT7QyyP5/RmDUnnO482ilrMJkztt27eTLK6yZHjxBfmYtXNOBJlGrYTkWhgtGPxswfarWnLs+I
yEjBeJl3szliC9l+1NXlH8gFR4hufGAdJLOZLiohBRIIZbA31mpux9HVICI2ZsTSWWzrQq8OOOyp
1IyfgZoSai7nYEI3NXczgyNM4Oxpn8HM/kKNdSrV9jss5aGGfcC6va4bYNVpNnjKgZ1IMtJl2ehb
9O471y+Ed2vQxx/pCG4H1RiwogZY2J1mgmcD4d6uQsCvdTEKNsiTBoZzRMe75BnSxJ84KOYP3DCK
FKo66RwZagTvhm/FeEJtMQpUymOcFRvqeSlf/7oJnDv1Sk60PeaDDRWLDTHZE16Z4FX2G98nVTgI
0MlZA76HXvqIsIoOAp6vvbA9aFiaDzB/5kCWY9SQu74u8juD+t5pRrvSCtX9Xu0G13YXpuL9hmdH
PzCD4WmV05UhDHlIuc28IlWGg8vcrQSNzj7dE/HKlnBQc6idkxUPdAPoSoDmMnzqz2z6l7HzoLbg
tn2Y4Gk7JrBHYmRwfu/6e+K/n0M8thXxSEPCd69R28VNPzQ5Q6/n5XG6fJqPYvzmh+0qc2+e3lh3
Yye+KTezMTBokEzETEQJ+2Vu1H8UU2EVfzN/Tn/mC5/UlcYEWmI7nyoqXwSLfO36JFXWUjFaj00e
hV0EnsZ86HNv5L1g+5sq4JHCH25X8PNUOW5l6VOaoubNH4XT2UJ6dWYCtTbiNSs7e3hl94dtHQM3
Z8lLSfxwspYAAdEr+m0DVrHVHILXi6Q+FiJlkJztV4aTHtk0PrbaYInXoYY+Y2s9KPxq98E8LTGj
iRBtDaneYXMwpF2+YIo4Da6jNs3sWhC/2W/NEJSJIE2UGf+/QJsES6rNqESm2e9J2VUwoQ4etznh
DAsndBvjjfBZnnxFtBMezVJkF6uMvwN/Q6ggXiSh/uMKGl4Gk3iTICOzJlbAKJwOo3V1FHrTdJep
pP/rRuhp4S96OgebMjeMut+6+FhzYuP0SmC4apYGs7ZZwO14L/9NUJ02xEOmEeiWq7J2xvL8OH2j
LqbNAGGQ8zW0mCVLY6Xy1YWFbwVRPslUmaHGdCNfg7C+My9d35AqOGlhMbHoh5R4NbWgKiduUfFh
0iGMugwo9A2LS5Pa5sI28XgRonJOHO4vq7mkA+Fqc8Af9dM4S+ILUR0JQzOF91kbaGPYNLk5Bdme
EAXkZFxqUW9GdCgJ4ieTcB0OIFGeYWGT+MVgxHT69QXYTXrO7IDv3GfcbvYxsAjiGz6+CYPeHF04
Ppgsp9q3yyQEWMdxHDx8NbwOnKc7AsuloenbQzMQSThD34Hy0k4+YdxjxaiMnOXkWCf8l8uBR7dy
jjsN2ZwAireYNYKeYBKpCKQbHfU4WwbTWIX9fpxRep2YePaY9bKbzaZEhHY0ceBSDmRPbwSG+zFT
b0AOTqqkkCl4ixraYxkZlO8vUvT8tezuNa5Kv6+uHeUNaefJh/4WkTfS6hUdF1PKVWTIHIleYgmU
lZU+ylwZdxRsG8IN9Q9yqUi5FSygBSNWkU9wZcllOqvDkcNJKbm7mz/rK05pBAWMTLzUsEc7mdSa
44aPyfAGYRdTBq893knGGNhuJFmyT+BuRWum4AePofVnHSeuIifiagYgHbKkic8ZMJnMSJtNDZ2M
N4YSILRx4vOUvGdDsnfsH/sH3RZdPy1S9DaHcSDo08e+6PKbvw/qO6XyHBAtVMEvc8yz7ArcYqhU
jIkanB8vn4yHZsAi7/oxp7sx7+wMoEkZnzD7IaEJTyKGqwBXd7XZWy1hzhmMM+/FT7H3TH95gxXQ
ZWkcGYi1qvdUGoSpi0jDL2jVWBi88byK9raauG/Iew4O2mxV18HTx7jAqBIxPjW2bupfUd9I7aIL
Cc6Pj8YdJXi/S5sduak80x4hQY7HC4UTigyAhQWh+4gK7tj66e/AO8YlzRe2wiCBcHT3v0PEv7Oh
gLXOAu7gM1Gnak+QxSQKAK3HdN4vlaplsdLVAmkwCQeJWVfD++2bnP+xlyNjbym20oCzGNTxBcFa
X7azsanElA+CUuG+/0ZTGkYMrAL+0fIzIgs77Xkp/7zSNwU4/WQYCWJ9twZjEdFw1YXWwYU0pPcJ
t0hhaUpgwq087okY92+A4wZ+ub79vdPsDa4uMmAN9nhldsK3mH0hEQxmgG9KoB8fxqC5TQ7hQfo3
aV/Dlf5b18DPwavMUzoIiLImhTzzvm/0a/8eR707S6A0M119bhnaVfHxi1dK4Sprvj1qzaDJJc93
DoTS0fICCoBsraaGedneba8vG1u44lc5vJLAB/5ednvPHnxmKpAP5w45N9hicEzoDf+Zy2a2x8rr
sEWFFlBpEIbgRc7mZUuAN6v84WasGZQnlYQcsUem+1SNnmvuD23mwojReuq4QPD0/9fEjR+3UpIQ
srwTnwbWO8cq3A4aE/+pAsse4gQ9XTHM55fTLcEVI13pIkIcDXYnwU/7LNsHE8Tz/lzhDLuLCbAP
YvwC5HyUlipVNzviNB+MmByhfx+5dPmkCUahIYZxYhkxW9I78aSHCH8Q8awVvLpevNVk4pMY+pKZ
rVd4UOHS+0EQY16NoiGdm0Cp0YXUTYDebhVBMqlHaJQAwGX6jkYXadTDMv528TLyc7L+BabqQFm9
AIxoCtcvlwn1irmRTYg0ndlOMbo6RlV6HVRVEGsa7ijUMJlBEFY3JyrevJMEbisASDU9mvZ6VIj3
SjylytG8KYTV+HZBM4ohIiIxqn7mJFWp4D/Pm/mYpyoWDvL3YW5R2QQzrhlioYwjEhRX/n0izTF9
sqdG4QV/dAxYBLvXzH4ZR1JaF/pGKPfcD/q5HTCoKhM77O4MT7454F2ErIg+vLXr62FQ1KE9McNB
4f10GbiPbJZEVRVzrOlfza1r8Lws8rhJ+SaUaj1nCOtG+GTyobCz7klkt90OBQhJ0YLadaROOTnK
uMM+lWf/5IQW9G80fwgwAL8dBRaFwbrBb6UQsMFsmHBbb1c3xGsKTB9o/EHi5L/iWZG2slhChblH
hj+EzhM2re7+0Y55/hwOGJKatZSd5AeKsawae1gZGS1r152UO/duPYB2qOTfPNCuvnvfHOm3u7au
Xxf+NX2ASoYomIVRPSvFgPlD2FLsamVd+h71EXnG95f0lzYUcsBUbN/O7YgG7LHohsPDre+JjnVC
r3zBj5g6HEFn8ZAHdxmvPZ7BT54KvNKbDAoWBqVscy9w74jgHKoLKZIiryund0O9zTk0UgmPjNL/
6H66g2LUGQNYqJd8DmHciVvVvvlWqQrCztUtstLHSzfz9xBJAaFUVT+WEqvUb3AccERoS+XO36iO
MGswP4VQ1NeiSWqyc/T40lTtZjaPkA21D/xK5y5lYC/7wIrN3iRkUCUq1vz4VEsY6wZftwak9zva
JgHpDnWnKHrKApgroGXobwZPkG2w/w8OQLiRHMGBLqJlZ/fLSbNwG4yRGHBHTRQKx+pu9F6sj4Mh
Fv0V4aGABttsMagEOUs9Tm2UiD8ICDhVMBkZikiaeHHwsPjsZTqUAMGsnvok+S3Y7k/WIcZxkA+w
6s7aENW6+ymOyAjVKs96F9rON7XeUD2Zc/PN12Bv5aSLI7N3S480f4dvFrZoP4Hw8osp8P0iCr6F
vafvKxk+8A95hXFp8ivtKlN0jaJF9k/6/w6sK8Rfa5k84CFqUD5Bl/peKx6RrMOCUdodD/HvFFJs
ML2Ay4HbyEmDaYOGyZ45t6xPceUWs3SBVxIMbE/he+T23hdvwrcDUp+eB+JN4T8K+s64+SUt2SkS
dN6Ytv9zIVjCHBKX4Nc6ZJJzUq9weY3iKbMG8+UDD6MzB08gKulFb7hzvA+IB5iq7NyiMV7kIfSs
K1EmMOLqF05A3rL2cMAwTaPqkByaeSaYJGZMIJVdpAKMjZnCUg5a7NyUfJvDZy+SQ7yfZcs43tS2
gufCjvmSN7KHH49vAfMoecSsP7iPlPH40oAgK4cP7MOvnfx00o7Cxbgfs+G090dNRPZdCeA882j8
kJT+aiELd0D2vx5uDcb12eyvp/3FSEwgKYxnkyOmbtbUFG/wPHPst7ZmUc4caPeDQjPHNAbQvCHq
4d0Zm6Wl4TlUodOKb6Fo0ujXxc/r+hQfr+R90Gxd61ldZYbz5LSEw7r7WoPZf8ZbDA/E1pP6ApTg
Huo40zupsM+nka8PG/wnTnz8H99VJbIexOPUs9BTf5QAFIbWozXYDYYR/LwuDvqLzXRu6lXbZcA3
YEG87XUfgwwcoN5klkm1got5S95ISXDKet8A4MNMRpwG2ZqsBh+KefOfBVLTFHezYxTfDF1sx3pB
nQME80xqvZauBkiiwz8509RjhQV5P1MepsUrlcwdkn2dYwBRd6OkDO5Tt33Gat+3Ra6BJg5risdd
MfQaLyrBCtsxtSDEScdwzjdcsZIdW8dLQ5zuvyiAm+h3zlr9PxNRlLrGMLAEGXEd+o3Cpbo3l0AT
Lj8l1F96QfYzgbgnNSh6Ccy5Jow5brgG7kVIqs+UlUQMlI/b4JRHOVKn1tIbyfyqKYNNwIxHpB1K
X9JIMXmtg1aW8L4x9FZ0VMPOd63Ql7S+TYfYreqL/EV5hGExx3pPN6+H2N9qup9sXIzpquwkiNVI
OyNjug2wa0V7gOhRSfkT53ntQa+ClNaUQCbtfuh6hjgutDsAhz5JQr2yKWUX+SPxcVPfBoWU8AWz
oM2jNbuBuXA51yh7hw3OofmbN63qRDgnwerWAzvSkAYBiiU8cFyvsnRp82UEO3ucxO9R7IatvHSD
OxjYzFpWYWJoj2MkFdUDVvpwF02zt3MSCxeJMUdgnPPHEWznmzDHyyyZ4jdKL+vdTjdL/TxFRrNt
+8N6U+obKzR/Wliz6b7D78aWEMtSpe43ER68MTkqQrinEzTb+5tx8R4TKMJpjYPzRq0UG97shwLl
sRw9Ab/qBG+iONgmphHNNjGSzIobsiJDFdRgN+m7GKPI3ckm0shQBqsPIT7D21PzdULDOO2xQQN7
c9dzg1czkWzy2Kf/2h//eHuDBPwHnwjsBIqVwbr0Lz5n2TfAagMcUMSA9b78sVKWRajttThcqmn8
i/u3a+9oJ9oOfIDRN26May4stRjhW5+7f1t2vg5A/6Pdfszp9ABYnqfwtp46D7ZUyrsMDd004e/E
9rCxhiwDj5mrLCuvXomziL849+vgVjxak33LJvTvQI5KBZ8HZ9UEgIAX/kFiHL0+qjAAInxDEcGl
UxpWcmg/N/VCby4+ms2Obpn0uw8jlI+xDMxMl5ZqlDRxF+SQqzePYEITR5HCk9YuFtIuYAVMFs24
0PcfK9mwrE6FuBKU7z9svqZcQSqi6y3K8wgSjMZ+LdnWrSz7sT23KRJ6vYZtfdpnggor3xCud5cs
e2Kr7Ii9VZcj3rNtjytDqU5n8hEwV1ba4gWMdb0VQXyj/+Zgb7ou5VjMKE2weT0nB+r2rYgfRjtQ
SV/NjZ/Bvxed5UarB5L1izZrok3knkq/43ZMKaKEKqSiIS7iB1TC26AJkprBFSKLnu2co9koPA6U
8C80wDsCwVCKNwNh0WAa2EPvUY1LmOEjBal2A6NpTMrqP7E9O8QI0xZfoyaiPN/sQTTN8XNCmYeC
S7e/znJBtKfs4HaHs1T9i0ldbyNmPHrrwlXpBBj4voKKBMiolQJxxTbPU/EUu6mdlKe6nWqSM4Sy
vwor5os87lNUHpbCbcPgLfbbkTkfX7+Vmfm2iWI0n2B3SBngA0APiax2EM6T2/IPA7/Y5qu0EjxB
yHDDEqD/UeqwnMWi1HvMkdgGLRJwxuDGq2hKCz3OnbevJ6A0c0n25R3kY4QQHW0zmT82mjXcxMAH
D6/BluiagP1ntf1Ae+ZEbXOulnOMJ8iPuK0bwr4bDFkZnlTZIgitgGl3LfSXiMlUKb6VwGihvr5L
LPf//62j4v04lzc49ClVR9G8WyY5cVKS6Zv3tUWRiEgL+3MSJhOa0VnOlJLWmcpmrGidjMLwwn9s
NjJ8RxM72M8F68goTE1kSp8YRPCff8dTaVwINudkx87uLAxf2U+tRwKAJ7KmjuwHbfy7jCqIUaKE
qZT5Eof+wuADoerCt2BfeZjnMwwzuezikW2/asVerXjTFlS45clBvTr7e/LxTtsQpyWdA2FJSsJj
2rqcgNc3NWbkLAT0MomTSMogUav7+FMRlVWG69roLMu0w8GbQsTxI9MWNvQ5rTjrwWY8su/r5Gsk
SYkF6jnD/YqMO3zbGxtE3Z8tXqc/uPK73UTRyVbz23OedlNAH5xXWkc1Lib/QzWXaGWjELQLLw4w
d1q0u8Gu173hCj+AMzPY4twHPAS8GZ8DBvp65oALb3OwrpMR5tE8av1u8cJvTVcNgzH6UAt/6/eO
1jkuV/9sCxx+fpRryQZG2M2LdeP3ZB1XkrLyYILwo/lIKZxYHYigEKI/KIXedf6mhlSyxJZcBrlC
RSrw6QfR7qpfp8bpHS9eu1/4nkK00iYaOM8psksAQeQ2ZnZK8JkY0XpzOTew8WRxCrDpbpop7V17
+VLAhx7ZJCRwyNPW3vi3T2LUweNLuhUdCvxoAM/dAZITr7pCINxFuH3aSsxND3Y0U35Fy6rvs5r7
zwHl0Y5PSQe4wr5cuaHjoPnhKqpiPvP2cIsqmQ+QrgYiqcGuf9KqMajE7ACDTqVlIWHUfcf7F0Qn
V3tQVDrIzgHsDqUWtWCATPPIHERTjTtI4BnxSv6dAb9StF22+SkDXHqzQcfha0bSeuNQR0XlZroL
5UuTOoWMG95pNzaBpPcvkQdm4eC7x4BNKtahVQJGywqJF1w14cOBut7MRyV6Ox25OWDtJn+EZXGu
CapPUrV4Xc3NirzsuxLit03kyDiveoXlgD7DOpec99ARELYPAH3aeLXB6l/y+aeAC7DCrsnM7pLf
COwDR6M9F2IkkiTO7EWOoMqqg0SBcztjQ2cYLoLaoAtzlOxHgSAwQPxOI9V+ouo97J/2dF+fOWR8
3wXYIwonv9k7gVjesrUOCsRtYzzkvw4XDSWW8FxcwlETc8umy/EP04bEKiUMyzDK5XRFwliWjFW3
mcoUTBkOEOqVB9D/BpdAhG9dFOFGU62tiQq9AkpWo/m/DBPKP5ToGqpYBIr20zAGlTVsxkMbsVGt
gweGHd15CZCViEiwmJjYCSe7H1+1L0wn1tyuoXv9n/fk8DcLZt0JP0oUqBC+2E2mzKAH/0kcPtoo
26Rg15dDM8bIzIyMeXqTQuEKgmgqDdS8IZlOk6R9t4daVvSYjWkY6ZV9Dwaq9DSdwzovzE0XrWsm
2qhWJOILvApnv3TXr1VorzKnjo2zVCOXa4OwTd3zLrwqjvTAv/RgMWlm6v9Bg/k4aiA1uqBYqDfP
NgS/EngSkAMrJuxvsqcreU0qLZusSz/7Bh4DFNJzJQot7Ga9u+Y4jZqQd5iPTSBldUA3Dqemf2HW
F1VcgjL7Ks7+6QefBi7weaijNM7Zl6Y2QqAF7KwANc3UfR9kEOoVVDz3SBAn9773YY2jRovFKvzr
NjvELmd8KJKmauwCsc9+Uvy/48LTumBMw4l7Vgw5mzsieHw9VvWRyN1tER7tzw5taI2dCw601b3L
pXsrj4M39zT5HKxcvrJRW6Ip6YiaKQxn//qCzY2ZjQp3XNxupkmGzZBwcsTFeyP40mLqfPbMB+z2
wZxKxdSdZ1LI2psOJqsVahBLN1xTmc/hv/DTu50bGjnPiXYeWNKeANxQy6t9hsHq9e9rIqkzRC+i
Vz2kLS5x3P55F4QW7MiGSaADaNAsILfYg30WjHZnO9DiT52OQ3Id5hDCIwxW/8LGlEETnnXOkYY9
n8LMqKtwIiwcppkVR6x2sw7xbMt/yihaKqVdDiRkMBhtd9jUI9OydAEbp4i9ybFni6pKuLEGXv6a
pSfts3TFWpWCutc/tN1a8wDrhabWUx6vt9xntaDUS1JkbnbMFpZ0kOXQuku5K90xF/oPeJOL2xYe
y7mgN2yJbBwoOyuTZWi1xEDAPYIGI0kW1XYrWE11p7x/nycJ5yh+rF2Cpwl61sJOHoyQqwCcPOvZ
60SGFyag3ORIXvQ9x9caVDLQhSK9mWiZiF3/9YdYR0faHMKPKOmU//jv6eV2uf1/i1oWtHxXPkL1
3BGBtPR4gFJrC+xaw6+T7qbd6IDsqlcJn5l42BWXSA8146eZtBGkIt9g4fbmZO0KGFuImMGph4rV
UCrvm4QxqYTUqEsOY+62bZtWCI/s/9aNdv3XMyH1Qp7qGsAuXtCZ8c3e1KMZCWwFKndYnais+T8h
s4n0N1zqmKTg7+vkBCiYL/BcRhfUiEAoNia4cjxoLd+FFWiJ3G7dngPOjtQaOOGd5GTHjouFBsQj
N7K09CeJnQUg66k9W+kHIrxnuhyYOjJQxsFlIOvebbrfi3+wteWV0fDRnSmgxeuMjEBF8XLTuF76
zQyv+/kysDj0SkSfGiwT4MYIwzGk5rhZkhUisQVhNrOvNO44mXw58ub3E1B1D8tn0C6hXL/0CjnF
ptcdhRAMV9++2dSSyXvuwnc4v2Y7o4IsgAHWL/f0p7djVQ5Z0hxoFjbyJgMxpYuRnWXApiAZGnIT
Kkq2nAgZPoFhr7VQVQNObortBxE2mSHC6RDPse4l7G0fNG7EmvKRP8qSAztkrFrp/TV59IXQ8aP2
oLDUMZ7Mesa1nwMyHP/OXCku0IcWHBFCQyahH3+HJ7CsWr3xkxU3rXvJKD1rPKdeEDEn3NDJaJ1k
c0i6OjLtOOWF2wJ/8x7MUxYRhs9OqNOuarqzm58WqWGgc4znB3KdyRcQavJQP7mvBEOzXOxTDmef
pOHcRcyo7+28OfCn9q1Jg9y+6Zo3h0ojXen1XarkQ3OE30i51WfxsVobonI1Iaa9c80FncrE4aVi
n2y8+/R0CriWrdDKAC5qUupfxcuSGUxtKdK4jxDA5JFgrJkBU76LhpULlehgHTNvg+bZUoOAQ7B3
dkKWzrQbb2nZ5kCVcrmP21+05DnljRlNbDIRlYxwMDic4fsxFaq/2LqqtJX9GRJtAmYnNMnzkTKN
t2av4yc4e+UNiELaYxAqAOfJvB1UG5MW1uFl4GrRlYt3trsRGb2M4xdFe5YVGU/A5gslflooC13n
m3Ll+tLqZZpMx/4A0sJJl2BxkfZre3hcAFqb9Yzik4+t4mABuKmdkPyL0MscqWz2K8omXhBsK4hR
1KBEja1FezK+0L9kYguJqCXeinRqhHTtcMzrwluTHEaD3dzLVQx90vwvH5n8D4niYfb4KTmvjSX0
xe0IK5IEUrqC6RgBzezp1n74nwd3CkYkuA43/Nyky8O11mJNFV0udi9Y9kJKx92t/x3VKkJzVLBB
FKm9JGCQeqcFxIpqxU8TJx/Yj46UpzLtlGViUu3Y6AQdSqENVZao+ujEFezKp12A9kNXcLInpfff
B3Eu6xUglDd9CjbYGDhSK5NpcRdDwvTtK/ne9wL51Gao4I+BZEF51ygxkxKCb9ETDZPOEm2AMS6X
QzsSO3Ei+mfbq7qoopjgFbZMvYYQYAboFeYQONKDwo5GpPMx2Er3f4BlNfzzlFKDVfoEkEwkU4m+
+bgZSGqZCLjU8Ds/fX/K02HknmSSzOeSmv5RcF90DNQrxTkGUw1nODK6/ix7JV2maV1qIneYrxfN
qPJoN3QSaJ8ivlwEIMQH4S1rYledr17wVqVtdNDsZMqVSffDU0tL3WzYnfJd/K0C0LHMPxicPyQ6
xFkm8g8m7lFCi3trr+cYBnNLcKmyvpgU0No8ZwLdAtNWPBGspKnLVms0QNUQ0HNX6qsJ4R/qQdKC
VtjFOdwpTN5bdTKHK8Wr7l0CSUcPCcvw91/MQgxr462+6M4nzt6g4PfbfYd7BZqvXAUmQe2tpKBg
oRBTPJnw+u+obi2Y1d4ZRGMVZWVM+zkH3U2WB6ARK5CaEQLUPf0mnFmo7BUx6jT4hUzCyftPeBk/
IJZHPchRW81AZzIIZFaAqaVHMWJjzTapepWLD5zjU7wb+JDqQ3a2lJExTUWjbBghg5MgWtJkb6Ts
EA/FPCAf6Yw2Y+DH7n1dVZbRC0w3vezBwPWW5Z6ompnMdN2fRfAAjQaf8HZ01tTZmm1VgjnLBMyV
Y1DcXk7WEDqExPXd0tGKU8qIP2+2W7NwskrW4x+z/B3Bj+ul0DaHUelzyJIJ5zIst4XcVHL46r1y
ZbfnI+vCuulEuzX2+xvhk6RNLs/SZmmSMDA2/iU54xgH0kpxZdaoy5//FFQ5t1lSqqlWxwkpZDaf
X05FIwfaOSHAPmFe1q8I19juM9H+Z0gSyith3vWkgyhC6AZi1GC3cWBGyz6e6XV1ZCXIRgCcfRnR
HQchtfzF5VgdItlU8OXmPPoxOa2CtSnZkauyXUkVkaOMbxLzIqkxmCaZT1U5X9ZrT0vdoNyNGao8
LtFtTkC7XLkyDHPmRTDvtUpw93DIrraC08UKMNrEYfOg5Pl0k1U3oT9Qbw+/DIwdw6zq/uqkN95W
6/+98Lwr7wC75hDBXvepfnrb3lLjt2hMA89woDXsaQ0BL8HX4K/tWGZtAUoZiFmPg9HvEIxx08uB
VHbVV6HpNX+RCwbWE5o4j6iVOoeI73uscEWE0SZQL8WduCPRqIiIszpYGK3DNSjR16eTy0fbKOXq
MPVbM+ciZs747VcXXJN0vUUWNNal+OyZH9eL3rzsPx6iAVaW6dEZWJ5jxmgMOcEHxoFaeibZdKwC
KJ+1qRhlA4EuWJk8zQde/4auvLbhif1vqTUEn+L9sIu3WVaZexVHbdAWdDlz7sHqLGj9NdJPqxe1
29L1N40i55Ieapp1uoVRP6q9oUhaVcAArRphcjybPbhShqM0o2/FBv1l7fenoGrkUFTafMbY+O+b
NHGI6D9t/zfnPlOsQWBOkr8T4sGiQy6XD+zE+h2yI5zdMF3Ma/wb1BOfFUL7S7nwxCLag33N2Okq
vjxeC0ouk6I0UcV7qJOsXwwKys86f1o54R2VFIzChx151YCmvjRi4XJp1FDM6DGcF1rE6Rp+Mwlj
RYXrVKE3Tw8epEcsczoBeoxzIW8Eht+1Cxs69RlgWCuFaLm57S15Dck6iH10b8Obzv2ltwJVGk3r
wVJvMvHDY/rhV3cNMpvLYlCqogRgzGY0JR7nYYinU8HXmpbTyINjCoYBvfz/mTPESDmX0g0e6xmE
P7WJzR81De0rdg1D4OqtUmzy2YK0N4EiTPF8FGYCGmU2AJMCn/ujvIBlOn1msYua5vgB+mjdEzSU
RXaiNzeqq7cJClknqgnNgpSs6rqTcQI9irf3D7mAr/UDBT7AHAK1gLUU/Q/yGt1jSP4xaQtzxUkW
ZEfrY+tjSAqosyQVeiTG9OkAeASMzJEkhT8nNMDIY1FpdXPj5nLxel/Gk5Zocepehxm1YuO0Yhe7
luQT5HifOEk7YMZC8qnAcx/etfg3l53YhNrSkrX5TdggHiW62Cy9y9IW04vyc6SO3RIjvLGq0Vwf
eQVpaqFXfH5Iqmuovl0LGnzppGYMDFtwraSQDNvV/E+dZnIPFB0ZnDOw2XC/3UrW8zAMeGpyTEYu
Rk0JeRAklIVNdDlZlYtTU59WvxgRuIWqfQUEGpE0cRY1ySroZmjgZFqxVIyFl7Vdizbm6QF6+UkM
F2iwZG8PRLxr2P0dwUifQ+LBgS1gGlv3aMapebKlCeU9Ue0cJwFNsJTgbkZ3nCZUr/o3hM2N5FU8
CIkakfY2ItSbnM3cVBJGkrWBHCr4t+OX/W49BQUabIT/s1LhTpOwgb3P53ONJ5pC7mdceRGhxo/C
IwOtYoQERAD1v1q+yRQpYQAKhoyThihum1hyfL9n4NbdZZIvh6/xJEIFuVjhZ5D6+x0whg8lOwYZ
0/7WB89KlLC5vqJzpXI3qtS0LpPG/4ECSSnCttJxIuq2Q2Hjdf9ctCEATgTPPvVZEq6Phhz9c39k
7iij52uWK6kXfaIuYuLqZxdH0K8wGZioc/SOOTpsVQGETyRiUIzttTSD1rlFujqB+94jNHQE3mu8
vZePW7y4qQHiqLEk6/v+vgNMo4pK8XL85YKmkbL1T4XWDTgyLRaJ6pEe3Dq6WEm8wrNlfSdtFeme
cGsv9yYnT0hhB+gb4uLLmtjG9cn1FjcJVtaVcs1bWG07f3iKxlrGXMzlGvskfNRaxyhrgP24voLl
ageU7dAEhTCRymckL0V6vA3rEdcKpZtrJcFvNBPcTSh8dnWBPX3ibJOKcBKkPH2wzPoKWeufpt0m
f97n/Sr0pvWKZFb16PYgnuN/tiXnt/Z4ddJ1YbpfQfW2OwHMXEMurhnXiHXiB94Xh2CL9Eq0eDQZ
zBPG8CRPcqzSbpZOA6RhFX2Edq2IRzT2Cb7ySZ/lkzrFfnFN4qJ6EjcI98EYVbqpBumMhL+lcS2z
4GyyYI+cC0OhmILD/MXEBdB/btHpqNjH+8wIq/DFCshz6AMsH+CLhfuJ3eX476AkRHL4VP+74ha5
htduLu7jm5uPVLjJS6DvINor1ISqJK5+N+2QVxQa+LayKSwiyhovOMObmvW7Y8+ndRHCgI4X5XMb
eY0y6e9UtjHt7+TLEiyr8CvFpKNOE2uMPPD4EFkcqMBeg4ZYUA53fPQs3B3y+TLhLakBxjI76W+w
CKQ0/cXrqSICWPYlc049e1HBwcp+awt19+8OMZSG4AQMiT4urO2eq9X6kLnSqY9ov5MVh09jz/7S
BRTG7EA0MnEXKqAO/zcUfaEiu1znpKNB30eE5tgK2zMGwLD9jLR2ia5JyNj7bdGcp/fdWf43WSp9
ebTI9NVDVaEgHvFhc38uzw3dDFXb+I8vK5KXdvN8l80sCjMs8p8X1mTmRWs0Y2QMifgCARAxi5Uv
SGoUojgzQUfu2rUufYyAntzaRMsGINpYukfygDAyvn09S4xzkVKbwC4lHbUqFHs07Vu710EYSMNY
NCDjWH6ia8hPyucdzAQbpaw8eVn5Slslwivncgdc/DTEIqIsKANOlsqYwKHhgcAlArwnzSFWslZU
FlJwW28yIwcRxbrSzhTUysSuL5F3tXTbgxIsShkCAmxwFrgXuacp6F1JzZ0Vlv7daK+8+3KhAK2V
VQ/zmUSd/XlPNN/Z290v9sy2HtU0BKSnXXorqhW90GafJdRiUzf+ZKMrP+AOuiK+CS1f9S/Ay0VK
86fMq4xOgsBb0V0AacL4SoBTifdOZqCwx9OYFbrKw4WApYSwySyod7dzaH7HJRY2pJcLuLJisL6W
5DRWkCLSwhjZv+ROWfjTh88J+ZQs5XEtSk71kl4jYrG0Oi7ftSkl1eJrjdhzJ1ysybFdIouy1j2p
GdVW2995bfP6N3MuBDz/6l50bAEhKmawxtVPVHt9teagR9ahNWRBccA771hO9zcG9VD8hUS9H5tG
a5Hk/IWF5uKkpC1hLKiFgEzfay7TWa2lH090M3pkM7wWq680dVCAnKXvFTqIpG3sZygYIf/NPwEM
pAhYCnBWK7owzyhV3MoPnGHRoTPqTPrU7K150j75NaDCFNYnKMkMzfeFi94eNwWBUtr+d8bfBdFl
iyfS0wbmiUCDUGWfekjY7IVl27nFxCACKhGGyPFosv8Oo+ohxdXKIucB/JM/IiPi0rH7qa1kBvmd
om6FBPB3cQT6LbIx1oI0h2WYdY7Yd4IUyVKOKXBZkWS7Nvm6TaL/SyjlHWJCBQT6jhkA5OuKrjh9
KLIXCNIIhcSLivLGhxe4P7hXgTa57+AUWZ2XfIpnSP6qwSKl6WEaIvN7QC0TUaOaDOSTNpbqG6oW
JXMie13xf6VFFPb9gheRkSohmMj40MM62eJwHefHh9Ji/sl6fJjSc3bqTCZ4pioolem3Xz9g2hBb
IV9beT4uvuenQMgXIHGvC9W/6VZ+QDVEbLyfUAITtH/a48yE0nq0bSgjcbuMSCCk+G2MyiQ+Rjtx
kLK52Z1lGT3r094u57ugftMcF2V8lD4s28IFBspSutH1aGXEMUfJd/tAfdbP1YZv1bOSVsCj0i0S
qthmpKoPaAalTyxDwF2/AJi2f39iUcR6nJT8zsyHakHEWXXlUXJ20RFabM0Ex9/yLBaB27GpMw5j
Cyg6z2ekZS05EOIuS1nadTf7FCGbIuY0GKvTB9jU2tbWdyXI/looTFoUCf9YqaMcs+hPk9bROiMU
q0LImziA2hFbI9qu6OsPLUCSJPVEkZxijI5S6AYHKAxPsuXOXMNFuObL2WrMcNTzreaSW7a1iO7T
eFq/tjAze+maQqPEfF0UxE2sHBxSts9EuC4WOlwlgRsBjkGlUUkDzibPIUCjH6NZfYjjbJkbD9c1
msCcJ2fBZC52HkapkbdNjfonWbI6JKLhIac1eLcEF33fBF2rbVRSHYiDzWvMajFamb2us6SMuE6K
TulaImpEQoNQalZGuqJ4qFoJ9q21h/D+ETtYIyk/DRN+jXN87FhzRYwS9YxCiZ/Ci6k6O9IluEvC
B3lFEyYFSL9jYDZky8AnxNaHgP3LPcrQICVMQ1gLTIjU6NWwKJV1+mLYoK2Rrr49TgJ+KG7I4Yfx
XMXO5mLaQpwynwgTH3xwubTU0tSW33Pin0J+v8g92XZIqI/DmkjNunC0oM3kydUV3w1vhKQaCbkd
MmLRcBUBCLKau9u5u7myrOlYhedYZ+zYOLkGzDwyPMoHj5h/aUnOJoAoigD6keNrYY7jilLJTdzc
WCZKAh2kjmC5QFDvN5bEQiALYrX80QWUV/IdmmQ+3CgzPXMdo+j9bqTySsu48DhD7x3BCUtuwZ/s
xVH+4/1ZJZGvdW3LGP3rYuUwic9m00VWZFzU+yYAXRiO5AXyW1EkgrO+49q5woITX3V9DSPz489V
bAuWO9dEI3etF48RK2SAIH+wfXjmYYori3R4/mAFQtoDuO8OmRF6RZ8S2PozrF2tBDh8BXOdXMa+
syoQj5oJD9I3DbSR/tQuM6HaVddWVIaqZfFEhEmXxg6wvINee2fCcA8yCg5QR/H1FUn9GPBbQVhN
Aa0a3yNEeYM8v4a8CF+baSOgd4VF0MWS47eP2lw7JlLn7mHiDI9lDD5m774rNTASFmOCiI45o24H
kER8N4nMb03GOZGmMI2LmQO52XhpX4yj+hnHjoLfIl7gUFjU+g0QsTxyDQHZgnohE39peXEZxB75
LzoLstT4XftVKnWZmh4EO/u7C1dYybzDgTyRvCzCjaF3b6EzIR2Lp/pb1uVeoTD3q4fXV+sfdQN6
XHN4M76IEkDww7zQZSocUFc4x1qyK5cukbnf5k/k2SX3hGHxpoDwilF0DDjEbg+p78xz7ImlEgJl
XwQ9D9s5yFEiYGjwYKVcm8DX77SvRxp/9Um89vnUDPPz/pPk6oWs95Gyl4lecewmCTSpBU+bxHl9
tXEJiv63TE5j1W4weK6t+nIoSAs9k1G8TKtsU8h4P+0tYIAGjRqGc5KvZ9bo7fhPgX/Zx6MOrdPq
7iPaLSeOKNq97VJnmqoNqXa2Hr7G73FlEGG7O8HdY161gCKcZbrgvHiQEypcBH0mLo33WPnWQfHd
N4zeQvFFbsqeeKcZ2ulMj5Wpyfx/Nw3kRKMot547044X950ZCVnLWLTSEBE5VadggGg3ttbgn0RQ
mmK7DT4n9Ubdvrib+uNjHW3EUrR4fyucOHv8eOSNo3VVvErhqTCF7oPeV8JTkMgJ04mF534Volwx
vD4TMaKhSpzTpB3POdLK/6KYwPttzLn7l+XAvyUBfYqphSpC3hjDDZ8m76R8pCt1ssXNyrfq0vWx
TzyyjIK6ObiUrLLltzxfoktbhbAsUUTxEXDPOdV1XIWrgmKEwchsjTJNg/Im24VdgtdzpcmXmTfM
EVUXgDtDaSdQ49q6QB0tQj2fpx9Lu3RnGazJjz3OsRzsHfDc7VgyHkq9gqsoLz+FQ+4b3Tp9iVtC
WOs+FP/SAXnY8Qj6wJdFDwkYhAeqOcqLrVvQgTVRAaenDQnAlK80GV8RpukML+xdBoUH2ZjzU7J0
QDRLvKLr6fhQKlZzNDNideewFHbQcqumZ1PbvgaibCWUjRS+h7rt0X1KYitAGgOVRhtNqWArTX5t
dcd7bBH+HqrW+XZT6U1l04qUQjesD7Lj25vKIXy6mymIQZ/sIL/WoG4AgNRacVMW7orH6UXgu/dT
M2wkzIBSQ1c4nhGQtTwctkw9r6QNywG3cnGpwpF3Djv5NrieTahHKwKJP+DKqqJwZBxcNlbCq4br
BbPOdZfFwbvE6zBLIKcc+REwP49mi1VYNK6PrBWWoEf/neYirmL0L+iOnqfR3abMuIef9ZMsWHX3
EJ6UN1DnlOvun+EbUR/Oj9VBq7SsN/z95xoiS08Hi6rk0ZLGY93guBL3FKfurCnrs2S1kWY5mCIF
d4k65jcJSrPfbUNKDjc8Cj7VTpHJv3JsdCGchFuXEw8w8zaIhdFCLdCzbw/mkqTR5KYVFpivwXVa
bIUFSFxteYu5xPteJ6+H9rhhWLqToWNJRrzDc1i3QvxoFQ3i5KtzFdC0GhhleesR7k1z+DRCmgwJ
XVfrps/pSH1q1THKwEBHDinudAyJZTtLgi8Xu/NappySFyerkaCqRoKuYi+BTkVNQmnUukZ8OEZL
719MPC9dwwr7NDgn2XQWeyw+D7F8XgW2mL9LhkMdvrNk6koBWpe8WI3Kea71yaCv4KIdgMOiUiF4
RuSRlGMLJcvQmaQ3f0ZFeOcdE61DlRAQrPWl+SA935pD51tH4MHf6AluQba59k6hTpXm6Q59NhwJ
1rBVBjrzSi4ONVBCbXFPkIPnGdbHl/M3ueiW0Nb8NWNxjVQAEkypFm7BGKaD1y3/HFt+YgkWKodq
Sd5M9En45pIAzCscTIw9DJi3DGiF/DRf7WrXD2RsthCHz2ic1tC0vgpO3j0IM5xwh6j7A8CB7htc
CfFxqp/hS4doXKVfUXdq+djnP5KL4xKgX4hn2smpW81wQJe1h+/gOmXc56rCYlSOVuepM8RFWiq/
cNWEF+zkeq2aa2SMbiS28DjIkwg5euarBpNgtIIQGjJuv330uwpUrTewL9/491alkki188wlYB6m
EJ/qwQn0j/geIfbmN8/noVvd7L4CPsSYrXNflbUHkfGbxMO1vnC3YjP1p+F8rhVh/KedDTKK9n/d
XaWiml55TOpNmkcMxEkED9XI3S9n1y6XEyCRTWuQ41MAs6gD2+GLuaBjzmFqE9siiuAXtpuTk0pi
FaC4V9kS11N0g6mqqyTIfJDrmTnHrUMpmJPPYxG+FwSNTD+PPsm+uW+TrKdyEJEB+mEG4tYbjC87
o72Jeg62unhUDR0WYl6f7ryRUGFWOUBaXR8WE8lMZm0UoRBS1BaVnlF/9xTLXC7lcdZZzn356HiE
TtjS48UMNNnmWV5aS9PxWFSTbvi6GModAPd6lLIpHkS68V8va2TbHOPc1OgVBXnCaf+L/nLcnkPh
IUiVOuUD+dDDBwlR836bh6fzw/FpCYLCm0LJVtEYs0Iq5bswKRAEJNT8DqPcC90ybwr72Yhf4cAi
n6J+i3OmH3t8YaudysmQKsJqKjP68uI9uhJ+iCLubjNDroXW4NrT8O7wCZv8J9rbgp8nH6qbSC64
NgyL8aPtwLLr0fRvMRu93mK8I5SFmC+vFqc+keq7KMJ2xxgQ4aiKPdY+RQ0Yz14WzBOZQ6lisFfa
OFC1alNKUy5zPIuY2zEeUB2+TtB8KYIo23RBP5GvKwARoBY+bT9dvUyF0H+U/vg+5HMO/Cf6mv43
jlxVqvRp2lbGyHrSz56LvK1RMKolRy8+EDNQxBX5KF7qwcn4yycb7pix0kXclyPse0xOELp7CwZM
2Zpsg/UdJaLIPh2NGOpdxjAX4YNxFBH7qCypO/FUQSbRHBpq3tBfqYRUcQZAhi57ZXbWFwRTQGuz
fXlJO5FXOR8bchs7M+FumKFysDlMka0HK7T7v7nDVqutgXJUoM+WT+Ecu61NVrR+6cLLjoCtRNrG
SoS8fhg7hJCwO6IQ3mgjqXtZC7ymvBQo33P+0NFe9wBKXsww9r6EwPZS4lofkMArLJ1NX2YN/xZN
v6F1wCBcTY/78LTwNouQdgTBOBAaNiTW0kbx1w6yiJjRVYYdIaWvVvzJCffXw8LE7eXRBKhvzJQD
Pax9di0NyqaxpLLVasqvFIO1Qg5vx5owy9D1lY9T/JJrS8FQAZt7AkAm105B/CFaNIcMAQQpq9ge
daMFz8k8vRJgXs3Hr57183Wl4tCLrq/sjsOKI2UFjGj9e7qfCBUkdwrfHPldD0pPcZsj7kKXxKjD
30weswJz7DcdvgCnVEBtbp2eLFzCkLvluP/u3T9/Y0YiJgGFFUbFbPa2912wHrztuugdD/3hlCXH
5IF/wmrNePM3Vp/vcBnHZBcweay8Kqr7v1fgSTLXJfNnJas8wcOvLAGseqlkyBn/jfuCwz2w6DVI
y0Jf4hI/68N3LF3XWHUJXPbpqVtTNvYN+hd7nomq0D2TV4cjrjDOFpbLWHk2yyxYCqx3QJz9n7fK
h3YKLY0Tg3xKm03BfPAYIDGk9hVVyN2b72iv3Ixt/KesdyiVTBOzPR+HXRU2szCtKH5ubRTn8QfG
xAoMqjSJgJPue4cvYL3XDVuQL4qIZPogAsm5w55zp5fG11qKg7t6EXjaqk65s5usntIFYN1XsriD
/PIWfjtD8YpXdbNCpMPgBsKOlewloyvVnS10aT9ziWH8tH0rkZ69FgYnMxfJ9yEUXKf7HYw6sh9v
48LwaYOJvryhGnMIN2iCAoM0JloON0lfIDe0kv56jbhv4sSyrJWMlLlLsOr0zJIvcRDDAzimrv4Q
oNZJmo+OQ0EAiqyWaJzUNLtsR20VeZyHzZAoa+Pe4V4RJTt4yfbmEToLWyWZbrit+IQOxNV/Aw3v
YA/TB+jgxiaBcXkhG3GcYe0+jhLdQUbjYUDpsbly1tqvxdtrzu4BuIBXH6jIGACowWStzdAsj7k4
AREEKJ1L4eaSzdtrNVwPWEqeknfhmjAjTFrzeNJ8hYLyKohyxR2my7jduIfUaFKggqvOxQoeBaWx
RR8UePeabfLIhXOy0Qd70mjgaxhS3945I90mCkXaqciRPhm2NOVFer0aZJjL0olcpK2irIx+F6X9
bEHOGxmcXMKPaISM05Uj3muxaQSmSH8K7pnuUIy/Dy/apWsH10iAglV0Fuyx2LK3keZlJKhRFW2n
cnKLc3oX8OjO3dStT39ZByw5zq1oKU6p2RShatP/7ERrpCTJBQTZ7Ov9QsrwXNSHUzVB5bROOSog
XqcqhaWOTmbsXUNu1Vy840hLJ4guBVqXl+l4Ey0nffBBRpK2y7Hbwc7/pdO5Vul0oLySN8ugF1h0
8Wie0pLmu29wl2YHp5htJGgxSnU/8bsgBRQRf2/0CpPxfDudJTYUTWyoG/VwIJW4PkYnC1VcPKPQ
+7eY+ayqjSWPNDEU92wMwfs131p595q/yMl6umh8Lkl2pRbz86tos6i1CcrAcpKT9lRyJerUS7U7
3X7Xivs1e6hvyvm4uj83YFkMV6T5sGF2o3/++VhzRPEii+wn36sqVkIAPt+WCKldY6KDHjx0M8nv
UOg9l3mm4lBqkGnQZg4Yt9k69HCXjK9f4sgbRauTZ2yUkzmrxnpKpBfGoKW0fbJVg5rMWOkusE1Y
0yCpngy/M9ZEnyZ+R/uzECHVREvVuOMR0F5ViEfmDckvIi04tF+EKXuGdYM+yJ1l1m1GSuYP6k/a
Soo5mnlVboweiWBCVIr/Wc9sLRwJ4xkxNuG+h1F4SXP0PHUZkh+5CavJD14ghHMOz/1X2Ojre8os
c5hSoud1OBkODmkhsBtB51ZlEOrNwiJnCAEpj7wscJEL6fdPHxVGr6kZ7gC1lpvrixYjsUc1gFtu
clHzQp6gMoNSjMhHs0JnvyDPM4ju2jrQ3/dljeKmiP6P/E+nf1Qw5v4fabaJcRuTvs5HH9odkESN
II3o7ss1w8y41hlX98inVWskJs5JXPyhqA71epuB5datyZ0BY6/RK7e3NV68/zdHG4kp9t3a+Hub
rWTyI2txFxTtIL+jdDjT99Tz/e0ahHnX04SgU3IjGGk0GQ2w24YE3K+ZOMEyGtvAY0aBkCj+/kM+
OGPqf8TnIy2zOroJt+nU9Ok1etxmsgAEl7ln7mZhjEt9RAkpha+VVdgLC8h39Fz9pk7mWFo4FXuM
HysQFg0skjVOU1CcPb7XkowxPVvlvosbc98Yx+zIShY/m43dKZpd5kk4+RtcALYn4xCs3WlLchWm
xyfFA78Pqyorrv7hqDGR/dSZb+OGMmPNFi53mMTNbLoCtHDe9GH9rE1ftIZpkqzZ+SDcZ5c4Dvf0
Y/ZgM3BySWc7P277UtVfaRhxyWHDIi9EL+6yEf8+8pmYEqevelBL7tSoXAxJcLJhlABeLaGCswkI
u75hZwJniGoc9NAe3PF1Ve0+/Mb2a8hBck9U0jQXJM3AxRx5c7gMq3dr7z9MPXZCwg2CA7ljHlEK
fiG05OCSvSGxJnZkfwgGBX0pU0t9sN8oFQ1hMeM6vUdj/30pAIKKKwxUAs2DXrh8U5HbaC1/LSdZ
DW432klzUW7ykJPS/ZGhA3kJ0QZ3Kvd8Rb3SKx3r+DeWDqrmAJpeh5EcCcZckIq5WmUYosRgdWuU
Asn1HVXHcoprlvy+DToLCqEpusHKgLy9adW8Z6zIvNh9ML14S8bsh/tdmYAsGWayVHwRd/Zl4ovQ
0OqsevOCcFuqY8e/hqAKfr45AZSMvwrz4ecs/SfPUEMpGf1qZl5hb5LueUrnI2u9yf/zYk4+knNM
OZKApXejZS1Pt1zDXPNB2s5kXeNM73CnvSfAm6kBaF+R0yx5XCek+h6GA6KBxn4z9frmpFZqwrtY
2gT4cCVhBflAVqjkRd7EoacR9Kt5QZWSUQ/IAFBQ92BiRTX1QAitJyWJ02UHhIb0t2dPN/Td3Zqm
RLvyxpUhus+vWFdr7bn9NKJpt/oaFr1G/zrQZlo2uRwpkQnqvEskjrwo1wPbIbiQshTIUHP7fTkC
75KKyvbKwsZ5DmaO+9bHtSVDaTxgm4/nrqOK7yMW+MSAP7liK5lI+C5Fhh7lPzH3De4CD89aUkHm
gqq0wjFcEhxdmsXLuqGGTDF0DFuAoQQzXoF5K7nJSt6W8BR/bfOQEQcuJEJwgZfsoDDy87KRRfSc
qNB7jwri07bcYF0F6Df/EIUtVc6RSQiju5SW+G/YwnU1eF4gH+2sK2l2QcadYovrdPP74XO89H3/
bwtBTQHzbdLMeZgRwmisHmfNMQdKgXe4N/BsQlWU+ifoYQXRaoYtXzX137aTp5h3gi2sCQZ6Mbua
S3M+R1zkEbPThEZV5b2TDEB4PJ+qZmLMlJMfNWjV36Lyyqclcv4tyFFV/1NVb7vOGViwWKo8KCzY
dx5TA+foKZQnn5Lk3M7ktCpL3z5ZEsylFm5s5fsQIp83DBRCE3ED1LmryRLT/JjLfsfRyXEiNlcU
YLhN1a2S3Yp8MtSeKUH0PFPNMEDK7O81bGJVQOXF3m7Dv5PhDnBv0u39+k7Sdiza9xuBYhIUIkA9
qFrklEZtca40yioGwpTfJw/stgvcJPV0HasN+0+5kW/gAoV+GMGFP/Oi9q0ZWejrKSMol9q0USHs
hNEZWFZw3YHWJln+O5qct0+Kt5+ooBHVN+/eK6TbqbawaMP9nOyw/I/vwlUSDM5ky1vNBEpmpYIf
pT2mgmkveqdRc0kpB9tuhHztVMwDgAFYWCuQLmC2IwGYcyzfmCQGTsEJRwfI3GhDPEkT8eGBunFZ
1PK+SbemKfB/o1OFq1fQXvFtK9SXi3IwiXcmxwECnNpai53SA6ZrHA2ITXvh2v6O7DEKN7jAi9nI
ZCjL8yRv4Q0nqnhpMVTr6YBN2SEqDz5rzEKQHTr4QNuQ6tYKMCnIkona4HFBQ9WrRpXr4prbLYRE
pGGtZ09Frke16vDOKaSpn44hhhb8AIz/ZcbvuLOs9xlRAO5J3ofiYuJP2wp0OgBZvsCNAe4gAEQh
0n5ZXWMsdoan5ad3wAFph1wI0hGFCrdRV4t7n3MEluP4AkCHZb07lWKOxsOE+n1INhDvCc78lTH7
iguFJVE0fLhPOT1/rWD+xTpM9zHSD0GTcRgXfRHu5tu43rBFQcRL4nyfSphlJtV1kD2AGgM1WgHv
gH6tp6vngoZCb+Yvw95x853m11ejxEXVBX0O6ozWTu29sndPKAsoaOz798QdX9MJQGFBjI12d4Xv
5VEQ9gEKuz8HKFx0sViQSNvUjrpR/+gNZ1Nr9gxp72zkhwECgi1lxN6PGLA3ihu/JdhAYSsSMkVv
8jVxwr9YUE9ry9vw5/6a2L0l+EDWbi69R084VMRQDWAqagcEMmxfp5yoSrpGU05arwQF8CWA/HKW
2FhHWROrOUAlh9MurThrMbAm/pI5jxZwpDozul7lLe2CNPJJ50tG+PP/8Vn7LsrItBRaDauZ+M/B
SYZBoSOSXjBGpatL3lAxJ3CRHmnT6+t3wkLP3VuCDDfkGzmds8Ptz0IpAIDa//oBQRImlX+dxPj3
payROEGBYeIpVviLtqJ72W4Xw40YfFpoJCnEvLInTFJlMIldylom4uglDXgI8ezqb7DHWuh6Ag+H
t6bY4nBxmVfU5HtqtTyomhJGhOmYihaP6LwOmlWppsGN7p3gXQdnd9N/CGOx5lGV9zTbK8TyvA8w
VTfiH7ROAselavBAtQBhVysl8+QAMh26BVAdy4CATs+p6Dr60Vney4J82ptHsuv5n5nHYBbQKiq2
06Y+4vpzGX4+JufWCP01U8boK5SYazvahIXRiEhkQGQY8ltLGSPiB47WNu6abWa9dRcKjMd2uUsE
pLSYeq44UGh4u/yWCVdz2mRkQH1WE6qjEuOiSVCurajEOLLs5u6HTea7ZWU9DY9T3iPShCin5P+H
5PNpz6k+d5ckw9YhWygX39mP21avBtLfcQFcH95XTj6iNIzz5UaMguEAneCtWPAPkGPvu4ucVOZk
eKM3AjoZ/qflBCsDF3ZsMEXV2u5Uvz3dK3adtrhI9ANLNeNi8KVdHjBjJmw6FI0NF4bj/j2NaNH4
7ioQN1gdn4+cS65rA5lEL5z3aFk0JpVk+NwE1iAvAVcn9DJ/g0GbyhzP6ADcwkaZ+B5S4v7wFbz/
YfnoPc5/Cd5TL3vlvWDw7morwgd6MbuF6peDoWpfvKsVltuTExH4lyV4do9ofzhv10ObN35UCTrw
JKAyXR4aBu91nFTdK20fSYtVHXsxfTIw4CUJzBZWtPz2gGSpkCKhrj+Up9GPQXkw8DGSXKWEml1A
CaC8wCrcwKfLzF7kfnLIbc6wz2jSO1g0qesf5MIIMT7UpMA0P1hcAJyaji7k+Zw1vXdXlKENT/cm
5A30VCQNu2XvYk9Oy/HcQ3C56yffatnYyeIOwTMc+POmc1/8zYs2Nr++xqtFOGBaT+ak0wF4efg2
7zM4qN4Mf9DwaFdHkpg9WW1REQdaKyRwPZCxkm6y0Kwc4mKsDnJ3RFFSwL5FLjEd1VKivyXR0cUB
+eOoUbobUKYfENo/Tqe7y8VJrPdYjkSbVWHtm5XlLxnWNGUMEypGFGDsouvE57e1mzOaQ3YaTU6Q
U26B3JhV6d4yOIUb3YmHMMEN96W/9gKW2pChrJ1QtF9WWYWNxoWTTNgsi/VNG6/p5NNHSBfkDV5h
pojFHxtevGLYCy2gRqA1He5UbsEbdZS2Eph7qPyfjWeqY+kxCu1HpX2QwmBsxCeVf3xMWklcsd4+
hOu89pSNL2pMi7kPyCkoNKzkpOTXdtvZ+FqXxvIVUiKjIf/TaxmfXvrX8b6nNdtkP/4AAVGyYzy5
R+6dKhrETH0fmJJmocOKi2Beah7WXrTytroRzN9KyO4fBITp0PeD5vpOKKtHZJJW0w1wm7kYIjHU
f5a5UoX+lo/fsaIJZaeHdvbQoBE6nylpWTMI4rElT/ETXiYQu6pzoFIyqutc3zvBQMg4oHJqgVbD
UFLCmOO2AEuyW/wjAe5OPUeAjIzsoOZOcoN9Tp3DPbbfbqiA2ioK+JRGue7+TQga44KecWZoqWNE
TmhJXToIXBybZaDAsSVZHA9wT0Cx6vzq9LLxAgCceUlUFVnPp4TitqGVv+fjBI2+z2axQNRozZzi
/WtxM//9y1DuqzQfdylNIEISO+cFSxHdFrXwTUWvoWgLfb+UryRReUaFcPTYtOXvjnNFkgCz47f8
pQZD4Qm8CKJbR/i5Xtcda9MBUzcKEBfLDx8IqxYx4h6V2rmpKjcFYGzOS2dv9H0u0XTSTGxzofCG
AGZZcAcpp2u1gFe8HTvAM3MeIFmpJNZYDNCo4dX1gfJQe7cuAeofji7AfVce3OTYdvxXNY38olTR
Cgpqr9Zut3JIo1nYutdZGeyEEa/rMfDrq0BIvupDq6jJNXcn9Ui6TYpKFJITlS+KTR+o4EN9Y5Gt
Q788g5qgmQ/jz0Usq034AZZ+s63b4ysw9f/zYerQiUwcgOCf+qfnX+3531oM+hHCuyJ0IbXbhJ/C
t3sTspIB1c02d5n8I+Lc44f6w+rZZHSh8KuwYMKpwzIG0nELNaavIQRIxShSoy1gDBVqWYpvA4ti
Y0Rk1IHcpgIbUa/sM2E2jEa/9VHbWRhA1KUJwKkN1kbxqUbIYVV3NGzkLAcFtAf1ffsjG3Fz/Pns
owxWJeywd3REckwd0cG/BNl3GhS+LG9gac4C9tBifMSqWCxyoxWF1Equ5V88hBanWj/f7qIpDfnx
ZyYXjQUoXUVhFMAxpzwVlptDmifMtIt5Nz7M9MXvcEexgPqnk8a36OJWw4Zz8PsCpYWyBOHARVjk
Q4hViH4Lh5gdTq/pUOUexTW84hPnTeVSinmybPID75TKJPs+DqzT4JW2hiM3kCgEMSLt7IWCh+5c
/nIEIJ9Eyco3nhe0JTt0zWMTWCIZRL9MhYgr34K/eUTnYwutgvKLrSioiFjxyiiC4I7+F8fDqIyO
IJC9jQlU7uq90YtrIzKKlqpoGOZbSRNJoIcluafiWUI70InHANdQxn6+mvsWfbXCPZFLWcBP1U22
CXBSIS49FIDuu9zHcDleiHPwE+o/DY4OjVC/t8fAsfLz153WgK/Uf0wI5OAU3/V0TykkFxntpKU7
nmWaFp9Y+uPvPULAr55k3pmzuiOlnf+vAkQ7gAtOVq9bonJiGcl0Vt4Rc7+iFj+iPV458iapuDln
aY/tYVEIK7qukDIL+yBKHauLeUe9jBlu2vNHdIr3OzL8to2i+zN/LSMAidEDjCMXqSfMXdaFD0Fo
sDbnppQ7tbacnWlv9es8gfJt9UKXcV3JOWxixkHrOuv7ZiJf3F1Q8E89t/NZUtlhR2ddwtq0gYtV
CQ54WhlPnnfndZ5l1l21i2kyEuEG+YATro8x0Up5F4eh3+fK4OT/34DKIVnIyPQiM/Eq6n2NA2/V
KN9d1J7QUqdVgl53bdAcKsgvIW6lgJNRUi/c9xmzmep5yvhO1zb/ELVrSJ67IEyQPrawbMMZSmHM
CPr9Dos2GpADWaRkJ+kIaeD3bkXjqWzGa11q4fFillNuVgvjrsVxJ/VfpIgj+iWuy4MXTeA1JQZo
MgHTa56MxbiuEKxK6l/XSWTfdBhQS3iBQjqtC63eZ2+M5qGYaDkegaeU4x1d9VZJ/UWNRINXLoaV
i8PsBcs6EhwPi2erS4g+C+tkj2RYRx/U7A/7SUDvXJhBMNXVEKQW8UQzMcAYc8E/vinX+k5nhXsp
V93MPhHBQpJE9AUaAk/GL4xnW4DHJOWIUQbXDJjzjht4GOwf7bZFimCVlx7EBUBipb5a05jHfmaL
CNoz6ZKS47WZwUSxPnOUhQtAvdHFrGQPwuqCPPSEo/DB8ZsrNsHVA4q9j/fgLZ8WtDaxcCKF3jEJ
byKjrMHwI0uzJqvwEOthI2djlMLuGDhICL6d2OVhQDIoLRSGtAcc6PPGqxvnuf4BTM9znnaPd3mT
f6llMSxiENMzwhAFTq45VMzj7cUaxVJ4uILGFZg6lYoKp/GpcfUyjWoJuSQxlSB/symmlERtEIWk
dewzPoTwN1F2t3UnJMLYH6M2U2v9nFcowPB6YcNHfxgRRa6FW0c6AhQE21VMwF/4Uflku7ruD1oz
x+7ze6q/LbDMD2eo1vfCYtzPJD9EYEPQbNjcK8zMobk7bWHm82IHVTufBatCp5g78nkB78mDvWBh
1pR6obZbQPuMyKm69LX59AaguRDgIXBB2so93k/04KJFXoLqSK+Lkxbe4DroAnZfpPhv+up6q+8/
uwiE4491C3i6WFAM8eenFNc4RnQWqB+Zo8yp7Slr9z9QKMJ40U6+JxmB4c86giIRIWxeScRZj4OU
Nf6Zb4bXoWi7WQ3nCFFw9obn+5Bcxa/1MvorPwXei2O6M7gBeqRLheu+HleyeHnqhnhFcupSue0E
dnambO4MEq/KpyvMS+NGis6iNLY7lFfYEU+8Jch07URwGui8D2sZCKWQdt+ChIVNXAJ2B768xax7
wyXMLTdxvEVXVSIk1Bb8OUrJ7xfeMxvHwaEzFPMquVqRMWpHo9Xdf7CyitCjEOCKdqJuBX6HPGr2
InCEUbUEVq1ugXQzkg3ON0ranqA1Z9nWmEq/ckIKtBCotxCN2ZppLp3VofWKVmVNGPCWE16rYNlH
QhW+AjpYmxbAL26/ENIP2nskzD3kG2Modfmmu1iM82sQdc/pZ5TE6GPcIj1R/Hj6C/JSrF3XTDjA
4E4Y80IJ8vRb22aa+uwmkSpGWh9ylWsV+CCfqrZcwatjJ6ra32m+jXRulhx0+PrbxZTpcfNOGdN9
ulrabsgkIppky81uoFhsyZoU/1FHuE8VQJRYn9EUuPim9mKp7FY7K/8aRN6L0Y7dbWu6s1OYo7Bf
G2ce/CynDFL0YX0JuxxNrIPe97BUMq7+zYPLJNLqjFVYp3xVi2yPx3sKjmXZalq/z8tir83PqBFT
MN6Ol6AnNWK7qajiLvxcn2krT/blRcjCd9H/LnyZQxRAVN6EAmKH7WnpjuZe080ddKJUP3yqkBsP
CAduSuJObA//mu83PQGFL0PTQUHTbZ4Z80nFfFe99CX2PKxutUoVnE5qIzsbTWi2sDxwQyGE3bNs
KKNPoh+sgWV5cU9Ly8SdN4TnWmx+wLDQ6pLfQgz5n6zxSu00V/bLuf2+Z8IS8E9CVUMQ366C0JL4
UiF55E4DvO7qQpw/H1xjRf/XNNit0JNCuQ5OWkJiIm5bT8/Fvl4hCP/82QRb0eUhnWneXN+FdJyC
DF8FDZyDv6e7IaUEV7LfsyxbBt57INa82dRpOIRo6JonOTpzrbhSH1qX0zERrbpW1DMN6A/Y82yn
A/YQ91sBl75YTVBcQsnXtC1Nlu/rjQtI+rOpvwzk5P1sTAYF2F7WPZHfsJV6vLr4bz6qF/pzq4tb
rbEY3LJZcVHLZd7D129WXrQJ8TKr1/8OFV60oo64dqXScFb7OimxArywEiQYn25Yyxw5n0LuJ6pW
XdflDO69yL2fz/QASy9c8C7DfHki1MfDAegyHJ+wlsCBWQokgIvT9NMRKofJIGcNecQz9PRrmvG3
xrRQwCPJPSOk9xTHpYxl8PIgZWDZvhBlCAw/N86hdiRyEBjvTb0mz4KsJh6ZjctpDgrv5E1WSZJ0
fOANb6hb0XdNxZDa2jYeweu2pMSGz3idPboqgD5ws+yZ3mocWcS9FlIHN+9zEwkAlO851Vy+DM1e
6PhWRdzLKJ2oDdwNatEvF1aP0CdyxMdUblpr5TrOwLb9MsTN0ZIcItPM/2IOC1aZk/RlI00NScu2
Gn0jSYMwYP9uErtOkhuOp2nY3sluanjtDxXazEIGmRmRlGzZCm7Nz6LvoU7skE9g1BVIg/cUq/mU
CJ/ZBy5poU96JJMLKYWG0ZXbdcH3vmwEJXgcwaRBeExLptCob05/J9OYE/XfxhHKc6aEKJ88aATS
ovF+A96kxmivpDiOXUcvCPw9Cecfi9aYsnG1bykeNARo3ewWkmZotD+538zmr2Yx7FZjc9n8NqMA
Rg/O88PN92RtUgXajlib9XG+5qwHdoJrGA85uGWzoYUgtv8f59/5sznmE1S6JQDGNiTLtin1jUf2
QMQ47u4OafrfkMqquQwjQ3HJrs754jtY8IWDtl26yCCax/cwhHBHKMwvgsMReIpmvZ8zOEFGPnIH
4SbiBNdyIju7s8l0TnSLJ2HndOehJ/8HQC6nX6fkVy4xL6TOJWm04OzOdMFC3H3Fi+iIZ/B/XVAg
nu8i+wSalrCgJ340dzx+fq9y86P3hZ1sp1X9IkR8yQEadQrlEPxQ6IKVMIhsqI0v9LtevafmU3uI
nmjl7ZaOxHtOppXcB4FSf7vPSDkFl+m7P0TZG2ODUaPvaYOiGJkA/6WH6rdAoyBKBaECQYVBYoPi
JkGdaN7dgJn9IQns3/e3n7QFoorPBqdgBiT2ye76nzCZHUuD+WngoYDO3ieR/1lS5PaSylqSPuMN
wDi8Y8JrHD+72nWb2CO1MFnHcOi1CWVz3XVHRE0Snn0tZJc561YR4QgXYzXwYbvnwlYI/dG8a+V+
aCo21FAJwnQqnH9r75FfJMrmEFIqEtQVH3UTHp/AL1UbCX5YMiLZFWqprRqY2P2xSm2owtLXQEYb
3b+QRnnlhmPBjBLILJ/ZUQ2a8xrN6f5nOyaiYr3iLXSliV6I0MO4/wIv67PpBRjJ1FUCTc3IXXby
dg5l1jiiioFSBLLhPKc35fRW6hpmcM7x/zNFSwHKV4t02RhfkcKppJe0ni1Z0y0KSPg6zh2gCLkX
k0ncc/B81uRU+y/1JZ113wST9snpXnGcGpAzxXCNvW3DDMrTnEAFoF2w9SM3HkoExjdD9mNfgfzX
RcgG0SgxCoR/Q3w/8IuakMx+WHW7V2NENvLk5x1cRMd+AB4BR8YRDEKcP/gLTNhn8/8bzV77sTxy
Zfcq7JwQj7oywzcBYPdrtBgjSQ3Jf1GTp/Gu6k1SYdXUYU+o3ls8UXu8wUqsLkZ+DzxvsJSW05Nt
Ioakv1tS2QJ6JNM4vTHjcUwEF2y4vxFt2RMdyOqpcuYPR5zfFyWpMNvfQYENGk0xLz+5Mgs6sIQ5
aUOUs/X3JRhpp9PNZhXlEp0pLfAiaOkjhEuOHkyxVOiPCmQvuqzMCIwxVVAGHhXnILPm39nAEzqe
1EZhO09RhICYz4aagtJnq+mnB4UgKosoRiGmn/oyjTJliPRBHbMoJVNAIlYqtKgXjpepM5c3Lmh/
q9J29/HbGaCifJcS3ZYhgx/24pyJZAZbVYeNO78UD7tEx1Q1ALZygDtu6SDvO54M4xVFYVqoGa5S
PbmKEOyPubTU3Gtbp6a0LNTj2gsN5fhAepuW4tP/KlNMfBpmKfyiXjYDemwoFTibE+snbrMpp0nj
8m8GknXJK5C5mFl7F/LowFwfQAQ6YVHEWIzaVLBmMoyb1Zmhm8X8Bcgq2n0PHHrImsP+C92TrhJo
yZkmulYz5E+dqYWbuoqZzGSA/pLADafOB5KJu6xVvuwoPpwg5ot62xpB7Rt7v7tgO+9FwyY8FVVq
pcMa3ISbWKuvPTOAwi3q46LwSe5X6yTS8idrL8lKqHmYaRloH1+umhtTQrbTlC2XQvBglzpqAoz4
sKGhOt2OxEcOgfK74UXTKCbA9RfWaUVie5be9Uott75IfsYQa5Tg9qgwyrfb2ISsc7d20l9QdDkx
hOckv73BLvd0hIPXjGdb1d//QNIygKfwvP5A+87ocC0b7q1NoJafDw39VAkzenZLVNfCDpsd2Sdw
oAxvocBjpWjxcdHyDXjGBD35VrZPn4hauT3R6RFHXjL3GxEzZ4raxtq8SyOPgf4ZytosRNNfBM43
+FV+nQ3tAS6UhWbIcwBzstu/v9gbbFIDbaHjoWIHfVE3kBqw9Qj+QdG2L4VoMCAb/rKpUQyioyA1
QbODbj6mNbu5kDKX2XFZsU8JWL0B1TZObta42O+7dwDrFokP91h6zytZxHdS3ExMYO3DrUwIOEH2
ODf++x220YQqKFRxVh5aNcBXDcs2b6PG2fwvUOSm9umgTbyjZEEuxrvt4JjII5c2EtPs3/jDQXjo
U1xDTw6cez8LowIP6YenR4nYi+8NDSACESwjcJhvLwOb2lMwBS9mGsAUtamkgYI4Buh7z5/Vpq+h
OOtHDt4PFgjxce4BaV1H8Lz2WxuYUCRVBIC9sBPAwrkSfq1Xhy2AHmYIQeZwb+p6lxEcJNZgERlK
cSB8gCnKekjZl1fy0OYoRjewlxdeM1Ow9tGSI+CnnFY1rZrFJ7GgQhf3mBRPpClI5+x/4kGvFcVZ
XnrDi6cT6xm67JpUCAfJntPD5ohgqDEtZqyRDn7zWxtV1FzHMxPexmMM5rd1cMOE77zixXkKQ2un
kkxZEXGHhMY18l5X22jmxTJoWmaA6f3uQHmUa+GEI0Vq+08HKdzgQ+rZdCne2eAAQbsyOLFWFMIZ
VY1ZfUcmOjaUBit94x+O2SywYZPV91mbBmNHRo8Lwtm8BkerMWkBPf4J6xQnKwWa/NwKUmsXBXhN
NEUbg6Dzz3zZCWz5lQZmBky/6cY/Ku2Hq7R5cffXWk/6iY/sDONQ6sCZ+1KjcKMozU2Bxtx+Ybef
nNZtGN6j3Na19P0ZmPzrjtcg6DkqmNoU7/bPKZ2IpiV8n063R9Ywdw+ZSzb+Io213curY6P3d0p8
z91xQ8kV/ZpchCuGGQxrHLT8bgXWfJtlXsRcdiUQ+FDlOyQof6nl4GutHNNdg6lnd1h3wyetgqx+
Jxf4FPHCA/4grq80/D/CIKCnDulnmCQlGX+7QF/VjEeHjnYpTrfI1FZoXYz9bYaep310KKB73ACV
sfw76qfj0CCSzqicGNx0lbU/9FsB8uc1hCfZNCKtyn82usd1s8QgFG1c9CoEpBy8qPXtv05i/5m4
RYF6FARwSS/VvnNmdrlUWPmzTjDVKBApeRmU2AA30rTjR8xbQ6u2z/1cZ31hQ+Ypv12W/9ohxwJ5
58jc3BhwvE6T9BnAEXLVAxgeFQKcZtI6ofzmoTdHDxcVw0WGnIXKrs4UhprDKZwq2pncSa4mK0cI
aitlUAVyvthPUZIcjm8APyBncHYMMpsaNgb9I+RQmlWFEoO70j7AcaEOiMTdPiXoWUg439gVl5pz
hNGUqXF9BL9HGTlC2IVrwfU28F1DM1L4lSpDBaivymwGqgdIUuLx7BT/wy/CsrdDhfsnzedy/FBg
n2n8SlTyOg6RRBxzDXb5EKyosBTTF6y0yA32a18YSXK96V6GH4A2a1wIa2enRVYDq2hkvNmJLY1A
iMA4UmqlAIwwdjAZpKUGFMG+W/87/hI8lHzV5JoJeQCX8fKEMtYoLK+dIq3gHdVRCGmfVn5ksmxV
SwtCm2ylDcJpA2mfGDoGvlT/RAKV2Rjq8h7gN3nuhF0rQRApmG2iPkFl2loraeWrMWKNxznZvs3W
zAOdsijNpIMW96ATWOcCrhj1mxZw7H70Tg90POO9W2ts8DayfwvvJm1d7bGy5NEVEkPe1lyFLrtO
4/Le0Ad2fG5Q2FVDoyt258OvTW9NT9Z067+8y8vuHDF7/xC3ljiiYwVm5fEgH6eltSjw2zmDpkVp
YcBwN+zuiFkpIFw7dk6bRwgaT+PYFwXG4PjjITzFEr3E1Zeqjz1cjPLL7Jo7vUFF9XJ4pDrc8dqy
YbS4DdgZQ/qRSn4IiXzuB4p6cy+4J3wGrIO704D2TxGe+0f5QijhoFXKqaN232ItSXjhFT8s3n5b
AHyMXez1itqtmWcpfXDIFG7cxcybHIcLTwQajdQ0cM/D2BrTfFtdn1YTwJ4MxbZxNH2/+kanLMC2
RSsRarh0Scg+eEjhRiRp7aPnNj3dreWhY7CKcNKAvCkaNWmb0PRINakNVK0fkv2GFlfZPm5icSxZ
sWoIwjpOKpEWpxRGHMzEEoMC+U/6+haLT4RKEMNqFAckETCxvwdIQYjr/7lQotCwINrfa+HE/F8r
HJQi0pjK1y0bb7xoOTxZCf9Xx/47R4fxSvIgoVsKOO7C96sC7EAKrT+Eg/nu4SAw5oGPCW0bi9b1
RQld8zROM14EIKICS7kMoOBK5qquBdh8ks48SBIE61IU/y5vaCYHfAu73c9lwK4DQsbP3qNduoU+
0ndHWYVbMr0+oz2hVkg4PpCpqlyuHiSWqflqOBXE9lvlZ9qRnRs4lI+znAx3yLFJzrjYRnXvA0gO
tjUT/5pQbloXtEDQOSLPGRBcLkxoSs4szbE23agkuOfYPbM3b4eHSH81I0ZzawHlslMcFLKBmu7p
cuXZMrKOMytlBZhG3CoXmzhYFqXOSgMQVVVLvlGtoQFCe2PCsQ93x7kyw6Iknzez+3vVR+JgCd9M
7hg06ATnvNsZEfPrPdGnUNcjQ5SwrU+vXOqQ78VxOdd6fVsTtHpgFVb3cTLD1dkwT0DGTCUH1DyF
iTREdP8MqMwDzfClUdL3AWwDVN60iDmpoefyl/5rx1OMm5rm+YhwpjGXgQccAG0O3R5rrNccec4Q
TBpVu83NZIM8i/Wn5wDaBxnRNlNe8tYulePLV69kJuLP9A6eXKyZQ78zxuZGWF9jtuntU5jWMP2E
aRS0425vPOG47yFKpSAmnTenLLLjjgRh3oHcieFbqDNz573HgzOzPS+/5wUEXGMung+XjoD4OgyP
5IUBiCkIvPxfnY9ndAJy817o1RHO94pLgryR765TlUsNlXJWOkC1UZwnFHoR2aF+mSnLThoIOuPu
8rpH+U4MlqKSEnfLpyvL3OUXnlcTcmRWk0eDsAf5Igg8Zwcq3L9EQk7m1LyIPqw7bpISySbtfU9s
gfULtOQJnNeXbYuSw0mUXttDETHmgbul0OAzAxf4q5BJGUDs0NwdWh8HCF4VRCyYO2QRVig9uxB1
jP4l+6KH+Xap0Aef03FlR4kFsvqmIF4boBra7pwj8MU3wNtHep2APCPvBEbz3WbGMLJ6rMnabcIT
sWFeGlZ714laHqx+m6qHllu0zpBJ8W2bQdaWrVqzFGXMaNRkdYsTNMA8ayLm2ZibEdYVAgzcvv+w
LDpZtQGG5ENLPcW3Vd5xxK6+5ZGpM7PiQmZ9Jhdru4SDI2JIOp2oqQGEO+VHq+CnV9kpV7WDpcMS
CZ2algocWyes+YZW2UcZoxqMNUBpJ890wyqmv30CsFtw7b4JYnZwjliYHs/lpd/cypTylU5V9G1q
9YlIA+R1vnbOcaEGokSwjQrTm/vDBNdL85l8YsnBTd9FXTnq/VN1oTN+kB+K+CVt2+DVRMl8UTPC
fYgJk8a0R/pkXbt18cjUAH1N4LyLBi9P88B2ZM91Zn8LiNWbshgtxqFpC/aUIA42QPOzUAQy/XAV
CGYx56KqDdR+33/HYfDPgqJsaH+GkS/oQR3bx8kBwgeLMUcr6nzQwbdPhiZe7rfqSfcUBQ5ObTke
PkmKLGCVpG3iTPp5rptmiB88R87iP3QDvZKMRJfC8eHTij1grz7Cv4OHPJW1fd1pTu8WSv1o6pcW
BJqFEkQamTV58shRizhtZ0iAzVaTDupbCTKWjKznvZluggx59Q31jHwBorSH8G1vuaMgN70nrFOW
GjZy4K1c/O10VFY+RXuyIfxyvmJljhkDM8h2WmFTwqnURL7lTRehBHqMZs3FqopH2zm9nf+w6+51
X1KgZnqL/E2zl4TmiDmDb5mrOjL/ulD2SA89zd+9AM6BFdur90cJP1fZTDmi/dwLiZMu8Rhl2uXq
QbAh68ChUvqLTOO6hOVx7YugwZEs3zlVVbmVwCCQqVf51/VYPnQfzGLrlur0Yqv/XHHFKil70fuh
vU3mlA0lnicvTDeXpWwfpmryXgkr6eRzc+ypY4V4kAG14r4EM8SVK3T3gwBJrzirkXs8IDJR8lEH
xSUDGGrUUg27cBWWfeapAmSXHjSMIjWh79CBM+R5ODdAuxgFVoaW6+cNb/7oIROuTR/lie7Paz9/
qaJxz5ddMdVJxwKEw1ZltziBCUOBPIUO+pw9rWtRXToeoSZxL6y6HED+Zw5xMI/ov1vR2NXUbT3t
lDNJAwvUhrYnGKKxMH63zaBjd2IsHBDjZJHBkszqEjTKo3na4n+CN5wu0jF48aPCHR4h+bPEnNIG
T1Xo7REmmlHwItOXUFyQZgIM2cpA8zOpBKxfsAEeUJmcqcdhf3JNI2Gh7I0FV10BZ/ykXHeh+P+r
JX+mpFQhvp3ibR/9w1HDaLZd3q5dJxIiECQv9N7s+JCkIihwf03HapDIbm8mu3OgyByRwzR36xv6
NqZ9dEspHHptCNyTQW9ZPllDz2aWgLUrArhQAJ3c+X/eoj9Vb4yhx5O4pAEgroc+jsiBmLaiqCrj
6Lgfyl9q6UW2+KAi9JzC368E0SFSarquOkfMZBuBmlZbno+wv5obz82oc7dZWMyy++Syy5j8xEFf
LgvdxmKGbR5eEMqhZaxB8PFygbieXdHXwNtXwoqCRTJoWBlL++sgPac3LziB6HU/b7CGRn3+qGtp
7p63CVNelHjvG81CJcZvTGIAtHfyIlTVZSyG6iaOQKWrksgLZBlXeR1wIK57UvrZgadY3Q4vz2Bs
nk67YxwEa17I2JjLcFvAnUWVVlBom529El2wwQhCtPRzlFsgK2cWDWMNqTKH0xYAWmk/caF4EbQm
3iIrUz1f0DQjyEo9VOU0XzlbpYzGwGGmTavVnezbn+pBlAuQafYIf6R00Qu2I+V423HLcbMR4qT2
zsPFDZt1bFxVRjVdGujQXBpy396TODVZWYs4vS9nzP1dtexGhLepGtDzaHeLqyoZvC1hgoj2kjch
Uxex1knvrj/xivRUTI0V7avULsJW4CEQHDOHqtWuvMv4fdfL0KgLygKKI0PlYJNhHorUlDm+ozwf
DzJ2570PrIRg07Vfilu5WFPTpnL4b3PATj4bBpLdJO5ZX4dHV6oBBrxCYy4D/7YtJyUbOPfalP1G
BijXsZrGeQWkMb3slzaVOjD/g4g1U7R6Y4oB7csxqM4HcgeCQj2IkvgSWNW0XYCjJELU88j1k7KY
tn57Xa+PEQn0JZqRvNgzi8sqG8HgxUhp8ZJFSf9Aw7wNoO+iD101+2hh8CCr95+E1OOoR6DzpFFN
od0CHhCTljtS1P+W8HzRr7FJ/1KJZhWTbjIv0HoxFqumsGtSikFZ52nnWBdlP3xhSLLvvzQ1GvL4
RW3i41mSD6dNzUcvUuS/KTkH5lr93Kb5s7sEes+rFCrxhNRnA9H7bd49yPPvVzraTHvhktOvkFuM
0Co1BBCMLORLsj/2YAClzvB3mWh/hS8K9CQkPRi8fLKvqbvdXbznWbPOH5Q5YlfQt+Jsob3825HA
b2CUFYn7s8ftJmMv4u2TpjbCvzMUD26Auf8xfurdxKzZTmdTXdUd/6MkIGw3Y22+tQJDAQRmGB1/
sZ3qJBC/zwl8Yt7Z7992O2ilRmJyBSvCrn8D+GCj9EfAwA5C7+vCaTi+yCMM3j/AnRPnwN2UMVDY
k2JNsxNwFamITHyrvjMQG3guZm3oDTNhcLdV8KOR73DqCmJLHl2g8Pnz9IBTtCoj19Ob8ijiH7qq
zTqxfM2asEX8ompBGCLlxUEWN9uImK6/uuzQkboHZVXaWx0NSom53zLx0bRo+JbXOisqYrFBFSjy
fiaEBmnXq73OxJPWBue/cr6e3Vwz+CHT4svBDQcG/v8SPSyWh2y9q7rPrZ65lC9kIYrB5cPsfVib
hrFcZLR944QyBcz1zFjRVN6B30Hj5Ms/AWiVOXc4hPxcv8jZe7s5H0zTkIy1qmUdq9xAIvFy9MmL
e5jzQbWlchcEmXwYn9HqjzX0O70HxoAASIEFX6neofSsRV4AJJ8/ABeJ8ndn4ta4uS8BXjgL2eYw
SuOpeUmlQX7hMGXvz3Wo9VtCij0A8q1P6LX11XUKJnnwmUKfWdNsmmgRPvN2YqMKbZlMQSdtN/m1
BZSfVL2kGmBGs8xPNoD5OTPWAEOO3qiQcopKLwsfCtPLzfFqInnJoaeMHw2doxX0jl10YucpMaNy
8lyqQAjY+BjEDYPbt942PmuYPEq/XyZ7IFvq+F3hgjh1k+SfNzxc6kPkqWBlXYtD1zUpFilbmdco
mMKwkE31IMHr3sykmhGUR2kxZvV5fAFd7ZIEeygL5vD6X5jVUopPqdkxhnnRUg1T79C27Ysm5u6v
GnZai5v3mr2B0dLdgJoTTP+Q5631mgGTsc2Km/7Vw/5YfwDxDP/ORaA5IvN6qIHesKsu/XoRLio9
vzWs9fvE65LR7QPKm3ZAq/v9qzSi9YkpdxpNAl58SW3t/q7xw/X/UM4UIhN1yYjPyhBADrRPb5M8
nv9V4NJTlJxcnzORDmvKvl8/bSxwoOkfzRwgSF50t6neeHGYwm064gwqb4UqRi1BRJStkDcmMRId
FI3paO8FAZSUZbqeWZBnmOi9B5G17NjHrqmEmrD+5T2Szt2JKJ8HvkFRJKPtVjoO7DilTvei3Mbm
kfb29voPTVp9aj/G4MbpO32DZQXKifiVkqWH2Du5IPysCnGhdhsmG5AXkKDpFqA3e38PG6QY2waQ
LXZnJDxfa6vZzrSRjBTba/8gabc7nf6MOTQwB/wjG9eOpMOlLrX4T+mBlCHsMJFvqOMq28hMfDum
YxhTYu8x4T1S+GnBNBdtNCxWMTmJQTG2O5/Zh2IDWy2g/ZwaDy1K/SCZP6/x0plM+FSxMhU+J+r+
DYOUoDl3r/Ht+rxs6d8gj6miXN8RjCSWT3N7X/jIpDeklCQIQdGv3+djgyXp5VcPzpEjRph7RjYp
vqxhTAPc2ra5RRh/PwFlXY/uGc4RbLD6CyySNRzuvmiqVUyrwQIjo5ITYCcapnrwhW8fBZ32V4i+
GtSLBmAM+gVNmvlkrsQ7HtTlLF5l5uBJKy+LiX2pelRxjT4ICUZ21+bUmbYSHA3GlBciuo53a3/Y
Tcx7iYZn+aVOPctma1SB5vFtIgbdtNq74S2ieKhclOUqaW4ZBX0zPnXBvviiiPEjd2fIoDvK3U0A
bz2wugdED9QU7K7qLQYxQbMIj0V7OawtY9zQuXVz1SC0O6cxWuxJssaa7M6YCAVwE7LhnwD8iGuC
LWk++a0KYsVgKv+P3G60VjIIX1vtJW1QFmeDQ7RMuQX84VbjcQsWwUtcmff+TK1ym6EHxcboDqry
qsnWHePSyaAL3PXuynhLlqFXbjNxhqD/ktm1vNNq7dEyQ3l2IwsQK/yGgB700uIZImx0CWII2V3+
oZd4qmUsi422qFm1oOPE8XE6CAsHMXJ9W+LvsdUiL4aL8Y84BUMdijACfOElFVEoFgmnnU8Sah/e
eIPSVlhOsk1/vhnpO+4GbtwP9XiVpZ+9xegknvfEgFsZteqDcw+OJujuPeBGlWHh6xjn8t6iPg7r
mrW/GqXbF5iQZqbcO+Wk0OU029jFTqCOeSeHl0bv2cV3uOx5PeQhVCPXXSyeGYTdtP4jyOi697oJ
mkthhbGqaJwYD+qrhyCGftKn1m7Aa+DkYn0GcB4Sm/VcS7olnzpGQFi/XK5rRuA+TSjnHRc8vJMw
dbUDGnfkHYQrOg9wR9JR2WXyRxqx1zFxs2ZTLrARYUH+BNlb4EuhoDld06qAdtHrD+ggAHGBYJbN
0XUr6olvxgMSJ46L5uSOkonZCQlSaX2YZcMWmxaModOW5+wal6a7tIRDml9cSDmpfm2pKvMedWC9
XS94Zo+sgl9EM7CqxqpS0wnLvKGvniv06Q8Ud4KIpsFs0M4F0VBwjSC1+LYxQEC24x5FRPyhkkcj
pmpaT2a9MqNaPJdhmcucG+YAsMJ5cV0aoBVht3tn1uTA4Ns6Isn0q1N1QTy6Q8XRpttH2J1EF6Kt
no3b+26Gumd5olaZ8HrmoSLMg3RPlbGOR3t3ZTe+gk12AfSyTfiMiXjksqgl75Htkt5/9Oh2uUam
4xDe5OOBrXopQnrtWQoz7LQwLyNjXtQRRqqTlarNFS69viV8VWQuzgu+Gobl4vdRewESIYxOVrYl
8ChHCHhUsYnBhntdQAYt+PpypwCZzojK+WzadKY1VLtOnst077rGLR2GNdAmIjBPYPANUBPcrSwb
Q6YYoOu82ONc1S4knVM3zZhZdZ0kyNWEwI9n6wvBCIl4yxPIj3tN6od4/xGgFbtALKgwETRbtk5L
ABmSpTAmaF/47wfOCY1Eqpd+A8ocx/b1dU8hq6PTPvy1KWVX793d2z+E64E39qwiFGd9rdaJSVK9
5AI6M7HK/ZaN7bXc9V/lOYcKrroCuCFXukfTbxqbbd12heR0s918PwlQqR1O+1I81r4cS8K0MxEJ
ovmXfL+1p4ZOW7mK+f0KC6IEfjcY/01c6Xw+bTioZBkvrsCPJ/a9qKMPhnwMJY7qTUoGPZFJJao9
1t70/g78DXv33r6DWSO6XKqbqHe1ZEE4IRLl6mDYcAz7PtYypwDF5deKzqSH55alciByMVZi49HH
K8ydsxPXcOwnIZDaG3w7l1aIvMy6X92O9ZvFUV6x8toHzgrMsmguZXqGwylrl62PYqTReuaRTxSd
fUKQaBTr9iSqqBop/GckYFn/ho/vFp26HaLixpjst/Muak8PmRMNNSkf+do753vkv95bzmurh6/k
xU+a6ZUcTUPQRYcvGDm8jLGwDzPAkBTcXFogC9lvYk/v7p3eqx3a2E15uYIg8p7j/aD8TmRA7eZq
5LI600nE+yz+fx9jyejSN4ajGJvPPng/5gkhpsZEHDhhm8oR4Q4+dhuqKOjDLucSzX+3w/KvR0Sk
Hcz9q5yCHQIY2oZJny+PZzlVcLxwZOxfqNyuk5XExhLxD30kb19mgWCirGRUHmVJvQQxEEq2wuKg
j6UgMJZVScZtLJhUhQxMsAlepltqHarglpAEBJJXY/gybfeJVepK/vfZWY9VWti/DG5z+JLVEuFT
8Der2j8enyendYn5pQZUkUjjrWKM4nSL5Uuj+voxuFOLIO6DQjM2R3ln/8HeTjrqgGedYHESv/WC
b1uUrUoR9mdvNaXampc+5FiE53dkfb70It+PlS5PDnIT8+GOV+oRp8jr5GBboxn40/ui1g8XUO/j
YBf28oJFhdq0oGM7IEr8cOJ8A7SVW2pC+aP4GpaF9U3pmEKC0IcQoyQkZU9pbgvVGUOQunk5SxGq
rshH/4bVfzUICIJJFi2DKEiKFuEZ1H63krXHeZZyD3ESXFByixILRME16rogzeFNxVucknKVj1L6
11nKr8abbL/a7gcZtP6bK/fWI4uIdJB6wqjH1Q/JxSV9pHoRPjt+b7470BTenqACq8cU4wwnbL46
HK5mekMg+k3aRR36tgGwWkI8pBHlM8baxZB7T3kkHrrNF+EE+mopNjxECVNXv2jVcQ3VfbJU+Oqy
L9rtfG1d40UT6qiVI9W2UDqWiUWUbbH/4Bd+JKWLnKsSHSt+4j9lKKSuSfI0Wh47AAumJhqs3XC8
Un2OR6821ui62szZU1enHbrxBi1yd8NoVPjaUDcX3OmIDup+KVED3ZbpJtR6qqX8D4JpvXuch9ud
0SBw+sZCpBfB48wvZW5pSwUiKrjVuByeO4f5MBJIURHKfYs0rgLBd89uK6Fkc5hBk/t+SStIpP9k
QaJyrkfCBhDUkqgAyBwM774MGAHhvkmz/64eXODVb/Ys3ZAeKnP4rqvZZcB5gB5ZcQeCq930RfKa
wETLS20erxL7IGj5iBO/EP9T0gEXbGalBQhUoIIX9JTJEalH2xaxppcldNKOvKkjZoEVVKOPi4FU
GawpESQGxK5+gBcF+95cvAktbpusjgUs1KQ+F7xg0Af98ytglKxm4jaeI8833owM132bVKl0/VK5
mKQN8JEsS3pPbnnKTZcoHQMp9x3g3B2Gpy+dZxZHpxNvVM9ngw4E5/jclvnhGpGJbNFovnXt6vr9
RGTnEVt7OcCZX9QIzg0ylDYFWtN8ND8KjlZ3WVIZjZ03nrgt6t8O8ZNoMN7QZ+G0ZDQBTvEFPdj8
0qiKmymczB3WfTsdRjhZ1oH3MVWVuG6SM7Y+R1TN98Z9JFvcIkupsLyxzSn/r8YfFAMiuCM5ieOA
tWZEjq5p5pjh9gG5etlWFzTIN5rC997CPfVSIP2fY7Yqm+BFMtpweQaqxGQ36iopzLDwjLEnVrwJ
jHtqNMZwj5DPYs5x9qK+CVSJ6jLfKzLiCeosgn2ColKSa3qiaZIyORS1pIGqM44mUtFdeOMxKFpq
dgp4drptft8OX8VkthF1dqoJtx54VjcBzuGr+Euo77Azrie2nhqjO2WExn/x+t2Rccgsc1dNO1Jm
xIn+Lo+iwijG/QmIUrJW/lTf+3NUBUJ4c/bljYPEdAqJDe5gTB11l5J1WJtEaXNW6DCGPQQszgkn
X2ryHU0gz4mPHLruno9ui15qt7ftFcBFcDRH4Vtsf05vcvST472qbwYqR360di9OjsNalcHvJg5g
3Do163b/4PGvDQOgTHsz3YDk16VNK4Iou66ObMzomslXG/br4dw+wAVtjuAPOJp7MneZ36EUbKU2
BbmakLl2oe0XGk5E4CJekxERj+CjYWzzLkMym/HD+eeZCHaE2EPG3ReeeOt4xv1dM0j84RMLpk90
J7pZxXN9bkkLWkbb4K2ogL2JSjbvHNdrpKAWxh3IiCyrseYO7nbFDb5EvexJx2sTqBzk3z+lY8F9
+119wkExhKuijvfBwkfAo+1SCFvx48zw5U597UkAhu994a4DardFhb8EOXmn62Y2xP7+xThV2klp
/6fVJMZq8+5gbTFZ+XOn6I3ILhJXSlE461FDbCNzSJ/bcHWACAJwzLbn/8iCa0a7xnvGtT/x5G7p
+ep5oknT9PK4glUVWb4b96J/CME7h+98QKVBh2noT2f2Ip3mNXm/Ujx0bzXTnldd9b+NJ+2W4l+n
w9c0rVfJZD2aQVeOpSCnXq3A1oRD9HQo9YmmzG8bgJ/DS20T2z+c7lHMPpthd1REV0drqwBJiBN9
o+Z+np3RfwzmZYvSvoElp0NIOR5cbCsOPMvCsfh5r5PUdY4RHiW2hiPUoczXeZqaMmLPOYl4Kw/r
aZpqPUsYim72v3MNuPf9HMsBXKe1iINVx+jqQYJMehplc8KnZotxLqEN1yKU+jKDOZpHj/vP+l4z
X7JvNAQhWW/VgiN6JRMrv2wAPCAASqz9Hsp87KAf8Y5o3Szjo9sk/SbIJcoAyEzKXyrBOgY0pinW
Jeh3bBBTgU005G3kWfk0VWqF5NIuzgxmZW0lKaZpU96MNTGaSTuM3zGhgff4wNcHKeRgVKF6ZtRG
MkxQK+wr4Y3XDoiMI/ma0oN+YzhmdAD97AMQw8H8qtfxzDe7DLiN7iKaF6Ac9rof5Z+83p/QLKpt
DlI7Lee4tUvDPlarCis/HHKZjIKUkwqOTwTsxpjleJYsibWwYB1YDSG4n5ORbMpxpZ3qyZdweXJ9
RMOAUiX/JjoUT8PkiZZBzOAw1EUxPcqi5212qTKcpH5XOwDMgoAfJdM+8Xysv/nsKlNa8J9hkmj/
qhXgLYTbvC6YUbCJ6Q/awqQ7wcoQozumMZas+FQ0xrMo297ofUHySM+YkK2S9BgkTBXFk7bZPOGq
oBiJaq2Cyj7H9DAjuPSAM0dK+zQeECPEoiNjqvnzyyjOddR39G/vzMzXGeI4GRJmKHfjbZq4YTeH
msC1eNllzVp/LGy90ZWwVM4bOZ7poen1Xa3SH0Nu27sDUv7wYUwEnFw4bg66WPpXtFnkIgyyPQNz
BG1vDidWm/bZhbCsJtFMLwZTyNjzyUN6Eb0Iu6SRnqK3T+WDXACsDBkOohkSwYGgmZNer4SMLZ15
kFuqEQsIx5RCXazfyne4pO9BwOnOoR62hT4sNpCsDQWmulrCAnwy4S5dJI/6bYKllKq3n2Eq4Z2M
QbCMevIybbtfQ0uf4mMy4p/ou21+BAcrAsao5ODXSxCTbVQVuDCaIjrcybLa7QG+daqbtWXvFqT1
Xq2jIH0w2OunsIXy9sDQeTrMjYHpj6MgyIAEpmumWS5de06zrqtmxCHUpf9lizbgmR3hM7g5kPlO
hiRiy6uZETnYsVaQG3at2CD/joeNtg1N+DoU7K9NMp/GTNzNnaIMbiFWnUf//CVYmVIq/pbc2H1Q
Y2i+sXqThWD2Xq9lccw4gmgVqSmEVDJTGJuC3gQwnDh4W7CospL5Fw3AHQlA+cE7xpMx7hrS6e2E
//dkAzG14lFoZUi4buTmnLnyK++gL9UkmvuhO30sMkvE4CtN993MuXlbXchijs4jTrNZBWxkcLzB
nP9b2p0mJ7bnpTFEHlZbbUy32dAdTzaiauJOZnXoG5HxndKPa0Y1pJXO/0rPC9HQBP14MdiSF3zB
7RpPt1KPxr72THyV8w4ACD9mTBLYbH0AdNcG8CHapIU6RqKOrrJakwN30UHpGqB7YemZ9N1bbiP5
GpoXppiEbpoiLtD25AzezkIgQpKLdhwxFZpUW0Sbh0M3nK1w9X289D71rFbfbLainaitOpDLiZqS
6U3ao2Jk9FNoEMt0x3ycB3M3PmZWTrfP+LizcdG9mG6TcYPTMJ5V7Fyn2YqJgoxbZxbtT8WF0ldB
ul0nkp8YOCZecv9EYV1MBNFQuPJaZICXgI1J5YYTU8oEdorPT3mYSS2rq5/ias+M89wMZnwH1i3b
qWjzXxvwWrlx/4rW/X0/z/FbXyuVOTE4lH7N/cmzLQRYOXypMndFy0ujvdUZb4Csx4i877a06wf0
5qCynvNCfqhGLYFJGw+VpHHrstVfqaqVeJ+3VTEfUHajehEIIFgCStp3HhdsiK+CTewAT+3KblQF
7JtBJicQkZx+SkQLMUtbnVIH9JX6KbdkaGibMFG6vMSHJG7fJmAdemeVumCEYtAcThrhGdyAOgs7
6S+Tn8pVTpSd8kHnRG6jSQzhtkzyWOWY1uAmX6I1zsYHQqeNAit4a60BsKkS1RYZ5ev08MH4bpZy
BeXLFzwtv+B3wPPMzhc8qnlfTZHLEOr1SOvAHavJTr1aVzWjFTqkJG957/bH0C6j3xpQDzOLfFWt
6bT/qgq5ZDbjY2m0KlsMlvUR8Zrvvla0JRl3I6WK6lceTgowQpeHc8kiRtk6hhmVD4n1oo7Zypge
Nz9E7+/5+EtAhG4RE+kvP0uNtM13kpXHxHtLrb4I+7HClw0aa8LuSpnkmSWW1sIAFNpmP4I83xx4
zlotnTtoxbp2MDzNIho2/3CkcElHEs+vhuVKQ4uTDJ43IBOkgO/uF3PTSOKdckrsoIpIGNdLYttG
lWFCcSUYWFSdqebjvpKjZVuLnEAbyGTEhc9VwXxrxojUoI6WsdGJx6nfhu6LTr30d6UnlRilbgGp
fKX/ZY0CET3jiCczLCL8NhgFHX1Z20DIhvQACa4F7D0opCvH4q2aZ0cW7YEGxYIvjcqIPWxVoQpE
Whu+udRuviWWehGeaBU4BcSfA2AYwZxce0bDqgC97gLYbsr6IZucDhtMCuQADX6NJnn+LrLl1HUd
qXDWoAReJXhiiEt9juLd7V8pAVWSgZE27rxfuLd7M69qPzdumAGKtKP/fEP2OadDcAB3v7JYyT96
e4Ltd2Am7j1t6KpX35USCebehS4/1McNU9P+0x64orZb/zlZaDSZCVRWndwdHMjerhH5N6ojP/xI
RgaSsFDpyKGbouQmMChO8rnoz0zFa1DWZezIgFeQTXS171rEBZtb1o4FCqOaUTF+fiMGgWY5Joya
qJUzzWsWOMEAQaMGsyPDF38faPYAYuA8BnDLz8gXz+yd/TSyLnD/aG5HmhJL0M5Ws+oxWp6LRAk0
P/1nsPX3mz5tABNBVHLp622Yf3/KrP5QV+R0eRNo0tB3dGApbvNK2ZkkhxPSaEl2u5ifhsnELxgY
i64dPhHzSwjJEkNs+cMv8JbWjcKFgPyfcrnul8sZh3M1tcESYMS2iZy0lVFIX62fdHAxVZPfZZGi
Mg4d63uumAxRgg3LRqOWNY8wbH/tyhxaJ7XnTkvNfj5Jl89jyLwdPsvxuknBQ10VV5u1SMOHqUuO
bxPp4PWRdmwzjcKX7Nf9ZO5CrXxRxBArXfduEk/FweJckQJ2csmh7JHUYjZTnV6ulJJQ/iB7h5FY
pZT992oB0mCH6qEZt8waS9Mc4ElC3ZbgNpTnMV/KMfrTPFXkYitkXiUdUHq1Cpw2II8tsM/Q6NaQ
P2k0lF7DEe/UqUVAhH+RXPneYfJjvqsoIch1CHzwYnpk9yLjXmy8eKQkLq0y3I8/+3qXF//eG2rN
P3GziSxTVRl7fuX7N/Wb0iz9DVkO2fcoKl/xN/4Qhdj1xQ5W/FCIIZDNcz3o9pmgqMWl11QZEiq9
9MpA+Wcq+2Vnn4UVNuPCgvOZlDwN2JeUIpBZFDWwJhxDG4VnrHHlllf++S/PyE4ycLpB7lRt2UZi
/385BzBhlBLYDmjks99SohDUeaC6V9mNVirgfG3shB5Yb2pNxuOaQRThjVC+d4Ckz1GDcaJxnUnq
01RXkhCVFOPTnsTDfPulz1vHNbHvNDmWEufwCgam3NZF+ClqGyknHt42vJ59deqcAgg9JE6RQoky
ul2XXM8wBfxa85yCmOG/vpNg3qgQCJJUMCbzSt4u/AKt9zcE8i9hK1FVldSDxwXDRzdoiE3ddsTa
gJSPawQMTqL3bWajcsoR+75BTjRSmW1h35CHifDGpLfiShL4gTgxIKI5zaScP7qyEXlZOAftqsui
/eZOb1qKYj7Qjbk8yhF7mdoAS/SJoUVqRzLGuZlCuPK3amYJ4/qB0GjtFasbqrLWX+2GmphhffFl
OrHwCyvIeRH2hOGPigZUmmLWCtnfyCe0E/FB/ngz7yY/XWXVQsAJ1nNE5zi3w+qsWC1hl7Ahb16W
LyrxIxQmlzzvvKQyzRjFGymSTUC8OzmBDoGL/qmOjhLO9ZJtvMvhB9wEMkj/60t+aJJNt58R2QwA
i7NONPHQ6Ye1EMriWar/qkHH2zM+7Blzjxhj9tAUzjo2K5dGu9F7JlgK99kgnl43pEfSqAFyOYQQ
G1lBs+kyn1qhwZUD8ecS01Bti2DX12Qg6hp8zfEWoyyhexdtC+0SS79nSvaqThMnw7yt/CRndPQs
UNBTVIe2Pb2VEKaH9D3K30GKeacKlGeYntS5ZxsLePbsFipDTdZAUxGu/o5/qk39sPUOnsZM+RKs
N/9zt2e5LqzwvE0RUQsdz3DSozeF18YcZOniOEKS6LquT+eg1fNSZ8l3b9/HBJt+dqiDzDXHbZNt
AUov+P3IX0egQEsMyqfeatABXtIY1lNO8FzvH7pFfKcOdjX0nZEiB/JWr0H3DpkNTPhMvXfXz4/6
rUZi/SJ8yZ0IBkBrHWaQ9fWJf86UFF+fJwPetNQkwYhEPozLuLt+r/G4fi9SC4vyX3FQYAScqr9U
x70J17w7wk8s9edW//saa/tWYsNNaD2kO4dXkA+rd8Pkp+h3Lq6FNR3hiJjsFmoN6aioUfTPQ2xv
bhTqun+sTCJQzWDw7uYDDI+XRoeBaXZ1IklJNcU6/qR3AmZkzkXDFm50VCgo2urFtBjGtYiV+8MC
Il0V7UrXYo/8n4BsWMStYsh9Gi/kbhzrlj389hpJ3Xun2/qfvt+9WruaC++5if5TgQVSg1BP8+US
dSNNdQd4tuWd9xOpRWXIgyHL59ZXHKwcoppwQuveS3F4Q3TvyyNL9ShlUIaCtBRduGfIKCYYQBoQ
i5AyziaSYaQtJdirMVAazn3qhMCFA0oiD8mntWA1fQCpDzUZCle2y2ZvBNhOAnykxGfrXP1M1ZlR
kTuz33WKBBTYXLGTPjHHeTeO5uOJQSUDdkatZ3A6T7mZc99+1hOJ5y7r9SrQCTkZvuR/gE81yGfd
k0MCV5TPyFm80WvxHAPd2dct/kNkvyykEm8dZr1lBOCFWGlYak3H/gG0oPba/XzC7CfQ0ZGnK+/q
j5kkyH2spR+iTg4IPT2TIffiJ/vPo1jLjVmpPesARvVKL34ftqO2dy2VGC4Mc7fp7aOQPqf1UXpU
WAx+fK6GaUguDp4FLkfrkNG/r0v7rk/qAuNhzBt49D2z6xOEQk4500nd1P53E/Gq+7GWsFf25CZ0
XeLLATHOijJFLSj6gAMqdBndFy/HN0z3n57a4L/1maLJO93isFPt7FJAgFdqNhEaMhNU7T98oasY
l6B/XCKJNXjAmVeU3/YxMTiDIaLZDNCXBI/SQxpFxZyXiIsREi1/68TogDznf2uJ5jzEjAdLJmoT
vRTd8J9cwanH3PqH+I8htSE3w7T6DAyddUbj4LC7n8EQX+vpXXS51KylB9Pe6gd2RaZU56JJUnvt
4In23uuqeSJCmi7Mlt3AUj9woM9eVkGB3gEPxtT5ouU7yZ12DxFZBZMf5HNuYEaUx5W5KLxEJKts
gwH7/IW01hXUv4O2EeNXgbdEdpjO+q46/6GXemgmOTL81AXVsKOduUYKaRYFJQUrdrn8D1bMyViv
IDSOHRa1q8hyItL5j36Ev1nL3mDoBvIDtsqEsceoEiNOWi0yqZKC7NROXC/Uqad1XbWjamo00SEA
eB4WhX5IClbYa4VizZKlwUStOUbrUSW+dXeZANGR5pUDyPfCyweQ6Rb2vnmTMSF9uGcBh4dFOWm/
ipZWg2kiOTuLhZpmspvqXXn6C0J7mifYRyNm/JUchotPvVhRymWh+mLrMDTvOtYZXS0ABsE6VMmn
w3I9u6/v62FD37qoaEdV+pE1vQbLZes44jnNYz0uezxdZkQ1YstjJh2HglksnJWuEPt9kniboFZO
atA5GsyDMQrHX0BpXOuWalyqKaWtFKDI6cF6krY/OfYBG2bj1eUk5FkeOPk3CmK31LWNULny9s1e
hamdqE7hEaXdqfbCYDAINcmJo4Rnxle/1Z8gxB0zcR1WtGfeRhwFKxY7/rmjOT6+xipdHzK5lTFc
jPNNs/LYv4NYRxbfte1NzQOmtFRJ8MblPM1ice6+gceb9T4j9Ax2I+yUdvFK97bZwniP0r/4XLol
8UQppeVbbwAZoUgVqMkuvOYuHvXSQhUf0Q49g4U+7PzuRXbYq5C/kc9cFPqIY7L6oqqxJqoE3LnK
cMiq01o8Ju/CxzXTlJJknrIn6hscr/TAQmfj/4es1FtlQQ3Xl0aPllJgue3rruUMbiVPR6TvX+RS
UNBv3iUz42K5VJrBSrXo2dFHqL6DAiLCMwL7N50zAM9ixyc0ZLpqpCl3t1+GXZUakiOEidlILN7i
IWdX9Unzqy5El8apy7JRPEfsZT/7V0oyhtuHEUYcovvpLDBaS7scvYwSPfSUMx1D9vSEywFeFooj
i0JrudD0g07xGpIuTrVrE8bhWHJ7AE0hijnVkJsl35no0twZENzhyzTf+lzButXs1mXWGTTHnmaA
cwS/xE3jWJmITDgba2MDY8riES7ckZcisnQm8c+wEq9ssKNRaKGu7nOahpa1PutkK1dDCV1PpgcI
yAcoET1deJxiRgwsoZvHZ7w4zRCd0+1l0qua3mI+9eXSQI7CrZCtkxgYiV5pTVseLBJedSsuw+w5
iiZl7iIWabeAEGDAHKTm+2ceUdgsPA7kCQ82Jiys92/T/9cDDJp8+XEmJCNEEoXO/+SUmDzGwRh4
oAyxbopuYj7aGwmbKpDRIMijF9Y8pDxEZ8l07uB5Sgf8tNOaNAczdY026iyEjy7K3/c5JaU+qjVJ
R4lGOHLqcmjf/ONqV2PS139fARgHNENkb/l4PZFTAlHnTvXx4NJBm2WpNA7DMD4hZDYBraThTepq
K1ilsHbTYUSYjGeTyczTyt43YZV/lYTbQw74VZ7zkZaEhs/z1ACP/slWzdyg00RCRGD2oku+ocSa
Dqeuh/DQT3+OCId0TT1ANC6TRpaQim0Z3FwxqKQXbnJBwn8vJEGyWipmkZt7S2H3a1m8LLGTgzD2
3IXvMGdYPum+A3MJWCEduIekowa7jKuLeIgt+nribmC4vBshNlpktJgjtR4fDceQjMi9CeQWIEgC
TfrM7R5WCZTaZPJfXhLKtqjmBl5EGh7z6r7TXC9pfLHl6ebL2irGs7TOdSmndRKBOeZ+I+JzkFrg
uqAnpnwf4sYGxx/8ZUExnqNjr3RNk3z36MO9rAg/iJffbhwaaIFH/6nGJBNAOlzcUAOYMA5JXe3O
6xeMR/OGXi4UGNChObt4nm0gttYv7RZm9kqtVf8UuSqFKq7MG841fZwunlBhmH3/AwVX4Tl6Y7ZD
tcsSs4VoMCwCF9fjI3+foDh4i9dibjbic8f4GqIwuE30boR1Oy1htO227ZSZxpirhJdIXplKcLO1
aY+61zcjSJGReVJ2c33ykAbFMp/jvsreSeA8lpo8r4auVUh7G5wJSynd9QWPhpw5UEe6A1wczna5
74Xac1i81TrW7S47ATAPcOKTaTIO7sfYAkROdHfmDRepjBrykfNsnnGj4rt7LiNxvze9TTrE+CCq
1dS68xEqo4sZ8kKTlT2dFd1drJjaoGGK6oe1HGskaSa7KvTEi0y95rq81pZQW5udK3Lh4tmjHvYq
wCT0dROzvSfQlwReRj6hv+4bcFPqkI4XFkj99Z6Z693KLRnzNrKhafbP15XI4G13KRwjOhJJ1Gsj
xTKRgHdvsYsDnrCePi3/GJPk8mdrv5WOP54uUYG/VgfCFaSqJET/Shj+B0ixiHUxXDQ1j34ABtma
VRYNpnC1X3GZuVymL7m9oOtIJe7g3mepj5PsIOI1fsW2zy2iCb1bK7zC/LxR0GASlkoZ7QC2Z5Hy
5Q1bp8ATXBfQ9COF8vRPqHVneP2Ldi3hLT3X6QA4y+G/dpIa0U51Vbs6P2LC6O688dk3ZMJOoFy3
tJ6FBosd1AigITPdivOVA93XzVs8guU7gMIS56FSr1vx1UihQMRblu5cVdApx7FwEbVUa5PM1F74
YLKdpCaJhj89Sge/KDC9K0N+yGjOq7D4+T0lwBelT/2gy/jGDg+yxZjrT32/e/01uGXTsniiDLim
yT/DjP92wCZjozKhaHCLwkKEIivNxdJ0YMSTAwLQcSKxyJpXlluBGcEO0C6G9iNUxkNCBq2vy3aD
4G4HSo9H+6VjpWceYVT/BcCuf8rIs+0JRPKSEyE3umlogwQynuNex9UpTSPuMCVU3leA/2ygvXIi
wIyb/iPEHUKFxHQc8nlA2M3NqcFa4K9vGOQjHt7kX2ugKTcpl6EzOe122cVKhJIJK4ksJ2hRNRZb
oMKMDw5wyrRffYs+PR4SxB+fOLqR5IY76NlAQh10fPwxPRC+s8giA/Cb1DhVsrjB/+1EdgfuIAGA
hlxWnJasxwyS/AJlwe9umw5rTDFUBOvLLbaLdieWlYxkDRcQzymC1TGJz023Hj1TxPfzocO+ub6A
Wa+/qZQYeTn9hbSMdh7zGzASYTZeX2EEmnz85vhTVdv7twTKqu9K1fPpRNrxWHPVbsJL+/O8J7nd
T4QVwFzLRkaKQVdlQ45qC/FxrV+WarPTjhPefBIkf5q+P8axu3DdT1a74yG/JBByiBxRCQF/1NHQ
lyPH6tRAJGSn1/zzl+GT2aMGkSNiRXQWpcfeYPEDpnfnbvVvxRz8L08nHyuGMBo4R+P923ziQPo8
4ZPhMMNcTYAoN/Nx5YOBcJWMAepA2waGmTQZCCvK8OhR4ynHGcKSduV0pTkERCQ3APJRK4pyGIkX
htyR4OcuhU3JiMmENFx0VgZXdDmlY9MvufyL1DsSjkDSvpxFl2vBJvQ04IhadZdUkIMZ92tXhn2s
WpzoOWUzwjFxL2tA102FY8U0lForPovp7mJNGkA/XktAQPKQ7SUSKo8hwRDso+Y15LmHV/TbQ2y6
JQ3Wku11sAjDdRh0Kpco+pFNpbSHBMwPrgQZRKvnVTszQt/OAyp4IULbVmdWq7harGLkJUn/PEJl
iQCIFpgIDeHKYLpVWvG5knlvCIu2WvLb33u7Kcceg4ZzSmsAwQDwoiJox+qxB/8q06gkMjxNp+B/
yhLWSrBa+QkhsjzyXw1/NiI0S8WwujMK5hh9SxwptBcWbJuWB2oPRhDpHr/eQPZk0i20LuM99pnN
Gk6jgYV4YNMQ6vFGLVXacPPdQJKTog3l/6/BOJmkOpTNYveqf2HVK77WSEExDM7nNptqP5N52LSO
faJghdFI7cMZ+zizguzV5fz+q3GMt9uAKAWnstwq/w902xvQCz54Paq7nrCkeJOTJ/BEsORz1YDe
ZuzhJpqMAT8F4mosBfuaSPtWqSwvwg3RlmXHym+kWsz6eQKnaop5vjgnN3bBhwnK+Fzeez9ZuN1/
UNSMw/6vNK6dUcVgpp+TLVPld+tK0xyRDceBb2TBKL8aMKsFm/M+q+ensActwbzmzUeilC+ldxFo
WdCnv6m5kmyIVlVRAS/3ibzojLKimQ9YtR77ICculLHvenkx+RuZS87yPMenqA6LwdW+HEqu3fyB
ZeWWxdbZItvsKEQHCFbTC0bk39XsZMSYpPztOGYW2XFDvwQAtYVGriLXEmUDpM+GpqfLP774wcG1
QhZcchDAPFn4bOrpZ3g7VS208VnhL3lBWAjqaH4dE5tGBPUJxhsZujsSZGsVJsWCrQ3Miuopy0Df
y7IvBlE5v7yWmSeQ3bq/m+SZqX9vUDhl52PATtHSttulGurUkVq8L9JKB6TCt3mG23z99D7rAokB
4xAScjo8+qm6c0uqPxea4chmrI5K9LimqRX1ZP9P9dmJgF8CYFrhe3vf0xNI8Lxe+5WrgfOqBoeh
3TEc7+EO48zXrSO50Ngfr6JSwgQSOFGzzJ+Ppnqgkik/djAAyO4k0Tt5Oj6mhIAcOKg52bvYwNe6
EQM1s52OiHcfdDRRGjwKeLscBYmYapTJE4UxeLyDUdElHBxtKKGaNc4VL+SdD5wU1OUQFwj9oe7O
s/owF27ic1epkN78AKQs0u7gnFDxqTFnh2clCgUTt0KleDPg/o7V4wWp0nurVR/Oxh1/IZjPOkUm
IDkC6kW4kY+0S8SlDtpT0WwFc/NcyUbWCZEWTH59VWw5zgDsXlTdCbu7V4yK4S4F+E9RFxUjDPRp
WXLPloy0o0QbYnwGLr3+WQnuBHltql0aKtdukO9dkZ/OEr2UlX24BTqDmYV9tTAU7P0W578q+Jv6
MFVYTUmcmSTFg6ieiyS5QXPUAI0Ci5snyL+f0si8WawrcgpzifDYELjMnVYOoc8m80Qw5G59s7+H
6h/MKrQ8GnbSmINIExLkiW04IyMeSrJVDNHisR1Bp/hFs+EszMUP1vM19XR9iPXCxpwJhTj9TjGe
3COzM99ac6j3CCqGmfYlcPfsXQ/Rv6AkG8ABlJQe+mHluqe0ImFOf9BvU9QzUrNpfvrQOTg91WGo
26jpUypD/V5Z1HqIox5sdSjij0Uzd5hEoBTFhu5WUYtmaspI2s2Ao2NUOc9YlslfNrXKug6O7MZz
FTnIYflsFaDVwuvEnY7zCBr/H4ZAG6wE95LxX3lTcAoJc817Bk/X/8VYNlQ8MJXPEno7O78KOcb1
gkkGycb+8QoFMEOTWRDpU8VAq+AKRPfUFzSqPMZzcAzfDqVomisRsRtb8Kz0pOdctKi8DiKQu/x1
duK1oWJrAwHBVEHxclGXGPKeH3FagYlvwTmIIRa7YjDO7L2l0BkYTXWiJRunlNHB0feaySZgQUd7
/V4di4Qj59dRLrobYAPQeqEQj7OTFoWmg43duNIISCSQmwo72lfKAJznSrxTYcwcTI4MJsDV4suG
8Q9jZRryON59Na3iQT15qkTfAPwEx0WbYEjxYEgE/RcPL3rcNg4sCjFo7yPiV114HWIIVFTErWLc
d4TCbuZV6uU0LyeeSLaxYkYPhZxXgj7MMOLBzbq1i/Zk33IwPzpX0iUeREEt5NZTsrhM91cDWlPH
s4uQZCYJOVd9bYJsiRIKGRgIeDfXBK5z/uIYnj+NLAL9Z7kP2OYba24a5rRsk5uAC60WJr40jULH
L3+cV5dFjSJlaj+42eFBTWGaUU9vDJx5EzqYOHAwqkqygPK4GqZlYKqpIKz6NFMk7ptMc1yWxYgf
kbXGo5xWmGDy1/wakrdadKRKOxvCqwAAbXxKyxtyqJtnhXNGLm56O/O18o9Go+QlBjx8rQqNQFCs
aszlIG+ZQ74250wJwduyIuZL2daTjYVD7XUVquC/DbEt+Z97e4/Vkb6DmaQVlbQ0yrdBja8ODdqc
9b0V0XEKVUfoMtQCWI+gA8KPGRXKzkKpjr4z3BAHivjnp3nOiL1Yd8THNCwuF1UDhJElCQl0f7Fh
0p0i7BzFeSR9pybXqL1QqEO7gqTXh2QIy6EXNW/TCx1ClPwwARy78H8/YnegGzJZSk3sBz9FJnmx
/nRoRuF6tiJiFy/X2kU/qLAc88/SJIlhFJ2useuuhwkUuwS5L+V8kqi6UjuT8AcUYCjLHO22Q4LS
46P8qDEfoqG/33IFitiZnb9GeWXQfk+OxnA+R7s6jC/Pnw6shjQfbNOQNsyHV1n7tOp26/PZZF4u
/A4aELYaOtxkQXqvJ4gVCcQEC5jXQvHy94o8f0VJV3a1eI4PyzS1edtDbWktEB2NzzouuIWMeMY+
8pBcpYkc6V4qE87350FIigfGlGwvJeJzAFgCZfo9AsqNIKuA/7jSaATMqXiDIeWTRVZotkURtaa7
1HlIgFnADmLS4faFF70oiq/69kyifOF+V1YqSGB3XBGEQOv/sjFlbcwPSNVeFv++u+S/CDdiBqYV
WNotfJTYkvf6WL236dRq8SJW8L5cOIa20B1FmcqfRxK6cJHnaBa/B7zOp0kldhBriyPRDEw3kijQ
MebwUnlIiw2hp4hrdOYz3C4Q50MrD45tHqtEM1EYEa0pr4tlLffgL7kM4JLGWUBazhV7Tq8hPPdI
YAS/8u0RW3Ai+rEahBwzVwyv1HqKw49iBo7nwwIccAEMwFwlRwMCKg9D0IfFgxu3lr1+Q5VLYU7S
QDF7I/dZbCXeBPJqVu3hVngyHNKCh3Ir5byDiXDWfULWYO3Vhgd+4QG180Dbim5/CdU20+zZEXGx
Zctz0NtUM304Wh8Aol+qXh0mcSmUyVJFRhYwraXJODq9Wp76IF4qHr3gbkokIJtGPGETt6WR7zF8
+torBYQV+YPEHXI5ANVr5S5HdpRV0mtgG9Dqv5XOok22wZ06KnD6h3VrPuymj+4YiRxz5mempA1p
6Yw0jFZwlmUnduItbjWedecboMRgEytKevbw7psB9qQBWz9raTW/KJtrgaRgGbcg6ebjNk6Pwo+Q
5SPs6WjZsQJVWzmqHq1CMWFdo4Xt5xndNBQDzpDLdO/6J2pbxMjundadoxy64wOO4sqTVKf0knfD
8+ljMxCXozipS+DKJXDCSDtcwAEdv32cZClA/8yY/uORysjXRVtuhlteU2qPrir/dEcgu11c1946
luV1G0/lF3j64AAECSO9RzZm8cgfDicEu5FkKMwhddFnoLs+HpgYHsaaCyOA3ngSdr9yxRf2/GdF
HEsaOJxIdF4VMeZxA6JhWIOeEpdOfcdvKcRK09mWdDBBvHZFgpC+xkyuNjzVXRYM674cGxOcFwGX
reR8ZqHsL50K2Wh5HhIPUHVl0LKiXd+Qw1w7wo7j1Kgh94jLG7mZLh6k44h4n90sy08W06EirHVf
jMYgBuUfRq8kQSpRuyWIO0v1ufGsqMsuPsFkbi3ModqvstCz6cGQNC3BU+jIOule1txMwlaUWz1h
sSw1u1xuqRLEQktg4ZhO75maUH61f0i+4uKFunvR3uZeNOlVYh1Q0O65iCIoxG+sNBr6Hvyz6134
Sxdf4SOVK38Z0B+4rFp1tajQrfoqZn5yM4P5+5KmopMn9DEdQKjXGkLyqNBA72TpdwdlUAovrmmy
7TG4stWhaouh6lTOBZHx2qUddmiFNeU6Sd/0DUnDtCv6aOcjSIvtd0pz65o9GDtu/6A3XC1BlbxN
D94Fu35TxA1QyN86X9ARNQyhPKUShlCVCU3j6dKczxShx1gu19Xn7Ozk3agWgReEJtBFy9J/+BOe
WYPZHS3QqZJ4CnTkrpy4+5OAOwXP840QBiKCz8yfWGihLPKNtzk9rIj8VxH996RX4e5egmyqOWmM
JaK9iOpNAnBUNrhDhXo48Y9dpjZ/UPpF+i0nzz/Hcsin/Y9i9TxL6mDy5C2JxiJUGLH1ys8+1GWe
C8Hp0k5nSbmhgXJucAqrcnHqEQq+7Ssfp99jGyWl71fmdwhlwCU6Z1qtwLF+SBFN/6bh5XxhKaka
RLUr6z2W7OUUzU2lpOpRhDffAtrD7Ck9gldfMbbU/VHEXA/vMMVD56rAksCWHGRLOoUep8QubNac
dtDtSlIrq0aCyfzxlwoqlrTsVHm/96ehAFKdBmZGR7BwSDerv3GGtM3Ysu7bppE8WaJLLhDlba+P
/GgBRRJu1CIqb+j/72RL/on4pazo53DQBzrabFS4CAPfkRYZb1Kram6nkPEbR723V3MDbqvFW7dJ
yhKG9uRXxyWLJA7uCwx9NR/Tz78sFQrI9gedzxh4OwRo8cEl0LRx2EqPBYC2An/8wtQ9Mfgix9Vt
Nv4k/rgWxxP4RAypTWd01rDlIGwadlqbVKzrWX421yq5eVHwjFpMp/QivI+DTaEVlJvH//LbuXGa
spvuFMnU7Tlc+NUXFAdY54IZmUFXSQ0XWqGSmFUASrPw/wG16jwhcITey0oCVwqXsg+ccSZAqprD
gUYKVX2KlQxCJvo77XhAYyAWCkmOHpKFDcQcTLAA/s1RzIKERJwV5/yRl20fFhQY4zZ4IWA0EcsK
gaWW3k8UZ3N3Het/44NuxvcbLpkLA9NmHaTrqbfmRsPQJrEkfjaN3wBrthhjSzkwsM43vB7WMGki
xpEnEJTs2eCnqxXP6wx0BT/ZQbKj9qzqdJEYR1HfuAGWRXFFoEnTnux2IA3lRC6U4V3XaGd5m8ul
oqfPm7yr6EKVXTcHda6XM579BxWqkn6Ca/en33/nOXIKEi29dJdJLBtT6W5Y5R6f9BAYDmYKiZz/
21Pe+L6OeUdMJLmmFSlCQ2ib7ILFmRBrwyyB9MEk4F9YOIoHI6Qc4/NscFId4GF4R173ir/TFgIW
FP9NqX/Y+I5i/XJAbG6wmEnAH43usuepAEjS8nrbbwgaLCISCQDjN6agI0CrQVzlSFMflncRSrz9
hSEhsHq2LRHGN98ZeJMVxIC9sVl90D7cXLB5hZgBVhIyIxG3y4P6BO5yQVDmodprbCrbSkb1pUH8
uJUhz2U+gEX8ERqS1MXTGl321+Dm0UQjhR7Lf7eBaqtemsxPxo94G2hCAMMS7cmv5whqVO23io7G
9LbJEcPlXRlypw9tDY1UVvQXqKmGapekb8J+Jo39XURUIzEIw0ghCbdVZ8/V9VqUEekRBHnvCfjl
Bdc/+X7BFlsB9XTTMNO9Fr0526aTyZra/wvioldsdQoym9ehDIT/p5J84gbYg+h8FNPokr2Dgus/
SSz3ZBnMdrCqvAvcMWh5WFZC3UDRYJ//FUNPwOVxwRmXbybUL3/h2SLG4fV3slnIcz6BLS9jIszT
smUQyw5Aqhh6bSZopVBqbjOThJf/GKA68kPhJ7PVAv7SPqwKGW7GnY3G9zm2U7+KCpWyznUBf0eF
AeQPHWllmI/w1pRExkd9xiIN5RIzVahkSrX0Xaas5aLg2cHHtX5K5szQ092gsYnRSwzlg/N2Yabl
suAKBUC55bQSTkmWxsQgdag/NWEBG0n/kRnwQyGA/PAkDhjwzAyuMJhCsqRUVIxOh+lbDfBWbN3E
UqWIjOQqK72+PMvhAooehbgFHtgxpmqBne5D0aq2Oe+nQ6krVZ+14TMqvXwBua3dxZiYXLfpJ+mg
SszPvQqy16bwG6nVywdqsVuUG6J2o0JTphjVx0N+oQaQ8uoNXB278Ik71NWHvqg6AtCfOi2VsMQr
YFbkUL7Ahh/hB8SoOGQbo04iXBGcgbbzTuNW5vdPep+oz9wz6pzHAu9KN4lKpb/rZDz9GJI9RLku
cMjad/zRtOdR7ocsraFIrZkfLd0YGaZ3MUPg+6pUy1HkoFEgqQibsnqxzrr39jNvI9+8ldh9DvBj
lCf8urOSawCuJvrCLNr5zWI174oXLm6StPBt7XUwPke0lYRVyRqSB206JuuxK8IoLAoh/L9sBlul
jd39B+BplvsbWMCEnMxUBA70X06iV4lO9AVbbi7VbKTYiY1SGXyBPeCiWV2mwUJsRx4ZorwaMY/K
66pV3NlQkirXSvg6T/RZSGN1PtvpY2bTsyEWMWhFRIBBfUSrpA6gGc44TXj2sjWDmkTnRH6DyXjt
xJEkyYZw16/ehHqGzWekIMn6QbgDGLWC+Kxe0UaVViOiI71FXC9C+T0x+5IRhyiv2YWq0mRhSkos
50Uifbyb18BY3QLIeOQ+kwnXxtROx0SuzVsLnNmJ3P4YrQUHxPLoYCHgSQWUy7dr9mJjHTPUWYqq
0UMy6UxzIXGBFdzO9l/FFaV3wqPvLKnXjZkhkkdJRCxhEzqE0PGaiqikvMbn0Q6hQ49ye5Izeep/
s3YY82oJ+IoUVCRyqpBtHXvK6Ktn8CKCzIu9Wb9aSyDnQWgOWa9ql33w09glQLEIN7D5Q7Afhs/r
sZNCz6EP3MQ9hCN0LH6tAseByzNrP18MzBwRpBlxAgfa/0W9Uu70hJ+oiLmCHSadpsJfc9TnwS63
53ZSMJG2i3p6rwregN97khAxJ6guYzL3H6R5cXX5etUPKdL65wDs7a2+7C4PaM5Lt9aeu25IsgK1
6CTUBTr8M3vqw8W01t1kwUKpY75JF0YNMiHbJnLME/zHQzOxFyhtIJaLppn13/c+mKjR9+fBC7ta
CvahZ65jASGDdhlxh2vvG+Ebg0wA4U08oMmkQ+Fv1Z5Ky/mBuZKvQFUd2DGWWaUz5l57nJq4vT9y
t31UZ30CF1tjUQec2YL/T+eNdmoAfhcXQNi6fevfV6xhRst2MFzsIFqhfxlJmbWNWNz9Y8s/iNRR
qlcgnXzoE3a0C9xr/2FxMwkxiO4FAmwjVuw3iIthAVKuRboKPu2fdG33o5Fy3f7G3y/kVXzeiUE0
vvf0fRfTA+9uRSGgq+oLcOIr2HcSqvaI881NYc3t8ybwt38ZZdhHpuFw3cLq8uoMPnZZVjQvOJ7o
3HxaD7IDndXrmvw6lX5Hh3i7zozIx0RMDw7HHGEJEXwZBEe+fAg5ksn9tiYxho8JQQOo3r/13jkR
od9h8uszi3j86WanbkkOZRWeKvwP6rId5x5eoPc2RBQVmlrtbj/SZuxvM2C4DSCnunZZSO9gDASR
9uHfBEcS4IA7R5TgxC0CYf/cjfPxtJSlxjoC1gIQX3Z+uaW0FX/fpYAYnM62JYXaNjr/M4dnBvCB
uji4+h1Dqz+Zx+hGMPCPe7G5AoDwtMaK7SnjRTKjEBpXDdOJOS34qvb9bkyU/UlYdHDDxz6H5zd2
jtHpsLVs3jWXgHbBjkvX58jqtMeATtrUmko/3iu7dhhvp6QNWcwtRS/VT4quT6Z039Syy3OinR97
/wwI37Ihi6g4ETVhVCdxWbfjdxJ5WdVGPfTnsqcL7qhxsZfdWmXgnFV+25cXgNE/yexYjRB3bgGi
lE4Tta9CxghOdxm+iNAbb3yXNoWDVMnZM95imIikmaqyLSuxhZJDP7aNmH1aS1OkjAAzR/12/VfQ
6R23ikz6MDnczRJXVhlZUP37l9TRCFcJJULFT9FFkwE9Fca9hbocM7OVgzjzcjuWdHQAwUgSAbKf
nOGzHNuW7ZyeXmvKuVvXlqW3rnF7l7joy2UxB+ouEfCvBuKugV1slbhQtA/eEUdcex2/86sg2RkL
Rj53OoutAYSEkXDZ5gB+DQpEHa9MLjq64cHn7hGG0OQYzEVRy/XBtzU2czjUQ5NHHUu+teDv7FiE
xeeWAPZv+WpMo0oYFVDt962pJip8pHhVLNioz+1kvj2lnxa+blKqq660HgTKmO+KxSZQA7dNl0Ib
45pTF9H68xrm+6MMbKCO253kYhUhOL/vSODqzmti8RPp7hMoWSyynfb2/ryMpqix+7N9USwU/YIF
1ct7w770wDQV4rMfWBnWqOSWl73VaDNXLJo//X1yfGDqUfPsqJEo/yZGxlhQG44dY2Q3kGrtDY9E
I19Ubhsbf7LgR6IcW+0xV6HCYg7guDp62rvZaF53uO6X6kCcRZCa6+qyGhnVWoOThAl/wvmtaU1p
9hlzAbvPY0Ek2l6DeamRTwmavlvrXoKImcHrhdG3sUN6N7V8u7URHVVih0H+TM0NcF+7jf/3Wtm+
guDWmeTo2z98taZZJ8SFB2QrtX0ZLGJf3smtTz1mcZDQsp7eyj10xsZVl59BEw6FJkljtYSfMjWu
jvsoZmIsu52wX12E+1iEUsfRnAFt4HwOWtNzQad7yS9AYbdzdBBRoNR7h25PCjEoSeAod0OSIE/Y
nDOp6rxrpoNJU7WQuL4KHxWkWTMtCtJvdAvAllZZSP6NIsp3ad7L05ytbOlk7eEW+cVQz9lJA1Us
VzuNEVFmoowsIMxXLGep59P/rG84fA0dNWsztFfpx+sNb+/jEFfaac5B7RDf8iDwe+1Qx6u78Y2v
mXWZHwutFVrVPyopmm3JPeMupx0t9w6pIpH6XkWpoZ10wkVTFF6WA/VGfVBRW61JBx4yGMDGPCCQ
XqzpDjEkTwg+VrGNAww0ctzQTEtz+L5yP663dAoIb+/ojz8TBKJKT+KelMVMWZ/XFbgPR8oo2JHh
ngpyvzCDgBuequvK+Qu0thRFtnr4naLCQWXvY2faC6FMIXRdKi9+mxzC2ztOYVQ8fL7l7mEUsfF+
Zffk4klatFpW5AeHyl7q97rAsWRlIYTpZ3Exd2uik7oSn/hGHLV9hGIPh6n7QVodPb+E3NraWS8d
buzkV3ph3oLQ2+1IIZFZYhr/ThT4cmuTx0bGNYso1dRVtKwZvsOcXSrkFPpQX5CAI21Sjh397lEG
8bVWpPqnPZzU80l3hE5KHxJ0FKNDXbWeMP6BS23rKxsxlHKKklJkOX7Swmg888yQSe0455WBOgMW
Gmb46G74Q/q4lN7R+Lo81gu7P2j11H7JcO7FoQPsadus6Y0CLOB5DpTpoJbJATRZnaJojC6yM6W2
7AOGlk+MZXix+8OSEJRcQIjuuH0TxZEwMyjRCjLsbfYsUr60RD3AyqxDmk85TnUHV5pzWNBM5rfY
pxaJYtNa+5/hWCxoXPw+3LyF8IgtyTr6nrpaGH2vc87lD2EO0zv3+qiRzeHmjw/kwGdQl4m36oEQ
7jaN2gjqP4SbNVGKa81mdhCL8v0gIkaJbuXF4m+47ak6iS8b+7OUqdRCgkJRqNwvKsrFExm9EHi7
CMm+GUzBV+MgVY7LbvRFS8U+TBuGQQh5+xYyJQkGBLttGv5xJJnQLve/h572rW3C3uszzl+Njhwe
dlWsV1JqOzJrSU6BPkgavrevLgfUt7SKy0uEIZeBmKBu12Wgx07W+wrv7/Zw+Ts+Ejn+nkiGzwHO
Gf21ocmWBr2jEyTqpTYnIXyDZ4ukL/tFwpgKEtJaxyzgFTZYtZOeBbE7DgEBUxOb2uNJMlAMz7K7
XIx+FGUMG+Critpb+/Mu5TtjPpa/CDoiYE19sgBU2aH6njQ+N6hJ9zP/oLkFalv3GgXu+jP8MNA1
F+kaBoTbAO2bepbqgY2M115Geicz6uNeXZaQybiXOuXgO/1LD04F85vYCDFERLOpoxhYdEEkcxwV
m6B4v2iFlp18jPCCE3JMN5dDDMHNE8giCapOWHmUc+KzgIZDEzpo9GEQ5FMcgXQJe0sCN3sTqk93
zqC4xvEmcAoiMHDh60ZP2uu+uWvTgAWk2P4LFXWCJQ192tZ5okjbyFJKVI1szs3bBFu7CoO4pFDT
S4BVcuckZgH18Z/FrRPranUX9QdVB/2caQdB6VeyuSwsiLzvH6dL3MIp/HQsj1QGv+KQ40A4wnkU
G98Fj/iIvjylquzFxv/KsPBGIX0nflS7cx5w8FVMjMs1JY3WbV7vRTcvNNlGtzRYCGhnt072Rdrj
/gVCcfqhQ/iaqD8b6HW4pnuwPEgn/2buC3oFt8V6T9Dc3tN6s2h8S9t0mO2emG7l+IiWNZTet6GD
/BnA+0cVKyTD5jLE5GQIKfHpjczvCo4rI4wBV8+q5MZq/IWHFeCvCi+hHvkwbpd/QZsauDbSbTDh
T0C4Ab/MZHBeV5wkrP5AU5RVC8mOUI/S43aM/swWu53TOidbRrLG27kwUF3C/zUQCtL8nfdmrtcO
tihGxCbjCc7Df8w3sACbAVQNR0Hl4YuhP1igyqP6afetppemzuf0CLCTy5YhwuiEBe9//GzRmm1N
qiDFTtMiiPdsgdqYOvEU8iA68GB5jyFmrxOmIIlSIzcty+Rx5H3WnJwrFxZTu1PK7lbyFNdId24X
meGYsvOoMbaDboxJTW6SapBEk9OTk09Y/2Ipcy7OBo2MKF0T8pfdAOnY0+rbfZ+sQeJlxPPQ7ay0
avMRTDD1UhrJ1bZgm9CXoJPfsOiy8l1x/M+T8nHrnVdlFFVfsNL2tK9tzrq0umX+qYZK6U5TOnH8
sXernQ+Q2xuNYFK3kYhLsE94/4m2bWIXwxFkYucNjX8rWGcwVJuuJ59f1vczW0caDzMA+ItA6JjG
gJoyKAWjgOBhf2aRLEfsFJxOsOEgOE1QZ6udMXCQfeGmULQMmZozt3YWvrVBXDQoZXaE+9kDpeNV
/KlOv0J67qesaqJh19V/UdFfUucBQ+Q3GdvcrlQ0nnv5miWDE5V0fs2La+EqUMjD6oxI0gI0jYc+
Bck4x2cExjCX00UpRtbMIh7SLLwjpjOq3jSD3HicHnALKnTl1e9FupChz9XsMUbLCQrg+uuRwxwL
jNpYqD9UXZMlQroTtpDj7HQZbChh1pXI3+hbbwrlHXRrz41EQzLLN4uFUKtncFWHv6/vyCqOoV6U
68Hra8IlAFj7CWPGeAhLZ/ZbmKWAygvtgc3njR+hSqi3CNOrRAB9aXvJ8hskNBdIRs4xdYEjIavC
U6Y4iHdcmF6XmVFVGL1EuZYRzdy56wkjn0VOy+MLTa3/uJyBWQHKqrkFWEHIcsSzffl07EX8GTLA
gsvnPwFyDEM4P/tCRiO/muS68WdlDPGQMVb8z9GpXg1l4q/jNh6xjYC5MbWw/rGOqjyaWPhWmS/Q
geTMsG19szVmwqL9cpj1hxSM0orLW+D3uWRPENsMYOdYaaw6v/MbPRxzH0j1QAGfKWRtU8DVjjdP
3xRA9zehLCvyM/W+v7FOkSeDi2sdqeMXlFCnXeuk4aNXnlsPcBY9nfBB69FtsrmuS/rxium9Ue/C
cSns0QfTeV1/o/FubCaYyBDDs0rWCs/P5fYx1g2MkXniFtn/xucEU/MYi8qsbWrK/VNa5aXfmIsp
aRcVP3kcTojl1j4FdCN8/NjU3Bc2lMvq1xft0XrjaV2RyYS+PMirU/dhEDdcOMpdypa5bmAs71n5
awUylWkxWPRgFy/FLFEuohz0gaweruOrMvAn14RA6fS7AFVa/iUwNKBuq/DiO/nIwFAMb03i0dbV
stdLGnnBCpkBzgqRsvR+EvtheF58UBQEVG3Sp2GfQWnVX8Lj83p+S0fseyQsVs94AhgHaMF433dr
gIUL94toU6UMiV4GhZoH/kN/m/gVwMBSCPnke3xOW4GBtVgBMWzVkXE+v6YtzdKkMJtzksx3p7Db
UF7w9eHPm0lxwGPN3Wb7zc7/Kk1p07Zbh2X+78BHK76jEVryRGW9JkN/NHNfUvTisRmw5qAkd2bA
H42ii7ICkE2OpsfV1HWneiBBqYDB2wXCJxRvOyJ3OizxkV/SIpChbDCiWkTiN3HBr3e+6KsEhh2A
bkVc8/+nMnrALFeIiIdsIsKmd5XTOK63DrzgcVTJBcZduXW8m30JVrMn3bgycSgLRgAlw0B/dqY/
1Hrhatgl6pgQT8r3d8hhxv+9m0ppks1sJMl/PiyxcbR3ATOY/Mx9L2TbcNyZ73sJa25h9x7sSydi
VzU3iUr8iIIG4TCRD4j0CWVQyrgjhbEoVI/MJASXR9wxgv7PIWXLDPXUjXX30T9gWKZfVnpGKMkY
wN+l4A1YPQndyrEm0M2cfcXg8QWimlM3aS5sGUmW/tuDF45G6i5nnT98rdSYhUSn+j71FgHCoyDC
d10u1koZF443N/ZzxX6cCJ08Xasy5arthwKRDEN0ZogD2I0IholZ0A+kEf8jL99mNNn0BwEReAii
WeP/MDWXWWX3QztWOLLz0oX7k4Q/fxagERBH4Mw1PN/E2gk0OdLqFcyQV3MAP2c5Sx0Y1lR96wbO
KgUmqq9VjP3yTnRIN36ksbdZJsftbiX8QZbE67FX7bMlHwOREYmxSe03GlJl8rIE/YaK0HPQ89yD
NbOpgDz+R4j7H/3Ri0Rm9PBv+iAWNHA/flnRQOUFdZZCtlAsOPejO+JM4MSBcxI6w3YWkwahKDL8
OX7cubZns9+evOuw/Xlrhul3RzkE7NRaVwaSUzvCgZhACWmzf4nqQ8XM4ST6fZij/t4kFoQdH2oJ
Wi83KMEEniTk+vXt6XggilxCJDCU00bei5r3CrHhuwIQy7EVnaAeREVQVuJFzgyw8e52exzWkrdG
ka/CaHnRb6fMSilOOVytuNXcQg+MYjpzITxRtQkl1XLXpT/0CfvdWcU/apy/R7PbkSdRPLyiMCQT
/v4LSp81Nvg1nuF3Pzfs7Jq5fFi7oiW9Oq9LcTiELcj3cfMfuTuYuUz3ajxm01LmZr+PVSdJibbY
fdgpz0b97pqt2JQvwVpCLhhrbe/0zI+Ey5e3VU8kW2NNlNxzDfGnconu5WfsUAns8vUzwOlEQV3T
6fBEmwciI4/QaVABB5YKEl/X+d3ziS7FnC68i45frT6HzXFPWTdKVK2Y8XvY9ZCGysdOzVd92b+j
kjy8v++TEHq7P1ccWwbr9TbIZseIETtJdUJl25tlXJxzB8Vzd9SFgkB57wPMaA5qethjTIzoo3aM
t8wt3RxvqtJiLlxV7hNFaM61FGc5iEYv2FToiFjNPF3pXACr8GNGb7atMuIvfXc3bQ5GZE6DfP8/
dPha6oS5s9d6GSH8+KFbUfcKeQxJqLODg7ZWe+oNVG4yv0mbhN1QLV1fBrWJQuOJCo4yTg6tr8wC
v/mVj5cbkv9e7upQtgM8yvXjkDgauW2O+dJMJaTGwq+KrJPXo4SAaDK7sYWscbksMq/DesDAQtKZ
4W+FmF7i8IvrWZ9GNWNbb07mFVnkHnHGMxDAXFkCOwGln5h/2/YFrSrv6k2cRU9IKDX7V5+FgVkp
aTg+djXFBrtnQlf0I4TZsMSArb4+yYbmdUJKTEJ8L5mVCkUtmUCvj1lFMKxpPQh5ya7N7XHKxlu6
EwbwJvoZTMfXayC+6wn914rqAqxnK0o5IbGXXYenKwEYtBua44vfTVWEvYf1oBmhSU6L1SHL6s0A
iIRmBWVvsM35VofiWebBleTfZkkk3ESaAe/9v+zBO+uUO2yEOeh+mp7hjFzpnZrs+Ljxj1d8stdD
2xmhmEJcEaMLA/MqvV4TGIAjKWXHemCQSOSahumPrLfoBu66n/LqJfM/kMrrEqyM11XX9+EVwtxn
//WttXzG5+CUKH4QQmCzQCkV74GJag9cSzSxmRpfv6G4GfOm+GsDYS6/EeKwDeu64fWtBuBkazty
G77TTR2l/dKhZI+UARQJeXpIfE5uzHcVGFw8tDZcVVV/5fVQCPVbydY14xSpIipRz1t6sIh102b5
mMQG23EzVdUIaGuma+iGry+uj8KHRDNXeMdoX9XtaKZ6XBCOoCMJE/XvDPL1g6xoxWSHrln66RWy
hJk8wqD/E/nS/5JFuG8cxGyjyWHXGzR+QW0cjf5MyGmB56N3ElwdKboU7QsFDEBchlkcwOLBBLBf
/ZUv7SGvXMfxyaaRTdrO1jHroqex048q/Rmv6by1e8bJVS7c4ji+/1SLOmQuTUZeMrIdQhmeJTep
6T3FOHqWu4adsPtk5V/4d7vH8uIMr41ldyc4oG5QDYjnZa0Z6+SxzqVg9ukUG3XxwGmC8ASI/0vG
3a4+9w+2LAK3JGGXHNyRcA6fGy0PtbKGQwqVQhNriQjSoVWF8VFyZdIGMtt+NDMrZK8X/h1MMhxb
qJpvWB4fS8UvF3ekplCNxaNXXmww2lOX6W979j4ZFScfU7PQ9g8krpWIkqoeeUvVB0vS3zbwGLkS
y80/+dCwHvd73ldC6BrCQ46ddBUv7d+dTKpoiMJOCmt2oDJfCXDSmYWxEEDmM9Wa/wCNoYtBRnod
X6qEDt/DIeBizujMqOjiwzmN/1sqfPl9h6qJSpX7JpDBCK8OkXxMXFM1itiFiL+piHUkU0sLih7N
iFjb2uPocKCR7kZ/nv1l/Xe48eBqpKpFnkWxxI/KxZ2T1fX/c5ypyP03AN+Ic1H/qeDW93EHkVE3
/R9eRLbJeIIQ/etZ6+dY8liFyUlIBz7nbUnR2kYsB2HRlwRaMBlBlBxk9GjbMNrunxBReZLewD/l
5Bqj15zm714xB8D1IeheENxiuhxSr2RkNRhn9IyQn7AgGJgHQzhXAwvn189jmS4PaR1cacErtZ22
Wv50bnzjbkyLypbxrURcv6HNbF1v23BGg8mseADwOLAg3OjH2PzarWZUSSSD5Tyx68Tm7/U0zhaM
tpWj3aktnHgDlms94Q+JfzvzU2lepIyIu0SYkdpPJaq9PXmAjjN5yefzjVVY8rvoLe6nIAoFBgZ7
BZK0rtK7lY4l6iSouxOLb8cgjfJ18RdcI7O+sHgu3K/eljIw6A2KuCAVGjQH/pY9emiXX3QFsJxp
XSKpofQnI2M758rXfI0oYtqwYJGcLhB0dMAv1beoK/pLwFZ8id7yNMRIWXdUGL96dGbEooSY1HcT
voMvpYLFLCMIQDx1GQea9W3qpW9pMVr93Wf7sKQ9cns5hni0mswUwG0LTQ6yprT9MMY9s9fsrOPk
zmlRpt4Mt4tn3bgB3DUgBltQ2xKwaT0Obf2Uc7CSacokBO1C44NviTddJ0mw+5Zj/RYCgFXGgxYG
ECHmAFbyNvOGhXD2NvX7D9KQyhgpWYNBZJ7Rq2M6VOoyVdoCyO9YSDWR531TCWeWSftRksbkS2EF
R0mzx2IcTlkA0ySnOmeklFhI75QpW+v7RDft+PKFHmU9a8fa0EKfJ/6ExN8F4Yx1OHnbBw1vYnAI
akFKRF5vnqoGpUbv0XyR3r3y+xgtVzrpCV2s/g2LpUqq9dEZlkT0Z/Ekl0m98fXXw6VuNIfCuf7p
dPRVH+x6E1ZCiVFckWeUtLJhiZsQRqp84iqbus1QoWXYJr/d2W1wyJCdTc6/xp60jacO78p4dlRv
yqhP9DSTSgYDNRps8Rkjzq/I81HZj7DJJWLp/5pnFDrVxCCwhB+CDHl5MFPBSs2Tv+QuQZSQRKIg
I+LyVRT3lg+WEP5pL26XW9fvGq3LnbZB8L2wKTosECKZSmKypdjmpNSLwe2qv+tAY+lpsMzH+Fyr
SN+sH9pquWZ0iB3P0Cxpzk99zDNfnhNLGMCk8Zso7QeaVv+RS6Rr1ue8oj0WGFjADlDGbV/z41Jn
h46/AF3sgA49b/D1rVHaR8Hw9wwe1HN6GOXjiK/2cft1pKe3AGDhn6j8KCmtC78la+spr0WsQoR9
m61f1Hhu7adIYyzfz2dZjMYVKw462STJcqQd6PTBwQuo5gAoz7qCyAT8/NEFEzpGxhi/Vn6UFB4r
5Epuf1ozDdEX2vBTpwCpqaPMETncCswvwTwUH0Z+u09tVR7qi1h43RfXsqnWC2VlBDd+Qhp8z73/
dQjUbPVlaWJv14pX6xEOS80q6uzy8sBdxSDcLe6BBuaTSVtKtZc/3bjJpb8o5dX72ms72kTX9NwZ
dZGGAvk+NUxZ43wc0SMKuFItmoQN7qzXAXA66wlpJKQtwAGo6qRp1K4QgqnH7o0XqeuWSYZI9VI0
WWYqGS8Nom94W51ssNxCybhRC8FMfA3PpfEk8EUbeFYb695P7BOtHIt1GHYCIkUuV9CYi0HYrdhX
WqMIBVnVtfWNZRmh1FwMA9vD4Fo2vWyKcpq4W0z7KTVNIRCMjsqeMAkx7RqNvUoM8ePZjB7Amzsq
mfA74+xJqqKtTkE8lVpWjA2bVYhb0Glm4o2m5R/wsyFWN3rfHxE+IJgZ1akSIxEW26fgakBl+Cmb
6O2W1F8AmoTFcqVsYnrq9QHE2mBPGL91fEJizUKYyMbxGdnEEazrMPiu+hM2g9INzJ+qtGkDtKey
5Qgzv4MxNWhzzTFVSTtY6+bmbC0uNm2hXvQE3SDYdNAOe5z7kwy5z9ZozRc2VFozkBpIFUw3LmLk
uuWJq/EI7PiU/N19M0p1aZtv6w3PP/5B8gM3SWtKwq+VMnxvPKkS44ShhYeSZa4zsSAHZGLeAvD5
Nx7EcAU7TAI7gWDZlzZUTsytLjUkU+7MkKyS0u7i3RFsqnB6eEz7veGajlsqbBPz8PT7X7+CqMxF
ATggzp3j04UJYTbZgpUiSCUNHFgU/+k0Vf5GRz9Rr4sm1EMFt2OtZuWBs5sa0G4ldgSw1YcFL08W
L7wWcqE176EdNZ2qrcD1E0dwetYw1ZLy90hJrj8kq5yHU2w8+Lo5U3ODjvGLjO6zpnn9NEp2ZQCw
a2trd6Q39evuEuaYfe97FcnaRj4ZY2gRKddlzXvwBOX2S/8FPPP+VmoQugfOnjQLn7R0qWDZvR65
CYBRRvAm7Oyb4Ka943YbnHDF50DoX8P7i11qsO7KX0M5izBgi2U97IW+gQvIeAssKHypvUxDmGjk
UDjI2qASEwgXdBqvJk5SfPEZivKKbCa9Yq9aOQZeygtTPKPTCh3Cng4u9j/Ub4En4b2xcoqFF13V
4uL+XYgqc3P0qzf9XWexwFr4rq2+gqQgCiAL3VKGWI1lTtlFWWGCaOisbUweoN4RMwUaxgXXivtL
66w+XiMSDBVnyyf2ScavSO4A/27Tikc+sUfUKTfyDXdQJ5W/YAyDjZuYWf66FjAFNgwYaLqjepo0
ZFpPPQAhXfY1Im5TYe76YTe+UQPWnyuVkTmyiE8/5JJvI7VDCAJfyfzOZZPXp0+iWZaT96u0sx4T
M9tf64bIVH7/6o05wI9Z8oUo493ttTkOkL4Yy81TN8a9cdzWxWYIZOpN2bYNIB/ajFpjqWvUP+ot
T6EYXSgXxNFSOFX+r39nb5WkryTfeEfuEnJvX0H+0K77DtXlXn33RLWagGRchznvir8q3vF4w1fg
BcdMC6wOye0o3SNQ2YmQ0i1bOvq3O6x7TM6nuFkg9LyzB522L6LuOrbu8YmRAAnKw1+DQM1FedqZ
1SuNTvzpsbWs+IZXtNtioJzkBv4NCWSz5sX4NVFeZ2jntZidZfeuiMm2eBtMs77HgCAXMuneCCEB
Al91uJL6GS/A+sysw1JgQllG9bWn4pco32QZxB7XZBpA4Z1Bbz1FDkljtBwlzmZmoUoHAG+3wYzU
D1QzmZyxR9QM1RIHmLLh33UlYmgYk9idzwHayCZeuAam77iU4sn36Zw3XMvs95AD1CZ2goJAVsMx
zBufNoAnoHEqeJhse7usjZYbh3COubqOp84LasK8FpKKZbqO6rcBwRL6RjJW1mhx3DIBsuYEyr7L
U3JhQgo3dZFlcJIqgLaJhBj0YoalbpCJRLFICbxkwPCbsG1gbPKoGN8JtN7e33aRAaZ06EFKWIv6
HG8o30TWaxQ6eP33I9h5l6B4cvTFAYV9kOjIyOpc3qdaAlvwkqrQ78SGKghDn8S0BdASzyaQm8gk
cEbxgaBmeXDPMsqMYdbj70VHh5q3soIeHK4qQzFlrL2DG0AhVysV5IA/597+Y4GTMYuNCAwl73pE
/TI48odzMIV0nGrsvZJ+PJ1LPg6x5PWQnxA3poDW97ok+tQik/vxK+BJoJmOPwcbJWX6D/VvyBXC
pqmWd70AlTkgnm6vDqZZQ7DkwH6aqqBNzwrENIx4B9o5w3vGOxvjtBW2y0k4xqIDtUdT0z6hjP7o
zJ+RHM/HnI7gAgFRp1yVI6BRLclE2+KUeVYmXksStG1DzV+JzD1BoEBDp42Kx+8w/VQtsfiHy42j
zgXEgP2ENnueKMOxetq7nrIdi4TndhHVqvTtQquOoriog1XLayWzPaZd8jJZNJGzdawVU1Pdau3y
Bg43zlEGUk4YAN0e6V3lGO6qNb05AMPDALbrcy+rTtPXHceAV3A1Y+E65vcwua1h7LXzY+zFZFCT
6ZdB5UPZH+8OUE0P2ilBj+/gTgxYFqib280nJr1AQxAbPoV0COmh7qmf1Qn/a8ZoU3TgkUBQRqHW
pTypqdsGOUaNPFUDIKZKBG8GuKBUAj4v0us3BDw1H9xnJjtbb4MkLt2TaXIA5ijTQs66xCGolpDj
CNvRyZRQtpUo4mZpB0UYmb0c/G9VVsri2o/1hipS5FS6ygh6wqw8rVv7g/RKA54aNqf/2VoHgcXO
QR2x8VUG4T7pRYvMQHNibRecnyqneO2CHrOTFyFf+td3g1IRy4IbFdNR98OXC/QOxul87vzAViij
2BmTEY0WTIvwZjevC/vmX9NUxXHFqdZ00K4yaff5yQrA/HQu1s0c9u/SYWKXxGE3Y6BRLHW6Zgob
cI61E+80zbr59P+p8yAC5OHJrxrCd+PYkdpVIIOd85H7XXOGLGx/YU3Ved7gogrOE41wGPZ04n7w
9Mb9kiZR/fxSULM+tWraRYoAScA5FpYk/LZKaBsD6U5KeS3PxH4o7Tv6+97OfmHyPSVm3NXiyqWm
NvXTCn3QvZmDJbIiPiJ8/6ofaRPn+0gELPnptLINvYdBz4YBeCD9bE/SvRLTa0dxCz4sjWKr+cE/
eDHPOxGHYHlJiJmAknPsP3r+fo5Vx7x9okvj6pfn1pCC5UAjYqE8QVfyGX7Ld//iXSVqmQJnCfJR
yY7yIJJyoJXYEYx9zz07C6hbflK4CihcCWq+wKWjKuvZQG7YbkLKB1ha/h7CIsVPyBcrkRjj710r
e3s2v1XArJuDth6ZTK5c8hGarJd8WqSVjyRJAFEBxtsq0jqYOyYSVsfFVjJEZZf41gX4tNJBndW8
ndy5zqtsFHf5C5EJw6fYnignNMCu4oSmVU05DcoO5aHyhUbsIf7OsSx976ARdEebABTcNB+btPy1
t/rVUCXpBFcbbr4mpFTIw7avO7niucFj+rVd+wy7PNNU4BdMTBSaOc8U2xJGV1c8sywcMZ0k5Y0H
ky8So+TN19GrIl9nBmNwDPgfcSCYWu/BfKJ45klyKd9SB6JY6R57sAvVmYxfo9A9dwfuZvbwXSlq
PMFS+Sy/MeBa6XgXuQwheVVeBfCV8fweX84ZSO4qOyKOw1gy4enDVyj13ZZFjB/koA1oebj6iUqv
L/NC5t7vR+8L2YpYFWJCSJ2LRSy5YGXaJgtJT/UEvH95L7TILfew2A+yGCDYxJtomyoijgD51NQl
rmh2uq7EPJK877zj+/a+inzVQtS1AFxr7eyaoQhDRlazAwiFjg6/o0U0eFQWzTJhq1FmbrddDZzt
4zlfaz+edIoDJGYr9r21zkZNp+dCdZHj209hFxI0f5rxt1FhKe1nj6W/w0pZ/XwNyjqyYCXbzQ6U
osj6t9WOZPq/hDHLyqaTT3MFEoyFcizYlx2QCn9hpVFTMWOtlFFLpzrOe1AhbQdQz6LtTQ2+UYYK
64ckFXtrLH6njOAmoM+1KTFhCZ1AD/UPZE/nDF5W0hnL8uvHSuurpD3XCTLQDps4yGZ7S0KwaR4h
lmAdFSCrmGeAZ6Vf2MgQPifjTa0fdLgY0RyEbwGD27VvVIHobIvfAiIvFYLl0WYGZecSirpvXsTK
AEVWgKpLNwPOogClcRF4+47I7SjW5Kdl4gW/QOf/pPjH80Gih9YbEsDc1tnVTufwqJqUfGFQQh1j
FVKr6tq5Qu/y9QLTBAKLkSkn62sswWh8bn3Tcex3zts2pJ8wrR8bdy2cr7duQcQP3xWuHYpkCWVm
SSmyKOo1w1CXrGgIQaRn+lNzIZNkvPwDqUVhAkrZAFY7hZNSRV/erPIhU5MTaqkPNcMrshCsTXuy
VY06sIBByP8H2af0L24lX6xV34bW0j6ecP0X1dl72WwEg33wCloLiidV5xml2aE4BZ0XdFXtNkFv
Ws8XJYeZyQjfZC4Z2gw2Q0KbeTKA6y08ug+mSslswJefPAadH4Fkiw5xu1ROnsRuTNOEtnxiauoo
jY3FskAKdwcFO4VJgC1j0lJq3tJSXVov7h2jbk/G1qOvCROaUn7dQkh6dlPnN6xEzaHJ4n5n1gET
gbv5/zSVvzYBTpmPYpPes2BFv9czzBUmA4+eiBNhdvsCze8VeI46sIF5pwLeqoL2yWMuCFW25+SM
zqSCOsXM2Czhl9/LcR4Nwt+hrRLhOQd6jWXBdRSmmAdbpyVE8doeYyt/lpzH6Az3R1PCmYP0u8rD
tX8C8fuCZEy9fBDuL3bFJXSlTintRZFLaa4d7NajkXRZeKBKsAF5W4PzOIgYHgOfwpOdBxJ1TqVO
cavR87hWZBN/r2Wky9iqlqdWNhNjnhPnzM1eoVkb93jUWo38F+EPQZzj4kRiQatydToeotvWkoqI
0JewjL/dj0IfnJx4KhApDgS2DApwPu9bOm+77/1ToIVtmrG+XTzenBjK0VyTH57ziTNDZUCei1xI
7KAMFZwSv0w//jmVtY99N6RvRMG5NDmpFImdXJWa/EURJekjeLAVM3EUGZAZRXZLmR2/3gf+WVKN
IgXWA7OB4ot6K+LHae7ImlBELGsa7tAStsgAc5ld/8SHHgmg8BHyNWOc6vZIZ3QgsHA0+hW1v9Nr
ASN4WWMQaiP68nq67zgm3GBGm84mo/pxAHR5V4NIxp76hIQ93YT7XuhoAt1PY4dXQw+Nhf2iIJL2
c6jWs1q/ywPviIa9V4cx5t5NL6hYX1EkQSki5H5qmHcrtq7SjeDBe2O/FaUdrOHYKQbXsBYQHalL
oX1t9dblGaqR5VS10CaSshbu2ymwB7CCrLuTNGzE2a1MWfyHJdDpjyDZpsfKPpT6BEbRJBSUlkDT
7m6EYAruBrVXLyFdDCsKobPIUa+KjTOCiaN5hUdEzL0JG5eJG0CTJo+38q9M4O3VzZyOsVL7hNSI
cQQomNisd5YgjAe8B/PmBcAkfQVuwubTKLJFJIhqj/h340iMCcmNajwgVLar3PjVb2rhYWC/Efgd
hRqttDVH0S8aC29jIcbndQmBrnH4/62qqELXzLTfVqnOOWzoM3cbB8nCJI4KhhmW2ychLFF64Nad
CwzPIfCrPw2AMnZPopEJRTDz/D/5bUZen9P18CFVWw27aubimmuPC0sHRjl/3Q2OliblO0L4lQVK
P9oHQNq1DGd8OK66eC8bdiUhJiGL7d/GJssYc4oir1hyoadf1gsQ+Y+aL9dqWNRLWd0rPP000IEf
uDtRAj15PvDNLVAi6523IQdJ0vdCAOtuV3t9eDi1V5wiKsx4yyUcd6l78qHuOstg8uz85NJbRuoT
3GsPKB+wS1i4guFat5FmJGcmEIoJO3XdNWgE3HJfzpQw4SXzEpWrR/xBTMa1GMODFh8PliWM+sIw
u79/wTD3w+ANYCtb5ak1qltlITvnjlGxMrc+EEJTFkdgtpcSgXnefN/fyQyEAU3JHQCl2ffy/loq
XLfkJRVtRNGImcSllFHTfCEWF82sdnjXafFX4RS0LmzhkLNSmLw0A5LdLhlUekhYS5Xbu2pqYFio
zDX5nCq/TaGuSGa1/sfeZbOPDWwDWA5mektBuYPG7mPLSaozaXdRYnCcxDeX1KI0EIZ2j7n8iYYh
9TPnHbOUkUpRPrRAT66mDZGtw1pxj7swOvGI8N+YoZyBvtbT1gRYqePJWX5T4r1MzCLIH9xqgELu
oFG7h03lWYOBPg8lsKTQ010yR1hsm+dyBXKXvz01yC6IqvrbAeJmp8Q6p1hAkCrAW0QVdV2DrPMa
78H5lvwpWF1hM+dOt/1Vta2HUeVbTkhxxZowYryoyqpr/yycfR0cA0uMkXQYzUMiqJnY2fvQ4pNL
Owjg9vwxXWL+1295xeTLd/SnHz384ZyGAyESWqUxrqmqQjwi2DVBIoalLNnQMGTvVZ2UXhxa9vV+
TQkJtOZolodav7UdKMXDQPDvWX5LdDVn7nj95n6TXIQUg2+VdAMlgpcQj1rgMjVMyTbSj8zq6l52
RpagewW5ckeYydH9dMqqL+1HH9LHmqXV9jmTtod8DhMzwT6Kwml4ODhpsWrRjyOEmsZnhn1bh4Pa
aYQ5Ccv8mRr0f0poaCfpW/N9LjPYx9HpF6RLPAVFyWTfNLVHSuMGKALZ91dMIprFIusR6YipWV99
doXAuwixsitbs8OSQ+kjpf6OTvI6WXtBSPo8jMg02HWtS65LeD1GYbtZ1O+Iw1AmCtJWhAyW9b7h
HknnroM9BIJGxFzavF9oJtIAGUSPHzUmq/RwLcDJe6XX4gRYp9KlZTS1eq74v2pXXQys4HySRlGa
YE6l44pGK+he+79Lp1D5nX/RApdB0rQAhEMvAragCVdtYqVxEJUC01KT4UeSmk+YKhRiPlPUia1d
sHCfENNz6xe7GiZbYR5E/DhkwW0dtxKUlT77VHn06/8Y5PTJcP+cytJ/HnfgEGlMJHDdJ65IPR2z
7ZgpQLz1aFWRRb823bGn9vOfo3JMDxgC91VcRkZbaxcSYCSoZtkRuVatzGUrfAVvGW8H5oShSkNe
S6IDbE/W+kCPPLmwkxYVMyKmtc2vegv+e9xzRTikVhA3RuI6KueGe4ikyQUt7nbZCPgtTVKIamTV
bsnf6UA+cI/LUIe+42lb7NF2JwKyncy/S+LQ3ZVMioBKz8fOFiGaInIXW+K502/67hIH5fdf25O6
KjE3NHE11yd5jyHcrKoyeOIfk69sN2h5uEJY+6oJpqEfKhlHIhAUqWd+8f1losQs9tVHTm505gsU
YP807z6ngRPmjb5yJQ05PmuQ5htw4xNhmOJ9I7jdN52aWhQj0hUZOlSiZld0kaRRUZxItjnWbKPN
gPj2DWfOuo1xqBsEBFbpccu5WHNfvCNKR0kbZsYhfinUJJXT5vmDPePZNDjPRFdO7J5GdllSg1jq
wdYCdpGuxYax+9oL6gKkTDYBw0wKaiR7GNkTblwJpJwa0ZX6Si/VYd9i7YIC8RtQIszvCLySFRQl
BwYqIIdTXIGu+pcqk/McdjN96xDd6bjKsbyimBv7JDWV0J9i4fBOiPlnqda0d2OsppEhMqA67ZwE
E89HT+u0808PR21FoT6GuFzbxfIyijN5BIVV5fKjqtrO5nYX9NLsEq1PwIFw5OljdKrfRNbFAbBl
XWUhIh7MBFz3yAAycRW2nKfl3KIwKuJ8lBh+b9hVrQH/kYVFkJ499eA43J8MqC3IK3qCFvH6CGZC
DmLJ/zo7IXur1K2PLNGTKX7Tb/8pkHcD6+EEC/dX4EURRS4V0jf31vOqx5CkPe+GfAX05BtjeQo7
40ygqAxbtzER1cn66mmFiDh7g4F0LDs0l/6pWfYOXE/oM8w5fL2M0pXadfWglHuz34ZuDrPFD6DO
tqC3JxLeS+Fa2C8wMPiVIIel0DvMJ5eSMWStltaiIv8URHsNDqkeIc/vc3lLBRjGIKYN3YUMFMZE
V2a9u0aJ0mL8dC98HTFsMOJox/iwpGmiMt+bku64A0rpeURjWgVMh15ZgxyIA9bRjPiRUW29vSq7
nJLu6Cs4fLdJVRK8UeEXz0Pom07o/WpEgcvDb33S1HjtGwDzWvFOmZEhAbeIkL+AjgBNI1leAoNP
6uH472sdt40io9CpUayEiJ+tkWiqK88d4QZJGdmwaLwzznepvsY7t3eojz7rGIjgjchZcv2BLmG3
CSiwwAoPFHotXIv9jtgdmyB4NldPqFLKz/s0sTfFJ786Q2JxC/M4YBvIhimtZtFSqo/s3E0Cwab3
vccfSIZUNKc5ZNELMecrBgYH19dObUeaaGHpHQFgkZOu6ndTRCeRushoPLmmMTp62hSbO/Sf5CXF
f1jeV+1PgT/f4JsSq0VLzpA6B9UAswIXXV3dLAl0/q5DAoILwkaUJBBzTNmlg1G7s5ideOI0WhJU
l6IduXujg68fz1V7CBFQXBlMb/XQ9YTkbs5qACWx+z0Shim1c1/wspkfmV4iG30biJDOwpnhBjua
YSDksEoNdG8Zt9RP8UDQzWQdBvIkgA5UelwkNE/N0n0skj9I9qmON3zVBsU5aV+da7cmlpTydJKI
tKfqgNtsqywy/WzDbxKmYAgXtT8p0ln5UY/i/T/tHzcan6cDpFQjLuTUE1L8VzBk7YCNrLEp5HXp
5XZIwcLeKjJLgBCzDje/Ad4giN/X/HuwHLcxDoGN0mka71aPJDb2ocldOH6AWvF3o0WISwutims3
nwVnM2qjoGdZw71TpAe5RtHZq0ljAFWpJmDeyPvUK3TE31DcD1J3M7dA4UvHui0S2oOyGQkw9CAM
x6ZUg8EMubbsMZn/3dwDkhMAyjfmw4hsOGae6BSuQF454D+j90EX0d2Et8vvXJRTmkDOzi+TKegW
Gfrn8PZUFoyPIEdsxZlioKlxqIzUi67vIA91141eqFkEY0RMFNCMD/D/BJ/WMltBMrrD3lxFJyJe
3j7N5FdmHGuizFSdTQUslZFMkzOdWuKZkdGv3xaE55CRzZZl8aaS5vRB86zpIfk6Qz9sYUXO0WZE
pW0j9ir9UHTPvJXmBe7Fe0H66q7WyjiU/Va8jB+Uryv0BfkFzmK0TFW0+Am+3Pj2LQiCZ9ChHurQ
q9uUFozJzqtDQrTNGuEBneTVQ4fvC7WPu3IPw3zTOwcv8pKrGjLTYJhvswr4YzzMDLkDOs6FCfI2
mbr7C9Z60fuF4FwKgf/p6OPkK6FrRId52D6peu3spbG3jUJjfjfJ1Zp6/yJyeQOYCghQj4QginOK
RYRpyKqDkTDX3TydhXkaenYYNEIplm3DHdcXEv9GBGcSz6Sz5cJLuS6AUshDFk6N3oFTIHw/vd6n
OrK4j31S33SdpPRoJmonDOQJvRLaXp6uGqTRsKIMoIW4afDySwkeqL1yPMJYgCR8aRN8CBphkOaW
ALpLPUqifO/5tSI8u3XXC6whJNrM0myUTcwkVREv0gH67zh6Q5cF5FsVSinrlc7dSDBAM1li2kRo
48scy5Ugg7N43HrDTXtHUTVKe2kMABZ7xoSdgcMY12reqKGn2UfrD7V8B9GhPwHI6NfR/rc3HdL8
52uVX30RuH89gd0U0rI8Tj2PuneWzYQYumBdPp6SmZZlZRw4fyL4zey/V9PzcXAP6Tg/d7+umZc7
Id/gcfWeriLAQJMW/PpnKD6DiDVVwfx7DaooZ01+OCEyxu8rN4+FBUB6kRssEJD5srZPqrPjUzhM
eZuWliGdMQSAyde0jWqkcuoyZ6dOP8ubhbkcyB7IdgWgH1NDDbRG09dUSIvjQnVnVdETpBFSa0cc
GPL7BBsWGf/1trxFKXPnwfbqHk801sqffXUN0upurwK+d3PeliIEQQqC8xcseoCEWOcCgZvafKev
jADcM4kzrC1N7uDqf6nQ0zfmEHAAWYlWCJzKPaw6CYFz23610ml0ej7Mw4zwUgtOsOTEuy+O/nnc
DZ+S/OdvSFXLJ+uTjRJ8JthbWgNNG7QxmIn3OfKp6jG7yc2Agg9OhMpLtvUG6Ip5nPpicb6tvSy2
aGCACVGoo9eYL9jssxZiofL53SIENHj1MPp02U31Shj9duBqJR8rKu5bDljIgGiyZ5cdGcIA+s/o
sW8NbzqmI0cjNiBodkPoMlsbhKNW9Huk7FfGli04YqWZl8fsyU4zC8//vGegdpITx9c64WdZUqms
Fuo9x4/+eWWj3/Jro+qDbqCrKMO8RREiAEFzDa64Sav0E/JS+KlW8rDZ/AhL4IK8Y1BAugytzj1B
BQdVmEnbP9sQBVjEwbRpb464vcusfRwIUXwmCOa/0WT3e+gtXKea/4odz6+IuHY0wnW/rQbRsesH
wMDNCqG5xMEWi/NBDrx5xzN6/PGzz/9Y0BDVFSy2LEnoLfsynmZw666xHWqd8385TBM95seUfTGX
8XVx/w9VShBOGHpOvlfOkj2JhvuqIPrA8PM1pBRPNbulDIBJi6ZyjU5i/o7btVPoS5ZwIgVn/952
u8ZXTghV8Hml7naT8EIs4z55pGEZfVKgLg+PWRWLX8YZn2HVkwXTDjJ2ed1tF/FsGkEzUo4RUjem
OUplLXQb0b42QO+219RKdeIc/MEF7V6OVe8D1r/4q5CzAgpGYAgHLW56yVde8b0v4kpFARMjYL4a
k+pItvIO79rxB76InXbR7C8eyR2wK9JvWyIWRv0iRonxzkRCBx7SFW72Mj0LFMUGUGmn9HqM/Xit
7o2wylPq77cZ5F4NDr8yxandFRfIuLEIngAV+pTr1IchSaAugr987SJ4GwQrHwViemfUqsKrW+Nf
NS5Mh9eVJpP/rpddwMJKpiJp+d5WG6TH2xG2DgAS7MNN9Wqx1iZI+Db5QmYNcU2sCgQX75BnsTsz
fatIADOdH6z5m6adChbm+lNCTxWyLMw8kEQS4joDFz8mqAtWbyCu4hv+dwJ/Ta6WV6F1ybTfIiqH
Hpn112VzyT6gcVseMEfIA+y+UX+sfzNrfXoGNNYHfNZO4YFWmEP93iDbJUpAEr+nm2asYph+NTjQ
LHtu7jFN030JAO+KVu/UkoHlBlovwGRepJWCrm8Q8+kWzdRtdZRxDtzB1HtMcKMizR02dRk71rNx
X3125GGdMDj9ZkQiZU6b1Fjick6VufereI9RUEix0nYGP/75urpyWu21EkK32EBZfw2ZAkxEfL4F
T18ATZFguX0pHJrLtBX/b/Zud2Ee3MBlWoKl5Er+29gEMdvYCPmYe1j+hIvdY1IJNNxAdGueqODF
LeneyU4WcZee4m5YBRtATJ1NytXQGoLhbL6Cu16SL+n4dhyfVltDxgBEQsV+bweBxDUA1KYZMwyg
xv6K2jIGra9253B+A/jbL5p57IEMlxNqOuNZ82Hn4lKE60sfyK76ICMPc90Jbjn0J4t3uEHjKZJl
N+2ST7AoWh2AnOdh5oEEtHeq+A2Eq3BuKt6XkTtEmimTVL8vib+ET0Wu13BfNk7vFQ0GyJeHo9Ss
EEXhDDUu5hXVUnedJ7Q31BGJ7wXDndmd65h+A2BQpOlxtmZVcLuHbX9+ZFSERt2Vos0e8qN4vAuh
DPNkkoUABOlQW2PAy+nHkFXg8uMFApfgEtmRszQOchUvfywl6xfK0gbv+j5fqwuTLPFi6ijSj0I8
S9wIEqRVUjxegZEqhrsbfwJ9kwnwHefEYqo1Sip5Ih43VBtpA8wt5w5/Vuk74pPt7Y7QH1+8DdDW
09Dd6lBjYOaoKnmnvcYRRwMioGC5msB3m6DFmEcHHIk7o5482lo22CsIQr1Q+8n5qMPSG58JRPPm
s8TzG4pT5xMTgJG24x5q7IglUMbsJ2JxOpYsqL1iAKN+LRwSU1QLBv0Qjn4waBxAwE7Gxk16auoB
gh9YuhahleSvT1e/9YN5n0bW02ot5siLSTpi/JsIBeC9hmfT+dp43KCpa6HXwDrQnYrHcSznYG+e
UJesy9/sBz43fxs/6AAVhRRdhGj3lXIom068x3TpigE9lyHUDEGc6qIdJwjNtRLgZDmJqxnPt7wl
FE5mmcB8JaOInN/mX8DIqO5uGEritUhKLARuChbqHRYY6mQEjpN0/7bctLvPYFSdTNelBBtmxUka
xtJHNI6iUtrydzhfpfZT7z7Fmm8ibnTn1VlMo/MOh+q4Xd+zD7EtAFgNXLtoy77GV+kigaTKrZ+X
09HxrxUNxSyB9cJCuifD3RITNFemqpmHLJtNYoIh8QGAor6sfN+KrMfmwrbf1Fil1eOGmA0/+I7H
q0OrYqOmunOIHFvro9BnkQxr4HIzGUBI2RWQLOaUnpi8GbFDArH3RNMk5D2tibwrRJOap1Dcbvuz
/wyJs6QxUSpXzqPFt9q80QaE7K96O3L1EDrrQKZ3eIYxsuxUcuwJt0pf1GqkSyRBBCKP8sjo9NpV
I1R1mFHqHcmgzujVt+WqoMrqfiq31sxYqmZ/mXXCMIZMKkGt2O6eYKFxznRHSXo4ARDnf8Qck+rB
uAOXCLzzpoJ9cj6AQlEMYv3nbPxMocTGhhQlb6fDryxcrqcEWL+SOoJ8IuZ1gJN2AcTiJDUQmwDZ
qRZfkmo0IauDjoYBbzgtf6g1uyWqYQSRgbeujoo0/wDg6kDOiM0Atgbwd1AeONDZgAy5CzqmEfmD
Ntv8SoSk/xb3/S+Pzq2SV3ur2xEibVJ1giLsfGXGn1zaxHWCzyqDg2p87n7HDUjP8GgE0IINlNL+
mfnIK0pxNxzDdQcivdFP5gNgrP7nu2Qz2GMep/OyDsZwURb3t58qhaHWxV1tcCepn8U9Z4a6qxBf
OxtDpBTeOstdCcHvz0gVB3prrooQGQ9jKkf8up2DQjuLTH2WBRR7sz04ozYUQcvFdD8dJ/C1HcNd
cm/GgrjRF6dYfGN4XwBC2P8rZXt2NA/pTItCMY+bdRmko+joRW/i1/DmaODCruLWPjuCnFBlzeYK
BofH99Wxo3aVE90Pl9PqF/PyKq9wBLxaiE0mZRrGOWTCF/fz+4m3rLEOW8g8bMyfJFFahU+gpq1C
0xeRkke0zMUV3zDFppZIZxfk0bDN7TWK/vViwav2GTweAaM4APKwR8dE2lhHfX6FQS97kI6SE7RO
KexSmu37XuHdjuy0At3aHhrBjDd37GrNpcBjoVg8y8zcxie49g1J/t/j79gDK1vZGiMW6IREGZuY
BC3GN0++hRex81MuJtP2MYwakak4HC74P4UfjDiQ7fjtL1dyUrUfXpGdc7bdT3dABUP9cCZs7iMp
+2fOTpjwfmv/aWMW61aKQWY+3fxqAR0hpE8rHMdB0h8yF5kGxZx7ouc+iPjijxHDbbTOn1sffIxy
IRG0ejofiluRTMVc+CBM0FM/L88YtLq+Q+7ckks3BXAyLa5CObSLaOgjt5JFnEFKJLSsQRJyPKR/
v4eUL32XMDMs9iO6E5s3+k6g+nAuGAn9595c6/oFiGABgQkHUgXuoBmg3QrWy6idlOFqXWaN0kWh
TYI6d4YEmqnz+85gyOkNr57X/LDo8kC98znslV8wPsuBVYpaWHGZ/5Fg2xoyK8JJqiRYKWJ50vZ8
zCVBMpAFCQ/JyIHMxbggnlJ2OYvnG5I/ug3ygVK0Cxw7+pBX3xFRxn7ovumyFUiJ2/ylaEbJmqWU
xxC8niNiQZG7DOtDKEx/6ccCAAANssed6l8SAgNyZXYcnG9w6ttIFfzS4T+/mX9CMUgiwNS8yMD4
1l6rztlTx8/GpdKxPUX6LB7uKAPWfL1OUe/opwt+9jPW9VwDAmXM0mb6qZH14jk7jdGpuCO/U7yi
s4IrYQyXqqyrNYCeZkXfZR672ndZ1XnsWrLJpXm8gVdtg/FUQbRRjg788mBNrmZ/bHWNWInsZTlf
2knTao7770Yc8LlAp4ueAtkohOmKZkYu95+m1tyq35a2FTedg2R8nIidcL/4i9JledPMIjPZGdIn
w6K00i8mnmZyINShHalikvxsne10LRIZiEdNdxAiM9OWAxfMjnSUKHqioTYNk8fhHPP8fgIWYO29
Oxs97QUazCV7B2dDAjsSnlf+qLbZr6qWf55y2cGPBoXxr6SCbhghqOOv7JB3juVP9wCKPrZI06eB
p3bjrrgUMlqj+baztlb1AAF1DZ4eIJAADY0ARKznsQ3+HPiwAkSC49NHimqKwSlNxTtVWRkLJZnB
rmxoSO1O55Niy61AZht6XDv6CrE1kRCKwg4qRDMqkLv1VMK4igXXO0tttTkony5WGa8HvmeFABX4
XBrfxUpa/UOMgwWrGjIH6vX1qWtARlP/CcxRD6jpiX5mw1qGSrsSE2X+zBvx/SSUBIDla6Tlhg8r
4oxOcO+y6dOARh4+n1aYaHJ+3O3KrDxCfIRTCWwtCcVzvGV5fIfRksufn1bhD0WsUq2GsMR3mdKB
2MxB6BHkRf7VJd0/7mL1O4bd7tF0FnxLsxlzzTsgSVNtRQJGGkUxj41nODsi/T7PZ0M7Z2jXp61y
nq/VQwKjzWrZ1Alij3GqeldWJ7u5HH1VAm0TdERqvvD6+AOydU/VxL4K5Hcwb1l+HKB5V6S1/zlh
nVnecdeeifevu7Ozrr2NuUQbIF6JgdMnuL+sQvAD6bp4B9HR42YKebyIhqUZPTzxOaduPHKG0+dZ
LsOAyQwfKKw+lx4HopV2IcfnnbboFdpfA6VXpFcbdxpF/H1DEiAFHZyp8sWaev8SnXC9dr9ejCfq
UTxnlIz8XI3cq9QvH6wVlQ3p4jctbuu2xEixfLQqg523BPn0KUpr2J2emCXT6mlwcjeEAtYLkEDq
hWlOAz6dwxgMdeC7k4G/iUVWzmquhRgWqZbXRsQbcb72simXpy85pFg+AXhL74Ka0P2c2GFaO4ur
aS24624GVLW+sZfuHIekL3rgawwc6VX9OyomShIh+uKLh7Z9UcW7bG0O5XnOZ6EYjGjqfkMBs7gG
enICqVHOPy3mjz4adaGinu1u19R14LgtUODU4n/QfBRa8NdVV8iGTKtNU9c2v6rPKuPNhWNacMiK
H4KG0X7ljDK7L7td+f1qs3cI6B6r+aemdVYAcv0fFtphYkJRdQZTtKgf0LtrTogkPYR02orcvJo6
fphM5F9T65IrKhG8D1uosxq7d8xvgMFln4Rtlmdm3HOxollscrGbDC5J97KanpjnQLS/OFa1BPIt
glBGVR3Rk7vSZk2VT0bZaPQ8eMDBsFMtsAkDI7xVjk5Szb144lldLIf3Ub+3IreatRS6vLfxjUIO
7BHePB+hZXVP4RHfHgwJAB1pHrU5/AxmVV8946GoJC4SD+AJ5s2Rgo+Wmp3qZTdNehnVgMvSBzFo
ZScfzrX5aas6gzs9qyZeoMN79E+Fyga3xemfXVNmhrI+0QtpIF864D+DRvdmIdgWr9GpeUQlioGW
a/rEWEB0uv7zElX0OREfpwyu+asEX9TSultt6HrUma8vNGj2vcXUp31jv9wHm8lpP0nHensgYSMV
4hkfKuAymlUHn6eN8xRc9kTJodLsvXiilt1jX+IOjjqF5RankQfLFHA0U5mDNtbwIjumItAGtnF2
JsGQyOD4g3BDvMIhY63yfscwmRQ5/dhwizxZbC7sE3a+VCkxkXFehLjURH5hG0zo9EMp8REO615C
P4NgmvG7HqA2yGn9pWd4yrPSm66m77h+aEw/l5BFiqlqSeG3Mn6pXuN0T1/etSAZ3d6dzBhz1Xlp
V9iwxsEBZjp0Nv1SIyqbBwEscC4HR6HRMPD0OUrCYOevuhtp16xpHdkE1XH82x+abVYnQXhKIhIO
56cwL6FdLHhi74yWBHaaKYlKqr7ZMbJPELiSmQxL2m33i6Zr1kkqaDDqYn1ZTKyFD5H15kh5tE1K
ZxdVoEd1IZKsI/DPMcw3V8U3G2fkW1oVd1c5CBEyMmu2MPKgvMaD7c8INH0BM8xFaoZ+y43dRsKm
YR9IXO8NuavEX8fybvyHC4KAfBtqTHDTj4fvhqO1GsTyA1cZUDE3MzeQpXK8DkrOoPejNCeQWpv0
fFxgel4uYaYe0yPTCaFSBMtwIAzerhebgy8RY2cjtXd3IHclfd26WbnruQBK1bBybO9cfm5IxbZ4
PPo5ytjOWqxZIFA8QA/mxe/jz+eCzE7H+0urTnfCVMjzLT/thTXydPmDySddY5KFpthwQnvlj20X
t/s8IPvu78NwTMpLPCpyD6RszIvZj0H7ZnqlkBvR9fiE+w2ftAvMzjZp/JieU9bLCu0AY8kv1lqx
22/Ai7JgSIHUVfNUnC/Gj8G/p69yZzCTARizzNlKUmipZ91r9vpE1RUOhrpF3Gv6MNGdWsaiNKpp
VulVt2ITDXLXo2e953lN7973gKKLb5UHRx8BPHQ50j3wkpfKh8MlYTtdKOJotsab4Q39BRMpcpDb
2CYnHJufdrMasOlsZukfw+EfjCtqWzt6oG1X1LeOReresv6EPulz0iz1sYTEM8xPJ6/M/XTPU8Nr
8CIGPuWEpdhClFERmvYGmyHsstXHW5tRWg4rrdiEvFHywHSucVT+SSwzfylhr1mvmIWaRQ9lRN1j
5ofnCkWqDw9hbOA0PvmcNBSXmQdaa4J+25vD+kotrTBw8I3PUO6Tg2RDIYVdnK9n6tVWrj3OLL9N
H/gDA9IDczs+NqC3GZWcwLbnASWaufqeSix3RIReB3x9/DADmvEUmVFUu5dXhC0SRss2EdQjyQSk
R4V/PWBxxbC2ir3UB0uUfxlae051i/MUWorEJqj6Vxrj5iMtnBfBQXKC4CJEelvkE4elxkL+KMrQ
nmXHsZPtNjMeiFhqkKx65IMLYJYEdbprReKGBNac+10ycK7O1xVfj/ZR8UgSTWThxaV3kQA7vKgr
+EfOPhc36a+lawKU6cAKS8eDk/+Rqbt4fnBnVDuKTSR6fANmDuIbNHBKkbRdzCXw8bGlYZlkxRgf
LctyURtY7pIVFfWV8rWhNf2OEMdZNtjvZ6kdkfvAccyNJ4hyxz5gYbi0qzCEUbYGxVQ43GhDTCfI
wd/VPwotCGcdc20+jlR6619DYiNKlyW0YGNZrbae+MHWPAmDxoTgKFcZQGv9vENa1v8ehcVkE6rt
NygRIvltqSWOSzvvFfxH+rw2oWXBzd/nf0z4UmfM3+WlQsQjxZq2nIzAwuwpg5U3wVMLC44tfy55
rE3qIGc2HKUXkOpgXkoduKusI7gsOGkuc3l+voZR2Xrb+UEgZS4lwRmo0POLvRTbWk3RR6fuywwb
V727/yn01DCYxWlcuda0QrZjXwIwIYAhV+qQu1iPpn1cwcEfK7/Ojt2wiqxxenBcjUQrRE7V4Ohc
NJhUyghQ5MRGSsVjBQRCY80lVZV5wWl3i9w9ZS/kkMEb9y62CJU/XgI4i2Q18XeF737ndUjBiGu1
StjmALP6otVFptz1YsOMtkjc789q38i9PL1mx7Usm8rR+DwLorMMQ6tkbquUGsZNS9Mv5KLGbE/P
em/6+bL7Z6fqh42eH8PgezmFEWY15Y6gXoH9T9XxVDouj7XGIPWK2MMBkkeVhbAF1DMWPzvQW1M/
R9MfMJvo2rmXMxzsa1Vz2np3O2Jlx+giJ1eCHI47RoW6XEcvqJqULSmt99gBBVzKnbmEGhnpdHvW
orHKr+iveqTNdyG8eR4IN22Z2JKO2QAvphiPyAvboq6SALk12tApnTQ/xUvEy91SWId85lMf0jA4
7vtP5KDByAa4nyBupCXZB6aM6nRIzO66eIp8RN5IRCbmqqec+q4JeaKsTdzRB8brkVSwsJONotZ/
N8f2c7FkCzBmAPBSOprDS07Ed2UMGYvSaJz/BAYGX+zBSoFxs68vU7GDdX9f/sCd3vbVqZ4smFOu
BDHXWPrp2AoynnUb8xRJZ2txbB9KubDKBhz/pvt6RSS5Iib5QGpnAUPftVRGbx0zOGVWrgaptwam
ghMJmufesRz1eyYlTubQ9aMn63ZoWf6SUR+uCSZvC98k3KMNvJrl2/B2pjwuRRSSXOYcHttPd9P+
mEqbvTQlsiFiGMoOt4Hp3rM7o4vbh8kyi9DrrCDYtrFr1pp3JApDtfL/mxa6KT/odmW9jZCPwAy1
oVhLUEXJLo5uYroMgy4MPPAfvMqhpwPcAkdq/P33cCVPstKLIawfrdE3wgTbodyI/ZZq3aWgDm35
t7crowLwrjwaZCqIeA/c7pVgAB0m3wkG+heo/96cU6sQIe8cFY1ofaoB9/Y+HIKzJf0e5Ia6GfXy
qwqTHCtQTFDlfOFbI1XzNoyZWlm4x6A15+ElsZPrU0fFzEjLHsEzgMp5sIgKoEAJTDc9i8NMCnk2
WMClcW8Lp8bjfzaCbdFSCA73zFO8CE9r4zPDwO/EjuJ5YdEe2uiG6b7UNH4kW7Dfm184X76QlxY1
5GnPBUgV320rx66wmlp62W8LANQHidA2o3GTQ2c5hYvq6c/T7ZK1jCmpLPqSbB/alPAOvZQT6u+l
tT5KVTyIkWHtcqbGZ81PxpXmesyRkiBeUi7uGXhuobEh0RDqSDrQwT7R25htcnHKhhz/tgZ/TVa+
hxDGfYExPhTErl4wLHcP6nahYaXHDdy04WUXzl6DWtYaiYALYGn6OpC2RiKxk+cEH4fHj8c/hnEv
I4kT0Y9phh4vVd+wMDBM4hiIdOlzzLBtGC6CsmAdbeIoxjAprU+CLaoPdilKHUK9JNwcbBvgT2wW
x40oJ6B8jeCq5zywC+lVW+i6bKyNRil1jb7rXXXE9O4RKb2mohpyllMOoZ+KMeI+SzxhK4YJ4etw
pJNw8L9ey8/rhKSANSESfMPeam6bck+rGYjnE7xl1MprupScTcPEW2vr0mKp7X6mnBxlkhYdh4/U
KsGjC0V0AOArosWbGGjbAUhWaRsau9lV1me/gUL9EoY3wW36Ppnxkgyxk2VbrxQ6iWaL/6CdHnpT
jKzosWi86Chdk6dK9ZFIHoGNbS9mX4THl+54faUm8nLsF+FsclkY9GaHR9/UCm/+xHtbS9Ls0HGo
srWF9df4YExdhr8dY2M9y6jqgQYJgsUXtxS+7tCZ81P6oUcow41Cb67IGtFczRpQKKQpAR4mNe3M
USBqH6rMjg1/XulgdFBF4F11isuSlY1jdSv0T/5a7DrqRcDmqJStTJQBInh7hSJGeSvuQuGlzng7
qPJAfjY49c6vp7ykQ/7HimgUu/5sZT9uikuy+8rzWwv1OFa0a1HBg0rdW0fBZ6Np8eWliqLNPAbJ
9YmEm8RsdK8o47vEQILkgmhpryhqL/pMAvoAMkONHRIXcoyV/Th6v+zRb0YjR0w3YyGUm9Xk6/ic
hCDT8rZqpChv9fKZrWL5eFWiQVO2ldSCtxfbEPXMG7EjWqUwSvfIPOvSER4NubQ+K391Hu22RQvt
x3WGtU3f3jbOE4cwn9oSyg84Vk5Vb2Ei367oLfT8381UuUnJ3b8qSg1GAwst6WfblMZ/vbc6VpnN
+PqBToA+QraxZiI1ww9BucpCs458fQjGeYSENDe0SfKKf8nlpZsgS8bmZXH+ifXZvC5MRw72aS0V
54GnhYIkgElSWDltAewfUX+TWHRZXGjcxfCmnrlgBrzDhJZslY30q2YoncK/p8oRuFx0rOQ3FnOk
D0r5E9/SjKb2pO66v6p4RTn902dSr1eoS/lVfVjesR3UIXQfixTmEjPqre6PvAWye0t5VajVykSv
Jn0Tr/RovLSOOE0xkFZWG4xBmWh/9EJitmPgHm1YuCZEopfEbc03FmeC5PMexhC3HicViEwflOED
EcbrRevEVqbgH/ZvEhT2RpwBMwf3XhngT8rn7Qn9AE5L5cSpjbORDweZ9mjHm74hmNXu8o1xUT60
W5Dk9X5OxnkLeFzfrp3Lx1vuP65KoljcTteJqmtv+92mepQtnIJpyNaMerogNua6XmYjUBQ9J/th
BRPoVKR8MznUq3IcHa7zzHgCkYUFoQE0evKGWvMWgtLIv8G546SPxTCRN66/wM9B7hvpRea9PJ8N
zPQ3UTQK57mZUqYsgWK0nJunUi3XQ92HyxdZPz6YNtmUAtE5Jlxsh98J7BswY2e5wmv2eXvX4j3J
YGHBMKKljN2CtbvQeVoh13QYXTq+VzvYR7rHBMLBmQpCVJUKRAu+Qjzd+Opyp8Ed8M4HmSuypuYP
8L3YqJh+pwwtR+xI8YA3yugduBkeF1vgFBm4iGUpT4s5bkPLMMhudEp2tgrjoDJoCJpSCIKGb36X
leLVndRzSknB1vRt8zaIPyy56RMPNoCK8CRioMIdlJFWPIkOWW2sIhQTIW1xrPhFv+KaBHEAVY1V
XcvhWqCJvb7X5LzGCn1Mo63nspYjeSB84h6jvGedogMan54hz5xBP4wcWNBXuVvAkDFumHGL7I/h
mtaMyLPRNtB0URdVVqDbKiL0z8DauotQzVoZm0w7+kgaWrzZ7QC6BEi/wKtTHDlJiZDCg1ntU2ln
j4fYjpF9vXqQPAfd6GwLF/rDCBxTKwiFwCw0ilK97WrEgpBsu5oV6fhJPMHJHUIH9MFpXweOPBvN
/r/jDv5Off8zFl0F320r9cGxKbB37Ba8y0u1yBQ2I00RpmWofiXSljKL789seZTZ0i0HIA9DYNXk
/9H8YpK8uCUf+a0LOuix/EWNcfeIZibW5MVPwksNFp7cqXFqI1uWdZNcfvmFiKBE70i6hmE+PD2h
6jgQS4PhQnnFwngjb5HPI9dlNEnrdvAIW1549QaWsi3rCSX8e87waVMlm0vmtQ1TkXC+fyZqUXW7
ALAM6d/D/JJ/ckS/duDjs0vf0xTT4jkdHOMc6cHIivf8teUVwBI4z8A7mczxc4XqResnl/qzFukh
pp5evIvI8w9DUu0AdG3p7OCt0vfH1W+6bhZNQi6GZ54aYH7D/6HYD472LNywZwsQqgfCWPHsiHIq
26JCOQDkuYJKRvTN83vdLTdWB4TuwK3fhnCylH5AatA6Unb3M09DHa+GexwlaCv7NYxHCSlxa+xX
e4ROGwkVhcbrp4+74Zmn5Qk+0chXbvy4pTjge/zwYMQX+E9cS/fqpgUqBIVAfhvu8OWZtP4x8HAS
Tl8sLbW9xPuJ/WsekJ9XgXos7fweOEKFPjq3Se7dOFcEG8tMie4XbMPyPGMXSp+5kQp/DanatrMZ
N3csTvYBk0N/MsWOa4Wo98Fjko/XnhmJyxSlRfmpmqAqP2j2YCwBRf1UHPyOzyK/JKwyhI/vWQE+
aruKPfu9rj5zTDvF+lRDEWi85PTuGvWyFoZ2xdvfi69c3Se496NZIea5pyvfc4/2eiHjd+3W7g3I
ZzEkrPCHvVxkDYCo59wheLA1xTgyfKTjB9nrc/D/jAbxbyN641NxDH4qNCiPSKEDR3a7EmvcU4LG
Y3Dj13juvXyeHoVOta6xo8VqkR7k07hm0bp7cvPHSHYcGggdmUZJh8Ig1REtNbtOx4ScnwsRFPHj
z7x51ChiFL4tJIupcU7LTVZt6EKmKngvgA4TQOdKZk2ioizHjj0593YQWCSgJXdYtkU2XpRHK6CP
G9P7bf6MsAMEitVeO3OZv+/NqieWFdCQWng0PZYW6JFZ/OeHsu3TBWXIFeSsprjkfVioFrRYdSgP
P68/HQjbsLdOp+OaCNq68vbCJF4T2h6/8lJhmPbgpJmnFqpOVaW+9OFY77XGDJHEZFsFS5Ue9llS
98Ib9JWCevY3UBWpPerZaxccNZZEqPwCxKJeYC8lM4+bPmX/EMlyR5raItOvxSg8EbxjE2PxB7Jk
Zt5PNGuLYuegPqp01rMyG/oUETOlG8TSisYENNhh/ScdXdN6NYfwvQbAWr5NI7kYhTJuLEXiosmn
Sni7iXVlgvYeOPQyTDl7s6AQv2ZbYOMastqjad8ZMu07ZkG+1m/GYJdypRR4RJi/tC9mRCJjalIE
ofFj1lPgApUIhpdujc4ocSCCDD8YHOTTLUWt5KWQx/OzytlCDJm2Du/JyCksQUVyu7WTAGrIpcy9
GXnkTrn7UHuTZLWLgCLUFg3/cAKjeqVhOcs/QqHKmHdXlOyp/GdoXsRkg5ylEKH0ZzPDSz/i2hbo
g7L1/6xuhshI9zeD46GQyFV/4K00fUtbjwqiBI63P34SCOcfw5H6LVCTjxrWuchn6EX2q//k0RaE
9QzSETRtn4NOYHvIRhrCWFs4AmGzPM4pZkQGZMlRUCf3JJ7jCoKrfhKhql9Z933uz2S3qVJp4uxj
iSZLYIE8iIGudoMwvhgKwPmhJYOuoXk13r7dHI/0BvX7pHh3vfebdDMz+gXVUnecEbTjM3vvkgJ0
b5myCFt6769xusF251res5qmBzpKcqTHlMk+RBcdRrmXBzGMYNZd3lwqfLG0EOOj3HodfkTGeErF
QfQ5ycLqAJnQ96kmhcy+A97JUQSxg6tlwyiMWtiX9ZXAnopN2B8sL80VMuKLblYkjgp6Xa0Wz3fT
5PDQLLJP00ae8byQ1pnfsW6wMqvNe7/SzbfE4im51lrhU9wHbNaoBuPFJxW4wuR4WHP0PdshVBxO
9GNjPfFTkyEDxIkoWiMHkRRN4K1QA9RZMUtk6TR/feYrCmpNRuhylfobXyKSVhxpsJ10/VjXhzF7
HRbonPXY9Y86MFuF3x98BdGdq5ITIfBrTS7RoMB3Ce8d3tuZM8P0Om2wkvs37U1+SkpIDyWUmONF
2FwXSJePYT2+2hADmvSckRvj1z2HCsSpjD1T1VjdLb61TXFshKGoEtytn6vOm9RXSWmh0SXTycoc
Z2iT3m3Ied92NVHa2xLTBHRvc/K+yzxUKx7wINndThc6rtAe6ep7Z7kw/SGqNHty7onmrPNAJRXE
BY4xsbFGr7t5S41cuQW/se0ihXT0Q3L6Z1yjNOxidvOxcZW3FRvofKKuH9r9Dy6yge4U9ptLIZnG
yNnL5KmdF04Dq6UxOyqmNEFzwhuPpn5n8ixXnxKNZnchYd5fB267iOp9WcbZNUdlpeJl52cwHIxl
569WuDBSLpSWdBdzJmMUaSu1+TW3aEJMoZeW5BQNXRAgZ6qqNOO8FEndUm2JbcdOGhnx8OBT56kR
4kg58mDW4J74HEF68vk+MBy8dhY/N2lbFcJmm5sM3mMGdVUFG5+5owoJL3RcmaJb25lyaj2fOnc7
sk+hdOnK7hN6csOGjcwfzCQw3HkBw5kVA8xUTBbzaHcVzAw7x+HcEujkBFWa27rAqPHTnp7ACLyU
qk7QJbEB9ZyzbyCcCRiE9UtuIEPSYPkFoeXyKQ8RDgAWTj5UoqP+gbDlHpngy9wgzbfra4kNv9UF
q4O1lqrhg77RADLbR3QtHDKHCK7SW+V6gu3Cv9JGHzlXa589GKtQ1sScFkg1WkABYSsbUNCTW9Ga
2370rIPXnxz5fEEFbC0d2dIpQPX/rNVS0i6OZsxIcJDXFoDlNT9J0gggL0cyIwC1yDMBzm6esJsE
TQzXM+8jj5+6Zjn+Dbl74BQtweglvCXqQ1X9rb+w7xSJ5B1pB7mXQEl0TNSnSkZZ9YIpIBYIlt8/
tHzsrInZWQRzROsEzoGokIyi9wry8nHyzTKwVDrcxgfS2oddySL5BCz827IDEMyTqgXodDO/PvlB
SPcBlvprQvvOyCeTAJD6CTTL+pdy/BqC5gXBZ9v1ufXYwW3mIJjZ7ozhm9H/lMudK/UleNPVuI8d
NUtYfqZtfNH/QGjas2324t3QOucog/HI4ukLWHz/MAh4h+C4EeJd71+Zopz9n8nmouuntRbYDiqF
qZh1T+HL4tl3gApFSYQttwTfx5Qj0Ocgst4hpb4NHsvakEZo5UDYN9Yqx2V0WnRWd18wc8EaC8z2
eeJv/2QzjWkLgopTBdprm1cju4zgj4MCooSEl1nYeMAUUaDnLy9DaSl/OfNbRVsGne9eKinHvEVx
GuunmbDk25LwTo/KxsAfMW75MDakfNYJHiw5M7/IgX8/HiBfI6jMzoLC+ug9K4lmZFhWT72u5KKv
I3djXgr+oA1QF2vaqFScp4cDeZUNoPV92hvjgaZwh0NCGUdkZwcsgDM1cnrMFFYizLjPtE0r/com
mkCbmRZ8SB+J7yXD2qfcDbxN8s7BWoQsjHsqlWkhBRsRgjah4UY7u2lcX99nV+ZlAzmcK4wE+qTF
kr0IFZoLiKdX2bt1cdXe08vRqvHzoIHzZsHguMur6kaLxKC7WeX1yuCp5PgJI9uMHYIM6s/A0DED
NQscyamSxzpdBgzkY12bXyOdhbieHkHPo+aMHiWiVKb+mqFLKRpzYndXzWISX33vcmvHx98pH6dd
/6JH7nB6Akr3raiQzTLwfPN1MZ4ZdBJm/6FPMf7l/SYhfFGDfZRwlxkRSu2uTcHEtL1af26pBiCl
MzASCuYCJBHm+SmTB0rMRpS+700+jy6VLCZwoHKPmm+gtiGgRuyZIDDkE9EnSWOgKaT53oi7fi5m
R8A8IUUG3mZJGNY/QYg5ecsz9tVNcCzQ2s96PZ5twmlQrJQYT2q5owUfdUZIMfuIqfoRq55TOQq1
t5oqMILfYdm/95wvOUJ3RUrYpGlMKfT2X9iAoULateJrbbRKxIAe3OJdfyp6jDimjcBq3ZB3KxpR
YnGmBuFdlbgzri0ESJ40fMs9J7xPLIx92XGx9J4gBRge8KD072BGikGxTUQwMblqIMJGxBdxHsGi
anQnE9rHmJ/bpwkvRUg2RyzrPNSkJ7woCDPs38T/rEi8h9dySPSwIcmgXOugILYxuTuRHL7N6Wcs
Y3NB5TxW5WQ4NRTqLmH+lAGmjH+mthcxnGythcqu34tVVbMV66xhoWAo5zfWYapvkyNYqraaHR3l
L3BiRuAjwYJ4Izr8jrvgZfgDtC776RDvHvK3PfXO2jFYkq9vV7xrnsCizqwaI/xCVmp48nY8Vvyr
zS/X1STDMGkLqOdGw/sO1rx9s5xj6/diMfhtAL6waECnyCAsK8KjK6Pn9fv3NIz13qFCRrS3WyEH
Gh5x2+DMtXidC5oXOFyyLtfjKQLBnGq6w7Gjf56CbUaMSfGshBonAxpQkLy00IGX1R+cqzPmGkcc
pNtrd3mZWLEcQABtpaoa0MnlKqU+NUH/3xvEklMVpPTc0J3+tYfH9bnt3+ikJZL1CXNiIAepBT1y
IHJH4YHD3r2TO0PKXve5LUa4nLufMC+Z1n7wydeKQesael3SMbhIYM7lG7m0yfruci/z39X8bTiO
HIzLydJk2Gx5lzwWUxCa3g2+jdLvtTOVWRUfOgP9f4RCII403zeXishNm95c6QxjamFkt8Fk6gA0
UvYirT0I8cykZ1weO+oznIIjKpn6lQ60BpFkZkVCeGLqyrZq+AePvkvjHjd/AxHTgG9CwPJwxUq+
7MjSxr8U/GMHfSfMge8a4GN0LNI7qgejOuybotReggNHSKq2Ntb6OTKzhQdqKM2pB5n7ZVXEUbXt
VD2YUAkM2YoHIV+UUsji5xtRMMTz38SU2eoZeYSSdgEpKYQelRj4IsaLX1F4HATu4XuRbr3muNzK
iy8T+cDZXP+BL3OEyS0sG6M0ywn1L7SqaF4W2BE6e5nUEhaLlrPalg+6YjzrouPVSJi/cT4ku9wa
h+HWyRj3xzkRI0e/fNZz7MZVaw82KRrKObf5OE21AoA0wnj1F3MdmVdFnt96DXeD1rsL/lstyQxu
x1keOC0bC3M3pYIgGzrMtEI0HKrCWQs+Q7cVCugLPeVAwx+0TIXz45U2rz/TEeNlJDXAglsaVr//
TTv9+MqUkXPHBpu1/jDzGDvLJT2wFLC3dKNdOzvAsXINaS0/pkAut7TlOYwFFhS/3DbVlOg1ecRs
QWvz4Lo0PCtE6YHRxbK4V1n4KOQLXO04YrHkOxP6ifsvM0ylQxYrA3WLigHp/T/RCr97nirw8Lum
CtuV5YDxh2UB8R1Lvl3pqTKb2nYhlRKn/9amynZgPmrVDEwDhhwkZhl3MXd7UD5r3S37TYuQ7LQ4
ugRkQwbLoMWzZ9dqot3wjmUhTR/Ea/V7vDs1UOGiw/sTYiECxF6P4+CwyYk7+Y9MZNYhdgOrsXDV
qfgJy2HhLAbP1zxX+f3n1TvIawaAxcGLpZt6lVmEBKHwHnc+SFObbg3iA4WQX3mmv1y1DMC/K2OS
zB4NFTUFL8D3oVE7Uk+4kEgUip/2HucgOH0Ctm+MzZlVkQAACrNrjKhy2qlVQqQruC4lRXP8hXTl
6cgvn+032bcHV+4luM4fvWRZlx33CkkUKj5ZFCF3XN3ZjM7mAIT+4iHssR0aueO+baQvuNiU5Csv
j5qTWM7ECi4F7YADZ0AUqrWtYiaLCnYvLN1K86n1BfWDuozdRBkXoPiM8BOtIKOEkdyo72YRcYtP
vI0GGTt9IwzLAh3AF+nFrmAc1EJeTwCddhQy5lC16cIWyjMmUgvjUK6hja8kMQrXXaHcgv21R6pW
Col8YLy5z5pRojW3360lXRb5Fc1N43eZva6lSDJl4hHmTP/VCOtVJmrmv+bM7jh2fZEnA8eggn5H
IcFER4zAYHQfOmaTdHPF94P3cUU/nxX+Ecr3FmSeflVsSbe43DisjN8Pk8/BhSfVc+GI5psG92cP
szbCAgYFQTtA4XMfqpxZT7VSZvrS9TRPsbmbBxwY0PIwoKPaIECMFJ51K2xN0IUc4r/sa+yvFdPh
gvsZgZhWZwmnNXN7xHiscAXbqxv6XJuRczm0fcOIqcZ5MK3MvwWAyzPre+fuSKSFpwwCZvKQTzQl
3XRNqjojwx9gTJH3xY2+bC+wAcovoxPXcoDas7QS53ohwMSHP40LiHAMthLqNgfRA00WKD44lHrO
mBuPAbtGSZNDE0BIIpQ+9S/RVH0rLIOzyEfpz5XOmU8CBT15a1ShW+Mlg+sXhK8dcsV9mBulsuze
KQlMdJraZUCGEW0CephhlyzX2gndn5HSzceU5Y684UWNz4AkcxsxTDugPjzsn76hjxR9O22MQx7t
mZkXPvLewqBuHCc6gHkFZ/ws/+hjrfadN2v3ViegnjAU0lcz3kWtBw0Ba4T2OZNh67tTtEVjM/Na
H0fcJgIZMJiBtFCYaXW7lzK8kT/fC6EQe8A/qRmVQ+73rPXGPiD6E0JQvyC3JFOWtCafR9gO2eZD
Sq4UuGBjG2fqrCRB5ViastI1BOz7x05kMFjBJ794SiwYg/tzfQJRADxiUsKtYSp7QK89J+xFf6XW
AiMdsEZKMmJoxM91mTLNc4BAZozfJjEkwthnCHTBXmy4fglhmzt/gRCkx8TQQ0OK2E308s+Q/Es6
GiBnY1SVB98FLuATHNM0UvyMSZ9qujhonWxymXy50tZTw1OOwze91w9AOh7P5wv5T5WC/EdjXbLL
fw3qEu06EyuAbAddKLUNxhsVpBf0hflYZCWBimsTC0RnQPKn9DkyLWLyF+S5SyStnigaKACPOusd
fW/lYeiEiXMhUxmGrh6ox0wwWUpnkcTW2cVm3zicE7qTP1sARobwJDbxFtK1Pr4+lLJCJZohOgvF
QkUtbTSRwriJyKtYq4wfvWxpnQ8/XorqP70BkdaVBGC4j2wT6fMeP7LrNClMvkaRUqWlgpVgJtQe
ARgztLziRhSA1TB5kG9RjYaG0A+I0DXujD85a/XlluvGC6XPekn4zqVNeGHrIE/YbOcHR3osgZFG
qOZ4mTe/tfX/lC4S/ekDlfoVr15CrEXhTmIbASJj2coiY1Gw+V5h7ZmybIZaquXb4Xm+wsEx8dEJ
afvbYKan2nVvI90b7UVpbPZJv4t2acDY9aX5UiiWSqSrA8CQPw2gezzJd1iv7Duh23N9ihLxWPhP
I1rsIp3PZTCfaGt8qkElYgoa+FttDYSc1btMYwvd4eaaTqqVrjDnF8ZoWVFJ7EXnWov1PAoD7Bjr
1f7EcXR3iWOPPjrpdDDrCho/BcGWGPM9gAHQanZ+HQaDyohLpOU1uqqajLUTiJ90gJ5A3SOxvvcz
Bp/4Q79Dw/4dc1Ay+0E5vgpTzungrePtPly0hsVCGC8efborBAF5mWfE244Ef0z82REG4mdTpHJL
vwWBD9QpboO7WA7yZOaneV436BWxeU1J/9kQJBzqxtdt6WNaAgty4IHe+4hzBixUQ57p1uCIUh/k
xZ+nuSR6a6nvAuP93sNU5FXeWkBx8Qt0uLMMctUBoEuxJv6X3wwEAlQQWIkcYUgHmr54N7jjWWdq
MAb++PLYvJ+1Ds/4dwbvAaIKxUsY8sl/m2Fz5TpKCJ7qqtYoVVUCnQrHUlKnjrtpjgjBi1mcxgp4
q2idqFX6PwQofvH1v4f+iNEV7Aj1wE8/6oR/BTeAmudVzwXY/2d0v3RZdH/ZtrTf/ecmsm8+6juK
YyvXWI79Gjk60eF4rOGwLX7S/YlTNTpcIhOjsvzhFN/bACmVlzq2ysaF61KSFRvKIPrNJUu70i//
BN5l52Rc6+UpPYhX+kEDijpq1IZcEgzbTc0cLYMocpbo1Q14ApYToHFs2C+2phLQWlGftZsNRQDl
sR3NoGFUI1vrQ6QvglG0XsUDRO7ijeM5ycN6VshfEsyJkeiQn02NRBNzfh09Qqb2ixqwlz1kNqEb
gfQ/eVAiX7B/gFCBX3//wjacAtbLF7F8xNkcPCRaVS9pejPxZtv3FVr4mDa6nPuwTf8BhuV2Zr93
/3hRsvZmDlKabpG9gpatzc9vXmAcJ4iDQiHphYOjc6NxuUfRWjFmXtoiFzp5Pf15ioInT6i2ocyv
7zfFTQs0S3HC2HDIhg5j+yVcvXxbiLLU5jcefhTwd3NdwmAvuo1o0vp0AyuAgXVOXl+ge+VMmwST
gPk7euYDbRQqlNOFg20bNTuJxL2Ha1UxLKB30dkiMdsjaC3oYcbtVYFJ2Gqg36Who0xkXYyPE4Li
62h0u+dMXl528UmWHL6EPORx1665tP+1rzOUKK0ahEf+uaQMUeKkwvi8Zd4SLWuXCBeQ51cuGf98
5bj2qOQYBGsqLJsthqKx9EufHKouIKQMYxznEeO7rGRmsx8QjigaInHrh2wSDIBt9PzoF/I1nSaT
yB1IgqhI+8EmFHK4Ex0ZATgHkolA0BdcsSKWbrqxbEh6MtbR0TMCwbDrYudDC9wW35IWlRf/hTEK
Rlm3rrM+xjxSNmLlWZVgdfqpaMT9/VJIgb96epztcs1GTDuFqBoeDATv7ewplTCpmIBWVYY5+poc
ZdnzSykgWTIFkpeThSzjE8VZ9TvP3aJlo3faSWHLXO/GyVu1nzmsnCPnlJbBPzc2Ul19YQBnpN1J
5umcmY0HYaCfHiGlV2NUyhcIGw8iu7jcxjbeQJngVSBKeAmOnwTfU1Kkvb0hIFjAe8E/IDhAlVhU
MS5pY7XrKS2r2nALoYw2SfW8kzKctqmOtlm5Y2sjwdFaXN2RtemXEPmGQOVkjTzkH6ONJLKcmzLg
mGZl1GhfipTfh1biig4+7wf4/ZY55CnTJHDpR0+I/bH0cfcMB3g5hAi9hsoMGWJ13M8y+nKtNNOh
rUZyI+0gjvKloc5B0ONeC87qN9rK5uw+0Ezf+3bGFMVKvl3H0PAeobotI8MKNXUrOkHKtzcFrcr5
xNSHaHUwAhYU5AP1QNgoHx4jRc17yFV4cKQTLAx77eQMjqX00ZtxJJVRkv2SY6mwgTAOYH2GToh+
pHZ4Xs1YyBSWVjG+/yGfNKpW0VZAvgbTdJZDcVtC5gmJcbz521tnRbSU2A39VTnSpL7WQxgqaTwG
yKX6+F6XK4J7qT635/mKdjjOqh4oRQ689RfhGQ2vgnZEQWeSXLOxzM5tOZRVcE4CRw12151fQpvu
dxYLG7Qj7XKhT30GH9Houogy34JzwU0wFjf8zVvFoMZJdt5zFxVPYmem/yD2PGYyQcLSRjsafkns
V0vIqOXT9VDJaaVT8fr85g3uOr+IJsjDjlw3LdPL2Fv7kZsEopIl9ESOoG3msGU9GLD5En3XvAu9
zGxJuAZb34fIW3SKOrsQh/B4KHIMNVBgP4CCyIpAaF22PAwfvX8/es2/54JrbqPpZCbmlddMXX7a
AYPa/khQpP9UOqMiKK4X2OYMB86aJ/3cmyzV6fTx2wERQu75hS5nc7nKEcdAr2XGv+PwSuYJMYZ0
ioSCQJSDHThjFjkAKHU6LrZChpC5WdNyG7EPfqQf8Wr+EYjyIVRPrEL9ocldb0anbk62FyLSqdhD
E2G6Rvt7iShzBkSIxdhHECcy+BA1L/olsPWwOMC+hdl8EISlMncu6taqZwy57FWecVND9NwhfrYi
p2IcQxFU3XYm5VLi5oQYUXJAUtLLGCg5gCvSro1BdZlc/33fCCrQ0r2paHnw8aYC+OXiuM6IAjcL
nuVFCUvN96zrNk7FZncAz1KwKkp+j2L1xeHVLyMaA6dRQ+kkffgqFNr7/nUCmslM0FBpBHLaMz3E
sua0EHupqcgYH4trYWGwmofNe/0F0F6bYUJcxtoU/y282RmpsLmY1+FT1cm3myAH+7/h+qtcFCh8
51UWe6TKJ+EBxcJKDrp46paTPOf26n1qBHhoXRLqXHCyHi5oXu0p6FjgRf1feYwuyyI+KFJS/QGN
BDZAfFeOHnnnCfhcL7El01PVhCD8n0uvv1ngpk9B0mksTD7RG27155HDEZOJUtCOdwBYNm5daegp
fhJco9AmC59t4mJYrFkIHk4fqdDJxdh3yQLnXzqAR2giYs884xxOkF10LgKw+DKLo9Be+11u7KY0
K1VtNPGGQW8mZzbXwghpThhpdhLqGXH4AWYWFCWQ+YlB8oyWfaIEIqtZdWNMfG2i5muSJmJHNsaG
Zh1StODefLifu4Cog3eSMSRsPmY+7hz4Nj7YnrYAKmmVTZgGPJgbPD7DGHvOCG7wO+VKBPlfsLHe
tSwct9uv9Udkwpm4xiqdCFbb/PUubZaSsXzFCsmIGa96ATJCQr1VGs6my/UuGswrXUMo3vOUPXbz
gAJ7DowObhWhya6KEG/e4RUtM3oxZDr80HedrVdG3DkR7kBhJV3REBVffLY8e+vZH3OxuHQJOSyu
vKYnBAOSKCfcKv71zq4jcWFdCmEjiWxjdj6Pi3eXTfvSV7KGxt4Xelu7YJ/H6hC1Ua8UAnGZVZMu
y0nasK66xkUwAu69zamRDuKrVoGPCzgctVSfFY3LmmMirJpP4DfwI4tXOEkS1/BRadcnuf1VddCK
GYlDIgHYUpvj+acu/LOScLddTT9B6cvq6lklkb88HBBhTe9KhvyQ5vYFKhdh1XjgUBrSfFwmk7iQ
BbhxiraG3wXmXu1AkJlrKVFX5MmgI2CT+kTeTGxnd7dtsdLDET9snaOLjM0MPPbjlPHLh34dgwjb
OeeggKhaTSJwjUb9q76CTzYgCwweyJk2Jaz7j0HyqXEMOFtL8gkwaM47mjGXcNL8cb+G6x+MVNrb
TYUYUwP8frlj9HKXq6WRF2Q9aRrUbO1Lu5IxkrOuDPgsJnpgX8EzrPDBaMfUaYSBlLv80qG6rjPh
e/vpu0plWTGBTI5krvoYRgefrY3h1YDGM6+oL1XAq0nnkHINLUyW6vYJBZ9b40Owvp94863eqMMR
mb2WxW9mFyZqli9ji0UfhSyIrmZfk4dinW8kSnaDIjZ6LRagVURH/I2IoScWVESLBY76oKuv4FKa
QfxlAX0oXdKqE4uvPyjocS1LnJPqKg+URlhvqPUMbVTIT8KeYz8NSOUnnUiH9DO47J8tmbANi70j
MKUMF4AIKcWkfKwAHj36oLjHUuyYTsJU0H4OzEarUJKoi5/rmjk0rMl/zlKbuPWearv1nErlypGp
zV73bT8tdMRCU3AEgVn/Mj6SGSCF8+6dZZtK5uoPmEv5ptQcnw6eUmCEAdJFgIpnMpAdeWKKkGv3
uVaYQVrbjqDCvNr2T92E3dmyrVpeUy0T8wWAyScXSJZKRmBlTRu3o9ItkM+ENEeloe3CPOyy1KD6
6XmfQ5Bc7ev5GcNLlKRbYBn9q4ewEDREE2NQM8adUFA0tPCGbvtjFZEZXg9zagGvkOackCgFyGdt
Ld4N3MOv8udfTNJNfwA6tadTO/FsP0sPV5Xw08vq6uf1NYW8oaetNtj6pqoSp6f8fJk4oc2CGTz6
R2C88ura1GcvyLKgtW716nWSCAoGeEcXnna3g4q7TBQmh38HxnsrWj3uxpQvjrxx4fvbbAINa848
+BmjgWtgD46dquIvtqBuAi4ZhbmrxfIBrfYLwl7f2Cpu+oyXppOGwWSfJQaAghP5iqmoStimWTlO
V3p0FptY9xNhrdq3hu4Gwsb0SCFaHYMszmZIHyGSrDM/Spd59gwRCp7wBNWHXY0qvDRlJ+4fqiQC
NgJODYCZaptGpyrYlVBWr+QVERfuuVO83MOc/F3XW+lbmFkfPJppvZ1Fi66B6cnDG+r/3TlkOKHh
ittRFCd361RhetDY9u/3SWJduKbrgLPujsuMapFqwhR1Fbdda+a/EJRz8jFDv2idPyhQU5IXWO7c
rZYYzYtdlLkkY7hi39JML33dPW/JsD0hdSjUbScCIlW/fjH37uzqONEaHuc3ow3B74XTTBgBHAiH
hONXUStYGp9UaKYNZJZHL39oy3ilhtz9YaRkG2cuWvq0CQzykUOf13WcFif9pDudlTSM2ukP66Mi
c5ybfXpwJ8Uapqi+7TwId3SDXIYK+gkIth3zzQizBwzbsOmv2im7QnQZhbvuL3twdl4iY1FClplV
+WhumFF4Dud58Xbn4XSMGMYVnIrSRB6zUzhzQo17hTG1VdQkOw+pZjcVEYl1/7LlIjY8qM6c8KiX
oauaxMPlfvbDLbc41EaJRRZsYUckn8ZS2TXiIzBfGgxX9uPDc2jDPxDp9OfRfPDnkgYGDZ9oqqqC
kza6f7aUzXMIFA5ruPHkVd4zePgZvjAx1tFeFPqGuMO7A8A92ng8JFmYOPELIqXOLRxy/MhyqqWl
LphMoETshcADU3WTf2V2rflpgC8U2GQx6B9KYVjUg2wnnaJEZrEwTv9m8l7YU0L7+yjDiuZ/diNT
8NCNsJ48DqunrDecmklJ09bxsEJdEK8Bcp4iSugCjkfnRh/h4PyXutueYqA4zu07yBmmzXx1TDdG
K+Q6OE94FDrhJ5i/nvxf/XsiDXiDyXolbLme6atR50rC5pPsWqNqITZu9ajCx+OJkhABixGdoFHj
XYJr47frtUqNUKd59jHPyKxncQ95kY2DfOjdts8WeUaGcHztVtaDL33VVWXU2LAYwv6lIMpWSExP
oFlkUwhR0KXEpPPLZ4kCq58D2YZpPDf8+/r+qxAuANXGK6UI78EeM1YI72g407DtkW9ytfr7yxUG
RoPOKSZY/qIPK2lNK/qJMSlPVQEzGiJHcxLqQOX+GwWmUcIx4Q9ledZBLnPwW7IPATIUJrc+MYUD
Bfa5Y+PMdHcdeO1atn6QMQdH5mDAscIA9XKgEbcxW/l0iRlTuxeN3/D0JtpZ534ftyzZo0rk+6t1
3AB5nLbbxqgT0rS0rN04KW1o8jPcUtlLC8Aaz97JzLeWgbV5ZeV/8yyfL7eRMUmtiDR0mXB4AHAQ
R+s+M9K3EtuVp4EBvwYpPGRSrh7SmHinGIkW0Z7rQpT3FcCMyzYkr+xd0TRLT9OGBeOlwXnqRjpj
X/yYj39qFHhKfcBvSP+YpqppTDLeqlx3VhMaZ+C1BKJQHXVmQdIALhdFaFXvfBQqBZWtd0ODFGuy
Oa+VuZ1peyx800sM89MwYrV5btlEJTg/fhoSeSHXSt2msU5xJ7rFpS8XeVXz7qMQWBY9v0003/YB
yoXgnLq250re5u/Mlg8P/kGyqm2g0gOieH0GlkS6vCA48L72xhfqgGYqoRSIesKOzanlkV9LLQcL
h199pjbAfoTgO73R78ktSOx+cFbvSQVGRVQq9I5OGPAG4e3wWq/RNs8krq1xQ/RZj9q3cGKxLruW
s5iNQM4mjdjfajYA+p9LvQC+E5IPxSHo9NiaLBrg3N08zjB73oep7xQwIZvwsu1Upwc2OMlNPrHm
B9KWLxdb2cpnzXyR49MuoiDpO70b4Fs3Y3yvbPNGoSGDQqpX0JU80ZEqYfopEkp3MOG9SosTeOe7
xOj7iHipY2Ad4GqhTSwg/gh4wll9fqhggc0GK0JB1iygBUJ0s/teKEdpZuAJg92H2u0JWKTM/yFo
SQq8edXBK27GmY3ITMypBP10jxEAvgC84al8FctSy63e1BNDlqx+p1Ghg9vPFJKUQrrhCbB10Q2c
xQj/h+UW38qySmd38UWdztliywUA3Ksdnxg1k58OsXeaK7rXUsIcNyXEYvjenTyzCVPM2yhwjiov
FOFnD/43KJdHE4alCurGzDatq1epXKx9+/+pkRZwj+6HhcoZHY8fMzW2RzNuHqt/eFkFWXa9Neia
zN0xmyt+l3AC5NI8AucGb/lf+Pq1Inp5X1Udq8tZjQk/vPeAzNHNcEkuqefVfmL2zJUm0mGLj3kB
ZvYtUkqiM5pDjh9ARn082Y+Wg2zcIY85T4+xZAB0bwQJ7aXjeqbL9/bkCDxMt1oa7r/NSaOKhECR
WMxvXJp0JAz+zb1uUoaB4Diz7LIL7GMIZ0njyv1P4l5pLZHAYmsnZg9c3cv8BtHu7EUEF/vDlb4z
hYWRZVioXLqLl377e6k6HF709eUGd31Sc+zELiM+x6suNMLbUQnz5/1kdJWbVRizKplf6NrGfbUq
9ygKd25VsxgpvyaikVbX/O5FqktZi1/3UcXX2j57vf3FztT7bZ9ss3LJf6P0+dQKVmoqEKGshC5a
tpinEy1lkOHd8FbfamHjC6dB3rcyJ+5DuiGEcgBfUdM+KeEB5luAQN+s/lbyjz7r54I2IKp3DbR7
YP6dMLYiZ/OeUJs9EaAXCDUVrmf2blyqgUnQd9u6kykZoiZfXoUE9MLZnP7rfwjKNRGzRR3Dy4jj
3MP1lxHx+jSCGblqRipZQ2fH+j+VOG4GE1ys+yxTqUf2tyH2gopS+J7PPvuMvkhWbltWBsiQIdcL
KyneS8nTCtYynxOC2BhbSBB/lOsm9r+jvRKPBsq3lKIjvwwNZst9FwLtx34xExWkT/tRiCRN+KpT
V55KzO4/SrfrqCJJIZwnSmiM7XmPfIrtsGPxu6nA9DxX9lhPKHIpKV9eLr7f7W7yM9DBwOfswnWE
9RI0HtrlsbKhc/G0Vcz1VofNPgQaFyHIKO+AjJfee5T1NIVldzZSNG5Y5ulo4rRt+0Tz+F2LnRZw
mVRy1VSPwfGk73A3MkkuoHokUwq+/CDtWKBaS00iQvKSKG96Cff1CMoXkXI1TANXQm778FVDsiA1
iu9SCJZ5gn19JJgyG7BS/PuOSkiVbN+Or9H0HpQyebfNRDaPzBqS1yrBWfD0ZfeB1b3hxrSgUy0P
dRZ6cHayx2zXY14Aiij7X7R3oqG8YXjU6ZA/MV6bJzeniK9wjugpFL0jWDP1WsFMvrGVFJM+snUI
+56UOPwKdvcIJColyo+n04rnftC9MbeqHyecfpRXyOU4uH7qLUurCfo407XG//40I+CsqzBtE7zi
jnvHVt3W5ZhBblN6TwedbtpmIrd52zpDqtpSbuUIneuh72IwIM035D2nLQbh1nKP14ykFXf3jno6
hjl+xIQA6ZWOUbAs/GJm6SBdASyc8nRnngWYujndpyRjuNwneAAGqWH9eRDewwVVUHwKEDkUcSUs
GjgKGpbDz5lT9WQ/RplTNg8lPEtDwyOAhIEOj9wKankVzj4WbTVgETWDEMyq1tSZZyXlN7YkAqxB
FqHKGCqyJOBHZVdeMkEyCYDfu4ZjGOSOflEMci+y55/1TjfAWsnZ5Io/gCFoVtw9/DY+kZAYegnr
jP7vOkC2xKMBGzxxb9uRzNUhn3vOEtR/pPLPwk9L8JbttFZRfIuZ1vqTDSuBfXgPrPJJnv3Dj6KT
FhAjBbKuXD5GP8SeZzd3DPOnsP86Gy8pUFoi0mPD0x20+KwXTiZqm2efdb+AswAQfj8M4Tw/TGnN
qY+uzGc9bGEFrTo9W/jNoZNXKzT1ApN//jb2nhcKMrg9Vn0UakzGWjwhUnSaMnoz+njQTMSXzFyi
Dvt5Wd6hwfWnmujrg5CkV6hMlbLZK/lrEPaXa6SrUwNwtfzXdby0svHHyX0vhsH4lMPQRGCKwoh1
ikzzFGO5j3BxD2WDRmybfrZU0KY71a3JAFQnemasLoUfvhHhQ7kPjWnxUj0jZsfDOpbvhF0KQHS7
Vwit0nYggyxkj99d8niZY4b/ZRD56dN6e0shCab5zDzLZgnXWoBkEZf4i2XOCyyNwZQEDIWWAI0g
aWLu4iQG2IjhlNG8rNxZFeSqdeVeVHcKkUf1ZFbNIW1GdwAIia3QSBK4SuclxqjMy48EWN90QsY2
1xUAYjGpKtY8rNpEoxvQrWjq2AccKEVx2xi1HuynXXZDDBEH67FLSLIOdnuqMhbyAgjQtxu6agJ8
s08sWJ3RabwKQk1DICKzREfutxrsW3prHXAttn8jVC3EL96k2DKi/GN6cIxk5VcUzuZDK2YcAy6u
E/t1mpdgTJTkH7G4aXRg4EP2Tv9VO0FjjQ/vJqxrbl4MtZUphhcTsTaNMfcXtA89Jx7Rw51xG4NK
LZMfpyn5TKATyeyLZNmazAXABRkF+9DaEz7qbVREcGpcTQZ0zz0clT5X9bs4G7XvFI1CcRFXPBY2
qW3gl0XpwzQJM1owZodbMhEu9UgbWScFgjChZ5BE7TEm+goZErub6naD67uPpZihlI8LqKtXF3WB
19nnomyNB5ouA0hFvVTw5oUevlNtM3v/RAyvUGM8/nPvPmbaV0NZ8Fy/UHTGPHgTQRsL7CS8+2k8
aD4YSJN7uyVV6jmnRNVVaa3Jbz4ikq/zKMmjeQ3JPFQmaRZWlZZJkcfYF6Km8Dwiya7NvlhDLXS+
XJUagQ5MUPuQCQzt8RZLYlLK7PO1AiCrh0Zm0HG+S6ZXCJkMDoYA5spXF4G5gy08jfSMfYt8KgQS
oZXvoiqgGMuuiqC/3xgquLEaLkI/mdoxXFLKLF0zpwlH74utE35u387w89M4rqUYGTHyVjd+dEH7
826aMGpclWfGQafZ0A7fDhkxR3nKbe5eoGmdXfYTdI40bnhR7caA9Y2IA4txg/ISsMPrbOZoB2gL
kk2sUGcKOVrSyvqBPpUvqdZHhEmfCm89Gt2Ps5ygvpyx1idqiwH+5PuvjdrNQySlmBcFNTcINGDY
4JN4rmhu08d5Z5dv6gy9nF254/0ge1a62klGoXmpG/TUoNYLg9dfelj8FZ1EOxVq3R2axump37MQ
OJz3iz9mK252lIF/Y6Hs965xxwJo7TTWjUjOuip6G4XXsmSj73iXg5HfOdekcSTptsjuuro3V/Un
5MuWDUxNGqn9BZeVsh6TDeA5I+W1VXO87A4CS8Rj0ZD4ZtnaV+WJ0EUnDcsStAtv1hgRgLAPva8G
/iFUQW7Ej2bRNqFtrIhuXhwF8MiEdPP3/747Q6D/o53Cpur9vkTDj0pPvrkqJnyGj8qNnI1oBwrC
GX/6MPdSUoMUOBMlg5RO8rqR1KZbFAiks7FkvxuuK0j6D7ZRbXzkjmLztStfPzGx388wXNJxJp35
A5HV46qSN90W0YZiWbSichhgu4n5FFbcjCEXvR2zCBFCm0A578ueg0jR4tOMjQGwxIn1gYBlF+Hf
u3opl/H3fASoEFdMjHWjxW0VoCqiAPc+4C2CRK4KzCv+LWhYsYCqwWWsXt3JgFj6bKQgRiJloEiG
XVFAliNx0sVFogL4snariOghtC6wQHT9Tm+zAjo7PqgcxJb3lk9z3pi/DJS28uvvnsoKA9TPpDpD
ktIfTRhuaC4/CEpuq7UhCJ9DumQQ0gdBW6R1Z+6zxrlq+T7bOEItInlD15J8G2D9bi8Hd8t+dgYw
XrCFGTviKEvIBJ5vvp7kRSjm+XFfMrTAU8uRkf+/I0LMScfRVsm7tuQEC2zMJje25imnazxSbIAQ
VuoozVSL7qigMLZi3F/1rtyLIrhmi/IXhTBKNrO5ZHOVyYfT8ZXygkpIn0UzWBVYM71QskAsxyBI
tT8d4AnXFBChNV4ny9nsecrC5LxnhXYllugBC8LfVGt3lwsfD3qyuAN831VvmyKspKH2SrtgG+vW
ooZD2Pi/KaEYQYdZ5CTLRruy+yvjd1Tz6nFYhKVgXtDmRoeVEg2ySeFMpodjiii9XpuGDGOgif3o
VsZmHNvNXyI1rRPCne2yRmGR73WsYEJflL1QTsD2mvQFmdGe0RmVz2d6f0+PYiUjBTU3ZKpeFrgs
Sf4T8ARB/+1pOrO883iRB2p/YVFxE5NWxiax8W/jEpQ+dWjiZCS3qclwmc0LllcxpJvZrtMWBh6/
VW+9TObC/dDMiilRU3B29fH+0TMQL0NKKa+DvpOp2LFzifsXVYatxf4K4vsunVMyk80GGSfJIiVV
7QS+ViElPev7PQjfLaDkp5FOUB3YIHRCc3LdRjSzjznalfCtcSm4P3OcjuebbNb4ACp5bBeih0BR
ivmRUMGWY/kiibTzdKcoNvy0lZSNT+jPaOg7jro2ifkAPxA7QyJ9yTsGCQfxtgDjBMa6EI6qmaN9
LFj8sPX14lrAyzQZkB8ZFWrqFNJPdtjnMnoqvKsQMZYgFmZDx8/UesZ0hRMUNtUxKj6iwMdH0Xyh
Gb9Od1AnpECNCvOEsuPe/ZucKEfK8gAnI+xiTFeFrLXuJzP6/4vYL1Q4jf4wgzXA6b/ry+1As8dA
LvR1sxfsZvIHJYk+Q9BSFP6hEvOZJQhhVzlWRAOSQA2WXRpyMQUQxTYBD7k0W2Ja58VXH7smUaPI
07oRkHyTgu+s9YJTZxtXvuHqvXdM0tBqzEwWw/FuvL6HzLcPLRQZETzRkWC5QUjs56Yr+8WCgeNg
LWxxEOyFcmSK/9Otq/P5CrZBX0PD66hxM7P5RvBavsOAkCfH+741j1DTrru9rrmVbIiGKKhHwCFe
JagrZvegH4j/BU5P1QP4Xbd0c1OLfjK2hVQP/xUdN6TJxDeCA/QtJLZQ87juyg7ADZzEyJLIv9M8
9xFWXfGOo7fLfj/hgV4vHIppImDp5SVHZw0+W7zDK4sHC0p0GaI1hamEO5dNn7SB0kew8roDpmFg
fi/9gguL0lXdlID+qM0A7Gar7w3GiOmjmq+/G9YPoAf4YIOAu9eQ5kiHU43ISEklJTke0YTtyehS
sXT+n7RH/MOhoRHUNZQIhSyF3JA4vuJL3j3OPf+Mw8GeZyxWrnbQolawPrxIiukoEfaytPBQe38A
YpgR+IZqyL3hyzgnzl+EbZ/n6vQVn9BiCeicEmRrFkMGOj5tBDP3/e5+JnjnpMiEJjId5NqPixkZ
sQtNCRBEEeRo447u13hasfowYQi9MnsKThcLM6g3nuVx7nj0QsqX1mh0weEmHh/Y76NudLfOy08F
V4pD9o0NHIOt3TBEsPSHUBb3xg3UhqiMnwSQltnAJr3Rhjv3+iIQOZitj0pobsSaSxJHR24fRYMh
lbuJd9VJeLcpUxpznytXdpCDkG+PThP0oMbuB9oZtQOUGk9KUKxMDiW/y3PTk8ioRInqOQZc4bH2
kbySLlZjZCWCvvE8fFjjf9IniXNCEG5VY3vDSMqpKEfjzYsKfuZt/RBLZcUC6S3ZaWTWXfSc6IJz
eMIVGWhE3S31JFqW0roGAwhoKdbRAkLSzhkDdadWyyJQH+r5/n7UpCpuBGwVEVS+5iM2lFghrIbz
/B63WxSSuMI/lrJ0w6o1lZmPxsyB+HUSvySr8F2OqXSvqwP+ohdlfXS3soKT95tZXJalc1bDGY1g
uDNzgDJ6OzFipJVds2MoKN9MbMsDYQsqfGo4rFZnHwZPChEF5JoO78bOSNe1aiFghBk1jPAcWQhW
8zIIoZOex6sLhbAw81LWThAH9nGa/I7r1RY8ya4+X6r92mLuSZYLwxsIR6U2/8kSZJzX0igaAxDq
iaP9A+K3o8jpyp6admQPZ5k64jNSkPc7ZHTKr61sz6Pjf0HKOtJumCxIGvEiTipYqkfyz0tGr6mm
zinpA5L+O4jp5gU5Lzu24wBpIHMcQdj/ggKeQTFvD4W8JOm0ZiGsMi4gIXbPQAZhXc73TZDzgzQF
wmj/4j4YijXjK81JHpF91QBJQSUjrZIIXiyBKWtE/TrkhfLe1XBJn4qbI4cGFCNG5ymTfVKQzNfn
KznDybwRQxPINx8Q8hmiDzfSLmIF6hyfkedTMBX+fCCo0e4fiHbQ2puH3rJ7eKjbLbUClWtTe+wL
g1Iie3OIIBtDK4ZmmDjD4OS3NZwYlIVP+J3r2XY8S6cSIbtMus1Pqp4pjvghPUbAq5wbfJLqUhph
65aRn9qmJPNX9KAtKbpbqnPhbTb3FWb0L2AcUmqsU5pb0H+xdSYRTqbLzJJRS0CgRlTnhjOtnabv
eLsXLR5mItpzUsipyWIHFs9jnhqovTCjkoMi1erL14ieBUby/Hy0K0KMPu7BGB08dxHQJOgjAWSo
4+YoQHAKzmW4fHM5OKroqNz2pjwR5FMhzAh0cZTvTsh6y94OK4Q0EvjuW+fwVTNd2ml4g8k/v3mX
F7ASp2oAEGfjrG1dceXJcebOb6pKXDkwanxXtrI7zFYCsc+cJJBzKkI/eS80oPDzrJO+cQnEh+AQ
9LX7JNdWyPZyvMK6OloUqEhuWW8jvGz9HwBoIuQ7ZE68EcmC4amFtuCAz3I1uxoJVzElzxQFFgUl
mIQ9KpXDB0gGeg2CKjeiDhxbn1ctqF5Y3e/bsDaYcgWS8uyLV+J9nFr2ulR4j4vTjMjN5w4XJMEp
1yI9Dy51N1t9YoFGVmti932MrtLnM93bLkgvcbhFlzn0+nYpKEbVGGEgJyej9eTXOVN/+7fQ+XAe
7M4R7/VtG/46xlQnwBYKFP8kXnbRizjM6cd6tsZgY8aZBTyPDCYUdthaEyA3hPnLkvQtOhTG7LwX
vluRO/wMZzf/4wnP0moWDhYBv6NNxhSEGNuxG1RAWB8z2W6wDZvkdYqEPSCuHHzCOCpAbZLMiI5b
091c/KTCwrl1+zdOgTxiSrb3KsApkXW9osLztocDBng/8yMMyDCCagjdUdEtntB7m9ROSNXsSNg7
qHbZyIZcqhDXKwFox0YJ2YgCXVyDoN7SAdLZLgKIgaYf326zOqZottoVEuzFbr68/eRpr8AnoG9i
Wxy4CQwJyH5c/hXYoyNC8xvu9zkIEv/TbBUTa/yppxyogmO6SpuRURwjijREnDfJj+a5E1Nxfs7D
6JGsAhfl17sd8ibbgn7wNNlXv0tB8ikSpud2ijTSW4pwA9AF4Wr5P3sASgwtQIyTpueTB7sXj1e/
Tyc9PQd3wxXKDBEoIsbo+Ddc5x+C1UzQ1wghu64lXK3PQsrQHYVWX+8/8vHSoACZOwVcqz+7UaEz
wD6dSVeoDZD8DKqukErIFvtsRhSaxLD4fGmSGIV/4peF3mIuQlkzbZD6BTt2PjTJbj85LZcgZ6jn
vDSiiQ+I3GPYAdPXhCaWf76AEJfAW0ve2Ui2YX1xKy7pG7H/nxNoQ7+XnBZMab/BRW082xGBlrFU
RzwKpgfbUV920tNe2FCzGp5tVBegRAmh7wb/mm5munX6cwZzS9dW66a8zAbMzHWibMpTpvY3NR2e
eZulMt2BOcMT6Mt3NDCZWbZ9c9vXq0jPJw0aWBNrbOuOGMRByi7YY5W1LyLzlSmH1kMfayIr8RPu
rCkzy7iOIMVenLxJYwT8ajq3kgO6WTHJydocEyqB8jNUBUvfngVh0woRELmq2mMPl+0b1vI/m6c2
TCLF3M5h98FoHoWF5bySCXdHFjB2hyR7k8a/pML68wkcScS9w8onj6zbIcxjRQmVKV54GCCnCFdQ
Ydz/gvpS7Wahh6rRfcp6sne+d2VfNHL6f2iFwh9AImX8IUOiW5Pmxk7TbiZWgBGzDMYkwLyPuIFa
Rsbp3W3gZ7ZQq+GAa+fX4GWzmPXC4UjSrSY09+BVtBsFYEzOrmmFcn8TXw80a1xiA6Qunf8LB+CD
PCu8LHEVThh1rNcsZs2Mtt4f4NV2t9um8bt+ia69/BgQFBk7kij9Ms454S86Gchrwd0oaoGiTXzS
lWcCKuBeXYnARzF1UKko5dX5w22UXWMg7OlZclnEK60VnBpUlAB1DgVcQDAwFxDg05GG99M+WWCl
W/JTVVnJXJcK25F+1YJRcEVuGLgLwGFJ1lg3XuRgbd4n8ozH0ObQs8N0BlEYTX8CsPCHOSKGIuri
CosmsTJdJ5j8GKznZu2DxwpvnFUS4PdAdE8lJTSb0bVpfLZWUgaFaC1oJVcwXcmfPFpQoHTGeOYQ
vRGqRCDuauB+fHliK0W8C8Qp/X1nOSnHM+LyzRadMKuc5cpE16HrJxg7on4O/M7CvJNBS9FkV0yT
O17C81En7UIsfIIjvHXIpDFP65KCvpBvngThEdl1d+web0GRpLkaTB0UZ67NiX+l6jIv+FiKMeO0
S+bArwgueKd57RuWR6LOwFaXQC/sY4hIj9GeE+9I7YSWTxw+vnHcqeG5c6k24vRr/w0DtOHIhcvo
VhTCd1jh1ovoUxCY5ePRg8RTdyqswsqo0rBuP4WIt6KopVAGcTlc2m+Qb4lixQTM+Bs/O0mUMDTG
75hf2apnMXZHp5ETFAisqY/w9+s+gnb2wNJvcpRH3S/1pi82cC+/U7MO/D6JVD5lkh8vvsm5Dn2u
T55xFbkpXvIUeG3KalleebSZqLyYGUVboyZ+ERNnsooNEL8iDg8OeE5qFK37TLcILlvgFTi5ELLR
76HMI8H+wQP/Llenyvk10WkM80rg+cctM1QZayZqeST2cKR/7uBTmZV0VGiGRclceGRl7AKd9S/K
FjXMGa+I2/s+bPIjKUh4dUL4ujs10vL6mlAqhcAm23EVnhFIVVDrPwypPTPf9wCq8E8ITTHydLGe
Y7JXyXJ/e1BDslLV3MDj/FI3a0pSEVZyr3q1VGd63sM3iCXdA8wkrf6vXoWx2fSxqCdQISoX2N/S
/LQv00Hjgp9KrpSvBVP8qqoZHj+F5kkzYvnNjCpQUwh/D+cWekUkJzOrBWkQ+AEG7yUIoMMxpdsG
EDEFzm4gFNcUWcsoX3anBRFHlpr5BczMrSrC9Hx7XQB2oI6zbjRHofTi0T+BVyQOLmAWB8VJf1YC
CAM1k3eicsvEMRzt10aFgm9qSasa/qfGFDkB0TNSGIzeyzNMqlmbDw30CSSQ6cWRCmIkIwJ4CHtv
l3hYwwS4XBmSxpiQ5n4kouodiH+Og9BMUaSFOxP/fuHuEk8cnXiKghWht/MEGdUh+24bpZHXU9ft
4yvwBgTJMc10rh+GnjyIvGw5X96Trk6Mb3kVoqpfotsD/hGRBxunT5F44L1AJWed92UqlLGXQeKn
qLGJqFIf68ZnIZsQyWi5sKKSoT0VxZzNv0jq3SLo4uWNMppX22vZ1adaEemsYs3vu5Wh/VhZeGM1
l1tMlq12plbH+/OsXLMssC3JShXPx43LuafhS0XHu7nglYRN3LSEEsLrtWBIvCL0Gdx0YF7P3QdL
H88Jn0Jte4S8PflIS7QT+JR09AvuR8dZP7fbIrnzaE0TSb+U1XdUy/QZbpV6cKQ2yt7jLZfXkTch
RSOpCep7RlnkakekhScsRytipWOE+slOoP6ISlVM+4Zz4tXPETpWwPebByWRG0hrmuvk+Zul5jI1
4zEc69JpCExL32Exo8SCuKAJTGDpUINhyo+tm+3pgrt3rYWiVmaU3Jzq5L13JG5rgcm7COM/7AD1
N6yVMg44LBcWAZ7K0yH3tIOrjO7D1e2Nh3ZrR1Gbh7I5Shk6F6UUHqIZGbtF+pbDumLoo5hlsYhj
ORCCbbUs/s+GfhOXPzC6BoAkNVlCs89pt3K0Yiecx+Nrqjl5OkrNffKz2txeXbxR8rKYCNrXGT50
hXsgf61ufimqPGffmcyZbruXCQr5vBibDToJQqtsgTKQTeZAygOlXq5YtViGgh3Qyy+TkS2XsVkd
r0l9nFRLqj9JG5S+7Ni9dkCFyRovZgTV8/zMEMP1NAuR/Lvvyj1MPPBRp5NtO+hUjXclfEeLJsFE
UKW4HvRfyAEF1GwPmiZz2YgnGejKjmIkWhD0Fq4r/CGDi5F1cSWPaJYK497EpMbwW/Xw51Z3fe1N
SUXMuJeymRTdumDE13yT/BiSfZ8XMP1u5ZD087mKa0cTqXJ3pRmGLJQ8FWeOxD1bvi7Ugff5OkbZ
jGOOkOr0X/uRCIK39Bq/axknFwwZXA65y936d/Ob1UZBAwlocd95w5POPvQafEE/mH6nvSDduE1Q
SlPWt4rZ6UZ4qI3tQeHh/Z2aWCm+uaMqR3nVYX5+TfKpoM3pkQl36BC5MZoMqsCRp4dY/kyfAcyP
ra2u7HuiDQx2nHIXfn6SKEA84Su5zrdnMl0KcQIu5guP1sDK3EBcdaVf7gycnRZ8thJ/IV3IB9ai
ikhExmUS0txLsDEDIpxRq/aFGCzxxnIyV0zrWgsPxl6LwsZiLGvV8UiDcdAKQFExCNSQ7O4uEkb7
G+NKd+xipM7OqQc1BQwvBKYZU9/KfRZKOpjIN/aWhPvipqsj9FDAdoEOKamPyWGHRtVkyuWRLVj+
o2V/zNux2jWkoUhoIl5TRltquxeZunvpTHAr5QNyPkrIw0oJZCpNyZGt9Hp8Zf+q2z56liskraXH
K2+yJzoaZXW9xj0eV6HXg5W7uczeb8grqQ4OGXNb4Nll21z42XpMmwZcrhaWcdWMGnXhoiS/I9U9
RElhiccD9Q9i6zAxf5R/52A3AVF8KIdGK8Og3e5WX9zGqAOPTA0+JY73TIv9aXp8OCBgjC00qLhz
/EkQzZrq5oMNODhp/B6yH2s005LSLevwBHyhxY2A98sKarJNNMx+rSF3cLNkYjD3f8b19y2cMpRc
4OXVmcK2B/ZzCOGQ0qhLK5Ua3KmhEkMcSkeb7nrBvPpKTtXWhfq9kpLtXH44ZICHAUtlc40DzaPA
QE7wcqXX3cX/EFOUvtEj7zPg74e1e2XuWF/aZdPLQ0KtfAkF7W/KmGMqMZ10baH0zXrkmP4D+oLp
XjjHjS5R0WANqaY2Yo3quQ1blntYjdNi3k6X5hWI4W5RBh9v//RknGfEZESILmTDwlME6Mh2Aw6W
+qtE5mSuqucMwmYRMo7BNSVQ9mRnp7h0YaRr6B0DDRq4dOxMsRA3vv7LzqVtfNgkd03Lpbec6let
YnZ4Sc29jpEHiiQyJmTX/1iZ9cYRvam+HjrhJ15OrzV5qzcyelFnd0BKF41Xg0ZPaIWM6K4ZJOEC
JRmyBd0nGTScAHfFiwEaO4VjYypknF5FlE/MiQ89mrTPJoh12Da6/IBRmTe1en2obx0Fii+oBoX8
JQzFnFWwwy2Wax2TrtBn0If5tIfnOAP/AR2p3BjDL5VPoAUic/UGLcyGEWDsnaYZXFiRyhLlTB0v
EpB0FhyDH5C6T7n2qKaJgS5a50y6MJKznTPBntXqz9wt9ruuIkHTT6WwypjhtQAsdiUwYLhb1ItZ
aWrJtuguDXnl1fLsTv6j/gktzmfSomhEzH9yKqs06zebOvdw5NlBdroZ8XlHUywmdcziOA8s16Wo
XbZgz33q8O13pGnnIllWERvZkP/3zD4A89JktplFxfoiqdTD9C+9J+m5RsRbCxlHAE2lBzdLShyQ
VRpV2ZG8eV/nqOMV5ORLXfNA28ua+koftZDjeTs1W66sXc5PkaVn5lvy61iYfVQ62u8VGVBi1kq/
EPoc9Iw+Ce69MZB91RvbFMIgdWNetoP7xcx6Ryht0beSeunU0hMuQVra2X1ZtGyIe0/NoLYGui6i
OGl1TgOdbK0EOqBje/PqlXTZaReo0ZCRXVDMx+L5lGVQqKTYPjREjKxccpndhlvRX7T4GvScCLex
V8gIsibFBb6OEbRBZrJvd9OIh31oP5Hy8dkIkk4+qrBgJXG76yPTU4cF/+Kq2v6M3x2qj/6Hq5bk
Qeq0GljI/H+iR8L0LP7B/UovM3ikvqA4Fu+edeAIngNhSd75Cw3C5Q02+igl/sTb2+RlVFqdpwRq
5NJBtUJgRIJNhCQCPYkpduRxV5uoBGmDr5J8AuTp0NKZQRYcChwN/QVow7tIPSNg+98XCwHpjPQY
DFGVXrJsyYNzBRsl39qmqzbnlQW3GwR1dAkyaCQKgFMbAzjPKrK86CVP2O8HoXmXxuYkxUd42Zi9
gyhGFQJ+5DoGFiW6tPvcp2kUKwkiR5ACEf3ykle2zMju9gTTDKHHsaGIJ9LIaxiEJnMbp1rT3I9X
cxwmLrIJKL9ncRsDnvZEqQ2ESc9tT5PIj5Ag6yALfkOfBrcVqWjSuJhTgFPEZzjFOJEUOUcam5xZ
E6ox6zkNXM4u0qOGmSUXem4UYakoDSdeGyT38O8yCWjKvaxRvdVbtuhdU4Of+70E4mHHEc4YYi8W
xYx7hqyZKu12vOmnBcaYsRNDHKKjXykeJihvHFZSqXEh/bfcAWPPRBiFjn1I3fIzIwLFn0zGCmC+
TL3QiK/Bi8p8gGxGn2ojThOV0uweVnt2adayuJkzHAlqqJLBpJTZRliboKmgwwC53tHiSsnXqs6p
08TByvq0EtqYllYdueKLW4igUH0Hv6WRDV46aRsGsSjh0WCRlRe/U+QkHX0ucXk6Voi5cHQty5J5
dCxl0Frnq0fEiPJgx+5YjcQ++liOwrT226LoskBcq6Mh/yZUus09eoxDkiqbvjHj5VkBoffMWlOl
YER2Hj8yiDeHNDe0ZYGioE4JFe+MJw6KelurRv0H60l9RQiTw1wDxKU6a6MjqKJ69YRiXRQYrJ3j
GeIMt+e8DUV5JzPLpbkpv4iXTKw6WRSn2wTUk8GtzizUH8+9Rboj9J/AV6iRDbZWOidxRVxVnLhw
AyGbF8q83WC5V59HA7p8r3c2Waz4PJbD9bQ/L7bGnyS/EOiUsbN270SIxLs5KpEAT/8oJIbfjiOR
9CnAlBnILoGq5G4Ms9RxbEtAejx7d4lkM8SmNA/3ocza6J67Gmj7X/VfIplJy3nVYNdcDeLalUjJ
ZYVTTAwyqzRx9swOxDxZ0xGrZWtSkDZg1+ngxbio8Gd0zvgU9iA5LsbT8pce53g4fYHhuV/R4dUS
htcN7J6zKZp/BM/rjPD0Xcbhqf9sTOuukj65Js+oBRmwV+tRk72XEsevDKbq2YaTntAfeZ1kAMEK
epdj+O6GJazB+m/X1hRPpq59boAYni3rM5ZR0MzMCsijeqNXuKS6/DH1DSSi0Sz2MTVAm/Sm6YkK
2j7kzGWtZkWJxhC/XwEoJx72Xy6enwEwrR6eBZacjCGhxYDOYcr8KlpLlo8WEEZjWp8pKWwUbFg/
RrexvUpbOtQFBZbPgoaYfDN0E062EdmKMtLNrImjHcFWWCHpBK/eqsp10GeRMHLdyEeEScOy1pu0
bKjxFB2UooA71mD9He+3toPTPLhFPYDvKW+R8EL8+a4H5O7NUDvEctTgfcjRlqRKv6YEBhyynNK6
lvT8BQqzpLVM+ImW8y6QRdRMoSV1UiTgz6YjxRfn4lBXnNcMirr3Bj1rmJrcfvPgAG2HYGmnRQPl
Fv2n9Y1A4uzpEZDceFmCYBh/8wYt+QKC5nDGDAy7iOq8Nyn60pjXV8NCp6bY+qyBvfyaVefzUey7
c6yI2WEgyf6yJ6bxK+YOi5uRGFquMPcP8Ah2b6MYBFPFmTqfjhh+1+zbTmIazuqbK+NGYLlgM2+E
DMuruxhPlEoPcc9eYsEYkfZXsUIcs32r3jnnOq9bAGDXBpitvmF5bz4iYh6NSmcJ8UJDN5wn5EKi
Hq0LhuVwrD14Wlb2Vil/2GXHq9G0KsN9opv5gIF4RCKFbTb83B4h5OzkL7hvkKUt26LDRJPnfhF3
I1+EmDu6/aYmOuOSu2MS1B/40Q2FMvy+D16fW6Fme7TzzgVQJihx778ihY7V2MioOqZDYlSfW8vz
2CH+PcZN9McaFqzpgMi2dWqFRdrm8GlguYLrL9G59y0eM0VhxqdOkKnkBEANxbW9T/NuFYnK/T7f
IJjdsb/BkIhabfFpiYFgm4n1y2K2iFLX1TgIH22a46ZVz2E+VpXtPhloEEW9dDRwpJvXl6G9dEhc
Nlet5EZZuCKYCqQl+Mm5hocmtmn2Vuez+Zw/8gctUo/6Tp+5UlW9DAaDPl82glyi1yqp42f01+JL
1d2XeW/Xx5Ka8SKqQPLkqq3sOIixDWgBOpj2FtKpI3I41Afkjyi6ObL6aqhZTPNpmqjL5H+pabym
irAMeMz7yGUqZMdt7F6YM5sD9LGk899ztwUl+cuGCqGo2zi4f34b/E8NJq6hTe2+SvXyz7eLMbm5
yl4kUM3Qrh/jgCLwIdsi9wZf+hQX0MOsDk1gThq4DvY1lV/h9dYEt6Ayg9T4I+EIIZnCCg2J8ZH9
vksocu65a1oLEe8AYoBfa6LIo9k+4Qo2MREMPIH6K8cuOXdxIIt0FSOqX50bY74OFCWZGX8H8cM/
T6bZrXdTmPC0ZOZCvClTIodR8eMlOlNmRHC+4lVIC+ypSPbuOFzOnOUikcD7q8RqCoITh+r83xqt
1Vwp+vCAuhAXJ06gKEFmTGI1EuCcIIBfqbl7eymccCVTcLfv2fGoE4SU935TFt2tF9OB3vpqpDE0
EgEAxOzcueLl+vb8X4Si/XJ76uM+BoPTOonjCSwVHsCatXIPxdGizoWEHSMi9I0QRMtMVdhJTa7z
MSyprS1vqBbRQ+lLlZ+3db1C2n3AtIhjl646cjXzoABxuJ0uiGqfZocnXTAKKnYKbFEOGKv6ue+q
Wglio6OEvhDs5ysazYpN/NRx4mS+oNq87H5excNplKdZzHf3YjXK9MAVNpBVneG4GweboJOLnq6i
Q6QW1lYN7oQkpEP+LiFOGAW0oBsKlFvGveK1Hs/1z3yfiLDRwecfQj7jDGtSBdV//3JG+QcHg1Sw
A5ptzR3bUUZ3Lgi1epE8dM4Vwaw/+hn8QnvxRhy1OLMaL614qshaIb4AW5r2QlJoYc4v0EfbnK7/
LxbTFE5TY3ngKe2g/nMdgOVwZUwdlgXdItj91xfLITDeJYZ6jYfTuDz1UHWgo1szjIHCcRTI8xyO
gtkCORHGTLYUzjRIQwuycSfuxVdZke6t7K9sANC57YMsJU04npjFGJBglcZCLYZ8hrxNTWJWOcVq
1n2jD+55JXFpI5FSRMaE0yabjeScJoZg20Grs1YEhrnqVx6f4vXmW44tSFRGTA6OOWwmiSFRLCF8
3WY3H8xW2oq/pu4qmKQX5D4hDM6GUN4z7NJ0/xuHnc+Yz6mewB0DRUyYC5Rzh89NEgSdal3+XOJp
jnCSUeHIu9jTuBRgSgoYgH5akuRNab7p6Ta/xcneZYIy+zvMQXdyhPx6Bm/xvPAUFCMWs9+ARezi
Ztn5dXW0wtPpSO7/dEpCVmDJXdk7FkxNjoA3zy3DNS9F1oxTwR1aucJw5k2OAQTA6vec1ZIX/Y+G
DGI5dNkwcnQ7Rn821zNqVct7XbBxZvsxsxymRXSYQfL+EofEnbTRj27WH5JMrpKbbeWaeM57wHDv
dPTy2hdbOKHPgorQQwbpEFmXq5VC2wOFhL6+d9GzUIdBj3gu3lpStMHTUpeY62uGuyN5MTyYd6bs
BXW6uJrotLskhMqK6AxGLgP+mQqJ5coe/vQtDuggd9mY9SNc7eL3UX6NIDaV21Qmbx7ZDPf6hZ6w
mbjFZeItW3VYb04mPye2rAy8IXganmOLH1X1ip3MRvUHcFLVQdS1eNlZdpgfHAGfB931S24oGtQT
x5ehR3lu/LzNJ00qt7ThClXgj2F0RPYuOMeu9XOfmOzbdqvB7v2YjgYXuHm5LmQ0KefwN/INoCFc
boyvJkBwidDxK2XLKJq9uxsajdF1+WYNGc8s7Htm+JBBhYKWGgEzwKML6awdJX0xQZLgj/As4ZgN
HxNYhEk7EPjQw9L9PP8opkBqnQSjRXFe67g/eLrxxcD8bE22iLN92rsbXFXuEq4d8u/jb6u61xv3
g4pWsk9zTdGYfYLHA0gPGC6sm+t95O/Hmt/NtvlVqkPycvJVzs93CRCxxrXrqV1QlmEvXXyCG6/I
h6f8cNYlc9IzTS6o8Uz7Hgu18yMYh7dS69AuWwW47RduL7jKxPN9f9DeTDH6AoyDKksne52RNHRG
ZBXY+Zm6tCwe7raMA/d/QfFvq8yRfP9fafSwKyf5y+fTZa6m4JXo/ApbQv1iamU4LpQO8Pdewa4P
g1+/Pmh6ZQLzLhjkLYvVwPVRJrz5Yiak09l+iDr3ghhkeiHQNrWlDLJMe1nIEGwKmx0vdANhwfbj
r3IZHaBmZYt97g/IpWLfSeaQmBby9xSpSoXOSYNjtcHSu2lYJEuptHASg8LRpO54wGdFA3vae86T
f0kG2jLQVRumTvMjoZ5SqgfX2Gbb2+QultSlCml/UwyIOSDviuFthtK26Z09wXtqN5U/lY5EdjYg
qZtWvqHUf+e2RLPPQAwS2D0vNzIq6tFweTenYrV6OY8XBfQVLamifqLb64rxQRjYZ3eBaC+Dupqa
yvdQlSuKoSToUgQVmkGtejsCBOhdyLseAawswYMwgqR28gq+1VnGdVZ3H0MpuWHd0CAm4DYpsL/9
d8LD4TLhtQGFDClEwWmYcbNmzrlz+r4IHCUiV3pc0BDv0Bt1qCIzqzFX0chkZ5FrbgnuMJ7KpHaX
VFkJQwfwDgsVkkImMkMivrzvShPWnlpoRP8BApeEfwfvL83VQiHrmsr7AVlzCSvChPyO8+Hd2R5I
mj+Z0lLe2wTwEGOc11hdRR/YlnOhzD3YLq5ZbX8AeeoFVAeqx1pXBHZbQ7J3gxv30GhgGr943fX6
DDdfBDSjbWuH2vs0sHVgBvXknoxKJLZ/LcLMn2ww/z7Pa5JASc/PhxuhZ/16Pc7WIFoA37ajiYyt
KCucq16m14PHokIYgT89oTZscLuUpcj7ftcCR/32z/DSn9N+05pb2j3By0bUdN/3QYmi/WkYpB8+
hVGI4EiwZSU3BZWo3n5kxhgJAEa2ar8pfEQRwgZiLQOJXsr8fLrptWNtJW5EDgH/Exyv2Da17P2m
NRHElgbjze6xNu+nJiz/K3sw79FEt+gGl9C/ElX19TjWlP4+2fNMvLtTZAh2skVc6JJHfF4ZW140
CspJAAYgAihzCADySB+SAqqbzyOYbEtuyPt/+/GBR9JpSRKlzYPkkU1eGdWVCpJaZGg9P/q4XJyM
CSDXXago6I1SNzYGeKunRheCS9FXWy7XbMVku6RU0sm5yjrOXOgiKqwdxLRWBL1lNMNYP+hdj3A5
2WmxtdwuCRZC7rtllRugzua/+4XjtPToMBjWLkHMT6EHvf5q97tDoe1jJsp10YIQkaALRkbm3D/b
4/K9koYE+xaLjCNuQD2q31lD3LDI0keIjWg19XZyPviY1/uvdLDGsSheAkauAeF2rdlyXOfAmmOW
bhzYzxrX+e6+SQIWadP32W7ryovc0FziuMRPBt/hyzd86XQD7FnUTeiX3HPGofKZW8HPlNzAdbsQ
PNXBx5jLYI/eRjcbra9fssv2X6oUFsciqGVZiJ8wTYQU1Y6PGgq1xpX0/kxRpDjWHuz/swXD86jx
qtqlBBH9dQXS5HM7YTIJue/t9Ct6p50FA7mmZHaIu4dWIi2gcJx8by9Ayfzekcbopi03rVzWWvnW
AxGEEyHDaR8B2qr3E1WARA1kNC0TxEem9iLOp44bJxh4rCymNnzAaWextX66lUJGMDsdsmMPun4P
w4746jrMgiSh0+XpKdKCTWhPjqkx1EtbY0IOyY29JFSgpSkryW+6N2Ls2TSYiI9PIEio+OzHPXoT
CH8C9ITB32cRG8091ct5/golWwM2e2N6a0/MU6htRIan4egEJJh/9R+I1siUl18LqK5htV9v+dCD
/oP330cFj1vNU/VgiEX8VrS/q7ZtsvOlxp/P+23/vufX/nSAiN50JfCkPN1kOuV6dplZ9HSShR7X
QTtUB7G41DsrqdxSdiTSVoAI+zCybQPS4k13YPeLaPKzPa98J1VF/O8zn5NgDNBir+sdwk/z+GOp
kWNZhPmCf3XjM3JbL89BT+wKKxSiEwBBQeP6mkFuRiRriY3yVUnDDpKYEddqdKrcjIxmofNtjw5k
Ks/iq81dRZFs9DTK3Ef4MNr4z++jBLb58bxUy19qHSQTz4XvsUpiVIhdj4V2qqMk65AquuT0oUhW
p0NqlY+2tb8oyYXjZDe5M7B6SIYeqa43SYS8cEKot4qgCVM9oJlvkJxTcaddugi6K2ugK3gKZNav
0U8wecY10vDAC3MmSN3lBJ01lQU+cf6D0JTsOOTC1zJpOiwqtILrL60h2y7cFK7L6uoMcD0hEhjk
Oz03QOEC2ih+EsRYTkTc8UlZJ785tZUcdFukGuK+fzczzQrBUTz5RRuyZ3i5y+On4p8AuboypWyN
Lwww1jnyIlv8ZBdvkuJQ+K/FhwGdS78RkPNyP4mxu8DhiYPo1l7UkoE5jBsvY5JnGoMjQoruomjm
zsxeoyMlcDxbkV+GOkGnnmJlVVlZaNPCP8SeM/wp2YoQSvon6ea5+VYdlNXkpCaNo1jDfimn38Sl
vXpoNt65CeW7N+oFHurkNrblIw+IWsmiBkup5ICAj/XVc2YbqRMi5TsFvpef1dxB5dmzLT3Hh2kV
wEcSDwGV8eWYngYgKp8q1OWOUtcLZym4sWVoSFDxNmAYqPUgRoPjmVULN3os+By3uSsL/tMj9hbo
6DRTAkUC8bYHionWduDl8whmmTD4OYgxtU+4N64k1vAaCLkyAAD1POJ23DPmMvh713vO9DUeQ4Kx
nUYTciH5JHmePKzSSRqe3KZ/j1dtlGuX4x9NGI1YBYm6sgyvhKLx6IQyGEbnjehTU8s0leZiO0L4
rceGqxX8WzhT64i1f9roR7igXvRcPAhd3fReO7g+sPjVrVeQ6BUHXQ21a6xN/IAmgvZiT6ABdIue
V000Y1/aYn4/igB1QC1Exv6ugDVoB+cADuo2P093tyEKf3lfaHf7jVhZNQejWj2tCKrjWPpukvcM
+7JMH52ROn9I0gB3LQrg3pX1wrHy1wUPpcOVubcJ9XX0gTm0rPH6anp/Qn5bJmC84nc1G2+Slvz+
Il3UCwjD2idMGH3DZUERA0AFKyf7hP+AByHCqAS2iDVSd0HEsuFYej82loSFAuBXKXMd6aZqWiY+
lxM8iTwopswIOFaYDHfrMNtyOXyJiNrWvewHnRCwjJqlUen+fDDiPt3X7FbB384GHikby1tnmSL9
uilcdkDQeNXg17DKNuw7bmEJeRScmWplHsXum1OYfvtmXGkpBYPRtOIF+uX+43QCrWxRtD3ilCST
Bs7ODmrGlbZeJ7yEPgfd2iscUjusxZHK+nEayh8vumMl66kpV8bs2SH6pOTLSMOCi+C7PWx5fC0G
Xv4pa3+25W1oWkaVeaFX+jU5rPemh5cmhbiiYwUfmqnGAZcWf6WZo39CorpMS5dPaF6LsrLZcfhC
WaO8GwHC8jmvlaTQ736CvFHl/ahtW4NRBUMdbEHBZzznTrBYJd+hicW8bpMu6SNcLW3HjmIvtMbk
iCgiXG64+2utWfNoFo/MAH5gCSQHa4x5lRwrE5KacIXEaJTknvuwi+wB6Xu1m6S/iCUrG5QKMxdx
OFp/l225FCRW3Z4xFlWucYmadcpeNbF+3CFSbxgsGO5eg5IwVjqLwpBTL3ZOPA7iBib4FsTm8m9p
54XLcJrhmdMujP7EVjAhIMmLeMrebUzFNSVHvJ4Q2nT6zHrkzGW5lI9lTvQcEQ3Yx0gIsGKKoIMD
uHo0+qtA1iylQQ/LAmrr3ClbNf4nhpFT+4Z9NDy0bdextE2AlBslvij8cZ66A3SxrmiZMVdkhjEx
zsdGd51CUmUIJ/lK7fEL4BbbPag3cbs5uXMiC9hXljUzroZH7VgI25hhRbSQ8ImSfKqeYcO/YXYq
lgfQ84FDq/E6twcX+T0T4FX7m/V22hWMPLBOwae8jOKOqlIJ2KuodTRYj6GPp/7Y0MHaVKlcFELI
Ax7EHwffIVatNjgGYWe70aWRn0VDxM6OS8bZd/yhX+wMh+zv307SXdaiP9wrEa/wPNAuMVpJDAdA
QZzQaYVtCiV/hmd/3xlyXOuH/pnYlftoyWjf2G6/v48z16M4Co2hCUnvLilOIWBrXHWfpRXUeimW
IPaMppYJZKXxiKS45fTvzR7bvZhslWkxYZw+gcwtuq74J/HimHwDe8ZMfRULOrUhOTCBT6NAdyC7
UfKuXDiWw0lPtsiiQlaMqO94+n0pb1+G5+XLaDzVIwvGSUSqbjoodEOrLzLq1WcXVEYBVQm+GqKI
swVnMx5lLalgHqxkqgK9wdu6IavxHGdOBJMeWbeKv4rSJnt2dGE84rcZIdzn9ojMC3r0f6WahOu6
K5HW0oiSgy0sVtMYICJC+0HI84Bh8aIOc9A1jys/SJkCsPwkUGJyF0c2rpdkWTCi+Ltm6oTYNuNb
3FWd/XE9gVB87vNEl9XG566UMa2h3s+tJNK5OiUAGqLpEPieyjFGjPzCRkuRX4akh2BtZxui3FTM
LDk6VwakAewFJeoLSy4O9eXyOlIZGKiuIGYlAh7Tv+/yy07sHFBKzO0OS7Ia1+lt+QZeKDOE+p/O
HuoXNZWRkiv6DHswaBM2vUA71ElA3Z//SZLaJOfTHR7eTz8wu9Bq0AVhRVD8CB7pUrEZ0VkmOLa/
XFLvIczmE6+LokikMH8fvGyUyq0+dTNWPT5HTSdXgHc1ZDfiblgNuNXbYgS+XoY7VojESNuMn4KV
Wa1jlhMCSfTiUarSN6mYxn24oSbAx50+qgr9bTKWntZCoSut0kKX4LfWbXXO8s1pZL4yvbaKUpJe
y3yDJFp1+9k8f2/oPv3dUUb9g8bPa2mVVnQufyKWyx4VxU7nWhpp87VhjkLouX7PuLZ6RFKht2n/
B09AoExSqhYVDbXWPMHkecL6s3IL9WxNqmRVSRyN6MxgfCaVB4D5DLtXS4gIzT75dhm6pBeOMLzp
xjMZxUCdUlwQPVSppMfL7/YrGQ1NDA3QSoCf1pckm54zomU47Fj2bmLAYHQI/kLl7Ujon7My9RvR
Ckw2N0QUDD/NxNnlhoXRbN/6YcYr7ir/6cbGS3zoXk6qYg4KeGRVEiulpvSVktLJnZas/k7VNKY7
KOadN6qdF8YV0/rm0HPZIJKYjYkqQAIQRDCudO76z2J4AzIjKgkDx7y119hpfJ7ra7L5/NqKWIgL
52WiNMQZignXr01GLDLOgXqmGfqEadyC4UF+mCMPJZIMR46pQBOMIHCXGJ5IigvVAAbozUv/FbrZ
U3CUedby9YKTCOhLvQn6YU1zfFKMr6gVW4nEAH1hazWx7ZN4rh0s6q1AoZgx+va62lPNRY4kUF+h
9JtmX0TpDq42oZdcJ1E7Mvxsn8zmMamtIjPEPzzeGhYzS725ZMCyxlha0iacqLMaHCZagirJXfqj
qFo3VC2BXUupJ38Lebb0LIpvT94RRRXITdUzSH7lgO5/cChICgFE4Vlw7raRn4Fs1uiUnv01C64x
V12hC21Da8hn4RBd2AsJ26RxZSIcsVwY8hrATnP4J6Evr54ilOny6HVVfnWY3kP3vnni2tVQOF1a
YzxRM8+3uaf5ATastZQOktNP7r6vZjW44srVUnkbrw0Fj7bMmd33VW9L/HrCWMP5wu0piVPugrLG
tTZbK2yALl0emcbZZWFyXBc7Pyr5y6Fqaq3dca5BzoT2Ekqkqk1f0oTgngqkgPI6aXUJf/zpyT50
wgZACErWt5yPiwO4YrPL4rEsAm5Ld4GMfkVt8THrFlNPKKUm++F0VMnABY7T3+n8sqDFT27gDF2a
caT+ObXYd+N+UqYWR8QLgoquPwFc5sbnLjdNro083lE0NMh4HUH0YeqlU4NpCYrCqQvpUbWutkVx
JGQOA4WAJ1KSNOic7ClbTI0AiEszl6b8FehMkA79AoGszTMiJ84eSIaXi7EPTwTM5UZu7VU9dglk
PCNmas19UO5ANedVkeH1PWI5dUtULxV5QiJYBLsoEJn2hEcc2ZtekRpkTH60OdYGKXpMm6hyh1t0
g9HpndGHMEcegdInmOHXV+v7WTgp2atF0/w3uAG9ijqo1B/7X7CGdZ029ZaDVXb7u7tY7QzdTPiD
RVUg8UVl5Q74Azm2tzZleZJf88KKh9HKe1X1Hm7hxR4N/X9vziLNGFsokHxOaqKC/Qd8NdZUVorr
oS1pMdjpTmxHUEhD0gqX7GhlQMdFi9XzIYksS+6CLOQWmPx+WmZiFqABew5dPifKLsILPNQV+Msn
Pehqhx8Y8/G+uXdLrr9mmh7uYaN3h+tzSKvmIlZ4H7JrTz+wiqXvYmW/x/dJggt6EaP7HCtibt3j
DyOqsFV7yk+urmY3P0hBP8PvfhCuVT5mVKfuRFf/ProicG4fWNU6JU7+Cuem12JcWsNl70fFUfcW
INTVpCbBvQZ8CNB5y2+jd/LnghywENDHjLG+ZGIyQ71WXUBBeRwLP6AFxKltsg2YFGKf6tK45FR+
xZxRWafMaA3IYFDO4UUC4mg0mWdrBZFL88gxAccoUabXBAaLjxnbQz+hNWYM6yIaQFdVndO85Sbj
XsEVGQMv6jGqiYSIq748gJV3J1Ta3lIsEUPN8cdLYr74dLbDg4OrxH/Qd0TmJVpAnoVWn5YksRm8
03MP1B0Jnj+JDyjgCSf1O8AltR1EcTVyMW8b62WuaFGG1aXmSgRvUxIEq1aPfho6cMxtr7/rDt+v
ZSaXwmQyoYMxm99oAe85e8GfBewQsGpgNPOuQd85wUq/F6lGJNQ8z+ufHfGbWc1+zr22ySyZfywR
UYhTMLY7I0RjSYUMDJOCb7LLWE5NblXjuTTZxDrKI0YGn3gmgatcfyDhmNWFjDclAKBn4GiWsuFj
FRf9twEJbPQ61DAKS4QMRQ7Jk7RDExLrrVU2Rnt90xC0n7jjMITARNeflW7vOyN4eJuYj0fVkwfP
eTqABr+OABqJ3PtL0/Zgnae85LrDqOZINbUWosZJGoROT6ohIXLyX/99fOIIx/2K6LZG0PpefPH5
E8eeNSdWfi9FmTBlfy0aRn7ZwBQRVXE9J39zak8KfSZvSJJfhfszj/6gMLPNZu4wN9mJhbhHu85J
cKZ3fGUz3TsOgwKXtv4lh+omhcXK8LknRoLFa3A7s3tKIdjDAOm4QB2XWsqjel+KWBUCvl3othqn
O/CW/Amp3eIixqJC69oHbLyDD68k/5DKSoRbmHUAlXYEuHgZ8rjvt/k88HRlPcFjxGuP0oQ274eT
+tkEIufl7Gx7fSgOAZzdDfeomSVEnc5IDvX/QlkEFLV/uo9le919DmTdqdhNUIT1OE39mFtji5nc
riRNUx54sov9e4uEuvDnCWukavbYHIKzoW/1/Mh+tFvfH3sQyEtvpytuWgHmj4w8zY9O1Wt9KuMc
GUotOaT/oC8Czw2XJovlzOS2WaZmU5buowv6LEfvHZRikk2pZcjK3IEtGh5nOXrKhIOgQD/rSJxy
9uTJWbqT0DHFwICD/FHahGvDd5SStB6w39eOquPF46RUO4q1U/qGv3I0JXxXceHOV+WMdEF6gvCh
S2XQFX/ixNyOoQ+xdSZHoKEes8pGRQx+DQASo4TbZ9amBkEiAS+vieP5nAbA5/fpjxb1/ml5No3E
Ifj3hjTkJNXmWd1ZsG3dsmnrEWpyCg9CaTDHjUdr9GuPINByzH1LoeXn4tmqhFlN0YpajHVqwtmB
ni/yW5T6KpSVtHCZQmEOsgBbgf2DIOa5LVStlR8q0NkcNg5YI/NwKhwC6liTARRF8o3thb49+QdU
lwKhY+x2tIc/lWlRDDvHjpvZ4O1VsqfsEIwrdAxsgzu8+gd4zWmiaxdkZocBdrXS5D9noRT4Zws6
dswAY6gQNPDjfz+Mp6jbkerLek5vcNruTDB7zi6VqWtwCFMVjC0xXXa9ZJx7otTeIfVDOaTcSMyN
+ZCFnMjMtYgUndkyhPQpm84w6jAHIcV8flwG0qPsc1jgBiGP6732tLZgo9JBDHxHQjxMH2bInCIG
No+VqxEIjBI1WSplT5l9IacVl4ASV/vKOeeby9+EcL3gAZaXnV5l8FJQ+hvBmAGmiudL1jgpf8ri
US8650/0dSbqBFapNJF+pd6zBm/NMCJoot2iJq5Gzfi9+d1NXQzFK7lbV9BEcSZ4+BYpdAwz2Bq1
TDOBJFh3ktjIRUnZWSX3X1+9JOgrvj8sDTxBzEeXG+vIbajG0jCcj9pv0Eo3K2lC7uEVAQ3uW7Eq
1/Pyt+bdDtmkJLRX0KXdubhtew4cPqyjdqXjfHu5gv9cTff++5l+cQteaYCT0GIPl+1eY3K5jlQq
h1L+EdXW/OrKqmW2jUp2nu0Db7luErrc9Tc8qNbJymgu/kcM4rmlK7gJ36mWOni4yw+XrdBEzQYp
Ge33fzXn4GsBaROQbivGb3LJiYsu+gV/vQSU4EpCbJYjHFqH+2GOwgYknyhUCUrROjqFaAqec7Xs
ic9bloZ1GqFn38yCyv9n+9e/dzs1ntlWBHRPk5UgO9ZRZwVVAtAu2uqnaBXu7POiSrhCo+0PQXbn
vsVKECEil7iM6zbeUquNaB+xhkYzhD7AEDSMI3IhHMmePE7F8Nbi6RMCRt8f0oTNQ5SDGZJxi1IJ
HIhSaXFyxCemFmsekrLGOibxskSIirjjcJEzsp5coVuDxsXE8UZKn28OAZbjgNVUpWrTxQc8y7E+
WxdYvbXvyPj9p5NuzepRVkfiUsvPBui1tWwFGsIU4ZBzuyhRCynhzjGVqq4XNJ4oO7OIA5iKie+h
HlLmv1pcUmBV5kYTPHFdfXgLDav9Dt8i1xbFg+kFSERA6g8yYd2AOmbMkCG9vcSmKxTXhUic6HnW
Wwme9/c2yr8eN78hnz83CVJ74nVhAkx3vqVHyHuwaksf1l934CHqZhq43yLuYZRGJ0SIyt8KcvDK
7H5tuAa5FAZZknGvObapKcDhVGjVd1o61brw+a0OZDQq0dzJDGtKhNe7vOxFErX9GpD3wRz1Bicp
qpNuBgc2aGFM5kvNs89pWhi/kyg28F68gEJ6I8sKykAswQHrftUXYVilcIJqXbzx3isTPj6iDh1+
zzYiGgX7nN8f2LVSWWgJZTDq7bdkluoD6GmjHqCgyAhIMPKqgoaDcIOMyTX2P5qFGILM2MSyiPqQ
KOGv9TXDgiLZjV1UjORFI9deAKob3/NRVYLp6g6l11Wz1Y7RdTXyv8MeYcaYutbZElU2H56KHL0t
tb5GEzo9mAdUz98o0nK6CQfTg4chYpZVpQ2Fc99o6iFAdsYxWMB2exXC5DSMBPg/ee3fzFwPQFoe
M/L73ZCY8eQebr+SEFtn4Unj7FDY3XidGW0qabZEVk+j3SicydloWbupg0I5tBAingVgFEX+MIT6
oA77HlFKO0iW+XXzsXGc7k05YQ3MAMcqfNjG/tZN0MVo2UmTzt7z9PHjnQsCrE1cP3I7Oz4jEtbf
n9/jz2ZJNcvx1oataIz1nrayOoY03nEfz0wSyPaYcGQj5AMNbiOyU+kRF3+dLsIU+OZiqCmm/NQu
2joMQC49OlI+bWDplC+KsjkuFwZSH+BU+WlE6MHWCk9nK7geik6NwejJU8jNuYrTOw9kilPYNz7P
4ORxdXZhyIS28Xvo9Bex5jfYiIHt9ZB2jI65+RO3rBapyH0MneBg1p0Nhh6CN6FO1qs/n8SnN4WB
fzf50nusuOQlDIbMj/UjN+P6UyzKU5/CxIyD27Ds9Kq8nkpOKwMtKdvFIu2dWhJL0YqAKPGhSZNe
ZAdpyqa5ah2CO8DnTvf0f5zjwZbvyvzWPZq26ugntvk/bs1tl2Ci+mhX3CsOdRB2osNzonBpkOiu
TXMs+YDfTq/NFnsCS0SMBoJLxkFiQ9WVw8XOyclLQzTr7v3QdDbXamUDBqGLZA75jL3FaHvhERfS
R/QmJAWAvdz1z8ASLM6mIjj8tSTfvvruJh+yr5s5cpogU7O3OAFyVNdESYQyHElYKQSIeHPbwM0Y
t+aPcxXqzCIbY1zaG8eNvNHRAsEO2m9TeCnIhp6mvYqIA3hA7u80JFCcKafjYwvMxLnFJUKoTK5l
3WFJzZFNmGw1Yk6vqX8DtRxkMx5ZJCv2ZwMlHLkX7MT+djkoXMaYP9hv+wCxXj8KAOmAHS93lAjb
hKw9InQx4Lx7gek05EkTh+TP7bDXeUHRWYm+yZ0TodUV0pP7l4yoJaFmQOAmJf4u9eeiiNBWl06w
5wGiZTbHm5UhZh+0/xHWUnaeHw5MqipUP521Fc3rwG8fBq8dcqKHuvxVJAIBcPkl/OSyQ4mAIT3R
+1NHeCFM/Cv9+0FRpGzjRseNT4ZdPyP3WntO532A5wBpen2UBh/3zbW1SLoJkeUC4zANwyGxGLLu
B9xc7TUhKDgB3i72kwNW/CTEgZEJlM8CQ0JN1ecHUskqsOGxQbS56VOD6cAN/GanvefxAM5JT82y
ynTPg2ry+gngg3lTHETAqctMnaQtHGNFzjqNiMXw2COfsGBh9eKDejAcf3jLkCm6/dLsOi+4mVPw
J9tW04S5QjnUPupQUji94h0uDRa8WnQfB02vcK5Q4pJPNcWUM0DoDRmlVJKi/jQbzPU9nDMz2cYP
iNT91H9WafP6OnpypgSbOoSTkFHxvTIMFyhB84vRx7t3rtQjHLBTXzN4tWtJ28IHyEoyT43/FmAY
cVJEiNiNVnCbazCMH/Vh1Ajh7OWPwRy2OeczT+D2ediHYIF23j49n0wcth9zAakbN3u7amVwRI6g
dEbL+vUV1aE93HhL0/Ca9rG+y7oDSQlVZ8GhJUTWjm/fVxKLfMSf7W1uVaxDgV24WC/7Ijz5f0qb
7W6EcoAc0SrsLDZkQTtdsp3JO1zRtHgRNrmZBpXz8NiInLLtN6as252g0JcrXdhQukxVTYnIB+a+
M1ZraH3/ZUJwXqzCac5PSSGj+1LgaiFppcAJMuyuR5iT2jfB7sSz8ZGWONQA4/prMEcmnctrNjOm
LDoqLGkGHGDD/wdZf3jc+QnVKJaVFbPJCiBG8afB1oNXGEEOyMPMOtxZWqRriBNbBOi+ZaiPPbFx
RNS6yOLOU47Vhj1/D3Mz6W9xGIR/jlh2S29K0MQVqt4XiPl+p+AMNqFHtB5HBcwRAM7O/qaZKHkZ
qiX76byy0Tc3Jg/1ii6PU5swGeX/yVqf2jjfC4kT3sCGT8+kA7q6+JFWmAjsNYjJZLm+obaz6FfF
QHNYndIk92nnqY0Xy1YLIQjm/Wd5hA6OZE7fik1J9tkFrXESumZRS3fpMY+QHk58E9TN3GXODPly
nmfUWhDLz5fFaY0dhpOh393taqw7GuTr0+FUtH+Gz6m1iTuZsckKQGMCHmC2Fq8Isupvoik9X2Y9
8qNXKugXLaxeUGi2GhpDBmI7Afb1sJjSekPXaiqfcMVZpiY1PrsegeAm3UPfNggvozLXzl57Srrf
ro05ZgkqMv6Gg+X/OjpXV5G2/d9ZC5dsUXld/ZbU77MnumZIX0aYrbvL0II2juxdKo3dasUuXBq7
9wewOHw/LRcJpwPbWYJxofmTJwMH1fUbxEIUZ+1LGr+EDWbhGfL5aoZg97B7KmsXkXL2oWfL9MdY
rNlfEtZp4HpadCQBXAiOPekEEeDFSMX0Ec++yZS/WpwpreHC1vKr37ANP2OmzYsg8iDIMIE8u0E3
6oJTQW7gOyMxajkyOP8u3yGVO4OWoG+szO2yqmYCUcXwMfsnlxuHudc8cXn0iichA22GnbZBUmua
x8EIT8n8uxPDpUAks2VT0KrqPE8Jlu4Ok9vZ4AD8TxjOqBNEyECfGfCSYmXsFSFNh9tbJT2lrPNZ
PuD8u7ztlHRtK+5wrE6k6rhLwJm0duH3fpxv/RWDMOzAw65i5QxvhKaj6OrjF2dJdJ2HVubGyEDJ
UTgzDQHNFc8ZDYK3TnMNeXc+yL9Aq5gZGguyUus/Zv1u9/Qp78MTsOA/jK/GU2ZMCfUw77fOiuxN
G39fUgPJSj/5DQbX3MKydEy/i54vQEC0XyLFirddDNFyQK/HSsBsZcR0P7XaXBaPzWcqbHfoDg1L
GzUQ4YBB934MZ8wGcldGccILW6uF7PkJYiIBIoVbD+L9f13wzyCy5N9JDp57X50z7oZj0pygUVNJ
kdBTQ0S4yRRVkS/ApgcImtd1huUyqIaLatxl8ljSiKswlDLeV7AibShSguvfVQro+GA0kQrcxzby
SIgZ5sgmkH5eAg5Osg0D+DNah6GrTfRRSJsc/ioJJQxoMi5hO7lg6n5Ef7dHd43U7jiSgliTpwbT
OR8YjbSBXqX7jFtsyA19iY1dpHu8DaV/fgC6S1W8q7jvBQQ7SkGXkRYWhu5kv2xj9S68JGeKNTMx
KKtWClYkJkhxJigmrxSDhcTzt82BZxTUcKReYwfcu2WivqKmYbl3MEwn+hOYweq/fK1ScO3quZEv
6qIJyZAK3Lfi9Ac72wRLgCmgZ1jIcYNAMpRtw9WNHVWXllIUDH0agMOK3jkVzHRNMyq1UFNVBJwI
u/4zfjtq6VWPc0qj/j+UN0o8IgQfG1INkUIdHza8LoCWJhzgB3639hAe/Krej8/DbbZGTXdtH4w3
ZgR753MGYAKwWb2ZfmpYbpkcg1E2nsavK9yrgfcgyOKI2GUypeRBkNhKrfusrCs6V+6VZPMjR9UY
5Z1KAkEnJ7eqXg0GmqQtBWbUTkzH1rsEv4VUldKJTl2w3yJcg9kVbk3utAS425RtlT0WLENC5NL4
vqRxlbKQqs/iMeU3B+vr8LchcoNMwrrUOWowsFD9y6cgrVjwbmCQfqC4IMbXsb3Qfd+nkkUcJ1Y6
NY4kFLOP5ZzkjImJ9EiEDMCHKc+gHOiiuSPgj8ndiJW3rCrkPc5KI/1oVUf7yv/e71WPGbYEwxUH
WBweqGcdHwmA/ZCARtzZWVKlWZQ/WvdI0K3h/lNiXk555n7XApTyzSh2N3QNhLnyhrXRoNOjcu4N
NpvSEEq/gFjk+ZDSlkFFFWYM3MWdKXubqE3p8pcfM8b4LXSBoBxfLukZu/bJ3kueEnJt2T2aIB5r
oZBNNhE/wWw2cqlVyUn+4Mqp7v8YSMVxz8x9mZFo5YQK0tw/flnCS311fVOq7ySAMYfMHsBezPCn
A/uaAAMOFwd4Nm90fh4xLg89VHL3Kp/ygoRhwrYlKMfvXFoSl2I/liylUf7t0emD3vBY1UvCy3Br
9iYPkz2dPphHNFY5xF0tXXopN1GnHUHlgK4rDf3ffCbCgWbfV2z4cv4Y4ZcJLSg/H8T2e/Iz35Cc
S6bYO8eqwxbhQZm5Ki562LVvvuG7iHev0MdOwDq2zkoTYoOxFzw+6x8MmWSDxFwZG+LNZINooCR6
LnNdNNWsMdomharDrPSaloKzJelbaFY/5Q1uEDtkCjeH1TKeBmuQJj445aYW7dGevvTphxMjcf1o
x0AIBz+13LYofG4G07NSJ8G02F9CcdEzvj/Vk+FKltmviT7eQCsV7AJypTzgNfppa+syprNh3MZd
u6Moe0g8FK/ELocoCev+CLMZKGZL0E4zsag38+m586r0pbvAJ68Fvf8Y4qmMOL2vcndQsDwwEKYY
1C0KXc1bjVyUxL0xV1wlQdBN/lDIBXP3M5Sh+4so/+raUGyeyKX8nZD3xUejvhODmQG0oeqpehN9
s7qeizm8jeIcOZmDfIxQTBKU0tM82e0Ej8YzC7b6DjksgvqQlhO/0r/6KmKAE5rxnVboL2SrPEp8
qJ8UCsYgGNZFH2mUxsxJw+tTMXxLpubIRvX1Ley9QsstxwsYAiQzJMUmIV0fKjvuImA2Ef3Sp9ue
iy+nkmlWbl+MQ4SXd7oPxkq+qUk+Lco4E+PAlnzT+AX1u2hxp9HCBKt15pkdYYReieTQ3Bq7aG4e
x+pYtEq1BGChpF3Bc+Ex6RWu9Q5jFtIcLe6SsEe6OGL4T7ZAiMO2qW3g1TMjSotxXxco1mCAPttV
dozTz3Zz6uMLqFMKhRqagPCO3IG7KnVR9MHpIXeNnXG3IfiDSIpIztfgtV7+2bX/x8Soi6/G9jWd
LD2jiuxU8f/+rd10L9ehnoTqrE7c93wweAoDTYuxPL7xnEULjTBNavlnLkskEv13h3u3959c4w7T
KTSGh1G/43FVh75we3+0ecs2UVUjahr08cuVhjKlR6e35amsI5Bj+naqCO+uafCo22Ic6QYkDO8b
FBvNQct2OOmce21DSZazGtuukSXyhbYCQPeR2rUahlaV1O3UWQClFRtdh1uJHhEPNO3kxdcegYSm
CIf7CcDfbB30Tw4ec5MuFHsOH+wn5neD38w1cBQrB+8ltillVR2XiePx5+kf8qm1XbZcszVxAknN
Os6wBU29mp2aGz2PO9XAmExoKjVLdtaIZJnqEA5+dL2BH+cnlMLJ/0jbcOaa9hvTQZqrLz9omnzn
5Q+qJWLmT/TvjLQ0i1B9b2HbBTaV7APK+zoQLEgev52J0J+l4zIrp2pXxwdtVxoB7rFCuXUKMW3B
I58Odh8fNc30n5Gapl19i/udIQ79dNWvrQfDCMTObWdgBviOkD+VHaHokh7fqwchEmC/8wlOx5Gq
yu2kXqWoaKfHJ7mUsWU3P97i9vBWz9NtZb6tlRBmBseGzM5FHJgbWEo36mlufRbp7FFAzCc4G5VC
2x6bFG84MQiDjza84VsM1QC6syUg21aslUL7iW+ZQ7b9qX4HkuCG8UoAukl9bNeDnaR09zzdtOjx
oEe5pIC0UbFG2A/ct9DM62eeV26j5NLSdS73PLeQ6kaaUxwLrN7G31c/7PNloKwKUgYp9OX+i+4w
bQC/Etfmc2o0E8kgzoTMaKD/vSsxdi9hGNTFzWfp7uSbrQFvcDw+Rn0JAuAchMU52lGqVpFolEk7
OHaPhCOHGRSv0rX/TxX/NDwh1ndJAPMJ5i9mm+YPhtw5CZvuWSO6MMdECjhobHJ2k4LRAd+F2plq
xX9qzZkVTGYSApRHkyndXEQknuOxMX/ujnUBAf702iBbS5A8ow04QC2lbO8T9oPmLcBZ6Ku5kzJk
pOoUyh/iUKkryy2YZ7buhZTiuhVyKa1xiJUF1BHsyldeVYRp1qYOa5ljhkxM70UszfIr2NOIdErb
7hG9Tg6kkuDQtLz7mOYF2EbZOVf954rlTazCF4ZX/LjgG6krkszLffheirJtYU/rar2Y3Y2S88t3
3QdgFvBO3go/ufXVWbvUghyFjsucSawIHOWPezdkXlIWX9amfSGkEgNvya9rfHuaAjx87JmeGVJk
ZRBVn6d/nL3L10ZKn1EH+4wGAdd0IKbAt0LYZWZC0NAO+YTJikJRirM2tKzsij/Gn56elN3MyRs6
g6Ufqx/Lyz28T7g9YBY1Srkmg2xbrK4aLFLHPLz9/bp5IwcsJUgOXSXKg3CjY0j2YgMn1HoZ7xEX
1scCSrDLfS9wUtUNUTVRMv78VX1u5n4gxNa/bxZ+a5GX+FHfTxil6vpVm8O8w1f43wl8U2u9+Z/O
u8VB3DcLOHN+fVdLS5iS7RXzGE09OdwZX/TXWgklqk9LGwMVvgnHPoMj8hnFp2KGABVJ4/lDgdH6
XAL4UGbn7tYwjIP6LtqgT+10/ekMT0vRSlcF/UWKOMu17/Ckkz2bLet2DD/MlvuJGUqIJhdwJs8W
K0hsaWdQNlFSHtqKTb6qakf54E5mmgG/79lqrRWaQwQLwoCm71SnPno7FQ20UKXKSPUEgiNGnHYX
cCRmSLlZ+GmyocQF5FwylX4s5VFbwKnvce9iiP3IjHOU5801mVkJWmDrcJfA8AfJ+GcVfT0/hBxB
/arBobjGOP49kI415fpcO3+rmHPMJ7F5/agKdSWFKyRSinh71tj6Cuvf8ojmihjpzFduq6nDIaZ4
TWjn8KZXPo1hngYShWV5VKqZ7YoBiSeAiTvOObp99ttzJgT5HUc9JMnRKAFoFETesoWOc5r5ENem
GAlo86YiBOtFOFsApL3AHx30zRhyqUJ8Pjb2OTSa29+f914VJrqMSXocMDMfVvQxx6uVWYUCT3sR
Dixz9N5MEUTYOiyAOo2u4VceRVsDrOzB4I2oD6eFJodrao8xkfLfZ+Pz5HIHS3rhH4sFrs7b5ma/
3kqdyI0N9ldUaXGeX/Yp+rUjjtMN5L4LgR227l3Pmgau1FAiynUupZwJmuZjUkEYsMozwlyM2h/o
GYY4eAnmQuMjDiSJ0Ub7/zVYgw/IcrFZ9GQ+MFDZxE9jmv0vrRQpFYf+UREcWzLGmTzPMvmvqNXR
pm0ZvweZf415292LzVIwKIa3auRnXn0hZ3w9EmZOA8Lr2DA2CqyHvCt91cnUwKemzy2cQLOpMyIt
C0VyaFpgLUiDkhDRdU/EPxh4j+nO6eeLSU9KZtF6BrF0OLhWSFg04AJ06b9TKAyU2SQomV9Mkhpt
x/2onnNiURiFSBlYDILehSDCcz56cN2re7oyEvxqj6QbiWgtpw/PRhdqUeEXU1a+hJw1X35CZKy/
n0MJ91mCiOjapaoYfXNM9pQ830koXCGitdAOVolSloLCqJqxzzn7WZhwCTUg+5Gsnp2SMW0LZW/H
+9LJFye1XmKAntq1VZzQDrynNTSLxxpqFanWBHy5TiE/jyBnMX5ddTtCX1Jy1kxDMighN7vSLHf2
OzZbkVq+NaFmsqwRLMcgmQGnlvgpBszDgy5kYT/j82fT5da0y+gOuKtprFN9a0N3kXPhPjvoNPst
/ZcrMHcAOnfwGd3/Xw4BedoSYsub64sgm9mIPdDGNjZbhSzfUOEgdvoQP8u0JDrCbvn7V8a4G7el
Do30WwdaKSvbYnaxNQJRf5cHfEde2E9bkNckSR+L8vIrhFA6kPXxlDFtkbPzaZcWDCobJy/AcrHx
YgWakm+mNzNo0rVjWaLhVkYCYdyvW6nVFtoPrjTpBS/wDQLt02jRl78LAaoNfLwUSKZOALESl74d
uKPh/io5EW8Ikz3tGSzgLBugH/cZmPM+9gRNnWcYIkGPu0ZPFlBYEWRWJ35GNLbr/7TqHXbTYYKT
MHALxV4cHJh2/f/zizRADrJ4qppiH6LSwDbgnMH/EQR1lTlKWQTBMnokMklruYxh21mviq5TFT+X
qX0bhVEJNT5VGdSFPImBUzstKksCe3mFyCE7YtARNtgKdWWraNg8K6p/EXdDJgdqls1olNbwdp96
9hI8AySBnYu+9PqGxdS7iZRlgYCAcLTf9Ba7zhdd0I5Z+SiVsj76NEhc+s0k1Gsyplv652aEg8R0
Ftbu6ftI9T9NIxKBjQaD11UqkODcaq/lh/V4oWGhUTE40LzESjj/ZZDrkdPadebpwEEeLnSxaPBa
dATm5i3mgH0KCquJ+CtvQa4SL/Nj87PfCZa0XYGHqWFQTkEsnlaYyAQHfd1V2sRVRxzx9onyza3Y
7sbrO6c/Dn9jd+BO7TN+p+axRzLB5eoHBywA5rVnQCrON+60OLwNpuL9ieJ47coKDPBwFXfhe8qG
Dh3oIU02tBWS6/SBsuPCviBxknlkBKv2S2oMNsV+J9IDGu/kgxeT/KIoTZ0g2X5gHmyvKYaVarQf
ABI2pLHVBVrHha34cAY3CvSfeV/8rdbyPaOHiB/dMB3V8Yr0xx1kGcYVLLKtJOmjanVcZy7bLc3o
SUWY+COMnA7PRYduCpJNRIOW8t1AE/9g+M29qjFY28rd67HCkfXu/THk8srccwkZoYpJ7viahMaU
1OmrGy9V/LX6A848qTLBGpuZy8mgR/D+ZDuYiChu3CbsTEmBRy4FztF6CQuBIksSN1vq4XwnAqCs
I4T5ywdUxq939oMLueVKMuFlYbCm+ei5WtwSzgJkNiX0jJEwFnUqPqhEGqyOQbfPuLRbO3CHxkmr
LbKsVUWh+b0UM0KTOUk0vYFVSl+LDpD+aNtIvBxZsvExkIcF8lksgYBDyp8Ot8MF2ckFOuwtJAkN
ifqQXbV2elkBNTtIK2GAlI949gW5sy3dgvmRbDnycKZaiGwXc7hrzt8NO7jL3D3VOl3hyb3i44jI
5m7Pw0QATgbiaTE0Y/wc119ERzy4cVqm/vlUBCXKA5M46Gj3v/n3ziv9eoXfhnZAtWsDkBjI7fXp
xsKlcRNli72kLmXVOBWcvup6TG78FPu1wZfDXiDf9U3k/N9YKSrltc3x7MPHkuqmhjZjj2Omet5m
bLXK0KN5FGJjDrLIdCxlAivXobEYqmaDcbABE2scbl84MfgCXmB62K2E7ino7xLAHMx6iqotxXON
3y1IgeLtTvHytqG4FOMpvgQMDa9YQutTgX+nJKvPoGI/qq1X2GNtPQY4zQ8acCSWcUSdT7jS6p+H
gc9JjeWZ4vWcnTuvNUecrR49f0EvWF7jYNQ9bPcarYQ5Q61ZXRSXNsPgsJxwtR5rksnUA2jM0UFC
Z9bqHBUoYcE8YomRSKg7mS53mm0qlDmS45/u5TaqTtGJQVQSt/MWDA4feGF+Z2sxjr7QSmMjFbIh
sSd9QcglBrRflg2ofk+GzFnUqduRLVi2j1h8DAPLfpXx8bbhmp7uBi8YU6KhZwCeGg+QsGl1oHZn
aQyfDwt+gKibgkRGYO+EjjWmpTp0zYUfGyO1anbO368PbD/Hrv5r37zsq1wfSzip3TSUnfbpkRB0
P6FfmIZBZ3FfO5vnVSl8k8CwLjtIwJCVQ9ZfqY9WnEsd7K1cLJPGLSq+hklomtA5ObsPESdZe4tq
+kwMssxgCgwP8vT0x35QCxhFaGj1AGYhpq0wrI66Vo/iTb7sSU0fGBFgH1YP5ohjz7nAsegzRtLq
CfST9pH9URWOUUD3kGSRoGnPPIna2doPNXsGy80CrkT2EzgTgZl0cUfKRp8DTheEJbNBvgSPQHna
kBT0us0EpA4UxqoEGaDoZw3rndNViNgG16mdauWWza9Q8NQ8dvoeDym1MnP00jtkPbTofbtdQryR
drzwkwvlonJZoa/7O897aRKH4juSIXFY4n7bMqA7u8FqcFKH43nuI2qv2HZB674aUeKzIeGO0tYJ
8NcKOuaAASjS5lVqSt2wAyEFrJY16hf7QmNiG9RGqVF89LMMYRQN9qCln1iDmqUJLsES0IyxA6YP
P645nHwXcjS2DIsTwJ5rSgN/m+XYgCvx1pOHDk42fZhu38rKEi4d8McaFW2OX3q/oe+1CyC/U+qo
veO3/ZyABuYbz07FiP4VCgsK8Iw7ZZ4v5TSsqHaznjKayPrUl4qaZHUjzmj+A/PnU9F2z/J8u/bH
fOcaQa6UaswtOVION0Ib6lWLbuVwHM9PE8dhUN9GIOjukb0ndd3YKWPGA65Q2tQ5cR/dH2gRa6EX
Hn3zwo34pKqzdZajGkyjs7TUwl41m8G+leVZxEKlq3ZecPkoYPlpP2gvxrXP2xBr6nrNHQYfwkGY
rC2YG6XYsObqHVGEN9HRTCjjYBAw3EFMjUqKDzfYcOvoL07sHb5Zw3OLgwKjqvSsjAksKuV3sSLu
LYqIAokDE7Ls4rDf0Zx+yeF27sL4OLYJInC3kKsAG3YjoMO0MciwoizXib+ZiJJ/mSoRHjdjs9o6
uTlH8IBdV802syDx24DaaSt+ZJnI8w/kHDpbjs2439yrHamcIO8wanfEf4UedstLxZ4vVqE8mx9E
gtbPpz40XbX+7R/lqZIFWXVuV1hqHZhS+g5aT7jZX5ob5svrc2dmKdFZCaMICoqyRsSKZXdZeMH8
/CEiQ30nPbV4NzYqhOkbFIwFIamph0/DpATRHCqtyf4yTSoFEjz7A9DLdoKePfanHP1HtG33MH6j
Zpcz4CZFrGdVSKQEujUr1CEOAyKzEefGrOWb8WfOMOyg+DFX2JITqHp5zgRtW7UatvxMD+gzEOeW
h5CbkT9E661CDfJRw2pG9HdFAFG7lzucdtt37IlvrQJ3YdcKekGXe4IyUN+ZQFL1Ef5laOjh605K
EoW4YHR5eY6X2Irq1Ogs/CnBe+VS9UyDBVUebcCtCdfRNFcmoyuy3uqVnBmtDj0E1lEYSnAQETGM
Y/LmcuB/wT+RcgakkkxCoelu29EY/wvIGtPC3bL/oi3wfGZmnirhZg4JF6d+zmea+w3cxzsgJCgO
5mgf4Pm+tM2K+AMtIjsvIsNLxAonDysPmwYGsIjw23+xpcccfXRUScAXW/BRvBKvVTYn4w/H/jTQ
//CRS+0x087eGUwKsf4rss9bLA80yZlMrOEIH9iNZ3dcDm9TexR5IIDJr768a3SwUkuKJPDoke2C
msZJsxFichxuOs4ohrlJ+vX+fyWGntbFhZsHMwp2NsJaxxwqjuFd70EJN2Zz85YTArr4OdFap+hh
TiyQMLwicHd5POjqCdva0CAznyNqKwX8j+RC4F6xhnIih/hKTa5g7K8aS3+cP+XJy4Z8g9PuOpeG
AEkHEXCNCXqGTzVIy1wkpZQEwdKcWrQX096pQa0KEchnWMQeoPjf5rpUnIO+SY26P0A6w5xh3eNv
ROBdSThic5S/sEx4rLsXi8H5irL5mzOnQam8lrtzpkTWTVbZxasmwAC2cMRzt5NOU2fLJrv+l/Ey
kUHmBg9z441tPiGzmu99DymOYGgm8FScIsswBhiDf1hlq3sN80nLE0Vo9NP0vGzye0Y/J5zRyljZ
lupXZSE/T44T6Ia5AN+wktLx94DgbYdNqAeQMoPK7BpAp41KM4LB6AHaAhk+Jr6xBfwaqBwAJoQt
Pok42ZvcpdzcFFOdbAK3riGYAR4+I3tYQ8PHXWocHVd0p3vIuf6LK/T10Bq+i8TsJ1NRvK9Rq1sZ
VqGcBKQ5TECo2R8t/6vgOCZEMWNsn3+t+rMcaieOiVAT1TAAI1NfwlAhMRsYPa8ENIPB67DCoMUK
gFOsdYos+p7M8HP0fHMrbgQzC4U9eiHVr+6LVogjL3imBBVEUTvy4VYvccITJccp1GAMBJQ2myW9
6uyqmW2L2QJNZtBDyIMPH/Z8huPGk9CkHcN5h1AaVbVA2o5aiAcLL5cfWR1+rnb1zKpQKmN5uGP/
cYXM3jA365gqZpnM92wwfZUYcQOdQqk+w6+AeqIJEsjaTyKReVBjlJxmR5emI3sm0ShoyvTMaMFd
krBqdncPadohEx8BbBZfFw+gGadQoisvjcGUxxV9/F9MXcsXRUoT5THnH83WWuoUTuw3OFn6uEKw
JHWbjNPIqN4CAje+EzZHe8veN1ERu9sVywZFrOERLlCY5r/Hxp5TV45KMg7Qno0Lv9Txph4Ffg1c
//25FYVfVPQr6W0GJd3/PcGLy9pOeQsEPAkAVzosM4pYklil0W7SeQ4vcRswfaFMtckdkh0J0Auc
k3kXdeT5qL6ajXGeT1qBuxOuRkuIV3xb7PeX5ri16P3xOHNRrbrd8ms1MNBnJ1WXE99muCD3yFaD
N8U44kCXwaCi8OtJGSiLk6ef1rnQBaekAWl4m4PnutQXuZBMYozP3EofcZvMib5RjtuA2KgQeSPp
0ntZRkjmRkKKNnmXpVQVbQBBUrDH188X0pleiKSHKZAs78PjaynzOsekmoBEvOEbT8kiDQh1GrTk
wUXce66UjwkTu+pgQZLwlee2uDFN29Xy2Q9nMrUEaBpL9JiIeW5i/RIMDFxp2C1NSQozxpf9EeYh
bNkQlrDHrTxeg77tLw3QA2TIqMOFF+DfJYrlphgWdSzml+zTv7zRPK2oAICuRz6EMlVX8FUHxx8+
dtTh0kChSnyeydjG7nt1rnPt7zHAR+uQmRKeWyvxQ0c5+jc5tFZIV6How/e1rejl5OPiGWtD4dxP
x/BqMjJSwny0wdKJdvBZ/ifW0xI5c/wrPJIU2iT2BdUCIrOIU0xO1eGTKOWXSWzcIu8tORR1wrn7
7n4LeCNWbO2kKD66lrYplADovx2mn2exp7GMCg/N2Q54G+R+tq9UOUBmGUoYiCrrJTnbwgoyrrXq
i2/r4vKHgHcVloZP0dM9pOFKntO7cqwlHGKCDtr1RZywHm9N0bVhSrQ7m+AiPMpoTUcX/9IKxEPe
6XhCGlj42FeIfC3MP0rPLQ3FuZAjI4MvRghpI3k8VKEpUkuQ6rMxLOuFOnM4nIWm0i4dx/fDuaW8
I53bqVIKs9EyRZyBGLkPhd7d4D+1dJ9wYWrPEo8BDVACScsPJWoQL0wZ39kWp2icTCcid3ZljrNc
TtVf5A/ZaveK7E3sN0l/y1Lv5g4JX2zyjwiFHAhGTLTWgmbt1D4YRRHJMeBSNnyrcf3Czvjrj5U0
Vuqa51FS6sDnYRdaVDz+iNsc3dLHPjMmdRofhUCh01RolRkLtzywmHcLD1Zoy5JuQgsleqq1COE6
UFwt0lwjLhnMQOq+nblgspZsPzjRX54bA8EisqJMP+QapSfK8Cf4SAlXNDDI41yg4BBP/RxBHu4n
zZaWfhPNx/NFL0gJjySke/1I8Wpt/t0L3RwO3czoCXY7njM3DD3xYlFX3j1QquvOlde+mpAmh+ii
M/rMV3S9X+ME7CgCQZQYieyE8noSyI6IABPIGFOOL7b0lID5oJM/kPZbZ/u0p6jcHbFEGcYwJyyL
8r6FAX8nTrm2bCwmnoB6rTU/JvSpwl3vDfYP2nv5QZchfjbBK8KNLQnVrp5bT7lX/GwqySFGl3Em
hKqvmkocokR1UEKeqael/R2h8qSiCJDMuH9Dh0kJQz+GqFk9qnW9mFJsgiSffDxtUtdLqaD9yuTq
OuWIpuocwEId0yHVrG49OFtbce+wEHRWoCQnQQ7fFBkj215O1Xo8M/L7KLq7H3mv+d41ZHUIumpm
LZQOLGzN4hpJ/judaSvHgDZbZLN+6ZUxtHzipQ+MY/gfCcR/WVga+vFtrK2YrKIIPrsNp2DrDLh7
7BnqshMha/FicAbUKfTg8umxSAfBl5UOkBUZwo2zgsXiLFCNGm6k3LFujkxI8rH7rM/4OfpLNvhA
Hx2pvkpdsK9L5PVcazJ8aWCtCN3ukslz8y6sz6Tg/PeNFGaDU8tNOhGkeyPshJikVjDmQgsGYxJn
+5+6XPD9a7k5QP7Ic+H0xvVe/9cfeOr/Avrj6SsZ5M+fhQUTqKzedXktAuGiKtVyo60h6boPS5Kz
r8vD1ZIjp9262HbARQU+8z20biKpB9AJsjSxf11vYd/zMm7r4kOqdhHFrCO7trD4hZJIYTmb9bLD
PZ0q7vSgAb5d7H36aX4DfX2ikYcXcirCqS86uKn59Suovcx8SzZRUrq+cAnguhCU9Ua6deEu1rQ3
UjfqKFintju7osn7tNz4G9ImlkCgjKW4+mWABzinLBpXj5VpyXtgW2FXNu8/evlXeFFvL1+G1nG0
BWFICLnJYwMQZ+8MGkgGz4Snt66F1drbeGQiiiTXfJ+xknbEPghL1819shSvwuC17hjwztJ42KwU
L7jScC34nx2HVSBZ6XW4b3a8D1Te2Nu+pCROWXjWVntdXswLeR52qKm9rXMgsdXqGJNKi9PjxGPs
g7quUC2YrKhPUSIw+DQbrzYIuCabxN6GEUtjTcHE/n4yZrzyMDr4BVNqScJ1Mlwp1jMvbj3kTC2U
WEAXfy8W5IXbow7Lxvoo5JmyDGy4UR/7X+8yLk3M/y1NEcDCCsBQP1qDbZ8yi4/e6MMEXdJ9IfmB
eunWqHp3R6YcAUlVdrprpz9qVwtHwL1yPPqCSnKzgCVam9mcMWU7iBp6JBJJRMFvwH9CC3cT1RI8
iHtuokMdwWSR9exWTrfMegnpSFbN+WpTOTkF3GKzp2k9itqYLy2w/BbFjHgXy8ll+9M5p8i8wp+h
GcX96mPSGu/7+YOEYZzGGoJSNdWFRKkYg9nozrA8bz3dlcFu5ELSjqS8nZ/f4L5QJu3iY6JXWiyJ
loV/+dE6Kr9C40mRifezYt6FCPoATJ+uOT4Qb0bz7iZENArOg0KS0yGNydmyGsYFAb+SG7A6bGb+
cdMyw+VvR/KCAWvoq+KGGvcJOMhUc0eYs5HPxHslbRmiAA63D+JnmDi7tec0inwUKUoKYf66lKdN
+owdRoHfnys2V5g97DEnztmw8PKc9a1BABls/Ohxu6jABtyWzJ9yhep7OsgrXivFQ6Fdoqg4zVyN
dRWMvQnoN5KrpV7+CSkiupDf8n6q4nFzZkhrr4meIMHFjQ2Q5CF1GkTGSzI5kUyXjYg4uZ0Cl/gr
U96XUoNfSlQlupoT3ze9xKpQ3brDZ+atCQ5OnBOWn2VXqiDV3LgglbHm4PjfTzEViE83EQaCVbSm
bVZmrser7uetj2Gey6OQz3jclZoqTiIjZ58nLlbJ2aVpV102fKxSIdfRWgYswQ3mHMIFkqgUIUvA
tVeNb+9MV1S+uyhLd9un99Xxg2nIxis5Tv/V5Hl5+3wmx/al7ZdRWTqFqY/aBx2b3zFGSK9fzZOU
yTS9P5vwObyvCfELw9SHjKMixW28CcS0QCkz4IvVSwHAX3JsRImi9+gpTbmbKejr3CSTGV16fQ7t
M0MfBbXY/j+Sy4zifzePjJDi+snifx68vbfTb6RaQLgLW8SFRCj8HuzaUnKDdFoQjWuABOp+IYWd
TWPjfHEsnmb/edw40MgwPd+bEIMNfTeTGT2yQMSD9JI0HLvvavLGuIbClZv9GWMHo2r7jNpFcI+o
XdxyZArqUdloY4FYRa66zB9brwILermTFbaNCEvYcY2Z2s+e98a8+QTAb/Lc2xyIf64EWyb3+TIx
Wbslu+rDpL7kd5a/lHNkJW/E2YKdeGspR/vxAJtNhCY7q+WNoH8BTiBNncJLkM5zWhCZMDA3qAM4
YV7mKb4vbjM8tUCaq/dfOrBOZ6csmr+zF5zCErlYXfWp3KaUzD4IfcRH0l2kfbdAlGWoYJKBHSzo
zivxLL14ksQFOWDSxYXiPYafdyI9/1c0TKVKaE9no3InkLBXyNGiis0Ljj0dwgcBYvRmW4iZ3Z3Q
FYMwZuHpoQ7a04M8DoBFSaGeDzQkr5rLTSC9BrpM7WUHpYw7Z2FLtI6zd0GWzgp4UQnDu3MvRPJR
AjhALZlLr/TeG9/NMuSYl9Nbbuf2EJpT6NsEv6TNVkmN6UZ/RRwbaFiW78S91ZVPDcSbf6ldlNeg
T7WexZ9VuXj0pzyP6nA5fON6Dk0o2ccMtp+3DOo3a/t81cdENGP9iiQMMfwksy0tCQ7yZIjjRHCo
co/Ls6Lgra35U4Qyu63bpgWW2AjknRQ8vQVKUgA+uR7cVlWX0V0fDTpmwG8Nk+6qDHxYnA8cf1E4
GSdI04ikt1cXQt1wY3eb4TPxehLG+bSlDxBqRBvlLKKsDTZ0coX7GwyoM4Z/9UOuroxVP05u7mvq
4PI8NPae2OAc1F6vVDIRIskng5psdSQxJ3BQUB6WK/77H2bC1+uj9HkUnAaE5/cjkdIkXpnLva+2
1H0CB5p/tA5EUI0+O+VBCSf/ztalI3MQRyKTV3xNcCsSSH4SugUJmj1yLUzDaht7DeLHSLyur3IP
cKIXOc4edSi/WfIx4IW5tanUC6oehbgBKIzxcOnTIYAw97SW8lZuqo7yiX5YF8k74uRW6Oleva65
MOVgJHuhwUmgfY97x8JLWMe/LOdRiSjwhopGE2Xo2QOrpPQh9Fyn7zXwgoWR/oJl1iFauVCLI/r7
1+HHTVz3YTwBtmRDh3DpXsR6wsO3iyHsf113AEBZgLPPT3OMH1R0F3aD01haNhzWwVLffUhVMGSo
X4XCPEJYTxRI2vfmiANtTL7erWVE+D2+j38ybbHrgYKG/Hc/jM77HRXQOCdXFI2i5nwtYArGtDBf
lgrQdyeh1eY05qOFHp86Syhe/zQ/bKPyvOuO/3kOEkY9gUd1PCrfyS/+Gabc3od2pBsNzvx8TZMZ
N0fckmDB7dNcxplGpHZF3sXhQQaEDiSzeAF4h92O09YKsDV+s1Vo5dv8slUDhUjBfCbcHmnzsiyi
qH7Gh+PhtrG5VnTYLlVWsqTd97bpQhmAYNuDVV1g6f6ExAhmqdDzfn+a8dCqSXqbpC47rqnvBLun
nApig3Gz4+zv0LKJxkzb8qFNV1N9cG15IWfWnqcDolYo+7cqzE5dnJvH+hSlE5LlGlusbuBOgI6e
RxpRC3GvCOKTa5dx1pjXUpWW/soluCHlM5WnOVZRIg3ox7tnIMhWOfX5wuGmP4yDlUwKPMlDmEIY
0Pxvm8DAhQM8sukrIWIWvebCoPAc8nS/zyGRk3OZKjbIY5ASxUb3rSYO2kR603H6RAmPsBiHSZSf
3X98lWen80GVYwtW0jNJDaY3IqSi6/bOQk9NLPqkXm48wBCpEi2u7VN2ObOvKoFfbXaW68tfc5Am
3o3pXUjUMqE4hcN6VL1aAj5s6/DXQ9KF2VB4lIAiUaOz2BDYmPkKq+/QGL4lCkvZlZLw5WYZ8gGG
O6oAiv3996P2A2wk0Y9nagFjA3vbjn3/GVDwnOJe/sDr0kCoEGNFLosHs/RE2CyNrR4vXMKzhNyL
NFLcugrk6nVdyco/1t+x+35bsHgfsZzzpk2t6XVmJwTZQryiUv29C8+GV61lqMeDqTvYgnSsW62B
K8+NlRUR5+/mtNm01Iiggb55cHAix+HuLCSTREGx3ihhkgD5eeAn+lLzzwBBAgGqSgIUHVqsTDtv
sGN42X1G4cyqYL+ffD7GmEVhsPFxBvrHHWQiYFpLBuYOGDEyTsdPTxsaaGAU42LvXp01MY3uOB+y
2+ASsocEW/+OptGMK58bHs+Aez3PLRyymJZuVkXYQQS2mcbEqV2UB1wUrUVVlO5S7p9ex1NoxooO
PIde5YDwVpOItFJfnlGyK7LYkWnvjASDhruFECVVOCjeHUKYg2pVfiwz/MkuKZxGQYWYRthSeAD7
smDDouj/QCjbDVFIxlkIaY1NuLbasDG9BSjiFw3x7guS/Dt+vn8hU8PW3mux+RRCgxQod+SYV5dz
t75VGL1i4/vu+PwD7bzJdoygGla/TOtqfFpi0SX3BMR/I4BtPhM9CJ46MgyE8AABpeL1YB77bb/J
151TENJhf4dz6nxc6HZenIPEkKxSf3Ee2gC0lm8Oo/CSIa8dVng7fG2ku04tlkeVvrH70X3WSis/
Mfp0fmabi3yn3c8r3ceHjCyMFAsvFlV9N75ogm7wLqNxyZeBJvx+PRiusv36U8a2Ck6q6Xkcji5l
b/wX0i83dcoidHbPof+xLtu3+1TXvBBBPV8vhgc13EGgknMqXEmbdJKeW5zGsAsYH2DUs2O7QLRu
+/88K9B2f3ryGrXaJwYcYpJDhzTrrwpT+aQUeYJf6N7+AT341aD3JzOBBLO1bLCUtDzS8AElpeQJ
8isH19vyXj10vvOvJx0NJkBHOEDxk2RQH33CSJ8Bl7lj9Wwgl04rRuLvP+CPm23DZ8cqA+53IoSg
NYDd/2wD5n0JyaIQp7dgX9R4ZReVdpNGm/ADHuuLGm7upxllGRpEkKrMSEHpt2ub/fvNxUU13txY
IJwIgkQapOSJThRtf73NHzUn7koo3FJxTI51R598icHxr9n8ak0rqdFeZA4cP42AYingIohPf/V+
a+qImoNBi4cZSVlEzyS5ijMmdashbv15FEgh5b/nFISBWUBS+BwIeEQsDw/R9tB+c/nLvCbNMHJu
KgEJxLx7cv+V9DeBvCuDT1d2EjYoG9kOJgwsIRiGi1eW1Wnl0L08ZIP7t+LaBriw7KS7sBYorHBX
M2c5jDBlOPxSACUhrlcV6P3sx3fntBcDTgc+nyZLlmq/iWFGfrxG++umTyIpfHN82yG9x3pK5ifo
G9w/L44bXyMLCgWfMEgch6+ghuK4KsESLXpP0agJwKiFdWJQ+CuSW4rG2l4xjV3q7/TS9xULS44n
i+MX4vAvNkglpRgiBCBn0q/UxLFSHihOnQ50tbXXBYoQ5KOmLwfwqwwe+afdRLl/kXyFRwD3cumv
2DR5KI/OLbwxozzmUXx2vqHsA4XJmn7J9YslkA0upv/bdxiTlRKMYSMBJiv0kEjOLxHm46uIUdmC
PD6Ev37pipbCRv19fpSy+uPhWHTEMeLSlchYxv8aQDY2MwMJziWEqufJ0LeccPS1hmRJzaMwJm1r
jLm6pb6l9z84tCrbuIU4rVwjfNsSmWY/cSqHQ8h2JURgiFSXuUIJTRN7WoObW3jIHKimgb1k6X/y
xJGmgUJfVSC2MCJEvBjvfqNUpVuAf2qkVUaoLaYVrpPBMan7Iew5fCr8C2690EGdpZ+nAsPFZi0i
Hk6Jqrs8MjIYBU9jlqJephIU7PvYCQSts9RufV6zKJojPNybSIEwulF5vgtnu5I0DxnnA6yj8sud
qo64DuGxtGst5jgIzJr8LZHaMNjrSxqx17PHA03b5TlWwAedEjzTJ/TkmlLgsFl/w7fhfT5UbP9F
1zoCyBJAt7rOpVwaSSHPqDNP6uYHIfLpAZB3x4UIio7q39sJGsr84GtPHuqNEN2wAYFgtaEyhchH
1b9YBjmiV749DZdeuyJUKS0P4RJuHEHEFD9Tih/k3/cIti++XrEZ40y2tlpdyJasLyJBNtoygpOV
9j+UODUfe1F49gKoQLYSFSTzglsXTuItVs3pT+pZINmj2vGfgr7vyQ66IJv8yAtfHNHvm40whaMb
kVZTfe9dH6Aqo6fLnV3ZcVzMAlzO3dWsQpAK8964XXBTlL5+Kao6oEqO8JptDCynippj9jdgeDnK
P1hHrhrHNlXQsM7BJO38Er7HkexqOpt+WVjGK9e6IKhVQRrhdzI1fS/GATZGq55D3yPsl7Lau17H
pt0CxPHsuobGZUJuMmMa1P7tbockRYE0EsDwasShtg7BJnXet8N9M/Lgu2CRcqWDcrkQYkEkhk+D
4pljcbxcnjIdwx0KLfKCV2ltZfQxiS39GGFjUHsCgaBeuToU21XkoMf9XA6dccyZXDdc9YeD9Ufe
k64iy5kesRxmsyXJd4CG8t5SaJ0p9W66sBI2Rju8X+oCvxiGfnoZ0TlkCkzZlOpDuQAIUqYVPsAB
sLyQ7YgsP9mQfGsx3efDNmhFH4jGPbBuyzgp7Z03dqQJcUPVidaHehOpiI+m2fX3k90EpSJTXNHu
QBAhkFgr7zDljN8ISvlt6d/vFqGdH9DUcE5qdXZ8Jmxx8hxWWDLdQR4z0a18X/Z0GhKfoGYMDQwi
YfRi+S+fdj/F3P61UYlPZaKWEjUk1lcMlTz0llgm1gbCMG+4l/JQ0lms3j84OvBcjhMjImBSfmUm
GlwaDuTbskbhAhM2rP14TQFgyJSaBUwfHLcfKk2c5JKHKUV0bVvUoYCeCaFXeslBNGfJj7ZGkXkf
vK59tL69TZ/z2h4vIvXUyh0bGJIndUN3xMR+XAftc1LaT/xGSyDG7iX8ZTpLbJyfx22m2RqUc7O7
Yb/2d98vxzICrRqLHFhIda6VvtKghbXXSUI/F2lY5Qxinb0O32As2O+c8n/JwzD/igPBCzwzlhxq
H7BaRzq1rklye/NnUpdG5Aos/LwNC3EonqTQ3NP046y+OzWca1v0+Eh0EkDLNcxblRFmieKS+UhG
yOfyVWRmIkkJ3aKxOuzGQ+w4KraocGm4ORehWtVee+jev9IAONGth3veEeBFXc5HYPGc+RRS63ga
G7ncxPlFB51Qlf72xl+xv9AcMtCrFHpub5+ibuC/SqA75VlwuZDGOuo/pVwSbIDxC61S4R8QgFl3
rEi31My/WXALvK427gML3m1CCY6lQKZOScKKqKdVpGSyHFWapRAWXExHKseI1arzUC+G+MbC/8o4
zG0xMJR04yu/44fzP0sRpGfUicXzF9wFmbVowFL9qxdk2KcyQ8690WOW/CvBzbw/cua+545f+ATw
cEymbfMxTyIsm1YD2AsWIoM3WVJ7uioxWuHt2ivenz7EKL+ZeeIkJUOLt+Ad55k4HqyKEtRxR/a0
va2CttqdwU3db4vVEaFhevSACamFopTKIlbbfFzgIYnItF1vgPTEwbKoKzXJe8tSEwMMT8NyGyfJ
LMNqBXSeZyetuJWFMoq8IlDmepw2q7OtFy9zGeITlF6WT8ZB2v+yUeGYkS5ngC3l7EBCp7JYuEIK
Ji97H0FIRGUZtpICPCA933htZo03Wpod/EJp3KGR2D7ruxvMLJ11/0x41ySckc+afmqviMZrPDhA
0cZzWbjOt1zEzvANxtiAqUAxbtpegN7uIV3agR9D5FbXH28uPicTmgvUDna4rzExa7RI15G6IzjW
ORqCq1ohq752zq9ugFwIuPBvTZASd5NkeV+Fl1HXtnQZ6gUjZCZyzeL7lYDTghQeNTf6joVcVUQA
mcLPrj34fxkwa/QaRNnqQz00MXj6zlj2/N6cPq6gVDFlZQkC9U8Xpvo9NsQF2B7GSUTaEtwRLO0v
Wtgibb4P9m8rA/3h6c9Zyq1r3T8QZhGFInIe3P1oOgRcTVLUFLyOkl7u0CSSQK1T/7QIqKVZIwEa
qp2OHDSQH3JLodeUCGM29U6jWZiS6tT59d/8ZvPOMglKic+BEd9YHS+T6A4YIXYOjb0jFyq5DVeh
USHP5xhu7NL5w9Fnv2rs1v422Xp4tnSlZl2HCEiKrVLqvHsrS9EBp9dHCGUtERTaILu8jwD61Yci
JZaLh4UimDlrJWLdMZs6ZRSmwLmj3ahZ8wYk5Nw90uTchD2zzD9rWRY3MNSzgUosCcap57y0uwIK
IQ0GM2B5nZQ70xmMnsOnAETB5gar4nEWx0ztOVYqYAWPNzx1xPyv8Pf4Jh2XGsoJr4pfDzwhRGFK
95Yd4XW8sU+Tro83zQWnDDJWjRW3AqC/f3Ncv/R+eneFUj+0PYictN9Dk5RZmC2Q5EE3B7W67h5c
1Z1TWUyvBvqMoIc+hTOv0/WY2EWMvm2gP+GqUwfm51sIuZZKXnFNzDjKiKTP0HvaQF5d7ECR+HnK
b6mKzeTENhjBaM5m1hVPKtFxpVqZeqw3EsSHYGGkKuH+Ph4BJgtfOpppTpW5iAstu1qtGM2zan3Z
fivMEAp9FyqUAflQ5yz7U828spQbcUrQil+0Z83na4i5z6Hy6i61io8BUjEcsOUl33xNNuYjT8AN
HWcI1ImeLVwLhDQ/rmYVNKTyPia26/1XQJ9raWucg2FL1BMUtypspSLhz/GOCZ3rU85CUi7/nwfV
02tcKYf8SH8Ey9O9E5slX86rPv44djsWQA37nwbt9c6nk1GWhlon/G04NkDcVa64iSB113k2Bckm
zuKcSYe62E6fGbsjMJiBJ0FY8zpqZTqPFwfFJSajal+9hPcUnhyAndgYbURZziev7/CnKB5M2t71
HW4RCyRDmZD1BwDPE6qUgXRLUtB933nlFSQE2MIaB9PMUR92DSdSJA1slSvHiiIn9y3uhnpwGHMU
Gg8ja9rsUPqV36Y7JdrgyGT4y/bq66MAMW2Sw/0vYJE4tkzzEguvGWm7Cez7f3qb+smXsYFN8Znw
sNlYj4ih4kOmeWsqIPMKqa86EGQ0kFXPBeuzo8vpr8o/z5PxDQu8BYWLnJA4JQal/cVpkplAJuCK
udw+c/uBUbqId9ieKPBzlGweU+6BwNqFqLcK8bf8aCWYlpurweCAfbIKGs1Jvm8mWYsB1EQdq8Uk
fIEc+2JU5gZSgswOuRI1PDQCjZZ6CODBYuZbsjHggltbE8YRAdVk8sIziEDDFjCAj64LYwdB678I
THcc7PbfdqEx03no9bdQDXjX6zltfO9klObYMBmwMkCFsUxkzEQ28iS3wxpVTerCZRZQatj5aLDi
zcEdRF8QYL4+VpNrU0JlrwhwmxuOu8QL65fo36i3mKg5mJOFL1NjBFM4I+ojt1PcHl+6T3C++sPg
m8CKBKNYe1wpuKwls8WrQPfjPeZCRpSzDU2Ufpjl8D8clk/18cxcfu8PIwKsPJ4bZKvIh8AVy5tV
UogHjB8i78dIy7pb5mAbwdz1nuvDlHTTwkH9+1pnoqTzTmIiVwD5YvbA/aRcqQ4hnGnJWhnjumyZ
4kLl6eWskwZgedzf7be7DBmqnwxTF6ZrPh578qakt1gf73feC3Wzhek9O3jxYnY4YTPGFYeElR46
rpWwxRaPAaOVVE2hxICZuaT2U2h1lGulXQAm6piLNM81wPnY5eiBjjvq4K88WomncauRVy2bdORC
gnnqj6zy7Cu0Pf10EUofESBuQ9FVyCwG4TBVtsld4TsHIJO+5oVAVLKxN4Q6gnr5Da7YcLlGp1d3
pit1OznNG3TE4ap2aYrBY+DLKgfByC2shwAscBz6fbTgb/8/LbSUWby4zAKqjpdp1/YLpLR9BJ2U
4jlJF/lD01yr9MihlsfLKr6yWwUilWDqOYebIgmYhRO9lKJtEssOmsB5AUT1uQb6I+73lEqynmRd
yE6nd+s6Q9g+TlnH1J8kvWxINnd2UgWpqHu7K8zDvmqSmOy5og6pxm+YP5SBMznLV2IaQGOULhZ2
eszK2uTWaXG/GZcBB+JqlqQpvfEQqwcSIp02U8iCHLivdiy9HxjJyiy//1mi3pzhnJTFUTJ3dxVL
hXHQVbtgPetX0yEiEEi6/NqqVg8uk1VDxZvjFKOHWNhmnHgt7hjiCSocPowf0lJg2PIArW5m8pwE
HRTcHiAUv4UkjZVPMvJXONglHrAbRB+BL8UMbqvId4UpiDgnIKCpiai5hB/UEc/ObiKuBlryKwvi
R5rO0Dj0fSnLjpoG2MaD3dxY+uVOIBVX5N3Ek9ewHEOT5WCmOjrI3koatBR4pAaa5ApzFyovWZJp
BXRT9ulDwAIZBxOA5b/W+CRPdMFHL176bY0SClWeT2Ktc5zX2T109JPD6Gtc2TLi/7sEJ2/Tqdcm
8bWVXpqUWvOS1nciyMcqp5y7zaewF9rLIuPqVcEfvSW8E/8tMpCWT9iDqIgG4on11IDtmiOp6jui
Xo+mpJRMKAVHr4HzqKveRfU+ctgZYsDZiaZ10vcY6dM3EEgwUOgWhs2AZsqIPTONzFv3esIvDNOc
j7+wrkkY3kxUYw4ootJgl/d5piKCr9MZNMc5V3z5B1X+looyo5xAqPSBnLp//JlNAr1xtOMfWa8O
IpTikSB2Tf8ST7VEsIBbsGuHNV0orMMdG5dPpDV9jk370igGjLV+SInPZmwEk1URwRow5jlw1sOR
3ESFVA0id4jKqyK978TKBGfoWB3GBRnmSnhszPFpTPC6ERQDV23pXh0mD9JelJz3v5WQs0bNE7U1
1hFVoGa3BfKTr0udFF0dXScQZO4AUKBzWGtfsXZQ486kuAWz63CoC1xLsHWDRBzu24OXKdxYny2O
RODicI3lY8I+O1JyDq2EGlDSDpgenOlSg4OWjhKXC9MXAnv9MFobZRxDUfsx4Yz+0J+hzfojeUET
MF3th3BUYBvf7zDeq3NfhvYKCEWki/23RlYuOkoUehgFK+HHOl5FYBcdN0aitQVxcu12HA4reFN0
KwWu9q/26adrkGq8DydXXY8YoEVt5mkNj8AoMNlGT0mRLCUuAO3dk3sEZGTcJ9RCY7gbUo8LAF9T
Q6yGWXKuuDf/mohLMtzxeuKzW54mJQK0V7Ufb+19VLKBEZgsPRM5fO45Cq6jkVNBqdb1IbB4Hc3Z
BP5vpOgSmb3kb7lfAwQ/84J+SN4dWhwKT3Utpc6zH2pDgTQv+sGbxBXapIHxafYMB9f/3ZHPw5Ai
nkbPadxhqT3N4N0MVNUwHfFernUCDFrWmioEg401sx9CxiQf39/u6KkWSH6WULudoH787mcU3f6G
GJxmQioStLKWKogRvcGxv9CXOiRevwDF0PQ3Um3Q8Quevp5xiPDkqr0z9v3Fk3UI8HsOzGrY2Cjr
2UqaPCukLmWH9O0E/CZch3XY3kRQwJD5t3mPk31gj+6VgGJwhXCbe1Qb6S3jV7XQvPOoO12hGhCH
VGMQUdeC7DKA9dQ3CaM0da5tdDFLxEJKrqh5+45zrwhV3AhruTpQFnKly2wez7Or5HEVaHTLvy6e
hTJlatQPxzZ409UoFbwzEaLtKdAxjRNhKDlu3sgeaNGyqN2Ul5Droxdo+f3GrFH3C/RRkA0zZ6zJ
xyxVWmKRFVXz2zjgIWsCXQ3Dx98N4HvBSRSBiBneV7/HE58u0Fn4Ht+1GAC6T1q1U0laCTAaAh8G
U5iiIM6xRMZ7wtWFSrofQvXkyi6NXjII3tV4gHYjsBiTqGuPHgx8y4YbsnF+4qyGKB7ZMUtoJjR7
m6XOFmVpnt7epWp7t/iQqMv/eGiR5QpcXvinejqeWan2/NLzvPZS1uc7klPN88ncZ25nt5Aqpy5v
zX63Ylh2oU9iMdVNWUV4CN12lOEhLyNBMuh3X1oPuq0pWyuYz+Rb6FCKDgMuoBSl/wIDVdes1KXC
UpvSfrqhAzXELlfYuJnGIfAZNwLGUbTGrvUohCRCIliJLwnlMBBjy5DZC4HeQW2wYmbiCYbGFD62
i3+C2G05GVkPRXRGTi82l610PwvzvHDg9ec4Ash/6Hg2y9EauBldcRmVr0ttmHeKKdIv4UFYMdJG
v6mwEr1tHF/o6mYE3iNIMalSrDwMwdfqlj3/yaXiFyvAZPAmw7UQi+twsbXgJWMMWmkAUiRlXsmH
749a+AmCbLvPkIMkFiUzC2Bs1QGXzg/oCY+JsX3fGX1/7eGy7LkrdYbxW90XtkB/CBDFcHmtU7Pn
4Kv9UEfBXWeisz5/6n0dYI0L2S0dNWl0zGQsXQ0paQKq2MKC39zNZuv68NDLxhuiJGlB0WFYPZbx
RvudDdqMz8TNVIwPNWZVezi8fnY8Tkwhruk0Ck3aHuHKBG0om7K30wqfABSQak4gXzaFz7EC+7NA
ocfGGDbz7z1ESPIZjvgx80pccwa9kdh6hZ57rT2SWQOJswPO7NzYFW5j30xYjrTireBFKjbOvjVA
KfLtj9sqlqs2dF3yss4HEKjUfyR9hUaw6jokJiWrZW1ZwmL2a6tLtM6Ras7McLvS0N5v17/309SZ
3MQTiE7/W0q/Cr7l8YR8B2tXr4rs5PCQWielzJ/H7otqmhLecaKoMu7z7TcFyrryfurCMb8ggZnY
aYfsOE88wSLXeyn+Nj8nc44QZdfpTplMWvgmTs0ib1d0iv517a4VEftzOfmO9o9XIG5vI2Qu0b4I
ZPpJdO6tNq76Lg02tY47dsaVW7j343EtTI2RUPnhLuTzR1yxGWt3GIyRXBfGjQuRCNqTVRPXsyK1
2D2AhMXTogKPxkxn6/HfXuOhpxqF8m4plHynfCmxL4pXKm/kKrf3gk11ES6g1eDwXo+l+iU8NF0h
Lq/gAhwTbNA/eveS15P+3aID8EMtC2hfOiwcZs7J34YwQQ17ddcRj1u0ihEX8toUHQOGga73W2jJ
Ib0Ygqn5lU/RvzP+ycYwvxh8qrrxnBvpAXzqjC9EKYMYvKSHy5v9mFiImvMknGlIQx0G/IrFnZRS
QSzi6CeI+P6nl1+5D+ef4dCsZVp5bPix1QPu09i4dpF2V1COo8tZ4g/gLMlc2lBqNrnUgR6f5m5v
vJ4lK9gEsnKyPHT6euNF4ewW4nBnMux7w4PQEt69IeWv5Z/FU9SyfSJOOcNbrkPo9O4kLHiAiM/A
wCQuMk5Nv7UkPxE5Uz0oQLGcof6WKycJibJCmFBFoVwTExNXTGO0Bt5BXZKez9ez9u823BNLNaJa
CJ7uXeyXNEIB3Nohpl2mG98vGKEWpbXYp32RXQhnUhBe4YDCWjVEnRvLG0c7gJDgrjw7O+XqsOV5
/9G8ko/GwoalMX/NanVHMTPe4Tz/OsRZ0Q4OG0z4ofIUOHVaeYanvWC79K3jCao7YIAH5UiMvZ7g
pfwcwC4jS5YGPXtZ4zAWoaYzyaVqo5hW6K1otHaTBDkzAAW9Cr90pEvEolEBt5hUXR47CcOdh89v
m4eaymjXK6jZM8pg9LXDWXYvDuxPBAS8A3T1KgkedT1tXEeVjGf1RUPHD8DJ7Vk8WGSOkMEy+jSM
Lfie79Zz2uLAIkTnJx5FK8LM2AV7eeWFCKB9vclDzNrDH/uPNs/ZOPMVitAiQHOqrKJr6REc9dGq
p0TpT9jqdJyXdDwB4L3N4PLsXccxvA8n1mutACcUFyqcXdlOSogbSDX7D7eTDg1DRHLPQ4nvRxe1
mSzU07Fv+2CTyvVgX89MS7SwmFUhZdanPpKVd4pTvNcUX/9tlEqNcy4uxnobqDn6Ynfvr5pyTIUh
ZHxVxWEqKQsB4psI5NbvWhUCajE7ljBqOPMEAKxIoydc5jzyzu5Tafrr1sm+XNWTID7qSSvJ/fLO
NjRmO31Py5T5/odjKC+8hBX9GAHa69Y90+etgAD3E9LDMF1sOoD/oPfENbz+7mZysratbrds27L3
1KoffkXD9NAQxsPtlLoXVzytCfi5+8cFyt/elGHjvX8sunVlTC0tOXfelbhBVOgbn8wlqpZ3fBy0
YC/x6BXjwDr1yQEFJJgTioxdw4us6CFGSXuynDJOObgSLwTFJGz0pSwL/9HubAUB8BoFQX4xsYdf
w7RGS+jS532tFkZF34Tsb53lWuu11Vxckvv9rkkKv4HUO66iWtOjO7mUN/nlDXbXEDqfoKFRDHhH
TmaAF/VSXJJglSwomqoHOW7PBRW5S0z34nRJ4Y5YjyOnCAlrQ6bOFBRZt8HFiGAOaTAXPVbwzpJv
qVR7fuMr92svBiHJrPrJ/7qBbQ+voYPeFuFFKCVOv5YfcbTUFc9rBxeTfo91YgzLi3+iRQQjJkUj
CGlspWS9qAONE2rqRW2U6P1vaCMnGCy7gwpMuvAVPZWOHk4eKVOhDv3Xy1Ye+NVWZrM2CgEA5ilD
i46x7NYSw4sOrVc47ZVWPp5E9SSWEdhuNw+Sl6sOqbdz0xE2P0xIPF4xiX3zp7yOkuzNC0g0e1cL
wwynRCDUp+fEssRtzFzFnXUdW4uSPI4HVJPEcL4v00mdmTJLx1jUrMLI9vLuiiamn3F0w+SE/BuN
KvDitPmCW5hP31Y3GsgoVyBc0WiLnIxibU/B65hZJPUPuDPONTs1rpqfYGwEjj6tGXATXq5/9lHa
ACjL53jMjB5Q4t1odqMqs7OevUCbPgomhfVXo6d3R3TfDnQG6/PIPWtFB9dOLqWFuzobw0QV3ewR
Rw1KdcPoyjGzvm5FxpWNbW6z0O2QqmY9Pkos/XbgeEFkRentpwaOA+ITsU7zZKlSP6bKuvTy43aX
QXcBwO45YuOMXTsEleyKcDt5gyZ/CBOd00oj+WkgA5f57pXQXk7Rna3TTgNiShe1+h/ICJuYxS7N
kIjyI6T9UkywZ2P1SEY3ZgCR01zve5x8y0ngvZusUfQRyclhTNZnG0eE6UKIeQ/nxvKZgk2Y4jER
NYiDZtrOv5hqFSnIgkEHF7dzdDKxGgKL24EZz3GvDLRwJcBNET5Jl1cdsUWqFKejrHQusf5btjlD
KWkKP5RnzZ98nMAZHh0Y6GlY15kb4roNXRAe/c4to/65uAfU2vh5G5JIg2lmNqBHtk1uSgW1wWWR
4315Nl+TQTYndw7lH4jVsU/yX51I/md9ptpMLa/O/KwfiSuqAm14aia4zs+HLnMolXiAzqZ8Anr+
XfZmYmHft+qByiMSQI2lo/JLQMmGzJTCCONLBtxaClrYpy6f0nvxkQuBfIyaFt0nGgD8KxocGT9H
orutG7TPijzmOkDApHvpR3as5XObLF7K1X5yf0zu3SUIdGXthlKnxSP9Tb38oO1tQxwe40pGqOQX
ihKaK9FoqES0LUs69CAkKjRvnfFUUDvS/2kExhM6VlTr0fHyzyq+IOjFfM8uzfUVoWrObBzKoz9s
AD+Ar37T5l3Ufps5uxGSvMG6JY88+FtTeEgwCFA6UzjFSdnBBqO0dNmoJ2MaFOshL62QperLrCYh
Gn5Mhh+V3te1HmxnlyWIj7AQerR7CCjU7lYDt5RtGBkYA5f54SIhsiRjX3YN65u990bKiQsSHCUw
EBTpgCQFjSDr/Hppbhte0nprO1bu1vBVd5/0N+e7H5cQlgWrdf4UFGXrCoGmqo1nqOWDQkOErDWw
TM8D0GExIN88+X7yyoo84mQQGYPFD3q4cGX0slkFKEgwn3KSQSCeZznpaV/LVvB59OeeBXD8drz3
ZUpZXNIUNnHYhtOWjwOgrAzrm3jd9rq87jsTQ+rsA1ELQMshGt3is9+4nnl31RxyCZmu1Qf3341Z
yDwrrGGoVFXSq927eVj+zfsayvEWGNr8v3zmtReTwaguBxGxREjSUiKlNLLO0vWE6bwUOnUm0S3a
PTXsEs+NEHILUtEB3UzuZo9Gv3Ap0HGKTIUNKKhe9nwWNCpYCVO/MxpUN2zVGPX74I1Cv3N8zBg3
QK6SOlV7+EQNVymem+fcJGwKQZxwzYb8omg25phRpEUavlWU46+sKyEF4A8kL3gG7JFKubpVCsaB
3DuFIaSiQX1X8X+lIL6e1hHFCMZ/VyoVAp986sbwaIzek3JJEUrC4vUlUwjX033V+LRMir90yduT
qkwBAtasfPEa2L9gcUdl+xnbQn8nRYaCbo0MuZZwakxcJXSigT/xKvgcHfiLL8u2yo7Rox1R2lRy
dbUfjlCSR4a2bHNqPCNYOScwglKXI4EHp3Dvc7J//ETYZEPhsdhZwYmCjVxW2QW70/0k0J8fKt7G
zZQeIdGWvzZ4vxgbMluJ6qInFq/Sr7KGDHvNts/DTC1suj3dlcbaSmK1XvyIC8yAeTc1DNa98ZJe
3jNxZKPNrkz1o0kBJQ76N1YvQcVcUIvwRPA5GyB+v70NC0kz/njWVK+HdwaaNoxcBShpqn9iVJhp
zLbHmDHl6v2MyjqMwoixeNxT55PXuOh0TIolVrPkaXv5RjWGVidw3aBJ03BJ7tudRa9mXaBYYdLY
wfKJ6Adue7ienF6fjjcpfXHoyrijnIgMAVBSXeYrN/JUELrpOZb8Vp0Gtp+RFlNAHqyeH7kPXITl
LdMlNt3167+BTrS6KnJAoct0XhIvRovZMcz2AU2ojECdgjSPNaTDMkez/bOJsNhsFNfFmdOyKrKd
m3F4IPUwrUxgf6qyOIyjX9RXNE22YwOmtbby3Q/PgpnKIPJklX2Y1/e4uJzMiU2evPPLmNkLnta1
fs+fvrSP6lOAmTfF1q86inUuyilpmC0ts9nGKIzkwE1KsWRjk7XuiQh0ljy4TCLFJCHe9L/IZksf
+gqcKffiGx+95CFwHb0NeSYZ86C/6IuqZT/Z9OGG2PI0bt49nC3uoR2XP4hzP95n2zcogjrKfigM
n971wT2J8cT/DGjy/YuJTWh5SGcLo7cPdklixM0w5HX5aR8sSLlNQi2ZCF6zlwJAe1NiulZmhWeB
WhcUpMjhFcyjkIyUScqbKWwEOf4WUkOg70o21XMiWrdCdjc6siw6f6PWZrMqm6kFi0tOsU6wqZhH
qtRAIIZ/q5Ld+Sic84Ot1KnnkwgFvoymOBWilyz9q3O5QqpW7xKeX1vKwtvv5U2YY+RGGFcQBMW0
jSVU4+4fj+urWVVjeZb85IHx0KS2zX7E8NNJcbvrV1zuVai0oYG20YxQ61H0MKMGmy1180WPoeEA
c+RlLsTwzhnOKQT+yQPqBOXu5l0Rx2M/mBt7kEcvI2rMXw8kAoHejeAr8XFvnCAN3Mw67Wcr42vf
sDVgDi7sBMY8yBI9iEsKtueAPUMCoU1F238IMdnWL5HjtB5Ooq23BUY1oce89ttcTL2U8AGe/bVn
lQu70vUsZWcobU0WV8lZ00f92MXK2ETdKyCiifmjGloCdgn//spkO7VTxiHTXz/DAyW8hyCM5icZ
pRE0m9eBj40LTsHUBSc9aKHqbqplgiRPgZFHL0MTDVpG8scBm5uYyJMEQft2LamZFTSpsTPlFoa9
YdGqmbsqTn4RVi047JcudY9fY1eOd71etEcj8EFohenwsR4MIZTEicZlGio8YaV9XcYhPaulIi0O
ZTIWfSICxDz5ghKO7qmjR56ljVbgFP/ZPpqP2UHBMtvhmMVpx2MTP6JXqlCqc1FkyO2nflIIOLWW
mXbZjdlL2xAgFyKHdWbY2BgzZCMJTAWD/cA1+8ErtZm/zMlZ5PCcG+I7gSvNnViv+J5hMkdzzVpz
2OjmvCnQsP+lS7JHKuI1Iv0NMVrnsiFHKaffFkX51A1iMi8bRvyMTYLyujVyZToBtRrUA68bwJ/j
8X+ljyq4dsgsoywjN72DoZlsByd8VjePJRAhbS5HVhMPcpQLGSZT8cwbDo3siuaBE4wtR/rtuGS/
1bOrgbKF3AivlrYk0yCiArNJy+rPXw7iA/1ApZmvn9iSy7ejULYD4X+PoH2bAwmb1tlFkhpiyF/d
6yPMWaTjSiSXVOmbVLYWpGmB9MdOzj5zNa+jcfgga6tc9GDqo/xEKR3Ng+vanhQDrJaL7OLcjAs8
AasbQpLERyDrInssiqLCEgWK9FdYTV5v03pFzjL17c6XY3qf0CIwO5oXOK7KTUZMtfttd8XAlwDE
m510PsiHW/Imwnai9Bg+/7DCExc+YRBMi0Jj2OvnQVbHFHBCFnN4tYmJlDKnPeMBdKuyrGTndBjJ
oAN9NUnseSqYrULeBHr+IsGpw+AWKnQ7Gk2rych8y54UWfO2zh1hn067X6G7bvZtSh2p8dkTho4p
iV2Q+pf6SHoGDZ/+foy9pZR47kEn3Jv7FU6fhvBi0QeJ6HwwZ9HI5/FEXwLd+Lvs+JKBJRP17nrE
xFG8OLVckOuM30bODEDJnkSAGldlwpZsjS1D+gDmZxhoRsRPoNQHyb0gJRB9bcNHJcUzk6TdyTuS
PHLZrJKKPnMCMuKWGXGAQZlkzZXQu7Joy+Qn0GRA+uLYjTgeJik+qP77LSgIMeZyOQXnXc+R4uW9
jdvsNnYW9X8HynqAnTcZg2xDrxeN7SkEc7xNhQxeFVa7pj8OqpU+V62jNjh0hlavyYkDac5qK7gw
tQMRMr6r7uDb2cePCqX2ilkNpujQkDcoFbgvD8fU0TX2BC00egmUa5IxVkppif9Nc0G3mvOU0t3x
vaWQkGIxQHMjmEUacK1/9TuaFeQcBpMjISkWUjV43xm0AZn+jqPiRGTAFLLjv9K8EX5Jcyv2R/7N
8/MnjTQtiunzACIlg/wfLj6ecBxhF9Cx6Y1t2xa6UCmYpS9a+p9c7GUEbJVItDKfqKYAaIgwg0mn
6FbNGASx7/L87rKSpfLfZ4u8Hr3Ad81qLYakzmmHlhZsV2TrhQrzW/gqJUzqHVCYcBoAyP88MgxT
W1WtreL7lZM62y36uL2G/S/8RQfIb825hwJVrPKx2htGubRpjsZ+AukYUcdXXn4TCAeBYLYiWbE+
/eLgE8xAwnyshpreUyHf5375UspCbFqihwGnjHsR7s6ngHII4anknAK2uRW7qpM7bQEecyaiKVtE
QPKMN/YS8iA4Aj7eUDqvcuB/FLKYGeBlMJoJSWAqpLUCO4zAu0K5hToWQ1ehlkw5nH+nqSnzdY7G
DoF7GYDVBkH61k13UaKmJxXw0CvEICcq1nPi2dmjiIAE4n7gjmIoTg9zfjmJEDXkuufnu1MHKkeN
rbcGNlhOMc5kafNlQy2G9hX3JjGSkO024T7UaCrAxw4uIGQJd4kIBvBTMkcGotbJJpxU7YKh5m76
+wfYCy4nuFMKM8FKKgK1GCbxPSzmM7OSbT9sDgBa+v7XZV+8y30IXW4HGniKBHNpLvcMCJ/fwKz9
pmeIODOEuuheqvBrDGrblxGwm0eUCG86BvmK1Y10DmgoPPiKrA4KyW23QdPlsT6UubeOd0dFHKlw
U7v052uAsyb4587e3ySzMp/K8xF8QDJ/WtK4Bn6XnNhYVhtfA6yO/ZmnrPHhQtWBhGBDnW+TXdfR
cKvzlevknGXLPxQ0LsmaebvHb37Pd19FOPcUwQRF6riEFlbfQ88AoEoGWTOMOQHhFZM/Bk33yvEp
+ALie645RdDzTjqr2wUQPo6k2m1ZclKUAcG0iOOU4OISL7tcFnAU/HJsNHE0U2G26Jz3Ftk7M22u
W0gk4CDAdvJKaQgOzDiH8tuTNrHu3i3xK4FHY67/JkN2q54fg6cUwFCi/LodhET4QnEEwdl1rYBu
A01i6ZQhm191FoVt0VtTKjgHt5e2P0SE/Zn2jKiYRzjUmfl7iVbADiaP3Rz699rg231Q1EH6CY/w
oGUFyaWZsbK0s8Pu+HWdASrNZFM4rxAY/uvTqrB7niH/Sfp/zbk/vs/ln4Rru89beoA9rZllRqqh
8/lF+03UBPUTQH47YcdQCEfCdWMcW32MAqXo6pWbguY5OA34kXMYM6BxHmVuTT56arwaLj0oT7i3
heaRTAiaCYhKsfHdEj6CFC7jnY0a5lp1rm4BDuQjWkThdw8NjOet9J0pKyuXPkQUv7RVZPKTj+Vr
YbnsutoL2YegyhE1T/2mRamG1srqpfgvqvO6GUz5cbIvyII30vIhcZ2DWIVJNy5W1tq3Z/3fz6mh
UMWjYk8n/edvwgapKb5WBnVCj8MiTAxXObnFRNPNRAVeFlRc4jyxPy9FowQ5Grtgdm7QXcdJgn96
IW2xJWnwHCqaXCgRFhAui0CucxeDLxe12AZ5+JbCGBQ91bwePOARdYNyeiM5Tncbag5YpRLeNIbT
FPc8FkhLbZBTd6N4jJbwIMBhCk3whCg3M6o+od/tQzN6ORiJ8zTLQGXhYNxu7HK9sweR+dgX5b4v
fqkJCMXUoh8lkXM4v4AFp2AjmIhliXqSfEDTF0R4wTkdFqMHkrjkwcpZ/9OzajDlPxalQSaCAGzF
Pvr9t497wZCHaDW/ulTudDCYk8cCXhaZVos0qlT/XKqHDMFiTfcD+gkHLMzEN1+IHa4xmJhEZlNU
JRIy046eIMcwqqgEelKrkSCI+/xTrMtoCkT8WmnSUdkwEzzYXABfHG+2yNtnZ6ZRROAHcPt24mHV
OkOisu/qu5ch8P50s9Pe77h+0g9qM34Pb6zmSj8Wd3FsACxBM0thCuLaDKT4ukfP5tcg573cRpzx
WKIqWeN7qOvPmq8UnnMeJA0bKoES5RNWqfpLcpTp4VhZTNl7+dIf68UibO3HePnG44x94N6e+k8C
20R99JgeNktAvWUMUg8u3QOtwoaLRLHJ70VqrYMkD13dTf0229z22wSROf+AQlv2/UcYeXVHUBfk
Tl2OQunckyqkAcWmuww6NkitKG1JCfT+ZnFf+hrPFbvbu6JqxGWMW7LdZxMrjz+DW4enRpx0QJgY
7FZrE87+6uUg3toKn2GDKaksIqvSM4AXD5HedrYBa+yNgdyfw/Pq6laCRFzSJ9gVBa5kmy7NOJSO
yt7AoDFcfPF9f7+/mAgW1M9B3ygO4MJis/FAXugsGZXyGkEZ3Ed/zw4R26myYZMDSRkKNIY1Va8O
KpUMDyI+2v+7fKHSQI5VxNQXhlE6frH+ik2t6ja5mV+SG8hhEquaQh9fD2qhospLF8GqdBt6bfri
yuxVgVCsV+g1wnKLjHNCXqwiviWSmSIzwmHyK4eqGzROPePw5kbpi9PXLQS+7wBbK2u5lT0lfmi7
ZDwswYsdp+ZHSjMTu0HnIjIuum5/DInlXCpTOtGVvcTRkfcTX8bYiInL4hn2jdT4VuOsBbpFuY/f
TEB908yTnSnzEzmQsnYLChHxWlw+HP0ZhkGLWikrTnr2oOKSLWaYwXCj8+S/ECeQ3MgmWZrsbNSf
sN2p6xcblfkx8zlOKch9Ige32PDiHAjWxa504OPUwSDW23vMuEQP688fvnV00jPsKwXewZ/amh5s
GUnLxO1ajGTgtIQyI0wNbhWjm5zgOj6xGTzflgDyQiKKb5qJRnBmF+11zNg9H5LKMw+lIugSqi/y
HNGoWXpAPZjjZK0sNuL+GNl9f/kCak8R3pztRMEpvjRk4/WgDMwVlxuDG8J3QLVxWk+mlZ+p8hDx
bYWe68oX8Ig4YB4EJAmCciNpbFNp6ZNwCmS/KCxeBA4rGwEKen3iFfJAI+w4oB9yPv1pQrYjla56
Ib931wEZ6dTCtMqPDK/i8T130Y6b03P6QBHWvJB80lQLgd2oL2wZK9YBKzssyfWCgzOinqO04VrK
IUXm06Ar0rT3K/2fie533fAH0WcmpOY5LD3nxwcAGtG71L4RNpb55aaf5xRoWWy2Axm6H9Si7TPt
bNvA/JfQuzJQjojZyfKPHa/GTUfHDP0DrCRYAr27aG0AWGyUT6sPAnq3Ap5ChkNDRfCCLSPPaDgO
REoa0ctMVvlIRwtk3yajnt2TF4HtTM2iPEt01ej6QPwyTbfgrHbit8Ahsmrqa9Mgwj+Z7jbh9UZx
JkEFoKPmM9Hs54lVHq+UhZ3hjn7TrqNkxr7KYue1ksy3zycLG5Qhx9AfuP/21Elm/FcTVPRNf6pH
+e7x/8we8ojkwbkcExv8fyEXHnwPbQE2HmTDtpg2uBSwkyw7q7aXKdvzlewISLcYJPfOzFkFcsaH
2ixVHz6L3ES9GG7OqKEOJqgEKQQ7WO2eCjyoZ6bSDllCibO03n9q2fCxAsSamSZlPVpKxNRE4MxJ
VRKbywGnOL6Mtr+4Jx2n5FDN+R5Amt4yQ2KiFqEW5RV8c6qXD9kP1spQ2aevO01QVubd4hvPLcQK
eyAFErZhS7YUklKhK25oKu/HYlROn+HKewc2GTfAiZ4pQ2q9Ef0vXFxee+l2A7fMddhArlI/OF9t
0w3mgWumihlQdM2ht973Kv8QsFxB1rrqyqVrjY+GB8sJiFfE8uGpS46u1RPXihxzg0s+NXwpeypm
WmiFu9w+8/uc9FmUMtb+QFoYb2glxoBXCHawfc0VfgHzZLD1Pc9uprDh3fobzGGg2M1tl+PMQ4rE
ILah775DAXc1nR18jqdOx7s5+4nmJ1wUBnwvoLCqXNXesYyK+/35VX7d7/q3EyIed1YVLQIEtr2F
X7LgEOsbU7VIhQFBQMHzMJlrrawGyPnEbazvDcM+4YToklDydYduGbQjOnZBFebpRZOrHt5UERBF
Jad00hgso45a5RH24gFb6Vwp9vq/j1JQ0T3wEHNN5lvT+MIMYwmLAoFGZ28tQtYfb+Ehhuas6pwr
Y/p/tgI7UQctaW+dUMC4kJnOS9/AQZhNbJqI8YvcBEIorLHCbUsALdVQNfeKlh7bkxs4L8k8pjUY
0mPibcqizyaHZx8RIAM7s4pYEoo74pHi80RqjiRI0HJp2ZwqpFUp/Y0y+Y7RYfjfSNPiJXlxX5Zb
/Vcn1HRyGkD04RFpsVjpx9Qibae38dU0wyvTXSLkIedH9r4aZM1tgpMsV8JyziHKnneZuiAkEl01
6+8AJZ1JxBJ8VHEjpAvNw+kJDouerGVgOSLDDxdVOwu794PHWVg3RTEhftFPfmIO8DrXW01K4t6D
7t2P4G66DCZVHxlrrqQ/o9xbKB4+50/EZqQmK9j59rvUWsVbLZXnNsa+RDEDG9ZD46PeB82Z2HoB
9kcFoRfkkgiAGMcbqgiLprn1eJqZm7LewEVwooxCiTQU40exR5H1kleqv9/7sMjvYpAAp4rCpWWl
S4XDTciljBafId90mdKOeXZncg89OPLFP5IGqhGIc/G+obLDOy77VAev509ZqFjkB7lh5ig3v2nN
lpr4rzw33eAPfpVBugzEncFip7gh/0mjDEHK7MPtectPINpynaX42P4KT01cvwqnHMH5EjpV3bj/
HO/EOIupQQcyKZ3WofLNREGMkmz1zz8NTI8Mo9rx25JYVqgXpb58jujLM32swvw3mrFsFmh0M7pB
sq8kSaGz9F7RhT7f8u4k27QkFobzpLs/CNZfta4T/LE0hqSaw/H6WRrdTWqIfNbnKM2dNFFodWVM
TNExrM151iooURs8w/Ap0WCd7G9MlypZg/klbLqC0TRQzT/zg+AELW9Wu+oe8DNB9jVc0qN5PjES
RB0wLzSN37Hj70gRKadAjIOMDJwofLwyqriRO2DarPQg+Mrzxvf1Z7dv/+c4+y24L5JhuvgT67th
5TS/842bM++VKxnaWema4kZABvkAFCEAj3XCt+7iYyf1C5Z2yKZlsODltLg4tPtL6V9Pg4GF+1Ar
vEMSdEE8aTjdlIe1Jp7enZamAMYR9gmUjsKTSk4U0eP9wOpgvKE0cSeaFbOAlrhqmKRyXYlPJ/ax
oV9fg71xmKKoojJsCTacdjpWZKnMo5OnUJcgVqgkZeeMqFNdqw3lm3kopo9hoS2mSwydMDMs2sky
z11KKnuZzBhsK79FACQYTCV/iT3BO2wT0eH/d41RTZzCCQKCEEGKF5blTlgWo071t7Yb3J4dW+FG
hOFKiPv9qiNxqzB7P1h8XVxcf8wtPiQTJXGB4yjv+9LCTp2Z7sSl/auPeF/npRdKfkOX+nKB/eDW
Nye+NE9J+pBxjUmN05a7ZBhjt8JDw5905b/MTyChUckbbuaCGVOW/nGLMkTvwahObt6mKToLxGZl
lrh6STfespvegRrGlxo12dGenQARanIfrImSezwq4VL2KoGI7dtBTcz1qk7MJ3po3c6sNomf9w1m
DL9ZE4AeSWUiea4y46nAF1f5iIL6dI4t2zyCsU6/4wH4Gt2jacPy8BQ6CC/oN2+apiOIydIAXCNf
mOCY4vpMSaqyJ9vY+9jkPpmqpt1FuRHpG5IFlCMsClyVkfgt213pggDDmGBAV1GxuDtnw9gDwQV3
sI4QYYb8FA4B3oRnV0ReSmluGhtxchyynWz3PKs7wWci1tEmI55uKKiKjKBolPzu3CZNrv+1vbLN
qh600hZ9vUohN2dCvRl7SNZkvtux9COfrM3ViLusxFs39ZzyWZJdRfuBeo9j5X80uOPSRrfwoEan
PqfMMYw4C0i10+o6uJG9LhYY1s89jlu2ZTZqR+hoHf2JvAKu2bZpb8IjiUbFTFXw6rjyyas4/2PE
iKK9uuImRzRI5DKfusY0t4RTGp7xdNMAPQcZBpvoXYi15QNSmgEnVpXQdhuC0TO/G7fGZ+3DMXER
OdU7vSRX/kgur+XHRSpL1Wgw+L3nq4exyRNnLnuLvM4/4wOfxQIxmmpzgLXunkx6pcTxavq7M8J0
Ay+jTRLhgfjTiUh9qZezaqA5CLYFBlhOuKn6sCjq5f/9tkJsjKj4ID92ToFoRup6s3LBT2rH94X7
OpXdf0d59a41hKAFbccEwW2A5at1opWw3HpmcFL96+zca4YVKJ9p7SBmW3zPkab8lQjOpnQ/2mP+
X+D26VPQfjCxY2YYhHIQNTYvq6LH+iHOk+33hzqISHg5IcMTqjRKQrWHGnbGT3bE3kWXfTYU9s/9
5ONj05d62cGl2Q6jnN8hBqnHD8LC+M2TmCmZkC1mzhyszckotwodUGINPmli8Qxz872ZtdOJHuZM
aFVZlYKMLgddn/L2zBvTUbZAwemEAyrrJQTCBdLaZdKRnui+kF1hygt4B2xG58byMGeFxMImIxwz
PaDdyU1Z7G3LKNX4/welOwTvfjq96002iSkbOjoxeKWOuiLuMIFr0kAJPsZrZ+NNTTVbT9nUQvs8
KUFdsJtth6fsQMSCsPSyjVCpPPNzQRjgQmpQoeuaqxakpoaHbHDIzMBxz8A4NOoDdjXZKJqxb0Ku
sXSQCJbQCARlIsigQw/DkouQeZFcbHr+jxdqw+QiuSs7xw0N9iuXzbgLkq5sonAm+j5Jh7r27qOG
fWXpgT7twLn3dxJ8VlBzvydTW5R3p89HRiMKlFSQjLVXHzNTvZA1guvjK+RHOap+VCnNd+7hm81g
PRTVacHgi4JHdobwCeUsbj6LAqTpbXEvqA57F/n4YJBdBUAsEfXJEyaDgluZ925vEJOPqj1KNRKI
3zHWsB/5XlQitaRN1X0XX2TIzE8cYFtmI9UolloxkqzICXGZxVdSZ6GkFdyIgkyOrr7Ze/Mko/6H
CtX4/1xLB3oUkTd8lR9u9O1lv5x8wRVEjD3twNNB47Ib+Y0wsBRT+9T7RxZXFHb/2m2S0y2vO9Sh
PAh3lvNgQdVNi3jCKGPEK11yVoGsmm5Zycwp4a5TFhxmM9BWRVjVHzk8QZTyfszqpuM6NZV6fR8K
h4dVmmY4cegnQBLLthoQjUzY91owwEl2MoFjidJy+phLLYGsZUR4mD7Xhu7aCt00PWn+ZD2krFbg
m/kLS3rDo5pHYnF+Se4H3MKOyfiGVKFqOGoZKhrMDJy0i3fk221KdixX6ZtRE6Wd3GNE1UkVPokX
3oNVkSHOxrxpA2mP0F0m2zfUFRTgXEqXHfJEqfIb8FQ5wQQAUtFFk5zd7Vq8jDauIgPKG7qObZ0r
VCVaRWfHFXfKVUv/EfePmKchhi1eXvfFAMsX9jTquYboprzveWFDXoeBM59Qol4Jlrw7U9RMFgTk
pPNxoC6TRNBXyEaMkruKsb4+9DCyfQTh2Ni2QrZ9zXQXZ45vWRJLhZ2TdblJ2B73HvxCLhDKy8bT
JZEYfLegLpNaJfUUZJZHwIL9xXR2h+J8iWOc1BCuK6b03a6n/KpPQekbIEgWadiimvmch6st97rA
uHo00F7J64WsivP7+MEwAd/C2nBKg6JPA/t0ubjXiG/NG7HABs+7MS3ww16K8shsoUlY997vyEMG
doS5JdPm2hQ9cOQQWSY4MymPM5jdgwxtyC9/i1Ibywj7N5vJ7USIwRsExTKuxrOAxIOJ7r9ksGPn
L7McqWu/VbXNreik/103yuVG0nJpeoTk/0N77H/sI6izPARkQQAzBo03+sT10aIAN4n0TmWfrmb1
7E631iXeCw87/LN7K7XepaFJhGpJ0YITyVHQKYE0KgJe+ECjWA8Cg9PKaEoqJ9yn+Uf+zFRDoqTo
2gPO3fCbKC+bPovuh+T7eQtt4tSQWc24UKlsiZ3gRxFdsxGSGxd4TXdbMx79aoPVd7mfVEOgfb9Q
UxLHrXd8GCAQ9B6uZh6/E/HI4CM4Ka5NN+OFa2iEdzBD0UDifv4bKK8p13vTWzvuXJLitn0voJAH
uVd8M2QsV/uFBycfoWMwgwuN1A2qqP6hnwkT0Z8/Ri5qopbEjiDWeGFFJYVSwxLRQYWPn9qvCepl
iCGYvVV4CDOYEWe73c5cH3hjn/zXmLSUQlEln7dQl9ObtsnPoSU4mf3A4JqurV8sqiV7gr849hqg
m0D4GduZK7ijx++l4p3zzy8eCYUiG2HT5SPjajV4O3Wna49xvgJf/9gVg/cGnRnc/gn+cbcw0bSc
a/4AC28m/U+xl2nhwnlOU1pPH/h7m4t0Vmq9RybYRpljPm/cRtWHqdHqM9f1425S94UyINb86DNq
pHDp+h7KzmP/xXwLcfNEXQtXxy5ODXBCZzi3+JMtLk8Gft7ybKpeyuO+bup1QaYiVVBBajE/TGCW
SySLHyxN2JKydO1N2nlgZzWF5n2I113oKKsOnDDVybW4CSK9707tPzKvK33Ub4rFz/aoBjnZQaMP
N9klFojHWdOomrkWUO/V4LrZQR3L5mCwdis1AhyGLgeiIoouioqToNXA36ATFaHuhgNo480jKsGh
3CikNbM1E6vkuQy6PQEK6ckE9dxbbhv+tgEWAJi6fxBaaxssWsWXvOGDYtoLgtgZZs4lUFJ0gSij
gkME8yuSqlYq3+kciFigegENzLZ6+84KBuYCBOYHdim9nyGxLFAj2BQ7wCFWXWZN5wB4KioG3hCj
Kg5OhswtT00uYaftqUNFbWFcSmyEHpiJ6gA3N3BbhTG9caLk3qFVva75jCuQY3z+qsZ47g0C9qKG
Q+XMnL8bVnKDX9GSfFv+4hbSAKvd2C31iE4K0MpilGIOliD4OTlqge6SK7WTrvHx2e6hxXK5umbA
eu3ZwBJBIDIsPzmUd41EkD4Ve0ENFnRDzLkuidpMCW9D/XAPC+ZaDS9a0FmJZbSAvm1lbbSM7trj
Eqi27iH/gMx4qnZGSRYtpNA+5Tt/fVSZyjZnXEZUwnQUwSaxXzYQdyDC+zP1Ho5lKx6MHB75cYCk
XB8XeHlBSYgLuinTswUri/2lj5jGcPTrlkXGy9S8P1jQ+9pZn+mnxkzzANvTllXejHU4HdW/uNBM
78FAm1FaGe3gl30b5HbxA9acduDRdlQAQiSfxZPKOc95hWPuzB/UtcD4gNiboDcwWGDEN1ss2pT/
pm2UJbDAiAg4m2WMkDSonNo/9yphgiKC/+6sJRUCb3lUIhgnfV25kPF6vDauRVxhKKZIdL8ZKG0L
ZNmqC82nzkUTlEAk2bU7fjmHURCHjKrv0iGrGlUaAUB/vT4jfDV1JYkcgKUHGvqguP9UikxepXPD
BHXUGUnUIamkUa1Rh4App1PXbyBs1vfWoT3ThawXLofaVRJSI8By7IayiytQ52zyYyrm2r797+yP
lWyh8FtpPydiXFp46QMzBEz1weZlgo95ShINNgymhcqrTKQkCNyh+RlQQyDv7K91zWr1SPtZvHsY
vTnuVpy3s34ugl7fG7jxB2lFQK0BQUkyRki2DKbXxuGeQUtLf74Sm3nNvj+KSN5soZWb8q4q5LUY
0n9DBFbqJ8uLJsNi1YZVKfraQcvPRcqHQzg+4T6wEoxnOulu886cTRfSfOWadF0+1wVICJ/sbAP3
m/2ZK4WQHVyhn7wkn5eR4QcvTvAm4gIi88jtGr5fLyDimX5eiDJNEOyA8KcuHyHfaHlDCRX94pGo
SqNVqAKRyIESjfUbidYGJbViImG3ZZ3gLd+SbEnnUEcH8x3wd4Dq3pavjZi6ZowE3T7xLe+APUhe
yIljANN+2sXt9y9LLkpNhl+Ke0Ofux81GB5T5maO7+l2ezqqHwJfZ0hEoGZ7cbmiYgWJJTA/NxUZ
tS/n8bL8L2NMPSQ2281SFYFrGLcTdK6tjzKithjoLZVU0+zQw2/VcGJ56DaS+u6iM/CPQ9AB7e7D
UUiMmsT3OYef8OMmE4J9OfidBDET3qW1m+BxOozkBonsGq0z7RqrpmbXa75GHf3ncAztQkvYDiW7
QBO4Wffz0CEqqkCLguusZbmC8xn+m6cWht3hPBMtZjwr+xJrL8j945CmUGrT57u0tU9peRiifjAw
DhxsNefEkBXDR/af3T1uCjBsoKMzgf2muG6bQYjY/Tlr8zRjU/WEEz0YMiYmUocoBH/XwYhHM8Rq
y8Zyambf7FaA3QlhMyqW+ZPRHZfRNOWfK53Q0Sp0ssiSoSErjYEaOuJ/N3r7BGimeomfjQCN/MLL
aIGp0lpaEtQuPZ1ygpSPW/UFTY2NzPwtnClwMigFBjC4VQq1V5Z8YrczDlvhm3PElVW7+NXs0ypC
ILdupvRjLmc9ZO8ro551TDm5KiTdGcQ6cdWUbpuexITXQc1jtW+4dieE3vInrDt9V1chzhH0wQHM
7m9iqUIXUauk0NDBvVoLeO0UPY3ab9kP+M8+LhHF2oCb4q5pLyFfH8XRfo+bsgy9gE4BLty/oilP
oVHK11C68X9oJI/6z5lEnRAwss88vYfyxZfC311dae0SjQKxBlVeNWFMvIkLJpLL8muT0te7ANac
T7YyhppxswRXogF7FLM4CgRutC9Adyn+KB4Vd+KfOnzM2HJ4IlSd8rICrSNVs1H34/6VHnT1odXl
sO7xytps8j83Ssw4NT+EKXvOIVBH+9p3jMWakCQG9+jzQvvhVs4ziVAVKCySArbBd27EVvbG1wiF
+cDcYC2EPpx9G2guSMLkHyiOG8dpBeQ//PrfhInCGsw5TRlBE0trB+RDUa6gGhy+W+0LnR3rOwAz
qG1Crm5cgmaAREH9rA3CEAEoxF5ijy1KkMAe3czB8QA4LksXd63/vklq6gymSIzcbyZTI8of/2jW
LNhABSX4MUpcDaqimObV6H4WaHw3PrtdBBfy0CLS9WNOouUCyc1pVruEWQaiJkBGqBPTbuzNiAkZ
DFRaebAGX0Ou9a3Hb3cPX0PDW2cf6cN8lo6E1eioR7oCBHNcg5WCeXdYOuI57gVJdQyqKyWf6uqv
9CvJJ8Dla9wK0q5fdhioFbca1WqTIq5/z4A/l/cipSt4lm7bG5sX04LcpChbWElmHHDQaDPmgddu
O3/7ZsEWH5lp6HVA681uLoQh8zz1xpgy+wzEZcQBrpoZaD5ioQNwlQN9i1ZGoxqu0ffxTFwNOkmW
SNOEDlZPK1wFGNe3yeJL0ka3qIajTESGlQvoxNEL44CPvQAnTpOUz7AnEPsM7tNYqr6GnuMb6iNY
qtgnz7Nq67x49CLP6PBXzP+lN6F0IVBRF4bVSN+bdvCv3borkScDRhOPVhrOVLuHkPeGJ7N45M2f
3moHv75zIxHoStahutA/gcd/nKUGnh89kq6zDrBk6+oS+XeWXu0EXUEtSFA6v8nYiiizaGI+a7Hu
0Jn2iaG3iLVW/v5Lb0ZQagK6DM8UzRlrpeNMnyybE0Utff1BSWXELdRaYcSPJD2jS++cUWMVEcBY
emF74MpuLkyk3ezqfRiuNUBEuoCSn/nAOUDJ620sqhIaJcHusEr7Sc21wQ4cdPfcJyPX8EYoMnYC
1qFAH6bxBjJgYltrpvzoG6A6BvwkLJI7AhENqcnoS/lTHtPAHNNA6gCIGRBLJ2zOfA3k0jaebgcm
kUY8HxaLKo4EBtG2o/mdmE6k5UqxMwUUAXq1f+X6ZbZHy7ajc8HSwLFGb5CYHDTl+MEmDJ7MRDhc
43qJrSmzMsNOQCGqYZn2OgCGfrl5VHXUhspY5jrQuF8NJw6JdioA4L1JrlvycDkvXeJHTMeOYx8x
/N9DKxdni7jW85sR6lK0JjboY91BS3bv9mHG6tex+clg/MsBvvvrwnC6tSQhkJADw2I7HmwNKP11
+fDuAix6qkHG1oBiDWqTpH1OQyVDQp0ytT4YLF0yHrAKZHT1PRJT7/4GOjGlbiK9HrWpoM6GKxZN
WhCkqnT7pJM7k6spXivK9PU5E1N5h8iHDWmiwWLuZPKt2FutEkU7cdef/Tr7OZMCo2lslABD0dFo
aWheJSvPb//IJnOQ/ND/N48tO8fxEDMHmjmt/nix1/lOGX9WQLg8Vto8F2Oe7XOyeS4aNyVRHug4
8jphxfH2ojIia3kGsGBOYjXseMmMi08BI0lIg8KD5Sx/+1SiOFqlbPA4finpRT8drfBHSXbW4G/2
EkqvY+j39+UY03CsqHdvdYY7PI2IojLDqzDMJx8jbm16VsW76wXG+e6jZ1gL/YXcc0XcNfLoDaOx
/q9/IQfG+ozc2oDmjRmWL/ssf/TwD+bR8pQuCTYOw5Rpgu2BUjP6YRRsuTlGh6lwPrW/W8xCikLR
nExKVtZLnQrXbgDhJpV6rdF4hfFgA7XpOnnvvnzIdYC1lT8leUhL/2UA1C7J2o60BJm2ykOpmGsN
Y+/aMS5gs36jetSVNiRwacf3Uwa0XZbbAdYRwNNinQC2wCCv3nX7CjMYuuDSTIy4gtzFZa/PgXEV
iP/cKy+BLv6R2uaVIgsmNUmPQFkp33Mc1NWMWqT8V0b9vE6S+pWazShlsLNmHu5fn+fx2cM9omdz
wSfCAu+AIFypqyw+qrilOXsjFyMesIWnaJvYwkytEZSAxHUfhA20TM4m/lbuCmngLZdKN12BMhVS
beAHgqMQJl1uk8MIk7eJiebzG5czj+jjo+aSzPHiOfbusa4D52mUBRSwx22Bw/ObGieXU1FhAMHG
wDOQHDzLx6wjPTP6Th/12mzmPYl7Fk1T+ouklpyjgFPTuP+3o/gElFibhuC4b/0iv7+eMiL326lw
Y+2xc9LM5ou0Iht0YSkmpNDXLWzefMY5Xzc1pf6ZLPoUkuD4dmxopht9Lbtz+F7R8ZJHzVkqccFG
dTWVZQt/XyUjS5kGqlX6C6GQXDBRKkXC/78IX1sQtdqE82lARbSa+jsnhQjzLQFhrqqTydwkBsn7
5csSedM+qVJ1vpb0F2IB9aPIwzd3GK6swq/AuvP4bFqwynaXUH0lVGGfRNsonE+fOT/I+/HqixZ4
vF/Rk2EEWtOcbubHfFodwMIyIDttQc16PE0Ggdw8IzCzL+oKUStmyzBMDyWnKRpA4yLEgSC/m24z
DCKaMuIORNvTts6ICkkvBd/kp8BtrNZ93lAiqwyHiBA7Xc78gwaCBx9dKM/4UVV/ziZ/sBR+4c3l
IeVO/XIogquLbZUUTCR7vgaHxyO1rcvIFGNROD/Ndri3mUiO+1R4HmhmGYedsv4iahJ9X65OmWU4
3Q2u0q2Rmf2jlP1nj2b091/OhFeZuwMU7ovyIWX+CWXfxvGCgeXzJtEcebJYRm6Ic4Aumws9nMYG
I2WFyH0kvthmyrQp1kHXc0+0np7uu10i18BL8xP/urx1nLhlXj1A5knitJ7xN1C1IE6qFxT6Q9cP
QbgIXsu1BGj0dz0MPbVbJukipBa/Bkz+ejrKFi4Sc4HLQAs1l2M2GMSv4XYCxq8DgMEirCv4UN5h
ICodvDWo+OXmbj/BP3q4e+G5xX73M6Mhy0NyOq5xuZAWGNWhn5svVel/hfnYRDBI6uoYSAKjpzWj
IEhcfjsa3wNm+uha46eZOCg5ld/hQR+Uu4jDRz48ENpuZRZvDRXpp2j5TTtJFzqm6ueRFvZiTLxZ
+CvfSO0SW8UIxzofGP88PKrpyE5U8dO/EM17N322G7mO7XtKckjIsEGkB+eHy6upxygapls8936F
Msieh9Mayf2KhH4c6P6uQvMrVwTZ6b3Gc33f5ygRhGO+UESFKqnEknwMFk6+Ub2sx1OhhEul1Ncq
2gAuvXZ/zUJ3Xk5o6bvw/5D8kTROTFdGN0XWx0xKgRZm6CNyQZm9T2isxe2B9UUb1eBhsON86zzx
oy5e/mUyFYrA+SmJa7qpp4ApPulOnouylme0oEIBr7B+SqRXJJsU7GgjOzpsGv83ilCFpZVLPTtB
sQx/PvemRvLfOqvuzeJ8WO//ko7aY48eR+6JXdNPU03KoYB358JBOY58viLA3V1XqnLlJTTf4UdB
t8bmO2yUOl+8SA/jQtPrNjGGxYVPFyeLEGirHRo6+WYOY42i9xLPH8V7ZyjT78gJ24n8FfZnvh4p
RzxvwO3UM6Cx0/h/IxIkp5WJ4nsv/uxor+Toy1OUTt8MvdYfW7Q7bx1O3/pCGn2W3PYyKu4heP6o
fge1wxpO1MsuKn6yXjxUpOUjOWxp5Sf+Houc3wDs31WWa3gAuyTK7KTsnOfePbYYC0gEDCfB4k4b
18PWnbA7nzy2rTTNV27CskAUwRKVUqE+fuyJS/E+WGzXOj0ZLwGBGnUCUL4O0fxJ+HbqirDUD0/i
E7nVaUNik+R5Qt+GE7ctQ5cCmPXMfgoEHd1qnXhLXBhfY/zBN1ijalNEo1F1jiQSMNW3cMF3rln3
p3oqEIoXs0y4vssVxaIc2OXsXHxLE0dal/3Io4v8TXYWx/pNTjIlcFI4lBJbc3t+6xWBn2k3nWgi
ehRFQZiU02Qvq3O6zAv6YOnIDrV2DiK8bcHXaJoHKs2PSuij9Or9o9NzHUizke1zJ3gGw884NuKG
WHq168dylBxVYvILasrRrutpSpoYFAEveNYf9OvlVGubPtNIljnwdWQ/YK//DEkXedIMQsn9CRX0
cl9YmzFfX1YPLdsePdyW/wzURfl1ZyJVKvx4HvXwoIkHkuCIrdPAKWsWrL/A8AzhdP2Bsy+f9m1S
fhc3RrjzwuPEXNYohH4Aj6vdILBXAlSgWkOi1pRfWKhfvKVgFh6WKRYifMSOsUp/MzXyn2GQNvOD
Iz+D/4ER8G1e4mlyJXSVCmEjYS3HwcH0ZIlLoMebeSEJrl+HgnU6oI/ghLxa1h7yks3Ko1jORLs2
B89fuwZpngBwIKaImNSUeNfWDx0OkPsuSB4o5w6vh6BpWOqySI/OPG50LuYcWIXS/iDTLgu8ov7D
EhtGL/2qCCFENh1+C1xp2c2jwLlLPlb4dt+t4Ga7O73I7SMVOKViKZbupRHKLAKizrr7ZLLabHBp
+Bad+XhvWmKSKF+J2vqw6hGibXConSlwJgx1yeV6l8jUzrzbxqKr4VoNnKu3J79zXCeNZqcqsVY4
cjgztHcJBz94AyXVtcT6zkMoCIygyIAIL9zJhiT4bfygL31RMMjz7EGqnUTRUkaK9Y71Wx90Kw7R
xo5RCoZvLOF2vyw/U7Hsy//scx6VSC6L7EFhjQUtcInid/7jjpiASfmjmP51oJ1rMKvwL29c062A
ubsn8pqbRFxmSlVcDXJm4wo3/GlE+OhLB39IqrxTh/KkW098WEa/TD+NeEvXcgAj+H19smSkC8rl
7GYOs+5GV1I8aAR6rh9iahFNAyHU8Xt3VoPzHSxL+XRBqwANwY/XXQJhQhTNwq69MvRoBAwwytwc
6mWESiTHg+MJ6PwpEcuKuQKy26FBzRvehN4YpwnwCrzZzGPYRyUnjv6GvvF0kjhTiau4j2rizQCp
h+oHxlapuIT9X9r9gzpJW2FGxrPjJLw0AKd8tyFyopQRPWNpZAwKo3/+ImyfAENEFTVU5zRHBWWN
AL8FbAEo0ilK1VKAnKieI+4mGK+4unThhRJIwxNhyGaHGPU4rV+oKqgWl9r4JR2Q5cB4QMmvE1eC
3xpPekHijAxfBse7r/BIEFqWUuNQwtF+YUurs1SGoEbQ3KMw41L0EadiAoUsag91UpiURpIGSvzF
0vJ4/WXcFFiuUcruJrZcKi7uHNjq2iDcJpD4B/4xsoO1ioE0ozdf1+vLqGCW9F4Rghyi7odncA19
fCmVHaTJCMRFNgtyHSBGX6hdu9+sLmPJ1nU9/VrSJKDp4fGlMYoxa8NpkV4Uughmgfj26n0T5cA0
B/UXcdV+QYdULdjPnIJx2FdfwlzPz7m36Oaxop7icQ5fPjytMLmJzMovFQMRsifnNkDU4LF/3kve
FCNIVlK11SPOgm1u9JtLgnzkls3SK0oi97piiVw9zTAPRbL3p6MU9+3Pwi2TYSEndy/eZY2+k4ef
AoqiL+8g/ie4L/G0RG/LiRNsyV4O2fXdimOsOGutbFVL2yANZSfb8LCcMcXf/P+8Tj1d3oH47zlj
Gdnb4T7qjL/hcxU1AUipUO3XDTnvQFOHSyJLQpeFi7x6ZTd+H4x4l9qRsfbuBpDy+Be09pooyjCa
MIi9gU0AWNWvEVaqy7LojHl32D4GZVHdHFDIZaNT4y04eDOtPv1wvNH+hxBh3wGyuOBg3cmUnBvU
ApX6ElUAepDqE+afaXiy88anLG8QPkRb8UZzM+AQpd5mWKh7TSMeM7xOva6X2AJO2juj4kKSLaQl
TTHDoJK5AMaaiSWmBWrYYjC2OaRaYJxiDwiPT7DTmvSXUCHx059i5rQlVoX0TF0Ao6l3kqoDMazK
8vrmv7JqREN9R47K4tM38q35wj5D9jtEw11gUkJ2qkZnkPMWoMI2E6476jAbIehASNIBwwQ0s/RN
JSuQL6zxZbp5QXTdt2h3QewGfoxpRcnEPK073UaAdMFeAniGfAyjq5XIayfcgZX/FMxDn/LT+Nlq
1NvB7CyJbwWDhWtzwOatEJOWk589ESjTCKSFLnMwK2aVpoyK4D9oIl97FpoJ47TBnyw1Wua49IrL
bavM4inhPcx26bU2nUU4ftRTPvU8JFSLYCzNmhOZMUaIXpjd+wNSddVBMKX1Gc8gUCfhCVPbJqAJ
YTkxyJdDwvAB16JubLLhmFjb6+co+1Yb65i8Aq2atzgxlsq0uyR9aysWkDSkl3MOJlTIb6leUSGf
otdysn44Ekq8lUAjs0y4qodMyF0SKIUu6GZ0BwO/FHVAfz0mNGC9iEoonWMP4Z8Du9LzG1BAg8VH
/qpCYMLYR87tpLSztr/75+0ogRAi5DRdfQdKYGcvxE4A263U6qgojpp36ym0CDbH+ncdHbI6pcLu
DhakJ4GEWZqsJdVsqG33d1sQvQV5ar8Dq5AsPvHmf98lR0r64SeqsBbkMSAoHkNh5AB4PJ5INvZQ
8kray/q4wDcp7zIwH/yNpOrMjbbY6hgB3sUUA+CSlIV7uHRD7kwDxRetbfVoH2SGRbjHvpxtkkId
e9P1DTIlWYR4yJIRvOxWVxi1Au+jZJPlUQL2nfuq8AcfAWO9Ad3lzhEyOgF9ltIzuqXwJ5nhvrP0
SGrLyBtaUEIpZAMbAGTwVh47NlOEYRINY4eTy4/svQRnhhjgyh5T3W+c1aauB4ZJbed/9eCu7Jcf
7tkcaM4WPgeD2DrKDbHdbK418lMYiHFzczX50X7NSYbwLt2graGeZj8I835+g6RRNopq6b9LQ2Iq
PWGiN4GQIfosWAp47AYErf545o4AO1yA5hREqYw7upgbH7jqD+LSnnfA5thz2QG3RLJVDve3xY0N
+7/5VMPSU/jv3HYSM2fgrXI2Q11XUGgZ8PG34a+J4uf9j3sP7LotX9to+Wa7iiOVw808EXlSirwz
/cZfu3tL61zcih6q3xHXGrWol0N2bXF+DQmKmAzZEZGw5Q6dHdmN20Dc3IE8sqKBxukw9zL+rnpU
IeyXIfWwOU8T5+Q0rQ8y8fRIm1NKlfP4Sj6cFEdS9Y0C+cB7DWvju1tiTfI0IX7nhEeTgRbSZP63
MfqWtCPzOQGH+Y8gvJTPrKuLV3wCjZQ7ERstun+5NGZSoVdvgLkiL9hCANTcfFedUd+Bnztdaj1Z
UmTtXUOHX45zxj2vPLRbGaTb3CJJC+H3Tr0GnLtrAg+oaITLO+rnNhfJhJsoDTZ2WwS9qRsIEx8F
69AbW1D2W6dwXvQUVwa6HYf4bEzIodGoTCqG5WagfV+pbIPeHiOU3Mv4QTX7JPMrblh8nN5kudXp
hQ5DAV3cpO0y0d3qPEg/PiVxUJ/nMVwGFOtZyMqqLCbBUHnYVznH5vhLNrTHqwj7R5sE22kIesi1
EDu7FJkcQTHBzmLhRDuM8VXda0v/PYgZ15+P3vLfRdy/khsfOvb8ZpYLAUPMbXGH7GyczaTinv1W
/PsunODP6khaQyzU3n4q7rLEAfpVVGaeA6OlMy8oJKAZpcS42iAZLUKoabtQs83dgciRzOY3I3xw
zxy54bXaI/N5xbD187OttlGMFhlGQwuv7PQuGmVT7443ueHC+SH6CRTIXLjDFYA6geG1Nmg7Wfwb
wsLwQd61APmjCAEkpB1KyUIBAx+buisuCJfx5qVg2PgQl66DiYjRJPB+MhzDxyIkF8cNXWExhgrl
y3DDJnc6/05nksLnXbsCwgHqEM09NlwRL39QdYIjRm63BMkk0Evg5gwdtquvwPWcEDX2aFth7fWX
+fD0/5XaDVkj8F1Vm1cUNONA9nFGrWjlydoyLjcInBsoySwKLoR5cVOkswGpZ64nvkSxe2ClcM/b
iUTRRY8KtPna7M8WQfL5Vn1BR3WBxa95cVCDYr94Rg8NQlbj9itO6iwdc1bskFrOfG7rVbqRpkAX
mnSELCYKGOUxF92fUypo3NaUxFWWt7GaJfQ6humU5NR0Qfpabs9JuSKa0BOjkObya37mu7Vx/6Yi
t37U6qdQbNYJ4yrP5FYS3Hb4Piet7nsNHLY94eJsCAyGjWjqfqCGPiisj1b7TWknnDmPgKasdk+M
NrysqpkxX8X6GBvsetAeHQLheXxVppN/QsckE7Tf2aKnR6Ou0GWYHNJtvfVrdf3oZg7/W37V6dx8
j29bWm1Uqsbxfk5ZcKgOUfecYAxufxxZ2qIZI0usTw8CobttX0c9bDqjfnL9OhL6ox3HuJFiAOTK
w2YDgcFvLxnDqLkP9RHirO0xwGgDVjuFjb1oTlPspyGr+Z0EDMSJWpZlUIackz8Wrsyx/WTg9skQ
bGd9l20+JCfUepoCBYdJ6npj0xlb0MMvmx2AWEZw8vAY7hH4SVNucSx/xqvONa23A9cUWiT/kUh+
R0a8GG7iWW8JDZ0sEwCt8IrglK1YxdClfhYHNHWOa8eR72yPz+A4jcQIq4Dc2Lxqt3EiYKDno2Sz
IuGNgnlFdoBLotmyEFzPmFU42hLB8HlsZYUDuVNXBp1LipJr0lnYFWrVoJoLGVrKmnEVBR8Xiben
xv7DWW6R2XPM7gG4wrfCRsGrbkzKuJtYzMdAXjGopVAPBTLy7UrVopqCZThPvdvsngoljw9U4te0
k1Ofl0HUQIbTXZXOrv36fsXQlSefyqhM3BK5f3jnmVqA34OceaJN7UvY6v4cfNM1Z1qeM7L0E3zG
Xj1uPq1AOynIBtdPafUbVxDne9Cc0a+Uv4D0L2wrODvptkFOzF93rqLaOV28scrWMTe9fJrpC1uO
rbATrOCEYu8eC/jDA7GxWMpRysgPLy0WhgJt+WOeFPakfJhS/su7heFNO4Fb3qiGVp0VmfOtp84Q
LJotbqPZOJpfbDi4aLBKk355uYPgMOEafuIkBkha+m2HDLYvJg4io7uV4rMJTF9uIVMq6CriCJxq
/hrI/I00Q98RULlQJE1q2IN1ACH7P8+i9p3TatXF0OPjwCqes5Z4FCucv11wYRl/Nk1Ji3IUV9uI
O9Bsrxn8RgjbTTcv/S5RybVAC1EPIqEgOFucwI1dNnx607ApX+cTd1EKlHARjlpqc5AZQC4kqAJ2
G8WsBuuVsPY3Vu8NX1q5cOQvGnCP6caT9pW34Ciwr2bWgVxODp++/R+sU64fbDwwDycFknMnhAZD
FZmxBudrAJ3kK8igMfSAmtGQpFMRGewcjQcqOUE8At6LzTMIadsKDwe+i/zaLKN8JBv7lhLFeDna
IJ5swSIjlIOQzmbyMvU7FhLwpuMRTmLojycUnOGdXwo9618DEZBwFyIDYiMjbyD0nJJnYIn27Q7b
nFBOUeueJuGVdG/TXgBs8GmvYj0Rfy3NNIbuPrN76fP+6aq+PrP7foxJJhiIp0mv+yfyxjtu05Tf
Kt2TvR+rJPOqkvnCvZ5Yg0cfk9VYAbk4oz5cPqiK/sII0krMq08ktUoE9Pn5Hp+WnQCB2QWnhTiD
WafBdmlkZdi9VPs5Yrr+HsaLGgmwp95wZaLMpy3sBbQ6lhqMCeH1ty/7AmDed3EoWTb0t6ZN3NGf
W/KodhWeWioDIAAOxXUvImMXI5RvTzCitMa1PoyVYSIobmEIH8mXOuaeZr4oDxFAAo/r7EIec5Jr
1gE0BGNYN3kAFDnhmvhVNvvLNI2mJIf5J8e5ZIyA2vWN8Ml7yj8u+6in12tlHAEPTVXGP2MOTsgE
hkT39yWZ7+AuNzPD5a+zwaZfAuXWRjQDGw7TTL/lXi/tc0eEXEKEHdFIWVgT3KyPtp/5eH4pLd+X
eF2icx8RU8j48oyKeti6ZTBd3oHKZZSgka07XTdVJu8dzQuFrWq0wadt/C8Mvl+CgTNAfhXVlv2d
cEnNPtCMcbDesqkpu+kfj1gYRQbMdrmvEllO92hRedCn5lg8DnCERTuscz9IBsrfMvZXWvLFPBrH
9oaJK7FKsOFsg32bygBZiErCR3/moFpPp+AIMlmgEJnVIARt/2lpm+b0o3mxch3FE4xGqk/etzyr
JGuJhIxq1X1iiackljf9AKzzoqgfQEzAY2hB3VVwdOtMlEXgkqgcUMJB7fTFBNpkN3MxOuvzhyGe
xSqOBmF9ZLWdrBZYAu+Bf/MZZjnp/5+US0SvnnqyEAiDSVv1aq04oxvihwrvro4T1ioRQWyMXRRp
G0LCnxt/oIA8aWZa9qu/h+85TpNXtSPnfZe+ja7vSNcSpUAKhWm1BUUOwSUvEoXeQaSUG1Cqz651
FRkJFxnyE+HgRYYbGjEyUTXvRLEdxRHpRfX/fcFJXVSrvs4XmdGRcBE3pv3nPxmc7pdL95MIpjfF
Q2zDQxyUzPSUte+ytHgR4MUHjTgzL4+7R6dvfD94Vec+/vIXmcGV4wke09MhkLqy/KkQ2RyJo8RO
BNYtftdjjCOmv8pkcLMlHpaa9evdo4WGUjScY7AgE7mgJj+sgpVDAb5JRHUwaK5pBh7mr7GYorEi
G04dtwOzf+VB5i0aCGIJzq2q6ddHpgpoY7lsZPU/8dUGZqjln94GMmKvds4RbryhC6r6WvnAbF/w
Q/xJRA8j4OnCrFvzJlS4rgDM21LpQWzqamZZ51AsesR8ZJCTbqTDDU/wRfuXeCdx6WVXGDAMYXFR
Wkstf6hKQwtB38gErlFlneNTAtsBXwCWT28VBGHR0kIcF5FduQLeYCbVVeNY2cVtnBih0TlVtSHb
OCVMdMabVqQaBY+9k60g33WMtdlxC1OdEYZg42K4ZD1bspUJfy3DICZUcEmaEsozKUEeBe4lBnPd
Xnfzb0QzvuRtCc1dwUDaN65ow8nEb9yyTdYbifiXzTVrDRYpWqkoRTrand0wQv1YEfc+Rm1yfhg4
B5WeYXL5WGOh7Er3yLwlYBMh/kIYmHFP6A4GbcOaynZZFc3ASV3gkbUcKx2sMSFn9L1eR5wpWgEn
OcJafYdoOuf/KU9XMdw5YkjMnZmtrLdpaf8junFHCCKesDdt24yjv+K03JkljEzrvvCSQLUK0T/3
eVVu82commk55zUT763/QE4hMpNYxmxQni0dPpnJ4/mRUv+nibueVIYo2mrdCjpqg+dXqFCFp20v
TRJT2ZLX3ZejweGYYQWPBitjrkFD46ZSkUxcxbVpHL9wo23Tr22qnP5AWAbIhsY7tQdIGT9tU+21
jvzOIjo5kQVkl/LOGWMyNz6HbyGxX9q0mq1bLA6FLcoANUQuPT6B7lw1NfBp+z879pLiJ6W3YM2q
AbZxrs4VLHDueIk3kpQnmYziM3zeHsgN2kR+me+6qtuBDohApfWCS4mRceCmIoqjeAeBK1bfinU6
1ZQ5g2PLyIeicpRQURyMkHY/VgCsgbS5t6OGa3xatIjko249OKxjsnNRsd8g3UBMxkbi/9p2wRTn
pEuZowXwT69AhXjOMUvuoKuWYcsV1kEFJBxxCSZPKVLk11MWRGOAe8Gy3GMZBEFAlnweboxV5K/3
VftGEuWMQAu0+hMl1WOPRX61bdJZFV5XTJD+qHuY4Tbnl1JR1nD/We5FlXeyPI5cH7VPgIpuzKBh
bvrcVQmB6DjGX5b58pAJATaUu1VDGulhtflGQlCZ422/NoIqvOVMRVbPwXk+Nmunr7scZp/Rgd5r
olVM0pjwWFR1CuL9dugGgTj0lL/jtXCL1751un34nQOUOUZ69ePfuGoaDNiVZ1TsfWQYv2mdvmWq
2xvIaAOYDgDQBvhcFruHJNDtehs9iY8HkgfKrIqTcXlr+K7gJoLHuxd8jlG1cTJUeNi3soNPRclL
jXRvuQTELa9K4/52gut+sEtz3Yb+pwq7E5qO8Xh8KTooGdEF+kwEFgiI1S6tZpi/a6+mk9A8QOEx
f4tHkPfAS9JABF60wzpW7x2AoS6ks7N5qG8o24xK6T5joRPhymIQbyZ1gpKE5AvEmaa19LPEv1bt
aKK4z5IYhBIzEOgud6mBhb+rQjfHYgGdse3cnzfDYuS8RoP8Y+f+MmYSMWgDTb9J6xQKeyw7MKmb
TSl9LFS5g4O1brgUP/4PNGeZ2ramDlR20ctVlMS/CkewNS5tqH1DHsfJvyPw5AHDYl7FH9JI4KwG
+4wt+TTSOT0R3APiKpkhktM5Svz3lLY+n8X+GWg+FlvDaFWIEYWly8y0j21g+SL8Vaae/Y3NOEct
LWvf4p0C2xnJvTpxumjBBz/H2wwafhmnGhVlUBC2MoPKLGoFZe96jEv2Ug+D+dUBx4hAJxIeiHXH
c+CSlPse015Dn538ECA+DxdjTf/mxFhblxO2Mz6kHKHU56Afej8dMu8NQH7XQUsd7MKmza4XdHa/
AxaAmAv3Zxu6dCXughkwoBC2TYF77eQ3A+Gb3nUz+EnVeFtF3nUSa2h9UdQ5qV5TmQxn3O50rSBt
7kZuxOaVcGEX+dqTHtZ/r7inVO9+iXGZ9aXlHHIlLPDSoqihom+o3kgpZjR0x0pPZEBABZzl7U2i
LH+qPyoZo+T4FMYpNYuLWZD5pHS4OGCwzCHdjt9Yj9KO6YZqRLDYzdG3F8t70hVGwNM6PVxCgFs8
MLu7PdAYCu2HBjNQz76lMGqLMrAgOTAIQ3+PkSSaNeGKEpOO6dnyN7GeIkg4amKBPsBHGud74rGF
/fJPbTV/ZW3jB1iDc6i9iyDpcpeQRq9EkC3fH6Pk0PXvc/7M+zvJ+OsFfVXff8jfFofo6Au/ChDN
gI97qLIXnOrsmmwQ9CZpF1uptVxkvDyszPUo0JRa8W6ZcCqQ/86i48kVlJidRHDkR/qN22VrhAjo
8T19KhA4YmfQASkmH7+dRjwboALUwqkObfIqRUbILPhlIHlhJvDFHs4wpjTqahlD+w3svZTWReWD
ZNYWbJQDY/hB2u6rHaSdxkcoGIO25Do7M52hpdbQHHmCsYLPlV0WihOqY5+2lrpd1dUeOqL+A9kc
hX5OD7O5Xgsog7Ky431Mg48N67WpoXY2kYGwl1uRDyEqxnKpOltlA5qo0ISFiAL9Ob7iz37Ktb5f
iULk8I927BdPu7WWmfAgi5Zq+PECpDEMIezgb3Vdz51LxFuMAfLoQQdm8MrxG3ptnxks5eTSmZwM
8qtp3jOv3Rw6WRtni3SlNmBSvr9EivLAO+1iqZDtfUzrMuIlDpJf5qbrcbc2D5AnNuWqkF40UIZl
VLCIh/BhmRMLDLoZq9qBbBp2wdgT087wrLBx6QXZ/v4L6xSclBwMSkfYL/tAqgNiisQ/AhzELsOY
xLfF0ZO7JzaFHZ0lWpJaKnNxudOxs17yaNidaFJzgQrVBU12qBViJM1auAE9WeLxvqhv1TTh5Ho1
Xv0rgc6WNTf4ocMVLJaYzFDn+sgL4uJhgY4Hsv1LQoPBp4VtJ1NXeAj0ZxIfVb9AGqBmydOvKp4B
hFpM0rWFS9bkkPvn2nMjb7gE8/25LSSGeHROoxX8U3DWFqsg+D5iGHqK1zRFnbKbQ+kdnWdm2reS
XU45Bf1ociuBB5d406tCSoG+zlgkm+zDohGs02fbPuka5P4WtBluJTsaMVRPyLptre75ZQrhEsPw
djVU8xgnkIpvDsENj5l0n8e9WXlgzqllz5OyFuRGRLqcfAPHDnlVPnC64JAc9SOO3HU9yIKwQSMR
LqhPhK+4kku/T6orqyacolBM43zIIxuTaTyAX/SYSEV5YjLkPHMZlEVTlrYSe02zxGjUCqlEnQDK
6ZKKtwN98i/Ua7PZY4j8C9h/Hkade9EkLc5FcGm6MoBE7r68/sG0VkGqXXpr08DLdYT2qUMQse3X
BFeRApFM0+F69WWFytTLlSwrc/1717IritPCp5nxALkudnTMxUk56nAhJv58E/ZZWV4TrW1Qr5wA
KDg+QVuSH7f/1w6iGmrtaXcuavJP1LbfDaFBl4zIdOeLIBXbj2UWaiKtY/+AdKARVzSpycJDUF7c
0Hz6m6uUODO5gtlPFbpDm3y+m4Svf36jImJPgHyf4/StV5GpqU4ZkpOI4uQWchexnN4RSFt1NZ+o
Cnn0EZkErAm3wiDdJlivP/Fyqc2ZlIgAXQkuB4lr/gbPzHULHc8evhRI8xp8FEcQ5KK6pA7hoEib
/BsdZPd+SAQpkdm39m5HUdiLgnmGiscin3H2HTan65hiHvDOoSBtKXmsB4QjggqbGAwyAmPUK8M+
fuWDFRfpovNJWiHlQAfN1uUP96mqw3c9U2V6euxPWI3HDSbu9WC1HmfRKH5ZA7YdQQ9mhDaBX2rg
NZ8859O9PbEdAL8f8adnIt8CLXJiqZGYv7XW4xgNj3sE3t/Xd+7JPoOdfffaeJzHxtlxtJEZsNfH
wFiVJgHrUlhzIYHTJ0d8xdRavMOi38vOUnOcG2mX6tC1warApU9x4Mzbr4DMEwT2DCTVVqPS3wAH
AvSIl8kiRqukZai2mbHg3RkRSTEyBWylSQ2FmEkTO6J6neP/YoPGtdu8K8inxBAZRLDvkwbTIcGG
UIP063OHVHPac7ADxAkzc/Vv9GM60lldw90qmxMjTICiHoMP6eYEPPI15/IUck6enWSvQxHWYpcb
0j3xBlmgJbCxDv78C5y3OHlnnf7sLTCKa69Mh4BAMcmiCQ7iT1nL/xeefOQejK2+FDtaagf3Tinn
uZjVx3+Fm0QZ+l3VKX2PO9Z1W5ejujOdxo9j1poTRcLQRgs1XwaGFdzKD5/x/Uh0CYsayaoOh3bB
mRLSEj5wAcR5z4SJhPZoNHdzdTkEWCbMXkZBBBsnhB87580IiNS3ExufBav6hsd4+4aj3XdIgcMA
gVATIpHoFmm/8qjZ9Dm7lT6pD9CTrYWksxbnTkb4+dr3CFORQ7DxmVIvWK+aXQgIvmBlDbvjeo3N
IQo+etD8k37pWhh07JTU2Px40gPrDk/oFtwpotzXXpfm6FsiwSoe/FRa5yz+Dzb/YW/YrNvCiSva
S7eSD0udFFW+Cu3wwCJxwbkngD7zS8RxMskGMDznOErzI9BZ+0aLRThT3ROIOUl0cb1xfMSbttJa
RrP/w1lmZi8+ZQivwZW39fX6DWqHCT8KfwuyGHpN7Iip8SwyjO1ThWqQKYgH6JDtWviHDutdW10F
dovk+wFzdLrl8yxhBCAEu59FqsLJxlKQ+lHtpLW0gBwdvtUF21+hF04tTCxx7IN3ZtFZF/jMV51l
tvvm08TXArf8J4SG7XTdGK7PUcteEga5KGGz6ibe8LC7CyLAIXLgHEaRAXWIkq++1r+sswLxra2H
2roMgyOFOPLWIeGQoN9IvrC5j1YcJ77T+UbMl4YU5vuyemAAjQk8za39o/hoCtTy3aDGd9aUzUx8
+Bzh43/dtkXMGtk27rgAogwgXy9DZW52YBd6gN/0MVN4FSlzqFPdpnCF+pNV6coKTb4t2fyXeQzD
Rn45Wz1ngV/+HCXZdaEGLRCCdcnIBnXgTiC9cgardtjo/sbyvTEDYZ6I+zK8Ou4cm910+sFQT66g
anvBNuRzwrC7eKVdojvMzVX0hTbXhXo+f4efUjMij1WMUU6AT8NULuL2E8B6C5uhwSo/ExAj9f8j
AKmb1KP6ttQH59NIXicPdOd/BiliHA5zqmb82cIh05+wauVXE5RX5b26DnNhuF7o5my6EKHjetIF
PKcnbi7dezd6Fh5quhOv7YAv8B4ysxdPlj0jRhEEQ65sAxXpfZb3ncvFq6V66Gsj+dywIQH5S5CY
Ly/xyJkMzycweXUm1oocDIATzwELhEC8ywcd/ynSmh+6mfwTtGRjUDOS3GkERo7wcIANotT4WqIr
TR+eIf3/OUGJ4O+awtP2Z5PQu8sO/4/qP+R87B7xNgwg8I92kTyKDvAxZEd9qqzIcsq5UAbGt86R
k07EgGzPT3Mtia3kWHnsiMHSGBfH2T9j6M87fQdB+QV2f8icaJB0qPHwETpQMfvRL6V4MvdMU5n4
vQEkcDW129IXgq4WPyGXI1F2Ljk25mnYoQABUg9+cwEYkOGi5oN/nrG84onA3sbXis4FyW/OWeQq
SQRSALUBOz47/aHQVRT17729kMZLZVURzzQ44hKmrLiRiAR/Bu3sPdE4wGLcKj1GIGyNUJGiHy0k
eOobYy3b0PFstV0zk8XG/gzivzpalqKZXopeED+TPb7wkTrv+rY2mmgtmWOiTvbSL4Dwbkl1Om71
O8QVRH87ILDqX348KW4C1avPaGAdVOogzfQpLIpARBiaBsosgP4EW/bYw0RyASZw73Qp4Bnp88jH
4bcM0Yf7bImbXYUWdyJ8/UzHShmEdyUHkwUUbEV1OwNWG4zeqo4js8gmYxIn7PxnF95kC5T9yPSu
txHCsVPAyMZxurBzIgu64Kw/IuirENB3ns9UFy2GdxIvjRrZrHQmOWblvQkb6VPJC4PuZoNaY7ol
WmBo7TRjR2u76RZ88P9etIWZ5T59JhR2vag6v/eePk599J+hl5HTm7WTiOcypyHni+pGrMgbdFue
8Y5XdaQfdR7TEdN16GLSGWGUMa5/1g+oV8GR3ZvAFwtY1yRzXwKPdZzLSPvlMZnU8V2RE5GlZMwL
d05suXkM1ICZ9VsQHvC+6yaSfBbAPlCjj8E6Yn5H8RSfUeilVuD4Wwlc2MrGXfuAOuWWwSGSqgNJ
a0OY8Y4erotQN9EnuUkbPELMpz/RYpkgzJEhTA0bFPeTmnMQ1C4z9afDYiB/k36s5N9aYYWVrJ3t
lxM6mqVFyGIUHAd6lwIx/kVpLXuP1KiTSD8xUaOXUHlJ5V00aT61h5MOQWwheT8vH1/a3AE8xb7c
zqwVtOLY4FRyduqau+3GTMff0RaeNG+h2ZIzTh1IV04X+AlePRFo8AofsLACvKrMmZLAh4JZnFuj
OM/AFTQn9eoMJylJgS8jyj0VkVogurF8wXOpSaYMoLG9bMhxLNdztWZkFFY6T+GEOtFiy6UKAe+a
SQOemuauwG3SK+1tlsfgxvrAqO1gKb9oxO2cGqAd1Tm25JhtMiNPhPG49r3O2CFdRygWXUlqVG03
z+mPivopp94FnpoSIi8Wp21bNi0QyzBGIRjB8Q3vbEvqxhhX11fFMk1Wds9nsUJ9yShWru/ysZan
1sAAfn4o6DZFdLhKGMVbCP0uYc7p9muy6i0oaGJ1CTdvL7VUIS8PGSeJOAPQ3GjBq0aD3q+BhPZN
vEUazgYXieV7djbma8tDJgyPqfveWfAqB+5vtOAhpJz+O/uuSUz9o63WlGUc24fhKi40LsX68xBG
hGi08hV2E+HiF7kCil7tpw8dMjUjCRHvvPnaPm8HZwcZKqUaID7t5zGtHHJD5WNPjlL3h1RoPvo/
6HVcTxQBqnBNLoy4bxaSj/bBtPzllG4Wwyh79UGvDOAmDLMK7rNkHdXuTKRXSmFnLpxTs8nGzqG9
z5SFl8+zS6Kp6LKWdPA6Hw70cIFqVArixCyYx4EJn0bARQGR4OrLNG+EJEZ18Xzipd7jek3k/bZD
0YH9zQl6DPeR6RW+He7Vc158b8KpedYYjNXUipaT3Wv+h9dc3FA38C+mdykKcqYooGTHqAwTFSVP
W+h/7wMdBNmHI/D9zDoAcpWzP8gzKByzxem/Nxn9ulU7AXRmIlLI4OoJBH1X0EopA1fLs5kUMbIR
Ajh5arC+UUc/u83KY2gY7IEc7dC71vfvuGfPxUz/wGFiUGixW9RfShhfEORjabZ5KrC09jQUq3zH
JzIS4qsKxxYzj9lzm361RhNBfdFqvOu1e905fi1oSiwWi9vdkjEBQy98d+MDsguRdadPKYAgrxKo
QYFKABF1gu4zzTbbMiW1WiBrP2SENvqeTMuZ4Aj1QvczDtdsfmQY5WUXf42oieezP5CbhLi3+MM2
IcuB/Ab3460tgPUucOK0kEaWdXv7KwJ+X5rMa7YtgOYO6VeLNoOG52mx9DQmELcbXBkVNyBp2Uvg
P/OBnPg/jbr9kMHpotd00wt74S+T+ybxJVWqgQSyIV9xUTODHW1qvBHOBumARNoX77IhI9mFAd1V
tiXaCLV8qmTJ9JBXulmoEqDbwcBUcdguCThpUpnre5tZGOImZTCCs6HiN51J0BbygUb8Lx7mrC63
AOP20UK5h+9yY4OfpgM4gArslYc1n7tk+T0mCiUI7KcBpnngTuk1yN522V8bhoBM/Jt4F86UgaFF
ii8CRAaKEJl+/pqzdhUvamEyyxIkRK7bsESCS3TLLsdwBuTRIYgk0VB56OT582+8oMniVcBDLDw6
brVDRyMvLjX1cvkDNNcY0I57JeevO5QsIoocihrDhCBA9+eJU8TpOeHdVBe3VJ6HWIG5cayuP4L5
QF4wb7ukAMun2cb8x1OcKobHfb4co1+8crIFvP7YFCARsgRJq772w44dMTjHWZJJIWaTlsj6dvKf
mXwQJLbiYWvPnD7GVbx3cUAbc7+vl3LLya7kgYrOw9FRtQsx0cr+uM0Tz6KahdxBf9UuTEMBipUW
uG3LUwYzEdmBEboHSwA3Zx/S7ebEM0teZu1VxB4j1fQBGih0m7JcNDFRPvjS1fixNVrgjtXXKCMD
MeL1KYVhcvDk6ZzhFQXp9Cz+s/btcVlbnew5iuUk/s95dcINaLo+d+oH8dH7n2p0DSXtuB8CHltS
bnaj4RbFqSuE0Mrw/p9hcrOko0NFDUwzrwIo/Ww/d40G9YB10TmEWtgRlBCvhOPWx5deNsmLE7vu
VdoE+F6pPfkZH6VeoxQ+j8xGEhpzMX3u3SfvlKlLL/rI1JgsrQb1SKhvFWHefDiYtJJwKBuAZImU
dZdt+tG1Oz40kCdlBc3q0f3Ns9zGY4c1D89X3kMLJo++bXuGZ3wLbrW0Uy4+KCTPyAfupPxbR4Hb
AHtWkrdvcpNsnTUOBZCt3XOYCdRsXJLlHqbJtucja/wKNaIYgrnEnQ4OyuFc08m6+qiIRUR2Pw1b
vaucV/A4ZeoYbAH21VfdAIZ12pT6/0CZPmgD1pghbvi0i+rqNyhC4H9P3Sw83QlSMDz717yG1g15
W+FosupCGS4I1wU1jBDKCDZ2+q1H4mNy2zXTsaEjar4hamBlcOx/MHCxBbbB6glCYk/zahaN5Grj
msFqU9VKZpYgDtDQ3Jg5MDg1JesZnMQy1EZmpAN5Xan5vJDIXkGHlIMZpx+kYGhkY+RBozcjfr9D
KhbD10K9mIoEtnlM4E2JDlTnn/OLBS5cQIkMoOQVMrV6os5SGEnj6rtoP96eC37X8JxPLR3WPEw1
y9fjuL8wEt3dq42cNALKCZqNLUO72zvNRYPw9Dl3Mw8bz48zI3vMW6g0ykTdZcZnn+ZXgFS+zjvZ
tH7n7asKI6DioX2Tzn8ZEZ9EssfXXbio5dKp7fNfSYF5lR+dreI29zQTC1unLJdmLHk1J5XUm3c3
bI6Xlsiaf3nRcxjo4cSzwMIkFx8kR+FoKjSoSx7tVxhrvcX28a2aJw6XK0kAd8+EpbbF5YGciWON
C/2sxwzTV9/Qq1Gp0knYMHgn1SuXLRAPTSP1FOQNLBmjev4KngECsuvTUel/uauJTRSaDgNWg19N
ppG+O6RlXzh8v4t61uydyOMZGTvqNVEvmgdMX0ApFWnwQTpKLA2ZcBF+ri9SEqr4d3c/+uQX2c1P
OuQtFVM+bCgWjPl26Ul7vXeE2BivMrKdE3cdgKzHBoCQlVhF9trMUIkAwh8ow/Sr5wPgKpTEW43u
vPK8aIFGssb761AS1ZhcrjBn0AI+Q3eDJvtxBdjbSFxpfGAc+iT8k1vmC5P0j9GE4TSwM5kJHzlg
Kgc7Rb19ouIIsuQc+boNohN6aJF95GrMkZbSqYYkzHVjIJf7uUgSF8iaJi+4SmLjxZWJwEB3ena4
ODibAf0jjRKEdibsU0CM1eM8IGRiKju5rZe8FJujpApyDUFc8BnkDUNfv6UfRa6UBoNhyxzFJqI/
RGkXsqpZ3njphCOL8m7qO4PuBWBON9mVE4bNE25bHadxXcX3Fw4EPEUsh3iiFyyPl8ZN3uiYhie/
lp63wUSOSmZMamyRAToexySTTcCz6jHNSKDt1BkIlrD5yNWmHiU7xz4utQ8X3Boivo2k+rM7kBiU
X711NZE+nady3VzzReNbO1k7jt/4hgV2B7aJZqBlwX6xR5FtS0UlGy+xl2NzDaEpPuxyJoDolfda
MXDhOqTKgs/mFOnkU3zW9CsDhcNTQVDXy8PgBxFsSAxkBILJGmNb6XeaO+FM8wcOz8nYGkPe7Xh2
HbWhij2OBIkDUJLajeMJCXWSPxQunulYEoUueXCXLDPfSM8AmwOjsizgYYm6I7O/rUSyDuBglMXr
HMh8RFYDqFnJymCpvY5K8y+eLKOXkV9Axy2aP5BAxPJSbDbF/aY+zl8wvkiI0RiBOHktVzXa+isL
5H+F2vfr+OOvJgSnyGfxhqR7DLPEm3OYt0+eIRIJq02ae7/FlPJTQbm++67LuwHChlvQnVvTFrF0
DklxVWE30YZjxK9652vQq79A84gwsDP9KHSne80Pn83RLXkDCSOCSTCb/wiKMoiMApLubpHIq0Rg
sOF65Bt0ZXlGSddSQaL+0W2EFFWxbNGWp13ljjaRnm5je2brt2oG5lW6UhLn+sQUMSxcvoi9fcQ+
TM2H84f84YiP4zbGSlkxad3IzGcSX1ImqaDNK5FaYA+jj9f3LScNGSKaeL1ZeDtOPeLHhomLbtBN
BLyKpa5j6uYkvh9Fh+blCHHTsG6R6/3Iol9LFgcePdWEX5gxU/HpZsXOc2xTy9GiABZmOAmhAP0Q
a2rXoWu26pP9GeBjdx/+xoWN3IWbs3nyu5Dp8ptKH96NQtAiWbSju5zcDXIPWX4o8+kYdUX/cbX1
RmJmtUnIPlnOzYYKC2Esp5SdBi5wavmchnMDVafbVREzxkLFQy5xjS56rsCoXyxjHNlCWMXRfE8q
xF4oc/Wal5M+H+Y9I+uH+YPSPWD5XlAkkKAacYOveNsjTiwyhjGWFoFp7fNPu7tNQjs3C0BP8TTd
gqV7JRT+m5C5ZuHeyLpI8IB6eGO431/97YpufggN1XbY08O4w69c86RYCIRSN7r9LhgDWb0etNIa
SjY3UM8czqjD/x5vwb0mhequUPK7VRu9tzC9qeo+g1S1RmRV+EthLyatOV294O/6x09BJtrrWMG1
4CWxMYu39Jx4LgZnoEnnYr+31TRkne64ArvLtq6MDy1LxbrIGXVqNMN8nBxX0QHgoA1vkT6elO0l
uk9KF9ViUxRSGdyBhG8mcNIrVjM1risJWLJTjTNdZKO4xngewXq2lsN7bKMAuZ/0UrxlgKdBWt1Y
J3WrZha+E6PB+n4T2mi502lbYfNMWXxuIe2gbKAZ34NhCWMqZ517q9vNxlmh7JcKs2Cszi9aT6OA
TOSPzmeFnxjpFX2yjBPi9+/T+uXAAZN+6Cn9hKhHoaJV3Z4jJzzci5kH+nAqf7y3Qpulne9Ra5yK
i7yEeuGHckO5DbvnATgGQv59sR/LHsBW/afIVfIbivp2vxpAnyDjPM+3UTMJFd3aMfbBOEntWDOb
A9mZ2Xi0CM3K3mqYF0T6lPboiBveZrznEfBTMVbj0gcZCrU9le1k6LGDXyzWuMbcogNVpeTUx1+e
V//PFTFxOGzUu+DXTjGlT+p3IDQSyBAwcOjw7+FWev8EcvhlLquYd1ZFAoE7y3PNcgE04Obl2JoD
2JCy227xOs5K3J7VxYzDQ6KmI2aJ9ZYRNr0VlHavSb+oo/j/KIoOnW6yoesBi6YU+SUIxCMXzDRM
VhoKHc0chacJn0oQOeBQow8tazTtFi0uUlqoG5QDnqNJn12qNsBqWPrDzQIBNuFJHWi761FoQCIw
LbuqgaVUqLpU656YnBmNM2IzMotRsBsvCCmbtkRwPwXhrK21f1EZw6zpupMTUlnz1M8SjlbLtf4U
+0uo+sl+n3SUPaQzWAZx1DmzC32FhU9LE0fgvV2/jqMUFfTgJFK+rsocEl586LEHCk/ywQmR3Nnz
+yS8y5SHzHjyeM2sjUugxotFGpS+mJ0WOX6HEjVLspaWfggiLVI7bvNP9YLa8wY1lvEAmFlay2V4
qK0iBmOLMnU66rcFVmNQdTvbofgoDlwD7AO2zQdS23JTD8p6lfV7upMbDO6+ILeI2+rCTR2DIcVX
/4Tc4rTjDyBIqsWKaTus3iaQcQSaDwF57JUr2bProeq1LY8fJlmSBHqu3Il3RmPcfy/JFKCUz44f
/wlJIm9aX/BwyJW3IxYW/C3LOOmsvE+D26DwHq+OAUGv1RN9qt66fbOkDQzYsdtJq10bSF7N8twD
RlPs7NX/upHlbUhjk49u4sj0m2dVURk5gipc5E/hl4Qm+jBudsGx9lVTXPllthdC0gbHKdCiinC0
pGybnM/qBqRRyX8xemX8mVuJ1jyichDbIy4AXerBDTjLJbNduD/AWiLiJbmoVpbr0igCrzocA58v
n/f3wGUlQEIqRbL14rjMR8HCCbkfE3wVU8qlaL2f45C9MXDgBKJee94J5KOhzeE9VwJL++EthcL2
jkb/GeOAOOXYUP+aGSroRmFpkQa+5oStiq1pyi9jCUYlTLbD5IlScNjN6P0OUUkgJp6uysQ7S7AY
AjsMKkO3vOtSjzpaVEUTfi0jbdKxAwC+NKPv/AZwJmSDRfxPJlvchGPq3Kx/RiOs4Oq9TSRd70Ax
XrI5Gh5hyK3xcquBD+gfEZmThpIpX8TYT2xlFQfmooaAM/P9sMAbg2C7XgyNbUWoYgmxY4NpNG/u
vlzZ2BO7eMY6RKXmTQCWqbgghgL1KpYpCDniA7899EM3hRWE/XRK1lyVcz6UYARXHHMLuaRHQiOS
aRGlJPbDnA11KpjBhF3x94y1Gha9INWPTUS0fpIFlewSDzh9I2q5Ae7f21qlR/DtAjum73hGo4I6
w3cyl9zNnq9qraDRh4Nm4WJVghHGgnW66+1mPb1/mgcuCL0MMFw0NAXlZVGjvl8lfUP0wQAcagHV
I2uF0lV6WNjMe/+MOG2TRM2Rl0uHqreQXkkK+Y771fmSGNYNOX/SjbfaJyJ30or7zIsEl7LhTPaz
+VkXAMG+wjd/tTOErEn6f5EQaJdUcrD7p/WP3BVSSW37tz+Zd2bfgbKOOZu0RFK18wTTwK3kTIbd
92H8n59/CCaisdba/pSUhYFMjWdJ6hv+EvJ2viebxRmbUnTaHO42RWAnm9tBfcnGWfBvxRYDeS97
6bXIBFW7PCivd8MA5RV/0flis49EiMoBLiKEpXiOKEDsCi+ktEGph27wp353AaLJi3ywnwHXu0kO
trMxdLGu9+nT460qZdEPDuUebWhdS7bsgLKJKzm/GATn5tBtbItW/3ux3w6uzQY8zgW7oJILG45m
8W0mVHaPwctCccBP0GF0OUQVQSFBONZRkpeoYfPFBwe4upe7Wu1gxr7XwPT7p9QHQGpGY0/VyS3v
MJ/Q/PCSRleaGdN/TTvXsMZ/jT+yukYvP+NvHeuNIvTjVrkolzk4C4AdxQjU5rD44AFMMwqJh6nm
+LzgdhfbNkXIWZglGEwcmb9yr6Meg4mYC4oj2bEbScd/H3qw+6EXXC8npXJe4fsOPpsNq22ngjw1
aeD2LQEbvJ8fWza6vdQxugl2ldxNS2W2dTrNZ1ejOByvRmeR217YF6zE8nYMoqce6X7iHveAZ9kN
TYk0D/+wVx7h26bOOwOfINSnEcdNEQNxmHpzt8ndCaXqkP18HHUf9vRBsp4cR/kPI/s9H/Gbxa1+
XLV0ntEQFey3YsSbJFcC1afCcar+jZBAc8rufWZKajuN8XmsPD6kXVupDYt3joYqjnq4j4+FbRH2
5f87+ndaicwe7vOtY+YSYczLA1bKnOCmLymOMfMhk/oK7VMIC2GRR02oF9ee2ikTe4zCkq6Zm5Pu
n50bkpibOJZ067PyzMI5+IpGcHlbueWrQXdHnrpxqolPC4NZ3mxoIYBr+yheihpjfNKjcxP8OecQ
g43TznGvZMNRmuAVJGGXgHMYPm+cF+Yib6JmWh8vnBHPCPS9jTpLsBOadaywY2iuGD0BDYMKdGWP
PeCV4cseWMXuukLvl4zbzy507LSDgLSy7h3NPpVLzWo9T2lgaIVpXmQkSsFjhAzMZ/4LdCdZ1a0A
0uLGClBMzSbgSbo2eYoyzDPfYKyJSFMDWMfZ5aIzZ9xhlSe0Be7nFGux+FL0DjJl2Rdn3AX5uxSX
pUPwUUolrJqyMuukrerIl9p2rZ8OJNFixmUUKrrhEwZL92MDABgodbmMumIZGDKzq1J1BaN0cCDR
96dGNHfpUqhiNMb0xe2V3+1tZRnbNxC4Zy7RKCi+EYHkJ8zUKRZkx/M+BFHbqlc0NwJ1ZxCar2Su
2RwYNN+lf8MOZ9VfTyub2UlSNtukQZreptiIxZGOXoSnHzsDheibcwJbPudbEdIf1gRgcngc2eoh
pZTkJpYKY+AgNIyyU1cGWFN98Pd+U2vLDuO3VlFqdOvHw9+O/X7unx6X5yZ9jODeVOlQzcvzL3kE
GatqSu6+/Ms17hVDsJbA831OJyRG1eo+pztGdMv2Iawr37rOui04zUsGWO1im5zRplZnxk1EyD9W
ahkNZKJHJ8TsXTbnqAXi9dQnvoVVAtxEs8b/9t6W5RQyng7uVrIDZaQFHN71m33M5BvM6KBS323Z
aX6uK+KIy2GJw8ds0kfk+oVypc/xsG6n2c06LHNk9DCfOy5xq69+82TDjn5639Km8uLF2qEu568p
FHUF8kKPgC5BcNuPULYe1V6UU42Ls6AMnosx6y4nNydKNDXt9zo+sR3exWVPIsGADRZuHufLqmDi
k5JbHzADs0pULRpEH0ibo+jG8rfCknLWi54dNMYb77gTrsC+ZVPIkMHU534ALY9ws2vK0HpXexc0
zbRqFFb9fK1011pdSI/PTueIFFYLLww5vIQfXU/kn+ZXD/OIKlq3BW6MuIWr7+WcxRil0x+/VANe
m3tggK64iH5TfrZwNnpt3uk4FlTZMdt5bHX7wEuEpKKz6oXDpv6V/sJ5OngMjCrqbbKtf/zvtBQ3
aIcKa/5hL3jKtTXKwkr/gJp7qNSglQ+CPZ6E/SzXQSTcy/p6cg7Z/FemSy5H7vz6mfgGWA+ON6lV
PLQru3qAWTLM4qyeKQ/kq72vwl2dF5S+j4Jn9ig8zC5Vy8spJuFoadoqFhhu697OjJuGyefEQha0
o20soRf+FBVndomGBNcuDJEM981xkTjLQ4WYZHoDjIRgfKfcaIXUtj1LRhrmLISQbEJUiNzVikJy
hJmnFzo+fnaI4dnIF8TLdGLfFMsI0eVVai4WPMlNnYWDGJw5K1n+vl++5L2zQxp0JGm6q5ah5O2m
tzEpJcb0jQegbshNFwf+4bMaxDjVm4wVNVHwtYG6Dp0JNAfoTRUEPICZV7TOMHHXFau+JwR1zp0N
tRQt43JBrQsRXnVox2VkxE286Tdeq+e6tNqRVRk2oRiwhqZ6BSKVQYNXDmRkQnM0+d00Oq9aSghM
dTbPEUKWo7if8plYaZGq95kJRrYrtiVAlpiejBUEReepND1n4Wrx7MACteXxziOylMJWk3YG6BgC
ludgr8UC8g4tD7ibwxq889Qv51zBMoGJazXlatMOh9HIkK6q9y/STNnxqpRK/afaycBsfCnjtwFl
Cp+Wx9HLW7K14W1llqcmcPCSRNjxVXIB+hCwY4YkUfLdwWe4Vsk++iH1Qy5h4fyLEB4YHrO9Itss
d1AcvL5W647lsux4CSKSXZ8Ua3Wk6TAbEUGAcqaSgTWZ+8GH1DtHRjeT2DmEuTrKqeROe4Sdrpco
i2OJWlK8votZ/JbpqXHb07xNqtEVeCffFEYnwHm2cGsiR4lHbyBb/iTCfpW0DqpEDNChWzOncaX6
Qn8uQ1gsuIZ+KPGWLH7EnZZuVTcZVRv40n41fB/h+QbngWHcpwRUVX8qIEr/YjH6+HuricwseCwW
DNywZF+3RTqFX6lqNOgqu2+MDO7TFZAQaFLufTYTi7YhWl5ndKj9dJA6uAaPC4lVCCzjIrTrw+JI
TeZtpnwCbquMt08vm5Zh/sIY9x19BdGcGX2cWX6IyINbJbnJ5XSHupCSAc8z1Fekkkb2A0gz9cAx
HCxqnIzqCNl071U+fV6DuwQDJY/6//DyaY12dgnXqsTSPdWTj7AbnRe4vXZYq65NTP98+NmRw1lP
bfrqfUGox1a7W3NJ3QP7+9zah0szL5O65YCf96505fyTjVFMMaSzqlujbNN/ysOtBzGEX/gphIA5
ho9Y44i4s47uGcpY3SppLd2hQtu2FlKKem0NGxbq8y3hcxzwzWLu+4P5gDp63ZX1TXuILvqVb/oA
nOKlAZPrwvs/Ul/870/Tl0DUR/30QKp1KthzPBQkdhxoltQFkZucXiUuumNDG4Iyv5lbq6osOAPr
RFPuPi9hE+RTI+KCMH6o5NLVTfJTHrHy5LRxoS8dXS2JIZ3VVJ4ovdt7cy9lcIm+ng3qWKi0NW81
n3O2HKJt11am0F264twASc6tpXLjbgUzRdTX58n1bZa1Y46IMhOakZDbrR2RtFRvscCpYXxKejDC
n07WMJsssZKQFpG+ONwCzlSsPsTDzTh6NBx237i67+aING18u+VN2rU+oP3JIV61pyB568H2M6mO
x3P9XT3dO+TtBrCUkxHa7xvZsdHyMlhsHZCLvUluzj3ycebyEAQUEnrfIE5uh3s6MjsxxYCPFwuo
tMo79KPJS75cfvStjUfNIUSqipqtbV/JDVohVNoNFEpTyRFt4o0eFoeF3V9iI+JVQP/QLGCbS725
4qbiAjy7TsElG2SmKZhsz3HI39OoVGayz07BbsKeuqT2+cy20KPcIxRb/w4/AnuBW6OPiIEIlEzz
VUIDF0LbraV0IMjfndP/xaQmeHoJW0t4pOSIj2sw02pNXYHcd+q0iteU1iO0UBXJA6AM4RuvUkQQ
J0CYhs4w7d/Lfo9UzdOJ/1/Z278Azc4g8AjciVmlgpw7Hc7j/Yzz6dSdRcqqRaEz/ciE0WlDwBce
k0KqyETAelyNNZA3bi3iuliYlHCkPIhIWbbrV8AkdtD+8HCseOCka7ZTgoUSMBIwYcU4JVcvlCXx
9uCTAarkEv1RiDZse2FKZBWwEBz3hG+uyPmm9EFHkYkZ6pFWXbxVwl60HDfuNVeNBndtvyZpGWmH
GlASokScrez23H+qhyRvCMB5dkF9vhFk1uhwbYuezhUgTzJAOdM24z4CVQKHyGD7uddymKcXRSp0
yjvczADxHJaQ8Yh5BNdS6Akuw4jLlk1eeqGwmzZZmA4g0aC2dklZmBSBl8AKohl7Tw7L44XYlEKJ
ZPmqxBImlSP/fRpGIHyvFDIjUpENM6lnmqTGBP061O/QbaJ7UvPanI2FASHxyU5eTynYdlDctEPb
IXFdwQX+4duWHqCQM669NSTtGPJNSJMVMxxljt2GWHXOp5MxULhxv5Pb+y3A9vmT7M8ktLTo0wl2
3Pj+wK6yGILDkIWksnLQwANyPGnKG/Pknc3r6r7rjmodK0CUPQ0jK4j+GVvf2xSrpZEif78bdoIG
4ircI4/Y/n5LOPUzuTreju7tUYI7YP3ivi6331Yc6dBLw9eurynEKFd9g3pN08182ZFgIntYD1aJ
k8fJW+fvRe3zN5Sbs6zf2+qIuvbGCaLgYNjhXj7yhseqbrJbGtdw5CtfaV8f/3J8gMEBpQ5g2A5s
bXEXgMQST1bMvJP2F698Zy4IzxOrLSenWl1JiL7ns2Yyicz4OZkYOqNW6MH7ERq24gLQ2gK9jjZg
P1TgSrHcZxCtbuP63Ypiny5jjRMTG8aLvWa8SrwghjllmEAqQ13jXyQ5x9KuQgLP8R/Ny4d4d06m
qPji/XwHbHu2aAWKgbhufXrDIqTL0T16NjpKU1gd6h4CY/1qy9sUl44FmclutK03KzFcWkUPBE4k
eDg89MSRHf/1zy16y65q8lUOh+6xjiOZ+4pRSn3FQImGKGp5BNNPpqg8+QjxbDLPjFosPOvJlK2K
UuJCrArC/dDeIPdKN7bGR5ogYeHaTWR34uwjkbKpS0jLCb8xsxya7aYnFuvQXXk41V6AmH0L4UeF
Y9QU/yJAdCVUM8FvPl/3YpvH7RSbCEOxqOcqren7MAhPhzgfiJYnyWm5feXTQevXCbG0oohl26/a
mNqCnEzNTPC+k2zaJqD0wFIoHANRwZuNlFTjw2mRVpeMbZIP97pxC4U9mgRHGwc/ZLluKxz+HCyp
gH5UHE0C7Yce0W7B1/Tx7w7ACPkt4Ot9dgC9Rak4QcRPBuzN9bxRk+5jsA6VoWV9IztF5Um5sFL/
0yUwHMDzGJNXuIQJAheAcB1vd+nKoNN55UjgeMwKDYVR5+HioT/krOw5jAPRJA5G2xr//ENHECKL
T9Wzc/iK859ZVpb+Ful1DWe+tOoURJZ/Bibn7cB27T7m+WS7dQZ2GF1SbIUJfc7Fv1nHCmdsJGH7
rju7TOefP/OSDjoiNkdk71Ru4g2vEiVMVSFI5Y5osudwuY8qo4fbSuMkgQRcasr1aWO1iZGal4Ib
1IJmjL1OGpA49qCfyDZ/VFEb5GLdJYIKVz0ACufL/tybNvZ5aFt4vP6RZ40equJYo1r7MtFRKx+Z
priQXxT2d/r3PzGIUapQqtmA2fQlEKwm8TPBNZTn5KXu6YvZFXkUufSz+P8yGBrO7IebAU2X23uJ
XNQxXJ6BU4r9QQox5TvA0qB38riI9UkHu/ktdB5cOf5L2usU6XWnICrVDsZY5v8WW8g+reZGHnWW
pVx7y9vOMkoM7w+yiUVYhB9EAuo6MXvEgHxdnY5WzxrW+NZAb6xrt3AmRzVQ6h493aSicUmSzzq3
yDjyobt41aZRk7lg7tZqUOWSwi6ZhRYOjeZzJSroIuVN/0QQKJQOmJVzvtaF/v/C8nDcJsSQSGMD
Xz2He2zPtKwgRY+FZBIlOP4FvN8/QvSH9brImged+HJY63x2LGNtIRz/+2XS+0w5KqikcXASsksZ
Z6/nEu9F6/Dsd3Xca5r5S4Lz8wSSbChpoYDZ6/K6bC3uWpEScj2nyn/zHgZrv31McRV3+MyRxbYK
B7KmrK292vKp/54V1pfGRnuLe1eVjalf62dwOguQHMd6PO6BMpwl/ENT/fqn6QlDaGEcfKG1cVKn
H4MsSHcBVTzoRyOS4y6ysEWOgO3njayZFcKtAwYBxwxyDsrBLkzjKeBscQXEAv2SjmNTJKZ1fV4f
wLR5imc8cuk3KwlCNwZgXVIafsqPnrmiyjsVLwIp4la/0mZcDtLmxjiAXRy4hjzUYqhfaeGjdsI1
iuDNDBAoE5MzWA6Q6GvTY3RrddBs8Tf4ZaY/6D7M9qRZIonHzPnau50DWVm1w8uVRnf2Qh+js91g
GHcuSKdF0bu1XjHRD1R/bV7eOGnstdNlNTMjDyWjP3d+aqNtWPhTTHcsGnrSJdloFoJTG3+uFg37
0btrX1anMLxl5OoFP4iiKorxg3icCupWtey9SbJMbFGIzSMoBDAdm3rcrGlsYS3JnNyxRoYqgweo
2Sqm4z9rkYKF3rhYt5+9vdkAF1UtApYzAlwX9b1KLWAVL6EFVBNxcIRx/jBb/YCyyglONCQA4IQQ
sSdsnoe0bjbyHZgJj8AsfCOQT2Qw2chvbfZ+f0tJfCuK8irgsy9n9sFM5VeQqFFbSsg+ZjUbYpNy
7EZ2htSQByARiY9NgseXOtinFavgKQarov2QSGm+zK0GcGug6X8+4aBTd31TaS4Ji4SbCetHFfoh
8d83XnpgUZ9OztSUhDthP6gQmPph1bOURY0kD+zekmK1SRYjWU0k2tR6IOsMVvRgCPhaXDjU9Y0i
PJ7fF5WU6OpoNP47+9jEihmfK3jYYdmfP2jK9QgyPAK+wD/FNkqrqbSg+P6BejdCOd+MxL73acRP
gtspKVvvjlD7Hkb5gyaY/zOLL4hEHHUYP3+8lOMgk1T4EjnzRmUKD//LBN8UjJQu415oOiiLM5kQ
tm3YKSfd1dZYlDgo7Er9+t8H0e+2dMApwzI7jxoNgVpLK/bv/vPpkZ/PSZS2949T/nGyw/bc8B8C
optrTuZ67LMWFp7UJdc1t+uBRaEjzfwY6RKM5KiTaQ50dGfvGkO+8JxjjuecLG4ieXRSfVqoefI+
Q+a0j1TGJEXifQCAd2DZhunB+MXKeUMRtiIm6ZCdGX4RKd6HoTWlGlOiPKTDm9Xz3jHF935PtwuM
sOXIwlhwgwqCWBzWLoEkJSSpCFgqI+aMsoK+2ecNToTd9haUKYPKJK/GzzvXDvOUvFUbyPYoxCCs
eg6RRpdIK4O9WPRRiHAob90Aw/gZNonU0Ute9mtSHTOtbG5rWTwKqs/6UXZwAIDxdiZhP2ScHgwL
abQlHYnUXZg9PdaGqIE/A+4xck6rOiocxtP5k8Gq82Df08/yuKpYNc1uYad7V1ubFz1yWa1IVh8O
WlE/07Kybe3xikGTN6MvXd2ABC65mJk2o4npoli2Kg7TjOdQDA4aujLAy5GdcBjOEpqahHwvFeuV
dyZQLwQj1sdrbpJ1RAyxPdx3Q+h1y9KZWZpx9RWbxqTIiTSiShvhJTPwffWhe1cZ5A8+a4O2QWfF
yvu8Xr+acCaCOU7+2GL4iBl8Ucp7qsylCfLCFny1Ka06e57YOafrBRyK7YX2MV+aPqT4osTivAE6
206B4G1T/gUvh1xlePsFHxabwTGRu8wMle8t7aWjM6crlZqMEu/59ydjYJn3SCoQMSFO1a3IU/62
hjETo1vj2Y4OF5LrFCsLgdbZt+HfDKCgvESx2vC85bx7REoBvuoBhM2YsJQTq+XuFXRGUCvzB9Nr
9yPRdXBbYAhQUdFRmLfr840ClW56UdVF45yy5H7B7H41vhcQGqUyEqQN6l00w1WOgmg7r8sdIMTN
xEu+FpP5TU4b6eb+Z8zvK1AoaxnGM7u9N+6D/nDBg8Dz3sPA73HCqcdF03drruJmP3/jOVGxrFBB
wV773LipZpdQ5YqfqkI6Gp2LbocSnK0cdFjs3iI/9m23OwQ2UrwHX0W2vxaF9qlav+IM7bZdzq9S
/opBx6Yo8QSrMvbSW7UUgEkNMDhryEtNFJsGhCVmfuHLfkuq4SCgpBS39S2qjF9FGicRND/wZd3K
JxMzP796wMz9DccIHlndKg7a6Lry/6sepbmZITe8OVYxiJPvZOisGPPPhWS0mHmyPX7cRzP8JVBd
yYGlA9VT41+c2AZ/FSy3nOuhAHli/5OuvnGRXMuUKPEikyGxiKsbnTM1l+nSuUEFGcQkZaFu5fMy
PLDLgxyN/AW02v5Gb2ONMLuk1AjFxGv+p+eG/d5e4/AWubLRjBpka2Me1WLxJPbf78Z4MXkrAQDx
pmMdTSD+P8+pKnRRXJuvzy9Wz53nnrfudGAPpE72hdvIUQZyWOr8sqd/z2Ga9BkUlmb61GYSXAAq
I5RxlRlWbd/COyD4amhoMf5Ifas5kkSBnXiELjmuRxcuja0RFN8ymvIlFFYC32TnwIs7BFh5nDmp
Mt/znyQEJ/w/JHP0tZkrK14evWyT5MoRedfPWrrF+vHvqmBbVEMu0M/kVCVMBDEP8GZ7PEDl1S3Y
8vnzWaDtdbZP+JiLTLd6ix8eSigfBe7u3ZJDnbfnb6RjDczeL9IuZLM71yMaj46PCthHyFtowlUw
7fFcn5es7FPIoX2LZQlb8XP4Hoe1Hnj5j4rUgShgexGbcu76LRoWtBij4iz/42tUfUOasbtC8DMq
Cj9MEGyD4NC1RPqhTlVOgh9VFM8kuZfxNIe+6VLa718YXj/ayp0KeB2CLsYkz+bbNBSkPNv24bWQ
AWOZTE5Lg0CoLWexwGuIXUGD0pcRqzcRLlEHK/Vx89WxPsHubCNEehqf7qNKjfWSTUzg8T+dcjzh
tjZXWYzB/aKE7YrL0H17ODo0nGQwOvpO7BeiHJFrHKyM9kCnydX5j7icAQqoeLZD+GhUIUScom8U
w7HHtdLBRkDLWawyUTG59feR6VMAkfclT7dDCB+ITybLa+laOOw4cVhWgZUtMvmgHh+ZvzFMhTQ2
Oymh7rM6tsZfZYW4TwP+q0wc2PtX8NkBVNmZ0LoUuHrDADhlGY/Veb3XQBWMvagFG5YDt3uIX28g
TEeMJrL6KqR49LferHenensg8sd08G5jldomH4QIuYiHX4wE1TOtxSuNpZEGM/nv3ArJ2dUlW/qi
XtSjK/6MAfe6NxxeghMNsmn8bcLJNn4efBzrJ4+zigKx1CyUSfj3F0vPav+vhiuluaI0SsCd+XsB
MpXDqXKQ31G8LY8aXtTfgME5HIhFO2RXKMKPPxfR3my8GnFuDkt08/QdFq7xzZHwCrcbi4U5LcKl
4d+fPvllgsbX/H1iFwZlT9NAZrkbwO2/rIOTB50ono7kqEOWytsymolpn7XOMTuNWUicGLYChSgP
4jthFbIGb0nyC+xIvC5U7Oe8l2AqZ7471gwiAVvnCEzA+TXHfP8hQ1QcnOXEjno3qp4a5HXcmaN0
bUHopGHu5mgWHMK2aMwYhMpA4f8P+TOy2AO+3HM0ShWXBS+0ahv4QAJb56SNQkBVwqflGBclhzw0
6odOfrBKy4MXBQVJFWGgdK7+b6WOf41XK6sh1knt1F9cP+ycD+yagvTs2RnvXrR3y9BdlwUpcaH/
9bAGPBsXaMddmPbz+k9cOlollX6Ch0rx9Fde2sUmO8XI/EWEEameiaNW/QU9IYvJljIU57jG5swO
coJnxarqgY11QXNCgdCI39assOUPyQVLQGCof/QWuZAdxNMWXB20z6+5HmppRflhD5EJSVvWFC6s
dV9D28BgKubrRJpe/axkMIEA4GWWia7QVKX7hszBg7Z6xVgpyOy0NqF0+SBuqcz+BYCmIFHH9PzP
J/PcOi1AUxozrmWKVhzl5nCDPQzJdAFJJBkdJiunG8ADP+H1+1zoCJ4VlEMQiNDo9SKiwh46D12a
XnkzJ5M8yw4icxKR+dZ2u2eKYCci1eYhw4rxSvK7WCXX5kBt64UpdzSJ0SGC8sSxKyXZUOQmtxV6
E/6i8RbG8pDAl9jPi8pE2pGg7oKUyoX7ferSkXWPNZwYTPoRrXDHgHymgvvcUoU7AWtYqUHQIgmE
Gxr7SsPvR93ncAUom/VFoAsypY6F/FVYGzN/CwbC2D/m2Tk1UaFpM3ldhRV+EJjWW1+B6Vh+Kx0m
WmodpOwQ2PNQ/DPwUpsQ3kSh6EvVI/CJg69nMxIq/asaqQY0ieTSmDSLZKS2ErEHalryinc4Ekg7
t6JyoU0mSAdeMaTrDhTZYTucmqaOXQ5Br4v/4y4bisrqPFGgdDpNjfHgSq/SfNr1RVWP5Jn9VXsB
I/z/X0RA+L6tZqfiNTgIT0HtPTXmoxkRyxofv4rOIIaRtZJ8gItLQtvqQXIUzk+clsur3yBVdBDP
1AtW1AdgnxDzmwcho9xXlsDidE3n1wb+azLKotr6oq9sLgXf4Ggw33LuLIxxirsoqPglc4yDrDA3
Zsn0UKyh0an1ZG7BAvgztGshLbjFpmFwirxGN040vcrot+aocN/wkMKgQ+DTAgSIs6HaE8CT/3JK
lp+DVbd1cghLMbd+SyIWlZ5yuMH6+isW1J1XqLF/uscznXCUK2/sSmEcbcWdL7XkVKipr7ERK7OD
Dd+O63TsGQNhmXHgs/oRTYMgn3krNzwcQ1cUu0kQNX9Y4W/0Fd46DzZO7rkPRftIN/D9jEYD+z9e
MFp4Jz58U1hVacf+SJaacnBJ5jvWZTu/5SASrBjcgJlmIxkIarRST8BH/KQJ26i7W90MnuQTASAO
AQ1IYVdIRlGpOK9XkXzvM+XHl/ycjVY/E9kVPjTH/F+6mxne1I7C5jJWNZ60SMy6ubqqfMgbk475
Yd6jmPcS755G9FAK/9BWeOeTaHOqztx7KIzwJ5b1pCNSf6JmPAcJv9Z1WbD0vB7mLOTCejU8od2R
TPsATpP+mEsye4jhOAaXIPh3JVUQBmrFDWKGF2Eaj/vFbMZjH/AI5agDdh8bDmyPwYaBN/xFG8yB
f7PoLGDyEYpQB+XMT8kBFOZaokPMb6nBNOtF5mUqJTNhtvcIvUzXdo5+BiO/fiSYJqdtPD42NlAw
BrYHSavp8OQRsxScujyZiHVCpaF2Q9IwCBBBsVzM/oh1PNSAGY15E1UAIxSlva6EcOHTmhsh0TPd
X3QyRYJV5+pRoG+jw6bcc15pa5j9OJXfaGkeyDorJRnCKKsZOM7p/+0MoobqYyLi4nMp/PHG8i/4
y+K+JXRoUY8oH9LYpmckfiS+SurjLcRiOMxVqMqbxcPmxtgglnXsVAjXZVGxRXFtdEDr/WtlYO20
pKk3nTGYVdak2/psCjwtoTHYWqNmYHAJKQjMBTv1jsMJO7odrbO126Ew2ksSzwUqKDSLEyHn9JR9
6gqBRau0umz1cOP1A061HZvROnFYzkn8sTLigriaqxjEMLcDwRX6NMBVUhHR1V63CPaRW2lQDIJR
8l+pEaiBYennZPRBc+/8pT4mNSbviSg7Yu7hVmSS2QeJhfatPyNaBCNVR0TUPs8+MFvPEN93GdVr
sZihLcSQZC8qWxRE2H5QofROo7G7Tp6IgRtqduOiofhw5rsL3xNz6SUgiV15qqkvjf/NRHP7dLpO
pJ9QFh19rkJaW/rAkHOz+SSfyMkaz8n33qSNe57qAGdqZBAapWu/d0h1R5EZ5GXWFADqg2QXvu3W
ITGbH4qrhhfjDCpL0WiX8Juw6YHz2MWpZBovEug9ThdyRzmfiloMX2zxaO14f2dhb8hakjWkquzr
kpmtBXvd6PiNHyKcZ8p+IhvLMZk/GLQPTJH3HS0Dr8LnBk8ppOTOxNIHe2JpezN1n5/h2VVg6WhA
ak88Q9vpp9b+IV7HfSaKbPggGOWzTC9R8Yx+OYkMvtjgX9uOSZplFwCGce8PPnVZLIO0yo3qg7mX
eZzuZIUOEKPlrS4MaJUkVSdAv7KezR0150raXHSidGXy8Pnw0URFnY4zzcD2b5XC7yi0wUCXb0f1
r2jAk5PJXT83V0H2+Iw2ARl04IB3HCNev3d8bsXMZobpLTGtejBBxIqTtz4+IqfWxNlLvMYjVk9P
cCkcybsGDjegPL3F49KMEm2pK/Xk2g9SboR1+RQHfdPArA6lXx76G/ADwpDbO4ZXtt/C466gaSid
cw9p9q54tfr6BKk0ldwzjY6p+HZctnsqD3+gchuRNVgW0AHyKJ3tgDkiBfvJbREaipIproINuPiQ
xuMS0jGDD2CjpA0Lmkmr6jd7HefN7SuIsIED7uJ88O3akj4GcTO6kc9zvEAqfOnpL0POjcp33U8r
WvaQO854reUjgLrTogfcqqAiMyqPMM9oR8GCvhGggV0wX1vWoAeiHbNrLuTUMK6hCv0zTj1iECoK
p2Y2/xvX04tTQABjx8SaCxr2KQkei7T2LhP6+Gt+IRHDFxHNb0xHeFXmJ+aGWBLSnz0OV4ycwqL+
Ic2kWXsn/0HrGdA5z7JiyLkO9nXZrxvHPcsyYLhSdW1w3e2wnTlzQNeN8u0eec1J/Eu5znChdlPH
6eONfkg5NxCQKbJAJl6uGiO8yPUcFo7j8xJRE/Xov3oxE9/PTZjG68TzK4/MbIQfBD9s4vBLyODW
7EQXG1WZTN2JPCOE5KccVcnoGo1IiHofiv8HtbhlRBU8iwrSYJOIs/1cGntoo2UFDuhgqmG+Kgim
iHLpqZGNd1YnLi9EgbiEWNkgUPQSP05oz/D1z6Or6qsrx28vdF4+sfrjS/3ACr6t6PnCU6HoQb44
YqWvx3ArtaqtR0Jn+Pizuzrf+DL62KZrjyt/UhAe76EfDDCnCas1y2mCcvCF2/+I2AJ8+YnXM45A
y9SQn437skzP/pYGZse8yeOD7suQUts8vlI9ymVBqv7e8UN5CbcKSMO6Mau4SCyoE70qNwkzBvxE
PrXUgpXwuWtmbA5h8584tGWJeUDuTTalm9LWcaqsoI39vwOacO0sX7OO6s6Rg3QpGh6MrT1RpGUN
gKZmfmRweOIPAnY0zdTxE8cvjpvtxPF259/I3PQpV1LLq7s8pIVaMSdm9isFbK7GFSzLt6Qqe2CL
037+e5uk21j0bLR3KqwOOjQX9fbc0HL3261O9iem9XTao5Nh6o9bqTruh4Wuwx/4YowG16Xwt7R2
7ezPkA34QdJs4eLO1+/E9SGLfwMxarlgVR4FFad0Cm+EicMeeSuBKX2gRHv9BeKIsJDxzkXS8IsJ
FwHf0zbNjoSAQkdNvcu/3Wruo/vDBopfk4Z7XUMAynJLSZ6caDSQZfbKHMGOci5QzruAL6fo1t0/
eIQonEwMjeRAyEGjOZWdmBqYUEh6avzrkhHgntN+jJ5Y22j7L+tpMmGISBI2e6Qn4uvsTRbkFeAX
3v2ZuPSRYnYmvNBjXHniXGLxSDvJZEC4RzicCJ21zVKOtbHsEuc9mG4V34V1/sltaWvESKICgdIb
aI9MW+CvRMFv1q6f9kVqJYNcRd9FCP9WViavquX1ZlY2fz/J43ba56ovoTY43AezuXDfc1yQQ90p
uGaMoqt3eEf+U2ETQn1TKSlDdEo6QYuujn5jAnsWT4oyC45CYPjk5j2rarT+isxGTsXDi61uoKGt
gV2gNEiLylv20rliCS66T2anlzMSVtVIbGOYTez28DxIt+8D0idUArsq/Z1citHQmx4sLwVgCQUr
gGgNrCegHZTduJyAPW4P5Ft/XH4TIqKgxm4dTYT0ROhTUaOoR99XsjpOIKe0ze7d2mA7kVuBEPeO
/gJKc+++dSEEpbBqs9fZhUzemE8C3sohlBI+lkjxHotdMCyONrg2ccjS6BDycnqE8ZJ+Bj09092x
hEKdr/hemvV4M6v5K7PyElgyMS9XYI9XrQu1nPO/SLmknSN+M4zVQoda+V6kAIM0estsfNQ7nzG/
KCZuovHleDS16mlNVNIytgQIo/qmu30EbqvBa74zMl5tv9tJjIKUjp/dXHQ8iX/H4oBdJ/NAQYwj
Bg0MRxaBj45sPufrx9M5WvMQRozyimiypZaS+HTLH0gDfgXcuBrAUakmDsLIogf5E7jSVZzY+vDr
SpoivMXIJ/EuVREbAdQZdKRlKAqtpS3SOk9u02tbkoBnNJSPNbeVUPhfjM8NqM6SNpjQlmVoaL7u
TcSPcODqKfNECsWvwrxzo7TkkiTby2oHqBqY+ArebnPB+7TWfWoeISBWDLK8Vtc02xNR+lH+Hx2S
psMgOqgVaiIjqZjKwaCGZmNYbbuCd6zjJt8STktax5eG2uQijKayqBta83TTyjwdNS9WrIebvgUo
ASLXFmNYcJK83L8zpCPDaq7x+6B3vy4C9EXrZl75RGbt/5/LPnm7WRcXezsIl6oa+LKm4qglW3ng
E0+2QIEclBaHyi46YcAyg39N4DbfVo4liIXl3jONpmpgGOKrbV9pIXg/FRQoHd92+ksciVbA6Sry
PlifOKqphcR5+mGZ0HFNOHJN9xIRiTIKX0M8QNwDH2Bx18gGigseT8SgtAS1WkiZNs8wqZ3DVSrt
TQ1BRXWsTpUn98fWFQ4oG535loexpIEYYpzmed6taEKXE/Fq/1T0t/eEHaO/WeseWQx5Peq0NyVf
dVI4InGUJgyTLJJDgejBVlJ2RzUbhXSAZOSDJt0rNbzj+A/7BJ/SBC0ls9zMwJSGB7H1FYR0CZbK
Yo+8XD8eWo3ec+vj7v+eyc4gf20PCrIX2MZUAqCmY1NraHrqskO0iryw6S73CRbMYVpL9StUIaDz
Al59Q5LEiup4MQ6JJqmZjwj3toW9v+2uTxR7gOuT6r13h3aLoTvsH9j/Ymnk1CrZBfKLns+w7Ihl
blv5V2hzn04MKZs0O1aBFLgvVhlObMEPGAxX7n1adsAlvvrxdK5q7UNmPKH71fxT5TOSI6tCv5Vk
cvFtd2sT7Z4+AnCWWFC+6alO99n2WlFBHQZebKbxDiGdrp45qwoEoWw5+kjtCp8Rb4zQqTCXqSDF
CnY0zIxKIFzu4gjsMcbegqwYGCh6/vd4slwPuBjeE9ZHMTIyKZQ7Ir3uHOMhKtKdkkbdgRCYmcL+
dmN7laldZKRlo47lUphGQSeVCFyLYt3JGwLb72hFUVvX8OlPmife2772Mjbh3sSsboiXRGXvL7EY
Es2Og/BmRQdevTPUDDgwXvagHSMdWN+M/GKdCoBeCb8DfJI0m4IxkzT2i8TD8conDK6batO64sgH
cF1AIr1rT1A/g5RKPkG3CssZ0NYX3rabNMfyCXYlSSKftSwChcy4PP6AMUX8p60jSUE6Lh1yc0gd
ko82+nSJMZSk9cDxWeHJIylHfX82FHUv6eOmMFPDpxXz1PGnlEX7tol+Whcmq/Bf8rprLvQUZlth
HOm1SiUj1Sc/y5UjxU/NaZu5timxnaNIFg9XYS3MVe3DU4xSZrjBv8A/KY3hGylVw8khVZ/Re3yM
urrNueWLag0mKCk9sdUXGe6UCVz7jgYj+bUOsCPYC6GpjSWswYKXha65ICTojuSoeuIg3hI6dzv0
+Xch3GIytdJRsHMqqC7Ri0OtzWlGgwZTj/Epxct/JZe19hvgCmBcJZzJooYchRpqDJdDRYxabR/B
KaTxcUaUU9nTNp3vYx98+XqsM4zCLXVj2HZYnZte5Ti3YsnUerODC7HaWhcpnIBNrQ8O+wHEupme
/XzEEyyIh6coKKfGId9j8DxLIDJABSB+XZjL0OjJOUL9JMyXfG5AjsHWyKEQnxJ3G1bgqqPvZbmo
WWwlheKgv20Sqo16JItSsE9ShdJax3Gj/A2NovNNgtzstnCTkInubjzGU9nBvPqV5eVpckaEcIBx
gwFzMYMaTlKeDxe1NV1Yhh181eKHwzTXbwVxqU57mfiAhWYQ46ZpKYAD6ESDqVtkMhaEKFcbEjJJ
16WO3ezume/vNyGefPo+bW575fX5Ijzivdp7R9mc06mnqB5qs527MeuWM9Ulo1dK5kq0z9nprHZ0
S5nNF/9tlEWEwmIbswKzQvkWdPyJE95FiJwBvu/kCuJSMV8Qf6+0C4bkuZLwguVciL9jZYa3oSJe
mRytYtWMz7u4JjZSXFx4u4RWor+ohXco/1KWBew//swvLujAKtvl/sAVR8W4mIC2N6PylFCyI+hK
B9YyBd9n6H18GcZ7JxRdK2Ohx0MJCuBDxSqkdVSrf86S9iQB1f8D2TojojTA/u39RejqxJrTbFMv
fHPJZY+fkV8sTQWqQpUyZVc/8BMGvt64ysH3eA1ss52Q19ZblGebi7YHvXgfW7Q5Kxi/kU2wnlMQ
dYr8+CqpznOAq0vY99aPNiokCEoM76A4tAHf5ufQjZBMLA0yYDkSXkX2mQvjofD6ssT9Yb8g8dyP
I6PbBKAwYRQfoLuGqs+po91zquemeQgoSF84fyH1f8cDzgGh9LDDXEZxlyEKWEfFNyFfFC0syApz
R4OCNIxrgkLFE8G0zIkmg+m+l32yq6nu2V+89YmvTivR5G497dKXtv5T3cBOSInEGuP5kA0gnpg4
O7tQCq0K+8Z62FyVVwQYtAVWVUN2aoy5pqStuui7xKSu1gECVh8jtCsv/dA5H2rGAVFvdu9aXNwu
NcT70y8r5PZHFbmuyUO7JT3SGFA4dhetBzjkABtRyPKmQSASDN78rPPbw73RWLQByjfh/cSnauZ8
zP/UlEkXcu5rTzvjiul7gjwUkDadJJMTzUHYj3CD7Q9u+3k0r8UfuVLeDdkV+3rD7kGXf4DvtIOh
/QtGcBIyf8WqrFK/CspF4P+fv9AUmRPYXxGAJnb3u1HRUPPNcyiHe5gQRQLMeanjhxdubDhtty2V
hSXGUVmTHmrki/phYKc5TgLqXvZxLzpKBA+HZWWbYf8p3wACi+HXG2PwHOcjIaC9AS7FaW6rMJ05
Z0uRXZgWLZZcdJNYOJ+ab3+IVZ8iBTR7o79uu02StLBGeOBb20JF70+lxRXrSW/Ee+mG3f58IYs+
6HTlICkeGcemGTyBw+bRR3UxLcrMf8C9bdFVUVdwlyBfvEwr6WQuoWdgVxaz/MV7+XppGXiIVkP2
xo2HWK/8w+3JlCzgH0XH55X2pdPVlIg8cUGiUjsq3Eeha18dPf1z4ymUlTJVIj/BSkUSHpWmNHAn
yQnJynNms8xDE2GHVeK3Eu3KBTZXQAZIi8STA35o3TvmNlxYP828dVY3Bhsy/ahvmOhL/env1B7g
Qik9Que6do2K35Eftfi7cdW5E9pvgrvB9fFsFo41qhgmOlqmsEMB7SCcPPxeZAG1Eia+IIYUpzmt
j7QoWnlQSF+a+m7EJ0duEVuY1HJNh/c9dTY13r4FFRVQReytiQ3vFGsZ9YuU37PH79Yu0CzJU8ij
0JKquYArJUjHAsfqmHJOGWq28DN+pfCL08B4xey3FHcoTtQ4QiSaEspD4akS/W5IPCP2jGAKOZsz
rt57SsorD/1OzcjRFo3T1NncWf7LlBFgZsSKCFfIYp0H0G5NSqpHJhAGizRkttN7RcJIRlskmSYd
NEZsCQLUOAVnGb1vD6Vcgc2FOu+wY8L78VC9duRYbVMnBgjwvYvO2FRSHmT2/7ovSoZ+arKJFM2q
pnwxPTAIUx0iwj86EFQyM23/Jyvi0f3MpMTxD53NnGCTCMQGYcTlN6qHSwOdtjfjOm3rWkOmLUsF
pFojpziFUnxCxhzsO51QLDJZATcnCEmSuBKaQ8o5JBExggQk61GpcHRlaT5ziDM1F6T+9ca8S2U/
zKeK3dUHELP8/hrRjfmS3ySNduSRo6zteN3IL+o7O3vi2bBfnauUztsS9aeEEPPsLSQ8jSAcBr2I
XJK7H5rbjUXJ1IXgVqxkpsPVxCBgxhU6sTPwVAUTOzge9OII6eTnqSSjodx3fFKMNUlWpjjwLgiK
b+WAJKXWJzzAguEUJ23bi4I5h2JT9KRFXaIV5Z6Vi8VbXkTlx2j3XfIRWI5JiFfbSTMIzn4FXj18
jrn5rF0kCDhTda8YMVkZcr3ENpeuvw0m2GZXl/Qxomt1jI1YW/L+LJ8G88rZT2WlcXq+Qp/3lE0Z
7pHwMvvPyzpLbmOf8TnP+5bjPYqMoKDhsjKdK1aaVSMswq/KCaQbGwcDmoAVzNRxGYp6HdgPCp4g
HvYYRNXWz0SKFZLtlGe/KYA1OXVNQ17eIf9sqbcnHshBBd4ARwUQ8xK4ZztOXlpm4sjRRs8iwdLs
eBrJiYMZdKivP2b72oJvPDzskSGw/FBzYlua+Odd9xAI2fTPrBWSbTj9BrfdOgwkMwL7CWVTv9yY
hTRqT7e/x0bYMybvCz15okOWDhSQW3ws8d/ENaN/y7k9YuS1YNyPWcm8wQPFeaVRs+Nkk7SW0ZYn
a1+r1+kIKXfB35+LW3dcJT1avxeP6lOQdBumHuPu6mXCtnfKVENaBmohjzyRkjydF5GHIZc/ZCBV
EcomLizBxGv50LcazMwdyfG/UXewwQnDHtF5t2Gj7NKS6ReF8M4S53XS2h1IOSGPNGFKJzRqZFos
TkDFV/ozY9Na2xIGi7gjsu4bSeW9G035bjg4I7PXAkLNhqJljvMjV5HyT7fKyp1l/Be9DEqN1X6/
d6i/uiibDadpT7PWzF2IVeokVB+RTrTr6X4Qa0u+OuOk8XuE3vhl5MUS7ZRv6jckZIB1APZSCDhL
iLVkGhgXYvMt35ThhPts0HOalIaltYWM4WrJAE3gGOxQHMPZboRci3CnANiQWqy17PyC23PtIa23
/naBE0NQWqoj60GzH8aopLAmano8FdYrvSLmG9edCeQZ840ocWEgMAzTmL7AVfxWOoniTEA6jF9E
+lVU91hk9Lzox3G9giBzN5psQCyL+zu7Yb+0qZALdJXCqIKr1rwwR/ANnr5hUbE6FKZYWbWuYWu/
Y1GtlitGiIkHYHEYVItfwLWv/WE00RVADDNKEY4RlErDKBkpFgmDzicSoGK8F5UNlIc39NZNHzLz
cFpqBcx6rt9aWoxvvbinLxUzaN3IY16fmDg6HfRBUFGAgUqZKlShiLZ2szRjEY8HHwiEMi3yx3dZ
VgrC1Y8emBQcpQuwM2etZZAi9vjxAyTV4cWIn/sNIk8cWdOKJ0gRGAUpjDbzDEdu0ZXj9ME8gl52
H+iYreKV2Nj7uf//uihmOno+jLMLdqVVqSns4xBEaM+wj0c8Ce/ie5CJcpTB0PqRXFmRb0iqkGTi
zbas2SP38vgwGfhPj28QMkapzYnH3u6IP50AJFlhwi8Ry/Zu8qxg3Wwm6+0an4KwddiSSvXTzSHk
s1pUKBfsLXceMRxvSjPdtcQ6kv8H+DmHZsYSVZzM7A7t9OGUUo0XoVCTIXdjBu0fMOfwlgqRb+vl
gMNeyPMEWBUV8X3XE8v4Yk7DNCOzkq5LcMKxHGiFcR1pooxG4W0XXL1nWThQzVKKOtuHHob7RLw2
QCf8TQbyUoz7K86anx1P4iIRHVJd/+Lg2PWLkDtGngmUYuan9troqfyuCp7ruGEQYsUg9/zKx3bA
r8UGOUxi2FoDNm5g6wzT6H2f3Jqs9FaA+j12ndp8XihvWOUKmr2EG+9iBNnSlSTaeyQ8rttPRNmC
F2q/gzZQy0QQuNXmhxJPYYudO8s0X0jcj5Svz4H3VZTEJPb4r34n4JeTblwkT0WhPJIgUjGAngnS
dK4p/5bb2bxbKC1pD3NfNQ1U+C8S6RESxC9D6rpIovEXBEZPf0beYdlpS8RYUi6tUgFbpFaTz1EY
RduE8le4br9xT56bFSmyJhiGr1Zu4TnWBd5NKdhRpAGobhuB454/VhXfTpqwlwWBw35cMqJOG4Bp
iqvh3loVGK6+xIvtGLdmoUxGoy1Cm+NOXGwNqSScfwq/M1vZ9t5PEUDSnSXA3pbUqgxgHAh9s1Dp
lqwUvvEO9AlJNsNNjaie05m7pljRpxOJ9BRRaUo6b92CPYoVXSZ3lRnzVAO0JZzXB4JtsLyLBMOF
F0aiMp469CQgFmHwOMnJXf5GV5QpSKOEMvHlQqIUEjTdAg9RVXOlVy/B30mqjjZ5fqvAx9QIRver
qFbQ92VMX7P9QeiD4RHLYaWxOtQQSWqZCuO/2YFlDReCceGAaG1dp4ibWFkfFy3OPGgDah2cj2N7
PPGPVEFAnxyR8jq+5OLG7S0jjyTDLhrxkqLQDC/5riXr4TparpwCjtCUputUGFOtOBY3xekqiXOu
/0hpkree0wCC/f7DCABQWonoXJklQdKVRwe/5yJrTNMj1T+bKv90bjx0Dev0chRyW1GfkoJka7EF
m9cYaI3nbjcqcPKLFfhxjEfUA2whPW2f0YNAJ9l6TOZoz6fXRBsZNwzsQQIHOfhrSVeX292NqVgK
oJJvXXRvv6Q1O1p1i0c+kO54SoPyamKo0D9VdqFWVgb9R32QL23LLkqWW2QQFANWNvZRbvvJq3is
lwBFDaaj+yj/WS5BUI6hNZngUkjOENvj0MYAXsD9EvoN9jqipb/S61U7zQ6rG7iffCg+Maakqfkr
i9TpS4v0Fcd51ZX5MrcMqPhAbwZwQnKV6G6P0VvgO6sXn3u3uCrhP+mEdp5//wBNA0KIOh3fyi4w
v0WwhGMxwFW9rnkXaHqnIoZFTFfU+yea4aTUPELlTHrSOYlQTkCZo63eZZhaw8btgIi3FFP0DENS
2noHJ4ZLRGhLaGAmUewQM2Q+97at4+MY1BhAjQQqhmFEcfV+HGKrfSM3c+fq+npCr4K2yhuAT2Cm
DUIJuUPEN/YQdOzSzS4RD/i+8Xw2gouyzHIGmo1TqgVC7cNPBhKtPhIayUhNLd7vRgAoTBcplNzv
vEmFLQsGc5PLB+2QkA2D0hMq3WpQaVCtleckY7u9mWtlUYSivMtSIsm4FA1XdLOPol9vf8vQNDZO
k4DnlTtruEOFo3x2jShMxCPNDD9hnqjvODV3abvOnYmNaNYARs7GDKzZanni8/IMEejoF5X1eG34
TZyideVVMfRwaxiaBDdtjkS61e8KAUfdxo4ens4PXInnLfaEoURI8fSKm1SqGml/XJcYv0xfjBcS
7o77NuJFCogN55CfmHt+YLf/h6+uD3PVH+AoZnnG+Xmi29ZBqnbVdiQGUX4djbbluWNqNJpJ5Zry
GO8ZqSUfCnRfcvYT+QS+p9EmI/Qv5Tu4tr5y8xDZKO8aVnhHYSZe3KoQQ5x4mMiVkD9qgt0v6gty
8LND4TBj+6NyfZMRsEbBrbFZl2zvA+aiUiWsRlW1D62pk0M3+megQvbqfiqf0cVVBKcJ6x7AOO9d
BRLMyxVjA+M7HAG9MWpShr4/U+j1Q2/aD7XxcEiwe/qpt7MWuBgzzOeXXN0FT2e9YvAlhjAIMgw3
vIEHV6SFP0lnJqaNdzxNiCcZvoWiNEu2lYqJLKW5U9ILOT9lc6pOR2Qit2V4YmHS9n9gvFHbP8GX
m8kqugDMnqPw7tGY0Otw4LvKJg86x0Q+1Etwis3a2whis3jvezl0SFB99wHsyFIvpX5nIcsrpVmj
kcD175cEyDLz5IsQpDy+SSrBjhIICmhtM1KWepBpoE0Ft4d0TpIPkJzDdPOvkxcGn+sM4vqz+A2H
Tggx0kQ+ZTPjCbNucseE9n13fGM2O9Y2Vtbx71syWdxIEqzzd5rXV7Vtwx+gouxxq2iTEunjvCDP
n1TW4vnZj7wpWlzrdQOj96WX4kePnmGHwAnkk/Bn3X6keOk7X7z6YrnNUTmpjTLIHLPen0Yx5BQp
PIZXAFEkAQoI/GkROaLa4x7uFzNhIawKgs19UJuqVmKqAEoEx4p6Yxt7dOYY3EB7jg75U3a9j6/H
JGd7tTBEl7F+ifKM3LN9+pyvIKwsEqc1+9siS7pUdNXwco7+f+Dw/YI66BBgNaiJkzkLsXm9J4kY
NeWHaoNOCc6Xi4hkKro4ChCrKOAN5C0WO0qYidoEcI+ndexpA+kf35ZxdGVHA2Nc4Rd9QxoRZ2P4
Giu2zKVw6jc/ig1rrODzQIKEDuqg/ZHFnZHXzeC0UmfcrCI0zhIdDBNyeFm4fzIJ65BYoUd5gTFe
cezSEkXdxPnmPLi9gv+td7SSSPLNd/AK97cLyL8yp8jN1eE7zvzRSsMQaU58KwL4X4/4EfkyCNFo
On98b0iYuXfxHGlx4dh5D/v+y7v05lKtaWKiICCHCEr9m2t4Npn9qdzeuGngVoEbQEypA3BKqXbd
BSgYAgybjmvgwvGtkcXiubIweKmi3QEtOHQWnTRXOd96EHXOxpUvfLdZgEvb8jyfEfBCQBtNAK+M
F3rYG7M1ssD4r1nietZWhgrdEEQklSOQbSe4NT+E7hG+IHaWhgJUsQd99WAWERI+KiL604Qar4Zk
K0jr4etlk4aLi5ctV3i0i/CnrMt8+W9y6u8wHi93lKr1DKEZFVZYAV9WQXBfo1l6N/AZI8RtYttT
zvcWNM4qx8N4s2mPokvP+ePb/QNxxKHF9/OIr0bkXtOghSvg2sbmQNtrevhUsL46yW5Pu9xPPjss
CDNvsy3CUC2ldg/8+dH++ttRtlnuBeFIC9a6CR1a7sRffFwzZoJwn9FX571kTV3CtL7mnwKyi5KE
Jbn2wsyJGAQzhoY+htPaI32+Ko/Tm6PJkRem3vYLBvTdm7zpNuAWyq5Mc8XjPhuNfur00JZ28fqM
SAvl2WBFq71xGgjzalHMDFdBZoms/c7ShZd156axQ03SIczZa9rP8YE2Iucwg+2CiE7kT3Yx4qRh
siwAKX3OTc+UebTaNRhmXUHIDOd4VsnXqtJA4naPjEhwgd3tHYHBfne80Z4bgCG00Hi2kqYggkzU
NRqkk2ibaGoUBDEw4Xoi19KaAivcibxM8zKVdqqJ4S+3z130oG8TCCp2A2l1GWMOBf63OZw98olx
CkNrmZgv7TINXUKHbeC0szcG7I52iyDoJ3BrkVWMVevhGZNj/pXUBEVvgijb477atzoPfWcGAceH
07TsyT4porxIVywdhThu6bDrZ9gMaQc/GSQfzGhxqFw1qCSI1aaAFPp1mXyfNabBsxItrBDa3NmY
rXRtC57ED4uGu9aAk8+kD7nL3KpRkPNfZu1SqXFehKsWIQasi/6Cg94IQzmg+iHjzRcCZAAoVLlL
B7bmP+BxzkDwW/s6bayFtN29huMXyyFUYFyqnwh7r4PTgPAtvnW0heE6E27n8N4aYKNt6DOgqsJ2
w6WMxpQzOiHA+2u/MS+zTX5sf8oIzRZzpk57sEkAWLCPraEAHDN7hJDi6q+fmT8yZ4dor2BLuWUQ
rAhUMws0tR5ro/xCGhwrO1KM2RNR4+OS4ek89f0J+krOtDJD8sMgA6M3pHnNpYVigG6PnPK6+Xhr
LmOYQNgHHjRqoi0QA+7queZh3oW+GYFVDAWWgrs1jJI4WJqSFP2cJDpGnpDpav5dHqcbO5Gwr5HZ
bb/A+IpgZAbQCDI6yaRLqOvDFGZ2jev9HPOsjylgu3QuoMNxNJqhpI6zV9dpa1wmJNavc5Pue1aP
noDpkc62BwZRqNKGbCQyYrClKthGgBRhHKE3XVVKhFOD1bNNM9LET58SW2a08H4mTKXNSreJ3ZvO
z0cYbUOjVr5zCYA01o14bD0ywsj9z4GjP/9+GDr0f+Z9DzJxy4etIksA2Anb0Xw86k5Lv4bObyu7
m2uCswWxfgcyFXJ3+Fn06uNnNWjZcvHZNC/ufRraMNFNImqmmt/GtBEKdbtccgUn4GVWs+hzQVPW
FMAVNkasckx6g+xPUFmTBMnHxniX/3hm09X4MraUzFM75uSwYGRHJbbv07NagTsceGGWndM3MOBL
99cJNSTUcZgM2YK5l2DYDdK36oDv1onBFfBHTg4Lt3C6cS7LNgPrdORY5mzM5YlZviG6A2E3+40u
pnpzLnKeVqhlFrZ4N0g2edMcNArR71VXxDav5pEhQy8vNGtZqiuh0le7gEO84AFhVbNuYRANNr7B
k37md+d31qTRg/cs4uKJiWQ7T0/QekhlbuuCfjP5cCW0XfKODnmbGRJCHjkTahqVT4vZzfwpVThL
Y8BldwqWl5S2XSDa9P3z+VRUQfWkPOZt7B5QYDt0npgblsMMf6uLgII+IkG+38hoxHzi4hHhGjJV
8qtAGkIEt5siD4pPFOVfttJ0HSDnXru0Dwl0/0rHlOjLvu+EzC5TtsChqmy9ER4+pqi69ctKoKbM
HybfVlHSmt7b31EH+SzyUWbeSdY8gHr1SR2H5U/Q77RUfaWb46trLloVr6/uKAjP3cFrFlqf0Bou
em0cfPPS7gn8hmV4XT/w6VF7pK5TWwT+pwNq5SD6TyRT5rZBwqRtFxSwtmOJX83uF8QP8STFTTgD
JvCjFp/HjInT3YDxM97Vp1exI0he2+bx0HnpTNkhiopbSDz1JP/nssxCp9HLOkkAi9TYVKxJvDJF
1lRtAA4lAon9UlkwYA6mCr4kwS53OtKpC4E7dMgyLoEgo/qyDk5OOhTsNPXkcrewNL8S4zorZDP8
aRBgPQFwtqcVSHFJM8Nvip6k09vY8s/av6JgEwwKA82kyOsFO9fb45oELcmCN0WxEjyzGHIJOmRn
f6wZON5WrKRyd3f/8yGXsYE0HcgfUvScBslZgSVvP/vl4a42gVA7Lrn33gGd8irq3fMHw8V5Wd7w
Wt0bqcQycexgW1Ys4DbxHzlJDH20VTGUYSdjMwU1wPfoDBv0kElfP0tbDPgitdAbNBIi5UB35gxN
8+j9ogVCytgpb9R3a11Oxot++mwzZwGr6V00k3m7X1mqh2NPbPDAuF3gPkAZt91cab2hrbs4CCVD
9x5jo+7PCWj+IjzJKzFbYDTtV53sGSjpMj+fhw2ZJrJp3zFm6ZY/pfljLxPPNlbYvJSMtaehtndU
0c23hjUBYbVFpNg8doK+w5mdu4WRr3Zi5fwfrJGnx9kXVIsYevYXVIILN79kej2qJJETh+/mmWqg
M73j6JDFb8Q4e0J/nIiXFO8ywGzzulKNVp8GqlqhxinkzyyZtjgOb6nbqOA+GP4TWm+MTZ7btng6
TYpjNQph5I6w2LtsBR+GHqrV3JvRsXYV6CKqmMLT5WdLhH2aQMZcwUTrYgbPdXzftUSzbvQEO9Kb
dOPYHa6OyoiVw9VLG3RSbtjsn+xn/taEY8qawjPdUPK14nZ3Ud8h/qKVn8obytMNQRgOqxxynvvZ
s+Z8Hdf2TbS6Exz/HziyTlEjLegBJCW0TeQhwY2JL+I0CRWvnpn3rTNf7sUoLY0nvfA4YfGu+ZAQ
zU3fjO4XUANgo0090Mm7F/R0Mj7hboyYjhUaThShUjc4V830JV8HrNvu38TmN3AsEBLySxfIlFGv
s/kdedRbYU87oNbgvYuMjHqRqhYZhAK/SkkUkAyr5+2tku+Qs2mxqZ8PZEdFZTIhrn3dbnMo1ciQ
BcvShMSuUIDYJLrTBp20tGGLQ+0YLMBTrJ9EI6g4BiV8vEQ5k745ZzghM81I9zKuDi+ngEH0u1t+
2xq3Kon3KG7Kkkdjxurbps7ICrHqR6IosjSRcb1AO8PQJsOX19aFWxR196awQZB+KgozHT8yu+Vh
j9ioHJRh9RJs7wDWAD8BeqLWEGDZZxejFdjlpgn15vRE9/WXdFB8qmAes7LGjiO0SfmxOVlbEQji
StoobKzATuSG40P0YEm5Np/b7RgPkmOyF8o7LyXxiczq0VQNgffaKUI7icLT3XpsTP4AXGhkC1gK
YJp4SKEQTJeXoiSZ8OsD1MRslegejkdL/u4fKlGGiSJjTl+QtaaSAj/oSXZfNpQIPvqMi/4vmrLY
p5JBvLpiRp15lsXn0M2fXxF++xp8SeMjZjX6vNFdaZjKt6CoASo354nC1hySFnJBPTu5V0T69Nla
OqdDjdF1bnxTM2ZJt+V/ZDLCQoQ+KFn/D0DsaPzh3Y8SzJPiIX5GMRehOSFPxcuWyanKDoEPZxLb
fC5rw24AJ506foVrReD7hQfVVB6cJY2w1BqDqKkeM0NwvtmZPvQxqjHbRY2hpw+x9fIFQqVmQ2UX
bZIQ/vDoyWZlbyWmrDHhJ+p5EuHeQXi581vQnXexxZBAI0NxGoje3gRmSlHRpPvASfcwjj+0c5JB
oXG49JENEsWobt3Jzd95PYUiXwbc+siLI053Z0r8Ehzj/DFK+qPLAb25uorjlO9VYryWFCHTfRCV
Ip/wekTTxJoElmz6xaP5G/gPqYInWmmiWd8tCPKrMWRpa4wa7Op1Y0+FgRIgMqyVWMvxxUD2xKzT
Be4c9myO7fTdefdD82rx+d4IXQqFGwpOyvun30ySXIQ1N7AQFnz6yjDlcvNMQdbsBd1cZxACXC3d
4S5fCI31oXc4FnT9xnnmAXVIXmJidAb37xGYNV5/A0HhVE+pYlKUlvZ4xzFnGkzmuFyf1JhH2ebs
7AsQAMAZqB4J2zaO9FE4VfyRfrwuYcwoTwLP0o9RS9rnvIznHMH7xpEFssjgOD4k4QbfCr30UNau
mUQkm8iv3Gy7d50ZE7oPVpA2crSsa3JwZvaq3mc2zVEJG11BtvtkejSM0W/siE0K4W57ane5BFLU
LszOfpXxqD0n3+3ZbQJ36x2SKZBiF1XUJKG7IFvI+5Bsfd/kcwEfYfCRvVlC9r4hSEgGXantoikm
hOsvoemfbOJOzVxypBM9FKT0TJynrRdSmfXXkoXgWVm+KyiaWzCuKNTEHu438OQhfQX2N3aSsGFx
41DqyATs9hsM9lQp/iheAx6TW9phuwjmx9WoF8i+mQxeIlcGYjtG3CritGtzGMIjO9at1mb+MORL
l9cldBlNhHfak+drtX2z2Dcaoh12/nmLn4RAy6o3RSV3zaeXnA7xTl177xaQXY+3G/oq6diMDH8B
FOKf2MdDXaOHcPUDQfl8X3d30baqooPL83YhI5hfsVrqSIMZ6LG+xFLC/bJ8hJkwvaavh021bocy
H71oBobmmnJbl+An/ZodXRe+7CTUixx0Ns9KALLS6hlexZbYYfoDKq0oe1rsM6rjeUAuyLvhwBNM
PllckbU8HG7xbIHgKK9RvCDnR1iZ/6LX5QKTKhM0a9+zxc5JlLZICkTq10SkaZKUD0t/B5crjkmG
JfCu/t2qdZ0Pb14sn7C1RFTIc5MYXEubAY2oNoE+y2kvWRbnrhLFQtLaZY6T0Av4KBFxo7idG7ps
tOsp5NLAnCyMUlusUDBGhSrrYhns18L62x92B8XerKBD7nqAUELHKg/hSQXlfRKVAb3z7NjfRwlK
eSodDJ1+D32p3xQqK9LfhU2Vq0wRIGAaLBOCIQJYwBL4XmROTBlxv7LePlByOqdEzLF4WAvLSdZr
mNB4mw7TCTvBvwBzKN3mGVQM1btx+Q1Og737UWw3QGzoK+pFtt8GYrogQQFbJ51J6Qupk+t+9RcV
FwQSwMlGBOVljVMMCAwtShhPrV8GIGsko5Cq/ZNfOfTNbnmrIgt5KBtNMFoKgZLiZglgtXFrpmtk
n0wHBSlXq7OmN2J05kiAyDBHwotztl7omRnRL1gWyeDksm/JfOKyZ7xNO5+ODTznk0iXR+kncWuR
NdS2CudQNmPBcWnUqOXSV0bTCYiaW41GXzz10HU2tO+eTcX2YBx0PX1vu3ZcY+8dXY9Z5VMu6zbh
lL7Vsc93Vk4RXHcZ2eMsPAiLWW1m3yBx7AT+4WZ/o+hmxp9gcuKwsnE9mjBq8iA5D8N0IxDQt0nW
bPLO6iSFFZikPQl4B7jk/eNQYLVdQgSfVnr/jMSTbOw0cnEy2BIBleQGAJr4rBS9KblfVOhKD+iq
lNiJqFfaQok4c4QB1ihMhgqQfvn0Io33ni8RdB8riTElmQcOsw5AxWzzGKqmagwdWTSEAKCorwf6
dFbaMBm6rf3iVKPhVag2TJ8m0+sjIDurdw6ZQnlP8PXvQNdubhwTPCFIF5sfTRuW2xb5PDqwGH4E
b0WeNawsXtgitiDLSmDscYH/ACpR4wZMcRQ7lOxndpKCipTGx8dQGEm4gD19O+7qVUmPYgisJxZP
xtuD29IBvikReH+uEzxN7ncT+0Hg5hquWYfYztAZWMoy0pmYmzHgF9gEfwRog0idP1uTF33V8UFb
O8kr9UvxCbaceEGruhgiRcZ6Em4P7tSiMMrELEuwf8gjumgCHDq3L7PfN3O8nKbrOerBMFrLYbqy
C9KCFRr8kp0OsvIwchCfn4l7NIOgi7hqocQiApQ54NQbx4TtpQvH6EbAMJ5m8U5CXXNKOInUBAeT
x9OWRT439SFyazhlllAH26YADCCEeQSUN1FS80/+q4UD7W0oOQVU/9QtaYT1JVJ70uOVp4prdzM7
7dAQ0uRRnWnxI9dz1dlyduAI4PRvfvyI6AL5sgZROGaH9MYnbdVaZeftsSmBHnWwuFfwYwSFs4ua
zMpA4jC0c+1O3Ci1BHtJkf6Ll4+ZLPR5jB3vFIhxJgzmePFemMaTPQsI6b44mpnn15YnzF7f2XCU
/TGg3azxUVHSJaUuvh9oofTSzz1FPPLPua5FKuseyob2iaGicB/bsmLovmiczmn0WW+o1NmFTnnW
r1/CL7GFUvk0Sbg8ylKStoelsYh7+PYuB+KBugHUWFnYaPE0BqS7W5GYW8aUuv1W8vj1c8Vr4ZIn
0MRJ4pXeUNRyCEE29Hvq8WBGtoi2MZ8PwfVm1oTFQnsxuEEpe2BY+dwCE1t0jTIYf76/u2mJaUUg
AelXmrVfO2g69ZKKDdwbEXl/KNm0GyZlvTWHeUbRa/Nrr0HSM5pC06u4rbSz362tRqWlgJryH2tz
I/pk4magiqgIqS8pgviAEFbavk94LlwhsK5zLqZr3LEge1oYBF1kk26tLZT8NL7jhOdrFQSQrrTK
bO6dR8A1vRakA915Z4PW8bUsyuyCtnhpAqAqs2CrawHcAVSNBCNNRTTXLCEeVcwQ5f46HoJOZP3P
PLCseWY20gHoxr+fsXDgmcybIjtPiQmSe2gCqpnEnLOsgmNps2fl/QCSrrLLXcVvRkYscXch/NHU
KB15TAnEXqlmXuzl3JYb4Q8PgtDZO3MhCwd/dZpvmkb+FuXNDDlRUdYEhggty8/2m/l5Sg/wlqGa
sQGyD3bEPCA5rEG3TJx+i+XyP7h78mSb1LYNcdWnrMp+GKoVdu30BVs3+J427EnncnGRKkxJm6U5
cC7lk2d/k/w2Uxm7JN3i21DVbVu6ak6NcVPnA/A+QngWe909c92/ID/OwrCm0FLy2n1rXIl5kvbN
JjtJOdARucmVKh4OfghTgur9T4ahEuz2Q/QIqmX+mKsUF6f9OVXoGAz2tENkNLmeWaHsshwE6BVv
diPTdgz1UINXldnR21LuiujhS76z/hISMxSIuMGL8IyVuf/ZJIYAOK12JMbwEFCkoJnXncolZvSX
CTwQxodv2AqIYNHaIqEl0pANzsAro4+sBPU3X2t5i7K5ggNFa9jbDroP4nLTuMlNWwY1l4Yxw+eg
O40pRazfmEw7X7ZUbPfBCuPR050epxhxZRMeAgvB030oWuxaS/7wV7h0ifs5iICSAEoBe/Qfmn1g
cSafPcG0rwSanY7yEnGjNR3mTOPO0YF7pb/MRvTedBOs1FgboLvArSC7awwWDLVnOoJjW1PU0GWA
w1zUo8fKfTCLqcwNsgDkdAL64AJ55uZNpBg4u/A7Y02BGDYwvNfoOcLOPYhH+GT8NXa/OYA3QIWV
RINLpeSm1C2VpiDRV91fBaxAweStVR5j4mXEURJQcqYu8CRs88mEAVYWV0KBP2z36lzihxE4SmP4
IqgpKZksEu7n7Q4F1TJBW9OYMPpCr09udOmtOYAtfPS7tbs2T/X48JGaUM7nSrTctAszDGB0JrpY
FJNrvg6zM3VJTcEuJmJZmLpvGsa0k4r16bYW/tqR7P381wiZWWm6acW80tN04j4NfRnNR4HQD9rp
ZXLv5w759bgluCJbNvZUcOXAJ1Mvru9a1fyoVXoFqm5//2k2RgD6LuEsE3taFvtzoWn7lq+UOZ8X
319xrxnw3EdZE2aWYn96QBE0A5GCy2E05Q8ephY/+gdFqAGeMPaM0BcIK8YsMhzIwTIYY0XQ4TIC
aqIW5Hpn6VrOrG0eyMbqjzjgDc0TovP2Nm61YFDy7oy2+8c0D00UpG0W8IDh/L+A38hgG83PM9FX
gaCbg8+9GtS2tr6mKBxDD+hl1kzpC1NGuoyLqcFV2txWq+ML9m2qWaS6wlIvOhYgO77S3QWWSsFt
OkhWa/DBNioG8D5OpD/sHdySgVR9sOwAKZDWwZeCjZLv0iOv750+0y1Bxq1dhEA2MbiPe2NoEd17
CEmdv60ZXqv7t+vg52WCB+rilLJXRs5nejsW8fR4xzaBoOQML4kLKssPgpdwFWR1y8MP+/wEvkAp
txtT9UcqVk9htZa6m4d+GsH8vrLpVii6HOPH2LvMUmtqUlG0GfGEhqWbnVqeFw+m9kBF3G2o04NH
VD0FSpUB7ZlZTt514Hf713frnLY8gtgo9+Exx/w0wV37OrNBzPEutyFXRWx771pzzHK8ycF3RFR6
oTOnJclYrjw+Fs14SvaWMW8EJtbnBrFi8UMM7YRL6nuzivZMI5/YGCFn4HelEOVcUM8AVaFTLKJC
QpdE6S4E6aZYBysuCnYDWW6woLzOo9cRVsPObGOLQTa0llusGEKeizEb8oxbgztEsB3Bdq06+KO5
YtLsujvLlELXeRrm+E3iNBQDkZ1h2WUjgjasteDAqyTrLclITK+DwG1OWle2OGAe/aif6QUEYF/b
xvQQSCrUj4O/LQIM3eiV+YEAgii1bURln22q4Co/GHyEgM8T3h94S5M4jX/2h8yh1PuBQAWVD1ZV
ycPJCW9uXX0pgS7kgDStqTTSNcFlWzihzbmpSSJyTcZ7EslT5SKFN4Xh3l3viQ2tK4ozspU70cve
nCIyz/WWKOZwVv+hee/KnM22LWVSu4FLdEXflDvdck1VI27y4aZMz7LtZUEQL+v6lsNs5ysapqr7
MVZzofihqPZxV2CKNGJ3pmZ5im0D4jUQdte8cf8yILrBv7HwSbiWLWTiPyWSFJkPtYNRZwUrfA/D
0mfMs4hMh4Q1lKatcDDTtx8ZE7O1tvfzvWhmxwUuVpafgoMCnq5uE7WtYts8zsSJWL+EYljljhxv
gKHrxqIAzi8AuhPnWIkJohVpw5HmkIqxIOfj8rzT1EZDxvs5N0yQ1YYKshkexeBVxAapIJKa1XjZ
uM+3lrCzojq1cz/DwCUeq/J9GMMNWfowzPPNRlQZJEWHqMuXa/yD/IUJmraA+17iSt8pclwRvCYD
Q9ErM7f9NGA57vHtC4Gxw1r8QEG//rXsnq48QcbSZ083T1gX50/PIlOZDOozvt/IYe72Mp7xMbWu
uZpCqeXCXCdZcVFoX5w0owIHRvvYdhZwyS7DGXJA64XwpiuYjZAC5g5GzobjwteHQL3lDzDh1GR7
t2BBJ7Hg9Pph+zLwrqXSE3jT+N3As/iF/r5YOkW5nwSVGGQAYZ6aCZvlU5r1Aq1woP/axj6PAuCD
2oo/qSL3vc/QrlZbUVC7IqRybiICpFCu8xGjc55nGWcRDAq16JQ5cGaa7PRO92pcvXyr3bVUd+U+
MWSAW1MFw3kSGQ2C1vI7uQb3MkDgNq1NmOWVD8I9jknPa3UiIe5W6pa8+tP6JADfYvOOFmBl6S+C
LhQu8ZLR3L6+BRO/LxS4bRtLNd8IjsLfUhzgMkrcMi4GA0M6KlIdlRkbucEmwNKTHjFevajjvE2W
aeIrprjNRVX9uAYFraeEnjU/E3I3wcgtiw4Z6m/lL9UfAkRLqvGGy/xVxkO5pvqF8RGMLZTqT3Bg
1ruv7OrhNuuUKl4AQcO5QOZZBWVZMiDzqJuGKm8Jb0KvaKnT57uajgj9w6ybet8zXb2fgaUerbSO
YWYVuamCjI7Sk9OMR6snUVABrQtFadUild1J+9H0vpfzDm13b04/CuS+/Kq5um3OIstauJmMYVX8
325VTVd04SarnevunjjwuPdqKQH2ngxI9NzNG8oJ188ekUIPxcCCrn+hpEO03V914lZ5f2smJ9so
6XsKqaQNRiVGxVtsTFr+H3w+OtfqarLBEGqkOTHNTehnijXC26ouzDrufVGxPaz1+iLvt/4dA6c1
0x5Qg0qwnAS5JyLj7dV6tQFwn5Q+W1Fe/E+Y+8nGCi0tMSCy9+qpa5YKp3E328AktvKJ5jQtH0Mx
QSxJV4aieHWdq65Y6s7iqKNlTuMLztcS0JBtvhiFEvDeNOi8DgaKmeCMaA8yHPdDWsjkhUNKqc6z
Jv9LbUaYn16Cfzu53nbsmsKXw5uSl8THVcFMfxS70lL+wuAsqYQUvvwUluFL1j5/prj6svQ91ah3
8aK2MRtHhrC+u/P/fHqJ8y2DLtG4SF1+PKPBaUEOhZGfF0tNJX/kywaOg+HS6FJFPQI0L2SlNPLd
sUyQHoWwZxE1i4gz7aHpdOrwEDYnvJBdcvuNHY9OkP2JkXwNCRagEwqDSFuwwmet7+F5Lntozqwi
Z88kELq/3bTQvw1vGWhh4YZk1V/Zak6rY8sP0D0ydDMZeCvCtMgSjERB6FPTBH0wAV07y4a07sOP
WxIKX5JQ8tpWnH2EbgmsB+CmPqHE3ROhJV9Lj9NHeukMu/Z2Yp27+oscGaGRMKoBKwfWqhKNa4Cg
87Y+KOjXXEsvoUm+HAr1kL2/SmLc1NhP6KMFJ3nA9V8b1A/UXelX1Wsr2gT/N93vcApG6UA80V6N
QI9VOMiOd3smM4SR6AMSTWwKBrPx1EWsQpy5X0kH4QYJ1JaNKdRw+znMTpxw5Ted75HUokI7gfMu
BKNskHG7QodDhO8ocseQCmp1Fv9pxkJ/9ELSYIPlD07kZHPDc9Uj2KAXi3UhL2BukBnt4yo4/KRI
xgqUT5RIBDeLqTfJgxA/Ezzae2gMLJxFkS+GuYmDKnl+QSEAAmFvLwjt38Mgz1ukV9R6sw3gOsZT
nqKwnzgRIiSFt59krIxlWZYOvc6zFDasdS+kYBocBkmSw0mJ12uuM53Tjq6gaD7f04ohDpO+JCwC
Bpw/lUFTWfCenOyPukXpFmQnc6Y3dU0KQI1msS8r/GvpF2Vou2K0ukEmwbiCXiuPfs/HvBQYHi/k
TzOEcn4Gd8wWNmgw/48p1o+1QjFNQ8wS7zP1bwyU4nHt0dj06jqj0tqTmlyB35d+VULMtb8ThJJe
cJuxW7km6f/uCWU4OK3OK/HQlkrM/BwShgwaTYVuO6j+82qdshYi3Z0Ip+rZDFQWkQIYgBr/oBIz
Q4dp2B1misg8gPwdMf6GqTQ6JXWsKZJTP9Ag0dKtmW3GFSt6tvp2NaTdieW98FIaz248va5ZW5jz
1vSb6Gt30mmgW7IyQVLqtQEcuV+p1crBDbq9ejltsVyC3jy1/Bnwu6mD8cIx7i6MmDkkNoPOGf7X
7yoQrFeNp/FSjL8Rr3jXKLM9FzuwwTnFO9rHkCo78ZcqnYrPw/GxB7HEK0+Mi3pChxQXr9nXoIHR
xvngoPJHCmoZ8xyqCu+ztsk5YRq9ady24br7HlImjicegZJ+K4QlCyTyNJLSQK/W+pmpgmOgzOC3
dZdu4cYJLmznomx5QuMcr4JZGEcn1Frj3G30+2kqyShmze9jnbgLhPsc2XX7JaZ3VxC+6t0qBkyq
yRyKw8/6Nb+IVhVdhBuPcRzQtasRY9B3C10H4Pb1jgnSfU36JKpLF4J8jMRnuxPInU67eVqMngeQ
SBdFKjuE2x4MZoc+0HiXD9k2c6M+hKMCMz5R5BOKmhrq1khrCgz7bBzpSPy+3Lsi7RweFHNGzBEe
WdBEDSYztB1jSiz+aPtGZH5Wcm6BcqUWWBVjmAdebFe6v/slEC1svxWeipwgZqAYoG2M1x1f5Hs/
M+jY/5dke7RzCRfyYQ7Gfe5fymh5+nsUNfLS9cKgbkB6fvtmDJRg1GL7kI/zxP7w7Nlnr4jWYfqf
ke8/PjMy1F/YG3mXmbLguFUxZVJcuRiR6vByCClHGgzF+M1v8Fa5GTCdDFHQE+39q2bvJioUY2O6
Wc0XArIJgXYi6i1dow0Oat383UWMg9VXYQaUvOXIKlFOdRj95/hseUzgnOiuUbc9UtQKSH9JhmGt
eGiG61wAoWRty5l4mi8vB4utcPQieB3MUJuDCF0zUjkzJ8d0kIZdEKEFokc+5B8OfnYoryrIfSJE
jUyl+uP7VCSnyCN8Xaqu/jTD06Jb+RsbexTb/0jIVa4LIt4OYngCJenwiWKYOFmbxeimmImzhK/M
4+3IJwYhVH5fo5Pupz5kljv67rM8bM59Mj+In/Vo4BYD14mTVJi5JL8qFq4X8k2XQUnZCRjVThOY
Pr4z9TJW4DsmejiPj0oeoA0phfiw9Rpt+ftefMeSFQUW86UxbD1TZwi8yRc1rWjlVocCHJqSYOrf
hPhdL92t3vv0jNS2XYOOufbl6I+DMa8aTPXB3K9nCf2nVepq+qkZ+jce9cjyPed89KjQswdHQ6Zh
l7KKC/jL6rFbPNNEBhMU1PYqNYExS2mQ762wZ5NAS72xR7NBt9J3OjAoMVQ7daqOARYLkdakxUVo
06/+MmbRJFNxSx7ni94iXHrDZL8PSpJRWpVL/+Ch70yL9B+RhcDeML7zGWbAbTKsNceDIBBWbKm/
9nSEZ5Guoeadgls2xeEAZrxa5ombQi6zjUgiGjpedHHcTHCqj4SgV5//RDoeVw8KAHHYk9KP48s9
JFTkSzAocZghpi3PInzw1g4xYyF22XuZQyoGFnB1dXpGTNCpspNJRig8OARRncwyuHz5ugDUesYZ
GIc8bp1RFBakbpd2POl0bfUnLMpLiVtVcqX5qGXcS5rVYIXCWglDgxu105wjcFi8Ice5zbucich7
7+ykWFOBKrvToxcicLQf9iEYMYgmOPGZiMvb4Vy6yEO9ix9/WFJ2NdDkXy4p0OLIloSP4Dhx5UZS
bItdURJJG4vPPu9JCEJ884bHtJivYoAdZ2nIocRixsX7VCMtAhn8I4dM6orN3xdTD9Q7yhR0eSKf
cygoGuOTbVjfOQi925c9QGyxLHanOPqIkNLoLL6SptgT6M/vEE/jOGK9+o2wJ1NZyG/h5VWePD7b
rlU/QYWFwfqHWwNm4BTFztX5LPbn4yFCNf9etYFcXYkS+/3vrRN5859ZXEKEKXuudfHX36mGPM9A
3nCQHGohOaNv+XzlQGPnzG2fUOrIy86F9WeniY1BfbJgdJOqSbIkblIHvRy6b3UOS0tcOA0GYD2K
7y8IV27rOGMloeySD1qVvBRzbPDavpRe56TeNp7RR123OVzO9XbVFoKhp/dPOz4e0THUMSeMoQTC
jYdoptDxHYJa+qvX5D0MPlIUdGgodbfCGvabl+kZIDr+U5FrPZxpcadV4DeB5dt1MTr4uw5QlfRs
FoxN3ybKv5JlXaW6Hrdi+8ioSMe2Wgy9GzNoL7qaKXSyXVQvK5ur5028WrE45xNUcxKoKijd4PH2
rUs3zagXCgZwDAK4HDxmlSMG9AfpAeJxXOD5TOXLFY2uHHUNv4MbHxKu2e0jUMlNlXczmdbF8gpa
7QsH+RUgvGFPgStCrhYCNixfaiQ983vAXG6RWEYPgpkOoleMLQ0jGMand1n1abiQV/RJSxOU8sz5
Evf+z6CZBHNIyBaTu3F4y+ojgY6LTXVqyZ5Bxcrf/B/tuEE9M5jqBIQjv9UcNC+MsPwlcKrP7aGB
aGn2xjBsUmW/LkTi1qQ6xngrdQSIcTu7PBNqU48FzjNxRx9fnwqxR6JmBQvgji0dDbYqwmIFhVEC
ZXtNrmbrwIrdOU+wmNy2va+kJFZ0dzFRfJQWjZKu8XslU+VxfDwLhhaWUsfI1ZYnSTgyFQ7YF2iN
U3xhJNy1lwJLfvITSBqWj6+XxIn2HUxT3pvGtKd+tWBercx+/LxF5HetT2J0shDSOr6FLLVQaUbc
U7/xirH52m2y03oHHP/lEn9K5sRshZe0t8xdCxJBAbl04nd6O2g9TkoJfb3hPre60353SVYj4HDw
PFOfE/uXcJHV0AP6J4C+b0MhAlpmtUZH33ndPFSk3dBgbBk6zEfy+G212JB/XkKc4cfTBhE0mVS5
SAmDKlUhQBqqzzT/CoIlMFFoF5TObddnG4XfcXu8QizOKRhgeI3Eem2YGh3x8mqYInoP6i49hCVl
t8L2ybQKzyBcnFvPdAdSWLNxy2ZJJpzGv6m2PY3BE8WNH3P21pY4jS0L+tO+SqYmzBASnRMYxs3A
MzgtgSIWfo79yQIZU+OLR2kI5vfvePw7vrHu/a2zbmp5c925ZLNKAkaNfKntrQX9I5LND7Y2ajCE
qr+kp5QtQ52eeUFj811+ppfIXD+cKx0CHexe4EzwQKJpjrrYKD1s1MDmJRrVIIEHeh7R0eM6eSR9
WEe9jwUou4HkorDvpBXl36/BwpDmyVNzFJYwDTOsWFUdnq2nY5fvT/gztQ88ZQv9OMp5aXJ42UUk
EuJvpPoOREUAsaeEoJ2Cjvy/jxFdh6ovgx4qvBi4xPHxlTV42I1Oqar0cmlD06jF4+qC1f8Mzy6I
hZUTvWfJ9g/8HGET8vTBInHeGkpIJw7pgqO7qda2DmeZ5rnNlsl08Qmsyx+DLPv/MmrfjifvmHuO
V+6dfwxHbhQW1ABCPrXJz+QbJNzE6aGm+OiDLqg9IC8ozsUEhegs2d10X7isLV1F+VL2pRZBU8c4
d+rWTyYCUoXpHjgcQES2TlzK6gfU8uTFFcmpVqRPB2Q06dHQWLVb56/ZqTng0u6l+hrm9xMAH+FZ
Eee3ipPFAQA0rMLeDcAQXAxMsQPEcnc0drjJfFT/Fspp2CankNRzYM46rWJae+Fi6NiDJI9E0Efa
2gQxt3Re2EsdDILMgRa/7Zg4DNCG7+mOSEKVMYl1cY/m7rhyrgOvfE3dwX9XhCKFCmKaFAfcQ1CI
h2mCrT8H+UcUCxILmTTF6kZiHTbXQExNW6f2H9sJ0uiAFOP09YuoTWrVjGbe7hyeooztDyEl461j
jkwhU/lvMa6mgmriXNrUpOCNVOy4NGNawiJQfWz6dSuSd8vlL2MdAEnc6S2J4S6EFEuBt/uUU1NJ
SZGaGjK9eNQcYenVcWOSp1mD+IyUyORueZhZpcDSTVGpkQm0bTuRcQTyxVBsjfCe8p2iMS/RaM5G
xdr1FVuB//nq5DXdH6OBWL7lU4YhJ+aGo39hndrHonVGgoTpcZah46XZEd27ZJWWAkAoO2zKlJwl
mxwa0wXNPsNpIa8AVhHbMHzNmZW1HUjfiufDp2WkL+0jno6uQWTCc1gNb2z23hnAnrn+RWdTb52p
ajc9P7MbBdBLVwYA0IhWhpC45JqWyl7iEI00GGhhgTOxcowiurbPq8FADTY7m5ersh2fyJxuIywe
IP9GOhMY7tNvGBgAKKXyFr+ZphjZGe3hxBpwOlAktFlx7CFEs/BJmkPWyGBUxafYBvyzw1iVIoBu
+U+q2Pr0z0oZc8juSSGV86P8NL9FkDZR2PXyu9YaJMEI/0zX8YpdH2EHreRUneAEnmJ825Y+eBjd
IOLFq5/mRIlB1FdaCt/vnF0VdyjXZDaYzm/FmO2fm4TRsTJZkQiS60J5vPOAt19IlHoAXHJ/b7k1
kO1ydBYf4r9LCw3Gaof/e2ReiOKmOo9q1gj87ZPOuH0J3iexxrZfYsVuwdgWkHw4cKVVVzwszv9W
fakQASxsoYYxDkpA7lBHktB5tfu4YP5rofQLKf08M4prso6erMBx5jQHZKvVGR3EZDNJVpnNq6nP
VTtVzbOolnoEpVY8YQZtwCsuMjd0I4vJ2+CehYgVXAvf4AMFZKB3fSI9jsPnFd3Oj3LPBh3WnVTk
F6Ud1ZmYo1K5NNLsiUvCxvArHX0xulFxjKTI78cVoo1ICz06XGdmF/eeZfi1CcFse9/dNZ1Hyr4E
9yIITyRyA+x26HlPdidzgp45VRvq5zTbBhzAj7TTqXpFMxnMW6kJmzGt+Iwr6G9D0MkO3Yp6aCcg
V48/FKNxdKbVlFe1P0g71MyzjxR9iksVxrtzylMylP/cHwWwpOJk1wy4ng2T+vIqvo9CJJUkF5HS
n/IPNrQ127zDXIRARxcD0QMzbeBv2/eCpQfWsWwW3lxRwZspgFPGkQUfPYbDrBNG80ov+NIRhpLj
6Gf5gdVCH1jhUFDZjtI5dxwH8OVkqrRGqg5gI6yYH5Uh1kkseBmqCGnkq0bkvuVz/QRDmLcnS4bY
ZEmaH8xyeg6fukLGnyucVZWDvxzdkXLF4FiWGpeaEWgjLpu9jGz/PM9RmFqgUs4DjfxZqsDc27H4
PcuocVSef46O4+jjtgTfVPU3mH9/bL3Ch4vKIXHeuwHse5stReQkRxTi1czDEwaq0eaTt6gz6pzW
z269VruXt1Y7vtLP04mZDWkqU0VXbz6exaSOr5RcqNz2Q+pj0lkyKXjEOYeahd2ixEzkc2Eji0ZL
90ooR8syhTLe30YsO77jqQcLDFnEgq+qIVudbRCrzmrmhiqwcw/e8sJKkWY9v/aBmoYdi1tlyfig
efYOwLFmoMePVvbXaH94GJndqqVUzKmLcwq3LqbtNFPuRR/YhExrSwJURmCIY0ZIl9Nut++lTejH
q+DSDnKdCDUd0rI2Z9nK/umWjye7AqRLpfQ6cbpI/fwymheUhApIktkxJDx2N35HZ/xRS7gKNLZW
O8PXx1jgm/lbKweiL37WkQFtlAgM1mrOSlAaviIYs+sG5DsS2r6bidZL6ro9Z9CycG8+fVQDXbEi
ryH0RG0xriUEfzFMC/WhUsh42IptuUzTiKY9TeMVpSIeLrzH4IXk88YoKc6BdWRr3RfwmSfC0Erv
EqUynNQ+qsmlJvzt9t2QnWP4xjYpxIhbx5cB1AX+EKy3W4EPD+qh9BJHHl6Ikp0X942nJd9h0zr1
ZN2mIDwSsG01bWTYrTqd/Euev+X/yvCnQ3gTlrNCqFLR4B2YrU01SsfvlFTWKHfAKk0hG5WH67FI
43suU3KLhpWF2HsD3l/VHdWgC2ChWk4ffNwd3C4f/cHnXIgfkBnGS8uFd/rX+hPl2wiXl2wNyz3W
k4dNdTE7uaRjaqz2Nif2+cx7VJhU4IY0dPWE7RG5zBhad4E6JEEziziqmBd6kXUeMC3aFIsBy+bl
LpPN/XUBxhO6BfIZDFiH1Jr6QSJNFCmTTJL7TYbr3Nmk7iGPqnQdPC8HSZvut0RUOWR4aQ2pv3jb
thQwf0R2c8JIp7lVbeqxH1NHmG9/QFrpgP2UbD2+HMoeqM5Wybp6ZPGaf5utrmf6FqLSQ2jFlRti
W8bfPbFP7nF1vfh5aC9pPHb6FfSgdeXVmeAhKMD6UHqLj9qiTvRVNb0H0folTYOorhf56Ql7j17b
w1QVs1MWFe8x+Odtb2DuTuKSfgn1i612eW/inXgkgWBU6O2Kii0yxvGygxXG6DhuUAQucz//Cxsx
5UcTmUChpS/omjLWEBQN5q2Sn/Np+yUs4GUnsK7wotlmdt8W4mLmQPNM6Svt8luQh+nO0iBy73l+
MOQhmoJR0yXQ12S5YhNCHGsVoYQr9fk4WjTJEe7/7EEmA5tKSDEzqrV7PVErd/gS/5raP2RGcbkG
HwNrY7oYkCsACqX5lS7VsabmURxYpob6E7f1MlKTAMMxTBKzlfkR20JNTH1BF39X+0Jd48ybWhjl
VCWj6Bp5XwcjS4CTy2FHljgQgdyjwLMt3lwUAgkUDSMn8EnfMJzSuQCNa+FAz8LccNhHBcJOhMlS
rJVCcAtX6XIEUvXm2uIPwoALBm8YokS2dOWbS6OX5Ribfn7/QKh7kcBbguxAAyFJZMECAW1QMcE+
BUjoripsnfa2WXRQjDv5irbJXV02RQ0klxy3YNW+sxxls/SY5R5IROUFKrRgv5jI7Tkopn2tSdg/
q8L4I/N1WDRZuQCfXAWZ4EG43I4B/pz34AD+k9OQ6YHBMASjVhHslzpkFL3s3ngv7de93CXUT3g+
cqUlV34+X4JlW7lXVmrZNiK6PlZgui6vrcBGZN7hb41gdWHRo2/poI9mg4sZhAmFvtmOp8Hx8F23
Qy4hX1mXfmXZQaWJHU3dqE6igeg33GX0OueotnVW65KDK1/BR4CwWRMy5HSZFT1aW94ReeyP0gl8
idkgagvyhPgjl+w05WP7eJ0yTfLoLTsGuzD6SM7s5i5PBMw3g5D8XJVCv26CbGKTlEqFeUs9WhTN
F3PzLqvGYu0b9++0jJWBBvLRZL0sNryihNY/VyK8aL7s2Zfud6/+KGNKYaY/mOULy5w54G2mCspo
VyNn4ZyPPhYBAarUmhXYqTi+UHgX8Q2vHTBqxMil8dGpHc/s7HLlXh5lY7kr8NALitF6Qx0T4Uh3
+7WJXuskYXlIvBOgZ8GZZ8qJNXb2Xe/o9D12syqGu9A05jZaNRX6yeNTD/RRDidJpLUB+byKIstW
JhTgHmiomY0Sl9nDWJcH0I+jfAztWP7xbprbyAoQP4nZR8Qh1A0dcQUiXG5vSjVCL/mAPxvbbNx+
1wJrL0HTGYacVyI7VR/FXQZTiyTzGscFhvxODVmpR042x1QFlVxf/zuR9TOYhPnQRAvppecMr15u
++v/KXrPNDqvwnkOp3eRFAAZSTcxMZRtwBDVG/d5hEWRkzcXXLHObIoZoil0/QqXM3947yHQ740I
JJYRJ4koi2u4uZmB4yQ5w2qfQQMnMu04GuLpFcXhyXQqCWvsFU9qnyeb6zUGUVLQNq68xOG0NLS5
K5fWEzhG4WDDVl+GtRRJvQPx+/mqLUqNqBDe2BIXAzZB8178RmUvFzi1ypZNj3RjaJsRAW4BstWj
KImVBGoitHs/d2uKULZ6OcWjnA2Xnf3bGM07aYmCaVl1h6MX7f8RaK12UlT3R1fM3WKFPq2DsUKK
CmBNpEYoge0T46Wop4zPdnlksUKp8yzH508qIyd4VrwLvy7rp4z8ooqCPh5/hYnaBMzuTBZdVhFS
3WPGM2CmXw7SnwZU/0k7XzNPT9390PXZ12105/It4dgnRpeTsW2EnXpxBKSkXg60g7CmBzGK16Yp
RSm9bXZ2XB6wUBY9VVUZhBWHjDe/VfJ+YnG1EDZC+4Uvc/uLh9XqtaATTMy3SZUoxFR5D4feFir1
lHbPsoh75w8MK72fz18c4jvrvtaswWcHM6ekT/XKuvTZw3hX7Jmo/7k46M+3bgM1Lq1hD/de5PpG
Byby8m6HJkLUvkpIolRmiemLj/v+IcJ7nzPZlzgKLPpVPExNlzev57aB5DcHgrtZxfZmVU9cvt/H
eK0OMoUexEsOAeDvobG+gngWMS3TrL9vUcv14TDZ022ouP/33JVbFSlGg16zLSlJSU6hwgE/Elx+
TfV0zle3/slNdmxKnL6MwOC1zIlLwS4fhNCdd2wOZdDqmFUa/41d06oDsdfNKRJbZzEQ5fM81gf7
fFCDOLya82EISemgXQGLBvo+dNTczH4RV6oWtP6bQVyRdVZNLpj5mPBgAQvBe2Fvxzcifb33hNFn
Juwo4Mn2DmA8g2xDDv+q5DmFgIr5WDESRTFmderQIqHYUihT5dpVNwEbW1FYxQeg5ITecS2XiMt1
yqNtjzd/WRDe4JjUqh2q0b3nhDdFK5qSV6fl7G27q/fzDw6cUvC/vF7V4P50MDoYjyxcTQw9Z7NM
0SIvCQIxWy5KrTSiwYxl878H52O11op3KTZd7xzWv8PN57GyS/P56Z57HcyBykfyogrXkRG9fUiB
clYRq0RGhAo69s+R5Lo1rliuomhkS3N24p+jXNDnFs5OHapW2Ysze/p2MN3Vq8beH7XIt9Pk7EZT
Z3HK6EbERtbycsnlrnp9c9lUbsekL246A/12PtInezNnnKwWv5es0n7XwQhsjXvrUVH/KSr8NjD7
4pIc/9pIb8Gl1q7qc7n0eQZSz/e1AxcKeME/DmEUqTxqXx/fOhwK8nfi1t6+yxtJiPMUyXivzePX
I0T14FPIMmZYg9xVVrgyiBwnDuvCZNxwKFwo//gq3JNe1196sSxlpJCMhk6sGO/B2HUEmsZLIRvh
9g2pYW7r/11Dh9u7TdkIZcJr7XVGq9ZgzTwjDuGTtie5b1xlHvFx5HZCZiOnM2W/8BJnjaVWTagi
c1xvonMQ0PiG9QsX1A+eC4E3i+OgrxaNlEvWOzGqA7E+eYAPeedNKppuXVsI6gKkK8U3kF0eech3
XjJnhNuwkD1pXvPqwZXo09TQdYIM6QcDjxrmIlMVq/jCvt2TPYhaWNy16kiNaWZJfAHrDbJeUdhq
yFcmVK40utWnxnmKZVbf5oLwYRa3400SD/vh3D0uYWpQMS38hMUo8y44dvA341tIEqZfPREr5Sgi
XxnsSY962aHWWMCQtmfmWdg4BDoa6HIzLrdB8lpSlGEowtsUhpwoSdOPxAc3UblMf97UzqqMxaon
S+fPgr/2oejHX717NL+rHLM4McmY4DpFi8NMCm+QWiOb2QXWWNXHumShqtzj9qe8JiOF50sKxSD6
y++12fRoB+WnfLVe8G/3EV1tf5Bw0huancav5r5FZaiCoScP6LrYO2V4iokAQmjTMzu/K7mOrsGD
/KTX8ZEU7elIPEmiVRzR6oJvyUs/5wW/TlnvO/Z7SwhcfLyzlc0aAHHscOoXbN+ojEORMjPoKicm
5AW3eTssO8Rz453/uG8e03yB4v8f6wkwFtH5VIi7zlHb68XEY+SEWU43B3fys0I4c5ZOe0iBzQF/
T1sQfXGv9Sa/KvioLSrNzjLepg0JrAQqZ0GkjTFTNBJTGGKF/GxkKNvTg1xmhi5iLzOOPVuXxH4L
vNZxT3n9vF/pQtgTFK/Tkw9iUApFVQjEByegPfcrhULhSlPgM/KylyubAaNbAkZ/MgAiKPAIZkk0
h+ZQdlDsHbBdNXrCH7AAdXiLdnIGJHoF2Wj4nFesdwucGTg+36pzIsf6bv4oiig1UsP14VpQv+pQ
rnxyzqZM/aOfd6nt12rfPFWRs0Jd+sSy2YB3HaWHt1qm4WwI7eN4Ud0VDqi1plp9nq7HbkhjV/2m
b+lPFiefn/tG8jZb1v9o0qbcd0yF7mn7G8FcEk+BOSBSauxR88IGLChLxllnewiTCoCFArxCTp6+
uztgu0cq2Le+Fl895cwwlchnsapvYBlJu5nyQy1yVnsBn6H5Yu5Mgu9RJy+aeC/0HMu30IWml67E
VadLw2au25AQQmQczfaCyt1VeX4q2b3o/AIM0AVrflTSkfn1zsAap5c9akVkkDIVZRXIe2htVDGs
tp53YmK8sP2HA8amFDKheNrnk6bh8HNZBoj2U3lhfCoQDwy1EE3w+tdHg/mL/Bs5xSil/oFB7Te4
O8hhmf3YAZ2YG6ddyTxuYhrEHyw8PuNLA7xhZgLKUYbwQzSooVUTiSgMvsthUzqC53osWimf7YZF
QFoOnIrm4mipuCXcYtmi51laC27tBl2S5wmGBrL1kZEbA0aYAkajuA4G1Lg2Bf/3FdAWiiOT7fjy
4L3AnfnyN0EaSBsbkQqzMFtVcYo7UBaoSrhuDEFGyarxTGL1xxk52mALPFIjfG9mRtOWjTqgnejZ
TNiX9YMYfBuCP01d5xanzfMZRjczVFXVxmVG12CqwIuKPupuyNsE5X5BcsDgzFehhdYQ0KBozuSN
LJnz9+ufOVhjbAZMm3g3GAp/wY+Cl8rkaFb3gu2DHsuwoawgPEegxrE1DskZt4QJdvspQ0zl8Ne6
TXmro8RhdS48xLrgzzbjtMwzibi1uqEFGqCfUpnH34Un9u7n80s336npBwE+XMiLvnv7bgh8j06m
rOJZ0c4UvReUP/RKOQnu5geXJDd1bDiqjT+w4DVmkAoL4xSzIIJm2xDexUJdRE0DVfV6+ETUfu0m
wl2f+v2qNxYjoUUApKkhbESrS17sJ7NmZ83Dtg6+l/nxljUGwcHI6gXob6ATdbcp2PGkiaZupTBL
oeLf0kRk7MJWfrxGyGCAvHEEE/d2MY3zezo1nXCHKgbRjr+PMwGrPD8e79qGWg5QlCVoGAwWOLNG
aBLsfFltIzVYAaQvPsmZA9Sd0pEPTCnfjQ+aRlqakOUCkPvvBzRKljJ9wjctptIL+bl+2wmrnkyG
c8JRwjJCPg9D5WIjHtdtlEq7MiM54vVf5/i4jus7fnaNq6XVvxcm3gbLLyOiCwoXtrI4Cl2hqebv
Vr2QyQU6s4DKIbAHx4MO4RC27/oqfGNbS3azKQkY9rwBAskQjg2Q2JPsr2cNLkCFXlOMADMDRnWE
T+yddug7ZZF9kyUz1NnWCHnSvApdoqif9dH4asY+NxNh5CwFff8qA21lXZuRY8DUYCO1+NJYz4dj
mby1b7YUx58ATOgPSsg7VLWUvc3PZqdpg9jl/dNBuTBtjWHKVrDQagOhTDouq/drpg7h7mb2Hglu
tpMNFUSlXIKJYCtnusjJuF4xKFMdorH+qNlz9qMfVIGffsFIZdQ8ADsY00cBX7qdeAeEt8Mu3zqh
u7ulg+inmwTZy7O17IuNwe1CZdbbHPeRS35KQUjQf8N5G2j9DjCrR1Tm+Btz1woU9TYSiltFd1KK
KQln1Kpe4KvNO1zzeQyw6GJ8TOS4ffwXk1rn7ibjUFNPQUh1WkwusFUslsdV56Q4SOSOPbfSlPnF
ihcNe33Q0BC45DslcpAKJq4zoJdEpbi8bsTEiua7QkOczmy71OPeIsj8pk6KBFMY0I2yGyAFtAiy
3YcdnzCU+ilQft5xJ8NUd404kGU+cw99wVDmAwJNAvrUrrmuVUFjVzKRd59iF/C90piAks+F0Aay
WDwc2BnYk8loyIHjfjRlGjQlEUkVlz72ucpgwhKUHDCo/52S4uCtXvI7dfh+41xDPIH+dxYb42kV
RCKk2nVhGkzUCQwApUXiRhRmIbLp9M54Y1KfU4ujMHGKm6FiMVRHKUCgjidW9rBU2TEHh0p48hrA
UYQu1I3rHdK7xdBoM04JFPVl5yZ9UX6Czaya92reGWGbFW5HVKd/mXdBrMU3vZMSJB4OBDfNMxc6
52eflrVTzylwQ8/ugHUF23AmK+LSKsxNRYevfJ7vmoSWbZTDtYlzXfNwj50YbujUOBhoKNjJpwPf
I7WsoE4u5vW6whh9aXReylFYNXO3AMMFr2+70nGxQzi3RJEMgf+ByVvsLNM+AypHMcpp93Ku5ZV3
ap1DZ2jVVWfSTgFABSSh30jqVGb1z4+5zCu4qASsZsNa2X+4B8zBtIA5jSsO8dHI9lgzbAgvKeP+
l7pf/WroYkIieiMaTZJkhbazsVyNQsQD+hBLOEWXi/8J5iuDz/ZrqecG+JpwjPnc+kTW/nOElG/i
3t5aIq6Vl4cjaWM8qR65eNNDVQSax3G+d3BYjqw9mPsWMh4ZLjX+IWV+pcngLIGX2yhTWBTVlEpq
YFJUvaNM6NWHgM/JPm51nYTrTq34NbbL6yp7HAdKgIAL+1yR2tY9r0jLcKQxHM4L66l8OIBDJUk0
todl3DpsLygvwTfRSoxOMtUwBIHL9A3iRWa+gDVFUqEJ1m45YvHp88fRtVRLObgLVRfCo0DZn4in
Nduf59mY8+iWtwlyrKhwmRJx3Hl9T676CslG2p3NAQYHJIwrtDO4YOeIaY4l2n2iOSDNSqxR7/wM
Lb9A0tTqep6SQJCoxGQIeZwoXhFuSl/m/o3Hx4CPec9b8U6Gr2ByY2wyfAC0ezEd+9joOBs9Eljd
KSFuKl5m5t3XUxM/EIM1LRavYHnj8IbNg/Ed35BmbA4LLhWVhd7VTNVS/Mjk2+RdttIGH8ejDnwM
SRBelITf9EUf8wShChBzZZoiF1jUmJfKeAhv89ftKABl1lBwedjPBnIcwhw94Is/YpHJ/uqreua1
dI6Jxa21IVrsp2JmD/i9MrbBbeNNv+RxJ496KG5N2UzSTeNyVd6i0Dx2WkfMpk2Uufp5jOCGdJA5
w+jIp7J8jgx/rnbPlhRu97tfsjsoIUAsfTCedmbmevRIYkhpMy/Ew8sTVNVQSJTV8WYA5A9kFGp1
BC0Jmtko+P2j2oL45HJCZZAKShvtE6AWeyzWbvuf6EOE9D9raTC+cPxO9kcMZ7r/Hrm6sbHWwpXo
Ntss5RqTJ47LiO7Dbml8N6oy1lEWMtwWCbWYDrISLKlHisXHDjjsV53A38h7HKjOLpFxYjAMV3kf
e21y5ZI66kDjQXtGOI7OQXISkUpZXGnx8HypqlEdHQRdGo4EP7AO6inMdCNvFB4LoksLXz8XGC4C
PvvBDTYR86b0YEF/+U4xdveueOgOjtIjGqleyUFBDTVY+NSTQeHJjtncUD9FvN0lquDtubjuNHsG
fli1brKMfiTy+H17kDBeX/7RGyD1Al+51C+cL8V0CwVL8DB+WHzpGj3N0Kn8HVVlF2hjB7GrONWJ
ubVwPqwbLgEjRInW+xjiywnwzzDz4NCUO8Axi+YEVYhHchf4FFXdkxclCJGpDhvXTtW3DBOpty6d
xfQXF7hRgqmTXO+IFP1We9JNY0hQ1fIX+/9/989eWF48yggNmkxECp7JfHGQyIBM7qzdzMvdmfID
96umzcLcZM6f+VBSaDHljOq5T4p4E2teZez0Ou90Z24U9lC6wJ+3C2kurrpPew23ar9VSvr1/Z3V
HiECpEksPfDdIIDOYg54tsF5bpwxW+ll7JwTajjvoxxoH9HeUt49wNJc+VPfnh0FgCxhkttQTNJs
Pnznuh3za4BAJs3u91QVG33bvnaC1y43FACbj3yeSRYmtDt51u/k/yVRqdPBmlIHJsrcG7gmJ0wQ
6y8hXpwSqWhkCi4ISemHZso8AV9oWUkDmZNF4eS07CgDObVJ8IiVhvXK8IsvA78Py8eUTkI1CauZ
/n57lHYIy6nGl7nG0X8WlZiEKgFiSPVzvrCkh7xju+lJrR3YPfPC9pD4csM1oUowhbs3ABrU7AYn
WWET3QNuOFzfc9d1xjFb5hDYQ8L7ZpvnBCRESsdqwZA59IF3woPkfOkPxh/V8WXfFB/nW4EBVLtq
gVdXRKU11ZbIqjQvHzq1vmi7+7nWpMMANAiZpajoz9WflDR3tFfF9fAq1nbeKJy19ifYwMdfNJRT
rfwYV0tW52MszwsF0GiMWM9vvel71ky7cN1dCztomAk9E74/3EUURJ80sMdVkerK/wnPPOdTt8xX
e6zJFqoQo1EE/a7rftoJkDPkhEt1qQ463dW2JKClGWZJfj0Svkiko9GO4WUFhjy6elj6BdpwSGU3
rG3OCej3URShuYabLYTwFmi9o0ietwFV6miMl+EEQuHUwuh4890VjpbFjhfL9CnNokuaPwr25Yrk
9OQBFmg2qbjQDXHCYT2RG4XWORXUfF+jVAwUXoeq/eoPtKn5QDDrxnNDdl3ARTQoJBVbp7ilri/S
Blvyy0La9t94XMeTEaXzZ07t6D4FWXf7AODwvskAVUIYeiYSdE0KFy7ryCCYtsChZ7eL4U18YrYX
/SbtD5URE5UyW2b1Aw+caOHjOKKCP9EBHv0uvUamTsHNaCld2nZiQHKZZ2nRCSpFV+a50S14hBJw
riTEgH2Dd9Q4/tpdq/pk4rUHUeDURFY1nVQbgZsimtj2vW38uq+0Viiv4RZgVPhq/gPRuUiRYZFe
Z02nuJKERKGlmMgI3jvfzotVbECOqLXqIJ32nkTqUaS547etxNh8ubcIE2dhLv2JzkXob4kFrJRt
yti7dsEBE/nK0foX5fX/h1w86i3VDnobyqRPFJcBoB67rLT5ZH51N1pq9UXSQZ4FkjR0Kg5ySz8n
6I9tlHIzyBt90V/KeCRyc8+BWtNUR8yoMVjTvaEfnyFiAv+Gj1SQ1+FO0itVtxzOQXd1umlGnV1X
qmnyX+Dt62JedwoIIyojAu5wNRPRtEbHEV/6oc/97l0p9tcU8qasO+tu6bEoUAKiCwyxESuf9NEu
+wfABgbW9KuLGRv/fwHFmXpFUzAHkeR2l/+3VBsHCUoZPwx4+J1bqIuyOKIp4v4DDmrgdyJwiTw9
CulB2lSTkKtcbgnWMQ+hHyDv29akTT5PhMhQIEcs0WZmnAb0Kln4yNq5AQOBRz4sWpB4GoXCUZ7K
7thu0PRCOKPl6UbffbhIAlryHXiHyEP62uV6RgKlysCnaiIsZCFHXEnd6QuLCdtRcxxVeB5ffQSN
tvmIrULQn+SitYXD0q6vtSualSw0rJZIC+MOXttgpJaJLVOdOMKS0cUyzXN6mTxAIAarGyTtmYnb
hup1lbnTjwHKMcEvQNPWZISzck2KA/h5AQ9tjrFGRN+c6W7s0dMpEMzgLuZraa//eAF726Bty/rK
/qjkop+8aMy2usbDrPSs2mRN4u+iseWps1Ww4e/LwsUj8BwLPOZja0aGI4p3IAgnHm20+m5CqRLY
A964WGxIhpVQa7bgK6U51ExDapptVYkUZ0m6XYWym/98YnnA6ou9Tfo4iskaZ6OrdgpycqL1gx2c
N62wr6Rpkyf6QgChbQr8WNzkTxQqdVOzsco6OQqv3Up7d4VeUeClkkDqNuVDjKft5XDrS6MoPkJZ
+OG5+2yko/FoWnQYY++wDijpu+JtvjH5c5IMy/L93slmS9C5btTaKVNtLcroSTUOTRzkYJZE+MLT
WLgoMiApVaTypXhcQ4oiijU2MLY04a9LeSoNWBYKON0iRAsJsmeK3mpyo1w62xVyTcQjJARPNNnD
ZRCsXVPqRChM9jNvTaMb7VYCZcepsbCQAnEZ6mj+M7QHpg3B27/zpmJNpg1PO1dYFpsaIjXFFTK1
Nxkef892WEK45OGwVw2S5Un9g0kbm23XPZ58fnxy+ivrVdrIta6m1O8mK4luWGzj/PCU4EJSdTgC
KI+IuOHJjGeRw7hNlMaq7LrAoqSSsF+fSPJ0bkJLp5nxsYiJIJK9AR7R3UquEbijcus37bhsEXcl
AjEDRjM7H/o0XtK6lBMbMNvVvauwCtpbZ8QtyJEG4ynKWvlXRXy8Qta4XsGUoHfDGmfvnbO4PKV/
zijfRHmUI+6tv07RoxgHcNdZMt/rlCrPZtiluGiigDmxZE3H7WKrrsvvXfhCG06ro7GqxRDb9cRs
C6U0p1HHEuznm6BiSBLVF+MDC0eT9SkmVmAsEpv4zKq/jt0LcTxvMxZVRj7+VgwlOsyMFcT778uE
J10aAlsh6/anjVMDevaCe4klDWcg0D4xpYAdXtcHbZdrcmBksYI67PSlInwSVFmGI9IlggmQi8gw
zrH304z20o/SYKE/CKzHEK96aeLTSOL9p5N38qJB/f6ZLvpmipDMxyodalBY39ZAIsjn3fvTH9/n
4iRPzPpCYv8CF75/4Cw14u0nukW/NOaGc2rH6nEZzR8rNDr0nwW1Yj5wI8jTwZkBfj/Fh1jAlFxn
kjlF/UQ1BpgRQmx1OhEYrKl9JaAvjde3pEZT0AUWCuXwPsqbqjA5CdjEwbISZOQ+uZbHiZ79Qm0X
eF48r6LzilFouDrMIthPZHH4TCiv3IQn3q0V3l8TvTccnKJp4jG6J5Oye2kYY6XP4ZdWqi5Q3Q0o
msCgARWgvyn6wa3rGF4XHlZRBDr42QNl3RB3atr/dSJxY68DMi3HupYEJ5MJej4eYhz/35c3ByX5
Wpm9m+qzA6ACyjvxDCQmKV3KmSZU76OD7N0osCrM2DoPEBQVF8T+2LYB3qtrLevsCusdu8dagD6f
l3IulR3Qnpvdz/mtgp8B7NtJ4d6TO5/dps87pg4AMkNa/3ikYO1Hz0GxH+fgb0YCkwixhCTHSR+1
IyszQPRTKguaezfn+9A6e/tqiDycJ1p+DrHeYRc891wXrTI76kuEfk1jSOLwxotlj77UvDCdmMfB
smA+3sZz6ArutNEKysub0/X6gj1nLvYn/3EpvXZL1/V6RfN7hJBMGiaLV5zyT8s13tDvueQYVBb8
uujZqSoETyXZecwFzcmCanE/YkLgjYK09XvtxUQmewea4iccL/HuJAsEzyqfov+QcBNeaj8JUUfW
wEvX0SGRysIV4eYsnfIOB47qUeDxZbdpz3ACSv2g28znLcbBiLlh4Ri5ewAOwIgFxaVxbM+WjK3y
DLRDaQrBTHNFqi2W7hfc0fv7HxOQ9xAO7RSS9Ga0zCcB0RrM8+uw8fm1apNVsEpYXNnAdzWgdeoW
f1xdCiciDKVApGkmxVZbFSoLA4qbxHBXXdjLo/d4adew8jfdCoJkUcbgJMNzGXoHP3QVhRhamwo5
iJoPbbLZApF1dOuk2BnUu2gtqglmUxhB7VPXiIoYmhqbBJs0m3gKKfy8xSmqW7qG+JbXpEYR+tIR
Rsu5Z4Ib2P3Wn5oT9tz9eUuaKCcAKttLHcN2R+Hf6MzJu8wAaQKWPJz+QNUAcUdTM/roLpk6kJBc
UMb6CyPICLGwa6zj7nG3iT2O72/bsF9RihlPu/4nSciVPrUf7fx6ECYoNvsvJJvP1hMnL0c0nQQp
3m5yn2IFq4shGOhnP7IAUWoPJVzKwuf3YAH7IJNPPNjuGCjrjmVhJLorJFBYWXozhHlUmEd85Jgq
WZMUMbLmIoW5tcjR4QWHtec6WjFCSHUaO0vVlcRDd6POWRR5EMZmsuEHzmUns8euyu+p6qVE4gMs
1nggdMtckJ6JauOOlc7MpcSc7tQ7UPForIrHQI20VGsLGEjrHh7qGXxd8ogYsjypFWfZ997EDjKU
YZZgMh7akXHnpcAVDkLAUooQq3aHHTdpr6N9+OMkfofXtV6SS7WBFD6ltzayqnJWD7+rP1osENfO
a/sGIbSAqPPALPWelUWxrcYrxPNuVUh7nZ8bHxveO/lR/8cB8Wr2BNGc0NKa//IFtojEnCl9XVBy
00Reca2UcHow7kkoSRqw2gEUpLjADcgwA8kniUdP/d/HpwglmLRhqK6N0dxOLvj/I/GHOAuAGqwn
cY0/E7R4BaFD0lf/I2lvm1ncW+1j370Sg/51pt0ptlxwJSgB7HvZp+wZ7l76zPvZzXT1wVvYD+ak
4uObIq6HedEQuvwSBcFu3aScUKiUTwdl7duh+orupnTgYNcO4dgI0AA8xW1oFDIVl2iwdz5Qaxs+
CYEJeCatDSpUR/WFXUsw7hP/wAEFixhyBb6c+N/GEpONC+AxKiLXxBrjxCEEQTuPlYCDMriAgLEE
Ag4UjFS32sqOhDbB7KirSfmxy7Q7VLuuZ2L/nnffn15A5JJUEYTJiQn2MVLZLa9VbvG5FP0YrrTf
BjhBLLzkpf4+z+qBegc0MJPySuBoCMeTM60JPYyC3WWXAjxjzrgqrwmc3hJQj15atYFx9C9QtM3M
gHdudLJ/EHoRvZ6IweASsDEVCxJ/oxZbOsA/LyjN1OVp3TLRXAZkPsQYCxzN0WgCLhD3usnw90ld
RFE1qoXXgQib8DRKcChfMwa29kIPVUx9pwpZMYWX2i9MbWehORS4qNiYhJorDcqL2rXBVXzpCWl6
YcvOkeuJ9Ycv6fvQIQmCAc90Xb9S1z/fEt+7/tZ3QylkKxGLN+qI1DXbGoDQnk0B8C1l9OK7QJi2
s//spFyDu18X5ypaW+Yav87K2j6YUgs1GiX+42wvLwkIj2MKkr+63ZbtAywN98lvfmllDgwKohUo
u5tvT4IMUEIuan9kyCjAgjOWXm/FKhDPL0orPTPVHIKZi7S2z6B9KoLm/QB4BEvAqJP+B/l/ssd+
emgLRBYQJpXwwpW0YQBnSSUhhhUticxDMMj9Sa6xM+uqhafOgpeQpKsNKDRBD3MsfUQEAfATpKFy
4UogaE1wJXNfXirsRTqvMLcV2lEHpuHmK2jUlkSZQ62ZNzb5T1jA1IXHURDh1JPmI38GoHM2Z3Kx
4mfucqXPlEmVAYX791gi2zKM52EV4IFoo2yP/onEc7Vkh8dI6RJvSNyJMoFaM8ipvwMG26Lefea9
wvJFf3tmri39sHaSe9vqqjnWh5JQ1UOzknMQ+JAqqrO+5pGNgFvGhhduPw2a+5jOJsiIstY3xkJt
8vfETDdZI0N4JkRps4y4bg37RBXRIhXhkBNNECyf/Y3aS+76PvbW+XbWO19cJsyzwROWCVaDjNCG
6kSD3EJysPUkY/51OjOVLCXKsvwe33k5kCHSCo2aFFsyg3d0UHRfMZwyJnDC/Fqabi03/5D2Kdti
fORrmXBDtnfJBNvt+pBmXID1E1IHI+5vt7CMOQjcOC85Sae+g2gmSK7JsbykZw4qVB4cnI5g3Tvg
6xxnyU8LQxOAaG84K52RKJRxDH1Mhu8790OSLCkAJ9nHI6VArgI+1Ac8UvOm5N/noIoKLQ3vltTC
oY0+5zJb7zZ0wgdh5/937fI85GzyuHzwYZet10a6KoFqgglAmb9B6iEqm8o1jNG6vN0QT83DD410
aEM+38pxfxuEWUrXmQ79xwMV6UpzLJp7vRUeeSe3lQf5NToxNAaOeUkN8XQMkC4PVremldrBjZP/
qX/IABIPHjdxEgb3HCRW7wEYDIkjH4aVFKOymcHqNBUrsUdsJqWxyva6nYsDu3+X37u/y8eI9q19
MDfLZDW8XAAl6m45grMLPJ9/jA46woUBlfpja/SZ30n83VJlnFBCTE/uL00cAoukWxakOZmuNFvN
wfYVmUY4kMtg/qXV8eR+GLCpVAcfUtEd9GAYJJs0vuZaed6V0sIm6ZHQ2U5iX3Jdy0qzcMR2jMLn
DO9dcg8bqn3uW+3i/437S6CJbw/yjTiHMP2HczOZrHiesBotrpZ0DgJ+9/QhFQzscF3JjgKva0zl
ymKw/OzeqFprHbkDVCgjZpU7J9cRUbLGSWqr8H01g5JczbNT2uaxLago6NylYe1IQa1e1eO8mrMw
grrN8hM6H6EckwjOACaQxJ6M6LMWUD2kBZUMVqOaA7Nz/2Vwx5tgOtXH8VBvX0+iYs8WWkoC3K0J
WU5/6lOWNApCXgkbQZiYcAPkW/hjsDZKT5whVxAwLZTvbrpLmg80ArlnvWuxnBMSz+Kl/96syuk8
pOtcs0DnJtx7TZGns+IAQJW0Vhk6l6Pn00bQuvyhniYOh7RjI3JuHkVnlkgRQN1DSSFXB+ub+hyO
4b2gUHRrZ6BSO0Ve2Krw35z28uyC2h9t/0JxwolYauFhI+acO1OtzTzzm7u0BEc2L6IU0PWQrLdU
epLbXN0Of9o3ILKCI2Gtn29llIP4KujogDw4Tv4mFEMVn+2KjGnOdgokXJm5PjZLBpJvTd4O3izc
VvSIsU5BGGaANal/V0FYXKnV0hmO+E/ldPXzjhQ2ZeOvBuy2gM059fdstthN7scnx2EFckLi8afF
LVU54NqpUD9V/fY3F8IpViseYgrVs/PoVKIxrGCBYYm6k+37n1krGkOwJCbV7GiTVW/CWn2tyJs5
CSzfoE3kJMWyCZdQn9CVorfuHhTlF9HK2w5LzMKz5MoZX5KHyxJ8dKBDmwQdQF7yb0L24tX5OmIY
FSnF432BSgdlzbKyf5LcWoxrPF1LwCLhoQ0d+jSjGPEhbffd0OAXOjP+OCTa8jvClEj4VAwhviYg
RJxvPgswEznJWLFG0sDLedMkxzmaQ9KBdtqgIcTLfDoLHD1w0DxXPs8Yb+mQT4BVEp+CzKmiTiES
CN/KOVqAJxoGLBWaZ2A9WJGHFn9MScZJE7yhGyRgddloF5yxZuXSP7W2Vyh04oP3q6ZSdu1NV513
mZPYX1zcJiiT5H24EIu60y68wGMuRGtUuUs6+Ei4dNltKl/4dsu/3qqDDOeE1yRMt/9zxNmcxvfP
09HFY3/SKU+fvKLLmQqLiN5KEfrDbJ5mJ89QZyAEHRlzxuznNvz4jCiSxqxna2CYZXjKrkLGkYsC
WOcPY00mzjn8BqsB64TSTsACSbKQORfrSr6PermdAv3D1+BBqph61V/LpKReOVfywaxXuoZ/LSCY
6lUDa1nwFZ10SQpg3iIL8Bketklzl24I7NcB4lFw3TXLi5afZyu02z0htyNRAI13JCXX4pykslS2
pit1DiGUEyyaxbDqePNbw3TPt7+M1ifB3gdMB5cgSfj850B3tBEsIwmQAuugU7ndBZkdZ21NIZLc
iigSkQPVBZnYOpddv+hPg0OybfixG1xqGLQm94LmAWBpHIbYETt26Gyjj3g1dGmLZ6VvZPvrg9il
31CszmI85Bnp1SoJeZrxG7Y+CcMqdSUrsz8BDtCvcCW3ep+/XQytmprxq6+/hgvfxPr/wdrrMAyW
kmKYahaSar9mgDJMtBsa1R0MLuJAGngZq0XTUA9p3+VPj9irL8AhV2ZzVK7MuuqnEEHIHDnhJn0/
GzEZVV5v07soBsAnxS5KYk0DoOwc5uaA6Fp6V+Kf6L6UWtyG6k5R+rsWfM0i9rXkv0UDStFp86DM
+sTbWSXu7UNNMyBYZLMVzTa2k4TMOjpuX+lZyxhDH40RDwWkFUMLIwraXinxVmtbud++hy0KaV1A
5mTL9RwuzR7pxiNCyxXLSIWYeYz0dFC0rZjhNz/eIEfB9U0ye3lHhvwS3nubG6N9t6MWtjxyiP8h
4rxZltxEkI25K8OOXMOWMszGDtO3usKsSxMMNo2VTGfUTRS0UT7VHDZyPQsCuVJt5QpBlwr05mUo
A2XU0eETyGFJt1Q9doEWC25MMrGGuq9QtwG/3e1kN5uKonttf78Qg6LPdthOwZZxfsx9sqF7Y/5V
2gRjoXMsS+iwDGW+2P3czvsGT3lATfAmPCEYicJp1eRncTxjsBTVjYhnu4sD/K5mHsA8RyuV0T+6
pjp9NanADYBnNC3vczY7PYvZhzdh3hAQurmgus9es4LihjtW+vi9+aXEaQVoU40YXkVaoHz3Bp/O
v/kW6ejQOBdOqUtvyTdPyoKd3nAAjaUEFSHk2geJSO6e4RH85w2rJ0HjEp80JsCZ68Y6FIH30wRB
NSaZ9tmMCU1VDwkneF2jdr2MWmH7V4VrOe2qH0tBir5njfE+fYYxU9DrHUplijef0rRokWYkhixx
e/GrVgpl8xIZFBiqCwwkEqDXkIWhc6t5PznE0s30jeh6kUbuqZkNN9yHYn0+g7ErxiMmFH1QZlvO
t5RK9JDGlJN8DQoZBRbzCu391AvNKssHGbn//YkRM3unzkXIiDneUGIGJNQ/XTNvBP64S3RrGV1R
zbhZMYEAPiIdOHUw0NUsIYdKTSwzRCi7L057aL2Lp7nCIr5UhmUdhEFU46P2obu/GxRgZvqS4t7p
nWJEpJSI0zyIk3MApsHMND4T9OgHIQSrQ6C7SmMz80PLUeAKhyvA+poNGaEFj8GqXzLUu+Zg+w9m
qo4yrp1mHXll9fjYjS/NadhZ6gZih4LRkmkZT6tZ2bh+kgzyXPUThx6LW07Vy3OJw/fSLmd1qE8o
IEW18B5YZn4EJh6u7ajUV+ORQvOF1SoPboiUE13vLwHNhxNgQyUhe/PT4aWyfNX4Jkwkk3ez5aGg
2IG8Q3L4FPBuxVR+fEBNLM3ZqEcEH4OnGULEvyLuNh5vk7iW06M0YT0813vMOOdOjpNah1v+HoTU
gPi4fqLc5orEAAng0D/V0bvZibKkE9bhGv7rsYErUEAHR3P4guyObC7d3x5wlsPZtusSP7Tc4ZIk
ZVT9RILZcxkGn2Z3mmXYRmjZgTznjidQjLWXjtlxvCC+XHK/kZj+NnRCfOeee9+GRfcv1IJDHSk+
YGGSv+kuNJgg/5SnOk9Ae07w3GqUoR3VD0OkDyYm/0K7el3tUnsU53C/T8P87h3FqtqX0S06dtWX
PC+v+15qavCEXQ8faZcK+zsYmb7N9OttbvEq3Iv5IxbkIbsIWN/aRSY8/u/CE5f58Bdgx3RqlF5Z
1eIzXWSFhfypxLvKUCRqG84qaPkOmJ8Ef5J7FeWhfIqxtY+29CWEgeCBks7bxWAfoxx9RwBkAv+J
FqTaEq2hXuC94v2dYZV3cRhvJnJ/14V1NZCRmSvCSdSn+4sMdl1bQXKr+00q5VI8jFDu8X2CEVCq
klWeANF+sZDvhlNMBovhXuQBRTQDPeK4kc2G/c0MmA1Wc/5BCC6Kold5vx9Xeu2BOnLFfGqBDcyy
TGsnwvAKZDhximfg7FJlUVADBIRM6keQm5JG1jjqaUQW7CeRcDLk9BlzRDubVNM5rBwysItcat3A
xeCk0ot8Ld5A0Xh/jl2vRbLLt85nIY9ylv32pR8/qTvDg3PY8uBvZIG4FhZaZ+xHypcZAildFu9h
LW1xpQRBYRbQKnhBftU0SNAv8VjXTbuD3dFg7eh4uhgVnXRFMlyZQkldWeEGgiBHR9SJ6mPzGdy5
wu3HecrIDw7RToAq8OSH998nMzvIqSvGST6zOu4s9b3ud27VsxFYE+sbHjJri5y6fIiPi4EVblV9
CX8ZwLqB+nCCEWTCi9W4Ah1OopfWdgHgwMfQkpl+DEVzlUxTlZjAFMJMYM/kMRUzFWy9Ij2vo0WK
4WW1IIzM3fl0jazjpTbNjYOZu6jp8Q7fAIFC0gtyKchZK+EpVNx7fn1Fqg5/30LtmWWUgdqgediw
fbD8eC4bZVYRLOorPc925znKvO/w1aDYjIHEqg/gPYT4zBhucfEp5CO1eOWcIBo4oZaG7N259EpU
uD+vM3Jz6HPy2NTs/bAflHlTjv0Pni9bJNb8OxUAchtnkO59G9MJkw9L59dl5PVLi43oAMLoNkG3
qX+8njpPXnGahTQqj8JEj2K/yDogrtgzEEkpwHaF/DGuQW/BmEtvi454knX3C236eVT1u08iIKjG
NySiyEbYWod8YYouXwCD5KxRDcEfelT+MV2q/a1Ni/5hcXGb5d9TFuoR+PRKFLvARypv6qNg9h5D
qmdm2SwfqwDmLPLz+kDK8pf+q6ESBa/sPTXT0QfxpdieccJO4nSQpx0mFB5jzRQqaagfcbti3Wql
KBJX8qVsspZhlmDs8PlSSBSN94oBlYNcF1O2ok6BjLk2cRPoeka3UcBArnlVpjZkzOzmfrfmJ9IR
I3mfc5YxNELS1Ova4eSuFuPVSWB7fy9ACZL/W26AEtAKL+8PePZJI4GsMx2RT8PvckeVma1dZHKW
2X1JPrbDhHYdBXiiCAJVnbq5fo4YecVbANGyRiAnk+IaDz5JsjOZGktx9ltRv42vC4ZYLabhF2xG
RgQ0T/TO23nNY5MVGz6Eb4GhQ7MLSW05xLUh1Sj/3J/+bjEXpq92ys8OCvrEC4SF3Koun6iiv1CH
4exszXeOt2gaPWsEUc31tixpOOiu6kjQ26uGZDhsOylzVonUN8U2BRpkgVD015La0JFUCxNCmoUd
fpm5QS+i8n5SNmZbP8epcVddibM5+XzKiGch9imTonjNRNYeQOwQKXPca3T57JLBAt1mubZtuXcs
w6o8ZL5UTbljtUJx3CbdIxByg0HaXuu4SAy5nVfdcoI1uvM+zCv7x1vVscrj+6FpXzfEGHNVsx0u
8dpr6cCcKP5N8T2e7UXYb9SlXSzUkzMgEubveB/FhrxaLsMQUsoD8XVyYSfNo54WqazBotuhoKR+
20IC0Wof+Y2urR5ntwZG9EYHAI3u+ldUPt7J+e4W55JmSZl06CvOnhvQoAnu6qu3IwqiVG81ykjz
X9uf/PVhPLNKx5Xp5Dnwbf5aYMS8KI5oMb6IyWNwnYtXhSZr01QDIboxZ9Qh6Fqk7XIv7wCwH+2V
93RUtV8RmdFSBztlRkVko9bkUByTwxbYfImHRuSIy8QpZaejHDeQhVuiiVzY18NwSVhCBU3NT4/Z
gzeS9lFdiNHVYuvVPVGKHrDLH8kvqcnFHUFixTjslWZoHk5LVwwnfUBbkGIyl2ZFf38N1QUXB/Tn
u813UacsF67X7qoeXqIReAsJcjXcfbIiLD0qkaJVDcuBiusLPViah9GMxzxKMk/Wv5yWNOkyjb4R
H1ljgiGti0gr+OLfaLyHAzUHZBFsA5JXH6q8l6LTJxABiB39opduFHA9TMCZNUVumkKyJ5CKvnAY
pJlH/0FRLvolqEPStMnFceR3oWegibCVjSpTIx17ETgoHRY7Ywm83EYDqWdfv06y6DO4KlH7bAIO
91p71rfFhMJnabPz1b/u57bE4XOZLt0Ul7CCnDcVFM96mq3iCSkEbsJgEaNORcoy2em54yx7Lu76
/OB1zmxj0b/tjg6p/zCRsHH+Nd2qmpO0L2Z5EMSAS3JVAXkLcA+y2tFEFFs3tPnY6OrrKmbXVWyU
LMPwjAtBMw74rezw60GNl72/WKBErQU7MBf4gq0Ro+Dyv4Q4awCD9vCfGpL48S4gYbT1HUTKLXyU
lrTUIkS0CH/da0P8KS3U0O2jLEI6kzfCU04tmB62/hjYtBsvLzc/NZQzhXnTwmAQmFM/cge0KdMV
KdUE1aLENTK6bX+ecWys0qKbJGMCJufcU+oflVXjQwR4OheT+CZkyRsnVakxXy/1IOLfrNtw0lH8
uUElVD2/J/hGvzYRX0y4m7Fc0fh38tlnutSx6j7K4CqtA11j/xLrIJKlYeoGRL4Jg9B+ltpSbZys
GGLd2ERdJGeCdcIuvhmgq1DaKWzcN/WwJbz3gOthyX8EhGhnrxf272nQ2ZLyELLgECfsX7AUkJmI
cv6wJ9EJhxveiqNA9K4Fej5SnJXNR5l8ySY6E5hOLOluC2bBhWeqM0Lkr52KVF36MU+inKP/288f
jxiVQSYlCSgVhocSMjqqNZ84/+SjLPwPbmlGeWCDLZXgEgRP8POZehvuuE7ws9t5xwBG9dSPD0Hi
7m2wgVxrIzyhD3AtaYFQBf03rJe2Vo0ktDvjxENgTdGlxrF4gWwLcgl6Dx9PaoxClxHdXlU8Mmb3
THlzb7MuKRsdCb6UED0LrzJgd9X017j/IrWWgmcyafRvzdkDLGjCjyrUaNkR8ZJs5DMAdNTS56X2
SA2Ef9uFyGYeKyxeqR6/9r4rodzM1wI6L0RE6E3a/SZV4oDEIxagXuZqPUg6XEHKTM/z5nsZPcz5
sLwr3sRfR5FnyVovtoCffCzkcbfhR+oqsL+3sdpDf302JsO0O7BGG6tBEGqiKQBLLlYJr6+QehhF
MimJ8J+aWsKfZ3cmgCn5uuH1GZIjp+OpPKCkBD11VQzons9Gd5QWgvGLc24Zyrea1HinBkFGj4wz
0LqogjWaz8a2WuhLoK22X7c6tayYGKkqF3c8Hq/AsbMShHTpsrwR+5Xz2RIy2xnc9jv4iPO1dSRj
OVEIhhAr/BcToK/l9HbCjQHbyTuKenXdb+HFr3IcbE+XE5qj8HuG9a/+oI4kHh6IAkXbrSjxJ7k3
UfaL11Nb594eAgZQWhGX/ataUAskrVu5a6Ctyd45zjhv9jBLi32hovIPGZTPobTbwnJpm5CQixrc
YEBcCfslQPsGSbiB7Kb1HKQBXZrd2l0ANUz4rdagYGVjENn1b4vJWO+eh6P9aiOja6DsJPNKIKmR
PWG40ucw2vHWm3iiUFvwb0GWPodhpzdTBtPEDF93s7n8jH3ee81FlBP98TDIMSrKPthhfm60MtrT
ZsYOctHBklAAMLzpnIfscMp16mDXudTL6T2UD+3nxYxR010uIdXAMoojWMYfuQfHJ8IJoJ8gCrV5
OTTrdUlKA0TdOV+x+B5/Y/LrNLMGShWPySWKgFdfCZoAjSxuyxf1NwGAwb7fFiVL1s6R8WtTsOj9
WSVKznYk6J2N4xd0lYcvBrKtwN1pPXaGhq1rQRh/lIVd7M6kGyabcyPRuGMHXCvyoXTkrdHXm3i/
hj2gcXGY3OkRUbgxmulMXb18LUMmTmka2QMlonOjvYNOi1ekRUDw1K9RPLHcvYZLvT3n7cxBK6/q
H28gPbHTE6EvO1P+O9QjxbRV7uIYoDlsIQ8rvlI7t+dchxvrtFhR619PUu4BvaOWBueS/RT55JLs
QB7Sm1YcD6oZEcPbxqHJrCnWA21GUcTz4INIjQW5C0BCU9RBM4Uu+y0z9C7uQPFEYPF9pO8LaBXx
T0Pg6SCTrh3AJC6PqaqHCE1NyoxdhTXydFEFn5hf25DQ8Ms4EZQN3+F4BF1j7HoxISGiOuzt650O
dKtgxGViL9NGULEv4MFoSe80JjhTvc52EBgfc7sjCuo6Ck+SSd/PBQLiMbckg7+AAP09pNOwQqz3
ur24lnVv1O924aUnmDotJ0CshkCCVwlX7+GiJU0I0J5Shfx9p6By2NrqDFnFfo2xza+NLTjc3gV6
YSe93c++LlWh7DzcQ6kh/AvN1eSNL2YsZEKRsGbP7X/bYQrIc3JNt4Wwok30q1IU9p/QTQ9Mv4CR
Gy4dwBahIeJurtinmaVs+Cf18CvypnB4/rtsjgohUv8lGz5+5LfJs8hLd+KMPNuMDiXWB58dYo9F
0V+CKHVRrD3GsAwVj2Mss/TXoRzD4qnFeBqXJS3IN1uKwJ6EqUxWX5yAcSrgr1+1tkMhR3UT5sqS
94MSGZxhSikrNvsjW2QPjr/06La8ArFBq71bsU+6CUrFAdcRDUCAsl5RQ8URFryN4/pV00eOcyfb
3LO6BgT0jY7BvbK4hM50i+XpH8NBgQGCE4sbV5x+NDGE11GAFnfCUCx1aI/ejiqQbCU6nfUDZahN
ByWeYC9fvUj9LkM9GI3BO4dYpJn5cTs5ik0mMZuwdMfA4VX9NbE70j0QFtknUuVy4UmjQkfLvvrg
GF6BKedJ3d5JM8SOa31lNP1R7MiAaaD4yGbAe6X4brar6lATbxl481zMMOH4NfIzsQBbE4yC0y+e
LNJmsnjk/XahHFqtwV4FL8KIz4Ilv+7af65BVloNQzYkpYPJA/rtL/dys75vYBFnjgOQ7cycCwUF
8K7wkJ7kqpsTVfknmLtGJczZ/Yf/36rxpaItD1unWSvyN+duxqNFIDRBRLVQPFLQe8Hzm8X22nIh
KwdFlqRiSqCBQuAiIqvpYkzn+hf+OIgJmux4JHFzTjwMFuLd+rl5KrkYqk4a397VROtkZUu8yPvy
T17kGuWtgNb+1VF/m7nWr8no90i3ulrYGJF4It6xxbf/c2kXIz594xkK/qvWOLlKg5rdvQQbGb5s
mMoWtHybYzgCbeYdKWbu37DXSU+crgNA+LMIyGC7ajrVfZDW4Qc0qIytU++muUxhltg6V6LiyebG
bab0hLGXaI26hZJBzKWPJgxNeRa/mzegkbDWhDJZWqSaYeoEiabUS0F0wFmzLS08Rk69K/+a24Pn
xlsH7pCRImNWuDrWFMgl3MAHJU4WKsuYLx3D8jVDQM6FVFY4lnAp2Ocirwsq4WgkXY08OY5boNYI
WdwL8Z24U5Od6AnPWmx/zdn5zQRmDuC1Bu28vEAntFME72wfZSVVWEpFRO739tbOGwC31LHGybE3
XU+mURDKtUGt/MhROFSIPn7bgYoVSPTHz49WOeWNfwBfX5TAQdpBxoj1yz5SZv/oNthQUnBiFxcP
yi21LWqn5T926m92QWkFNAucTefVTohH2uB9ng/a/1pQuHJCRwI2u1W1xopAUT2yP98ES0bKQLBd
y3P11k2RS88a71izzbtrNjoHZwjYCqyi5Zk3PNIh5cryC3gLDep2cpb6cJWhrsaHf1GHKATeIov9
YdjgMtEkTt2xlA7bOW5lcLP/CYkTtRUMCdGZXFhHqjzG+JkLNkOD7VrtKWkPT1hTSrWfd5hvsT+q
EWm/Cy8w+vGfAaVY/snfDBDPS9DovZps5NJ/6fv2lvR3s4Jvg9a2paqcdtTof+05TFHw/ooXUx//
xQPgXnZKp8jF9JhmjgEjB91/P4oiULbX4qYe/PO86ClvFJxtZkvrCBPZ23Nbu7sSKFzvDbkCF8bG
ko0QLW0U1uwqW3UbeG8nSi/rKjH0oH/BNE3DOTpOyHupFX5uoEAMXD9J/su+YmWASLRVYeXWYN9E
Jk97wKQAF7hR5I35854TJc6S4cH+w5CaGfei8+49B7DnzoTyubZnK9eGbkkcb67yhips7ou6qh2c
j3ktK3GQmYpqNpQDSLNMsiuwQemQ4wxzYkdXt8vQ1lpqUNt2bH/5h14qHDnaKsaAkzXkrGGN1jUt
Of0Aezy5wmFZELUtrxetpBg+acb6surYX2k8n3lJUbHaTxONhwUHbOq5da6vfIdSCKwGWiAmmgC9
o96PWizlEHeg3xb+mgf1onxoIr3jpmz3XFtsuovQ+vKf0eeMFDvCAv9zKpD6zZREb8TnqWBx7UMi
IvT1BHO6/wWszPbOuN2t3tn5ShxJOHs0YmqJ89/rLbGwMGqcoeIomPDHV0zs08bDsOqXDU/w2+Qn
OO7Pci1pZ+5Y8U8QfzKUHNLTUs/u3XAt/0lrlLmlrXpEMaWtKI0stF0BaYeIb41f4clkpGbWjSDb
z9+QpHxh6q5Yn/vGznaaJH/F+CUY5z83vbs6uFkDg1hreW7WzrHrhABWzy5oyG8qxoJh6i708gEy
D44afeZAH01I1sH/4S89sBVxzEt7slGvYyTyd0IZw7vwwf7wqIP/PBziQymYZZxXSTo47VrhbXUg
gb0FMEdJXmcXjabgM0SBfGldGc++5dr139aCugthzl+W3Xp2N6n8UF1ZQgCg7ZGN2dl5FIknZWCj
TcMte+/NVcxlJJk8QNFJufguGOBXmAj6t3Iia34cPNZEbJtnB9kVtGhIcUewvy9fMMKWZRlZsVOk
Ol09NSDSdxmR/VBejNLMCT6ZusLKtlKpaQTnMib91QIpY90OijmNdcVP6OMnaE1BaA+pSi+gEBtq
eikoPlVqzAbObUvZwLXdxC56lUPS9pJhU0tflHvc3P5MRmtsZKj1AqzznWGHhTO/bhNOqwRWMtD7
REIHo28J6sf+VV4MKL87b74w8QeM134oDamWGy1ilCxWhCvPPKWdb3C+yBB0cVez4kKaNKeHJDhw
TMfmRUOqK0Yhp+GrPEvqscxca84P+8BHg554QxqDlbO7MbuvIsTQ+z83oIlZLtJzP0mDSMQ6fx2W
QL75IWyIcJK6tU/G6VMxHkchr9451uacGUQHUtVn2DY5Ep+07jO621mE3AeeJHLe2mfWTiKWvvxa
1JeInj5W8uBAGxVE6w3ar0zxM2wkDMSXI0B6xW/pxMeV4JRiDcSjAuoQg8CiW1a5uoQuL9nBQ1s9
+mkKHfglykp5Lpo4tBIFLXPTfaqE8nOm43avLH3m0Tp8YPlrpTf89TyZhN25mMNvULktEsReHZw4
eGP7PjKre1JCeFsckllWDwvf7QrVe2Ku97zWcjVDsscCyS6Vjp6Fm7I2AAnzuW5BSyZo6lRvSdA+
d6jdo+B2eXKIaCsoB3mxOhR2TcbgesMKW7AJYeBMDi0O7PHAyDHp9EKRN8uAWekiSRg8a7G6lSpW
gzOMFYZgJgh38lvosTTkZkWhD01B6JeEdRRaU3DJeXjbCPJcMZYFZZ4Om5qFYxKdfRzaIA5iHjMB
yIcScKlOi+fn+Vk+bknrkat9+hutSPjOzpkWl1nDyqBSeu6QeVe/5x6Pslk1uM0Xs0YziUP4z4zx
3ECOdfn89ShXc9wRIV33erDYeTnic0ycxqU7/ZQPvr5RP6eQK16XnyacRZkE1fI5cqXWebKRwzh6
oWVlHnR7pua+E50Yx9+KSohHLG8rYO1IBXoYDJ8sQ9SYJmUXVksrjyU+bOHRXRILDDDShqadOtqF
FFCj8EbUuW3NXlgskWH7rQrKY2xqg1vqTPhb49CBHT1CJDB2AI8+sWx4D0aRUjyXxbsX6iUz7oHT
9gjELqCbs9ONfUGwuvFReIhcqeNXhkLZV03D5MqA6nVvVEaNsbobgjvcnJfk7pcw/nZcp6i5ehmo
uYbhKMFDDZ73gTPnW8qRRmWSMTGg+HsHlmJCTwNrG4tPGk/sJxDtn6hmP8s3+tQ8260hWLHv+N/w
tVQkJU2gzzdTSsqgAHEK3g+FZ94wjBAxrfk0mzua7OW/mhNM73aLhRWs3QoIA1aCvAWQh/oXy0sJ
hfd1p/JfD8x2ePV4gKtfsvFMb8obLMJy3bqgPSMyc1utPQCp3pFWBKWgq8cy/tcyv5OHa78ZDTnA
j3ujv1V+PMjsZjkpZJIWo9oJCOKEShS/Q7l41Y5VZAtDSN0arvrcaqD29Xsu1lJQ45dY/n47ljZA
aS8TzXCT9h295IC9kp+YFtw9puQG+KErQ933XgopiRWHhGpt4IxxfyxNoVgx713KPErgEJ8wg6N3
e+HowAHaWMMos8IcnSrRFc6gZYzk8IHAA7qzWQ6pNnd+l39UJW364U/U2L+ae/KmoHg3nY/kcY0l
YkFCSeejCk0fY16Q6ZWyIHis3k7dQAqZbf+jQy+nDRpZD0hrkAnEEoaG4Iy+nqnFIpLwF2KFev+1
ruNWxVj8xD8XFF80cLvimSPUSVKOT8HEatLZmWqzBsRhabI8aeiSgwWQ9kB22Zs4NIPRiz6WWF8s
oRRXmHn3vAOC+V4Ys+NSmzQDT4MXsA3qX5dUoYgsWUOKnkalpLvA8Ubb/o7/YTTytRDughvsAgNl
DYsqUo6Z6JhoC4+Xq7NkXTcBOPo0QLJyISQZhEzAAs2V5qAudfUyV6AvM625xN/3PbUGrUMq7lvT
l3c8AezrfSICR6B45yWMKpX+swROXT2sPR8lNuES43I821eklZOUbrUAWS9hpfAUMAjv/xZ+ihCp
sfiOsim/pex3ea4fVidYOkcbfbY9s+BNPf60+zuYovObdkkQbhn1DdMx4DG7oE7HLnMUlDtLCmlW
08R/oKy+D5mlHFQC648BFZZnl4HlOCYSAK23kWfhiqBkuu7bEAODXFxZ8yBNzxyYjPVOpuKk9pgd
b5rFU8O3yY+puXBGJfQSUlOmxosZ/GAj5bGR3wBAjLHwACWtcxVoLNLDUSkzqIRbEpJYG1BOXN3m
sE/JZTltJ67IxgNjMFJ2/KS/2WdoiGGvKjHAvf2NdoyYjPSIw1MrzuuQPeIWmHjqxxYtsph+vgNE
7uT6eGuAtm1zeN7VMHwFgiZetOyg3w+kXXkRHV2Fj1Km8BZDD0ilrp5FiXRCLyBXmhJo6MLW/ojo
5q/G5VTFXZL+0RmtdDP+hUMF0vPj6BStqY+DXgvnmqu/SS7joE3lHzmdQZMRoOX0hAbgHAvDed9Q
kgAzFW1vxyCWUKvv/AtB+M/MmC4wVRYpm9wa9a/+Mn6HtsQjMePukGgvDiYKjKVRzNVLUJic5z9p
grJl9pTpn7DDlS0d4kxmujDZLzRt8DsVwrlwMOx/levOHpO5Dcli1cRiZ3OPiUZxRWvqRSs6OdMw
efBctW84ZZNqNx+FAdXenFQMDEBk9kOz2PuOe6Gc1sS9kyXtnV4r6MBmS87dLnl7LA9xhU41OqY3
aXVa2nLoAg77H68+nLsnnt1u5DEOgQewd/7c0ZuXOxJUZwfL2buzQMuhgXtm2a7R9jnHy3Q/A3Us
JN4OjSviIz8zlIxNIWUEKejVMrAUZtoL4TIogCwbAmU59MUkcdw53WkBU1RaKiOvFcCG4CtCr922
7Zx+bzkyYhRCHojsSJNGtKQ35cWrKIRAaTL2cCgqjYqkN/HXn5vpuCXZ/71qED9XqX1qW4bUSAxt
YU/4UZ+lIRDIiNV5HDji5I5TICyF/7MonAO1Dm4DMf2+E30Q81FOi5zdpmZL6yGNRDS7gsxj/bV0
X47g848XvWRJrnXglIgEhfBBcbmZj8EuICEkqLsrvrl957jErOQzzB/OGLSfXsJ9p55SLUM0NV3h
YevXMpPz3Psg6FB/tBf8eK3YHuz5OhM+NZJSCKJhWOVreieUL4JxSM1Q8/LLqoU6iQ0q/Fp3m2RZ
wIXQ3a/kmKhcM9MjFLGvB4wkvWti32MLv5gBcP6ZPTxiEJ4dIkVhsn5cYd070g7atsIqdHXze2eG
b43arF1JTzzQsiaYdi3YyiExwJIPolrP0GFoS6meyxg+5bjHD1J0JhKvcfGQJi0vEyIyKhZVB4XN
l0cUu+lbQpTSXMZnfLPDNMPTB8nc7KRKQg6Q2q1WKDjADg03aHjFfBZrHfQ7lHYsLfuOGPw7jhcH
MGxz/yu/1BoIzDB82tiNNOgmQX19AMvZkVk4hdVZkkEQyjqNyyHmYEyMm4qeCKyWrT6kM9Tqy9XP
KClAlXXYL3vd9lkRIZX/99A1XqSfDr3flvlEwtdFeVDamwb4GhgYIIjoFO6cdkB71M67DabZz8KZ
Z6Dfw3LY9eMm/rQC86LLO5OXwuIIZl10dOYQdpZIDhxTCaQMptJMoKw5J/Q26tqME6wl92qt8kHr
nXcNBzNYvQtf/jqHJ0KawGjLQ0N8x84jSjezXhp3cpyzK0Rl2OQoKPppPIOvaPYEQE1sytc4vgCy
QdHr1QKqEGQkN9X+t8cUG20stIfJjlnFc2mo+vsR3m9Z8SHIav4dUZ91JwuHD/vOSNzJA8POaICj
YPEQvHHmdAfko1gA1tmVp/RfQB2k3W3v8SbiR2tRrHwAXUogQb27Iuw+mbjPpxVAlTf+F7wyuxvl
chw6rUrU5WoLKynm3vzhPMKg/zDgehW0DeBw5E/FKbuto52QHgRrvpACT9UmWlJPf5ljdYNbNEMC
sFuQNIQmwpb/yOXjr1zIzmlRoJsGJygCSaAILreYryIFvc+PCObwZY1vaUajHPzgfaiYkZT7mBXA
yJHpMvmhC6V5XUA/2GSt/AzfFNVvxjsEsueyAFRpd4GCxhc5/YYWTZXk13k3uNQ3MSz2ZH1djdjK
A6iNeK4AAi/dKYQ7qeceErsEuvpNV6qsBZqLRXGzEe1U4kEMlVooTr70tPCXo6X1cFSdk8H4ozvI
F7/xNhBiykcGPFTpI3hbPY41Oys+E2pXoLaS5js0ZozPw0W3zcKMUDqPminz+wropibsmytswU4r
tuZ8pQbYTn6yW2ud9zMQlUAASI7rJ9fGNg/lrDfJtfX7lXgd3HeTp7VKqmfoUdwlN1fsay0qcfit
IvHRlBwHLJ/OSvMcBsV3vtrCZr8gXD8bKXp8cmEAh183uhcHukrTlgHueFxGO/+ITfw9ygvx237Q
25XmAq3a1aBJ8s4Dx0PYq5ZPBP+aHVzbYX1croW0/rSN7ajm8SABmjW7nzSbc4uOQ6OVauXHpftY
Vm0XWlMrsalJi4VRA2pX/jEDkcCVO5sZT0GPSLhlIP/26d9HFNSJXOwO/vRNKI9gB+c+gkxAmpgJ
c/xXuotOyryQRvrEpox51vVnBetrznbBH5LHTQBlb2uZTWDDZbJyF9acYemp22kGQYX/a5nSjpyW
q1HN6rgdIXrpkUmKJ55M9YTWx8rJagn/qUluEwkNQVVTQfCL0YZb17ZMQIccAJ73uVKEfiWagdys
wjALxIQhUcAPFQQib9eEKf+rJ+DA+7v4Iimlhmb9DL5xKhC1OhCLlog/mpyNpirj6tXu3jH01pz2
kxHfAyhxgNHlQN8ZRBs0sWjBymS5n5JJVgiWBj4Sa+hjHTp2s45apAHCzALn5OaJc83dxsYUdwH1
MfmdlGdF3JmW6vEPzo2yWa907EcnuzwvZ+BETWRLNxYqrnqlVi71PUA1v+vHDZ5bC0f3eLNAOFQ1
N7y/vOUeSos1xKWRiSEWB+FQFEM5t7egbpz/oh31683AKYPnuuvKzVWPPYQ2FKDX/AO0fj3Na1KV
tg7fJHL9lNZNZYX8WCikq1cKry0hrCsC+xrnll6h65KCXAjol7jf50No1s9LVUQJj+L48v4W5i/z
0/+5nGfkHHx+LUitb77w5t+3yUqlEL5KMS5Zzzb8l2of3ZtY8/wLkjaqH5oUlAfbCVTYaesHC8c8
LKMAVowfuWDz+zJ2W9tXy1tNCcxCJ6A9geYOqi/i9YkV4H/NQSGAv1PLBOfR41SFYL/qpFUzBPka
SHqYwxH7ahnaQE2z5i/qWtaL7Oqvgv4dnmIrxU7LEjfdvM5Ty5suscGq7+xzhIqu5tg8uwUuLPFC
Jzs8EdtNB+OGZOPWp91wl2+378IXIMhoQqRfOx5zRvnUHmfmtk+K6bs3yPSFYIS84Fmh0Nc9KNd4
zs4q7f8Ne5lFWvzDxSI90QuhmHKrPeFeJ+Arj1DQB8LR6SvAf2O9Yqpn/RPepPu5laYu0FAgbbMg
a8M+ABZn+DI3Y1L/T5EiLictAPNQl7YJecaoU+gA/kiHrQo8dKos9FWaUPQVdvLMQQHzeAVN2HhW
JqEn/5vTzJxwzCRHlxTSLDSh7FSClmREqkTfaFfG4nh7KC/oz8ZhMIDS4T8SR6chXMxPAsQXj77n
IXrePeRk4wa5g0d1GtR5E8U7G0GO2vMewvPlFOsevmr3AC1ONeQYZLfxLFBbvpsU5owuX0WfSk+i
JTg91RWOBIZqG5eyu6YnPG0vffOB7/oQPOti9UD3wVFPnYKZ7Psai+7abKM2TmRVh33IoyikMUo0
u/ps1R1fg6+1n+yQPCupi7cnK/ybiuOw3zQCMDtSNa/4P5f30Nef4hH3yAw8E9/6+DkXvIRmauVz
P4sjhagt1Io+AYinFfz+wsSj1Nf86IjWrwFr9XZxqCMT8N5BClFhNiWWyURoySbGFgKIg4pR3V7+
f1oYUGLljNcVPHLMBD/yECeaTdKm+QbhS1hpnmWG4BepS1zO/BQwKfgDvFcRTu7/X4Q5cR5TdiPi
msS22xbsOv9qlBIJx/pudWEu6wFYKrSg3bEO/aIIH8KlR0gWSUUe+o1QhzaldktwwrrU5ovDB3kn
mewKkyCzqUYthBHmm7DTwK58D/b/YTvjDzlCThiMZezAXq03Saalq+1s6oetorWLzRhRGy7AbAjR
k42ByHQNQCWpAr5g76MvXBqoy71aU5sp9tn7mQ5xBmEp4HxJU0OSB9tYsVp+DmgbYhZ+E1WDoUEH
S5mBEIbF7Fai2plM8qPEFV4PlYDi46mMuvTUPkIIWIefr/mbWtPYn2jhen8GQrvCTLWHS6ftJWdy
nn/nWdgH7IySxEfQa93yGYLZ+A1PMTGmsO5iu4o4Kanj3K0akQwa563jB3XxD+HvYZ8UFsaYvXv7
8QYSGbk/3gsGRuQvFerz7hPtki9/jNLgZbA2Xm5Fzx0GL3UDXYCO9r+755bxz5r3QU5mg9BTJ6qz
7XxPNW2++2pmzeBuIGwN0xaBb5ge33zB/KOA1xmDwFU/3Y5ilGZY8aAP2aw2m1mXfIcqd51peVcF
hk+g5Lgo7wk+N2pnUFItSyBMYYU3VSR315o1F78cI0M92p0/yJX4dwI48gH+QQZF0ZYT722bs9Qv
NG0rKRZW48bhJOc9hzNFrFdXGQnxaKUZ69FJfMtQwVgg/Yv1rXQ7qXAMPPjs47Jqk8CaUFU+NDzf
fQt1zBAqOscHWP+WW+gfzmQQte1c3Oez+bbAOt/qxPnrcY5/Q4Duxt6cpVbz57QY3EJV1XaGbRUk
9DIlm0h/s6XPY0yc7DCMJcPv3vu35us14noKLeaA/v+HQwcUJegAik3ghsv8saVUTkqh6STzQ0XT
cV1F4LyHU0xlxWiW1YANZDUtlEycYtfCpO78PxVzTHNUHOYyOKEjH2gTyDEYAhn766SQa8h7qk/j
GnAqs7+TnaNJZFrwr0uBfAjKOvhTqu3q1dgW13O0e4Q3OcmXXgL1FBqYGbn7PW53EP0wKBJcbQkG
IZx1Giy7vCgYIJOJRC9MbkzZgSsZXqytwkXZRu+L9u00Mfwg5GUAlGPKO/jVxTEP0vi0XTuJdpd4
4boENETFXyL26mxpI3HsF8O1dQwdcQsZWxnBy1lzQ83wnvcz9y2/f8MAeKLOuK7oJfQzghVQbTA9
EpDW9IdTlthG8qtRM8ftV3HM0CLwZ+gWr/IfVixOvDVYUDN5zvOQWGPOzojMa96e5nMMduK6DDYk
jIOm6dehbUIQiK+nXrkaV2dB5wMLdJFr1tekUkG8fLoneSmfhpMZvlIfnEzupxmUZISNlRCtJmXX
JsJaTKJ2Rt5TsOJZsVbi7sl9FX1E8A4yYysXAffSg329+Idx/nqQQkMRHyEJIY/CRd1n9vQp5bFr
675PZmlYSuAvGFTTqC0gNkIoc4FkcsLX5aUYI8ZQI6JIXB6t8luhG5pV7OdxfuglHpzWlgzqjnVN
6bt/apHeiZsL34UXfIzoZFkutwl0H5JPJj9fCQBLrEr4zn4dwzuCpb/uAjR56TflfofFvjiYkORL
GP53ww8x88o2k8hypThY4rXe+SpXcWX/9LXM5ubwO0BGHi36itxy7WvouSCmt11XYIkbss+YHozS
R2DkAUQc1HZftkyQ2q3kEYrKUmr6dp7anxEoBvU1XUUwl5J86bIMXM7FR8JIwPjJglVkcF2IhTOc
8UduxcrNzpkMwqPw7UbhzvhWtCxfHAe/dYU5STUg+un6k+ONyCyz6O/PiZ0ImeXXs7byikS22hm2
L8bMnDlR4NJizDAnjQqOnNe7hgEx6LeOa7nDhE/j/AP6qJjV+xAjRgoKQBPN1gCsr+5KY4MqBbRy
zPOGmmQ6YUtY17L8EkPCMtY4LgV39YuHLmoXKlHzjNqF/4gDE1DoFAdvWZouknSfiQBdP2jMFNbI
5Xh6sD5NpihvtnHlVqUrriLYI3CSffgYWDvjr2qTb+JZDJ8AYpBG0EAqDyoKGcSDosFcRpwhfUxa
WOke6nb7ppPCAJ+7G7FJ4XtKoKnTs5NtRs7HlBiA4+2BFmAnKoRqvqr16n7b2a7TLe9fmrrH3mlY
uYF7JTH0pZmaXwKH1KirUEUBsvGpGMnrrzt0Wa0LNwoSFlTMsNc4S2TPV1e6agsZleIWfXf5TG7i
Caaaxa0Fzbp5EFiUvJNDPRoy7i6NTeZDG1cn3Tt5i38YPvAxjSThq103cjz84BU4GM+cOvbY7VUP
oluU7kTpoNKUe3+wS8UUnnJSI5ZRTcSmZNupyN/Pr/SC4owcN56uIa+4PQNeB+9Dj2wVvo6DitL/
+4MbWm1SoILNrKdJkchcv+eLvIHag+F2CkRzNfYkVKJXvCMKQE5H5XChsWlBi4UZizzrrkj5WzSm
jfMQOIHjMPqL+aAg0vZ1fXpGXtddoquOjo3sMwo7u1qiKthnBBTdKx4dhx14lRm2uuLwvl6HVYqm
rS/dkD/WtPOhlWQNE2GkNJCrkLSv/hI3GFKb3T6TvXEjrIyp3bOerWvDDuuXdbkR24t/1GOXLhp2
JxiTNzJwGLWXK/AlXOe4Ne5FXsNfK23XX8UmZ/Y6OfFr4Jdt4iw6GRWUd+gusk2FWQyFyPKvoLu3
wlv4+771fIL0EsaiRYPLl3PoHLe2PZNG8sz5CZDwB6LsTzdPA3M4WRBOGyKTZhq3/Rzu5F3PPy+1
cYxti0AoGSieKtl6v/4J0jBtheq0Ayx9WMLpqrwb2BwtGqiuraZVJuHZprKdDnpFXTwuQfniA/v9
+gx7o5K5eLnnaz1A/uZOvmKJQMhbdbKrG5ajFwiRImfQhZ/Z4uFMpyMuOoWAcZIyZhyxXrkEihja
nu+RSv/SojVbbtgI/Tt5fgUSMIO06w2PJT7qhLkwYVy2PWAkKjHO1KWxu1FhY6ywMcV3MAtDxYTj
iZ0HvewFA004J6ymKuGm1SI6zGLshV9QG8wRcXE+mTN/WGyy5J3ewwJ5Ued+lO1BciEL1hv4oWh4
gnG5m6ZK1GkWhfhHDLl6Fvid9hUBtvC3EnUFyAToQTtncn4tRUONWBJFUtWtckxkcrbLaM4lNIuB
s4cBwM1OXsD5EDvgFZMmU1pJyILtcfKOo5aPLvDSIPHE6YBypxFo8RQSmv7Frrqe4FfzXLUgtcel
887jS96UxsJArxbV/NkqS672XKtbFezVJiJIHKT1elYvBjlmllAbnxlQ7Ya3iitoHVMTzKVfToH5
3ATlg6n/t5rlgARJee9EorYfdg361W8xhX478n9tL38BeVt56W4qzA9kQq+h4eugvuGUbvVqL78n
WXraK7TnpbFAsCgH9rTkTITll/TY758gTGi9GO1xYagU4fGAGv3Yj8wBkrVZBdYy70I0Juk+Kq24
ojwhtxrcZ5aSxkXBv2TODk47s9QQobzm5o3fe2tyYtb9DnLozAIRQCgEoOFbpcum0YPNOHAxcjtU
e4FxSoZpPnTFyruPwWFx1MtWNI0I+9+Ew3g5tlDX1RHxiGwcBk+81v5Trhas+vTwHp7EPkW3LY8l
3zWvxN9KDSfoug7MwsnOslBhGtqkneGyWVXL0ta4YflGORTRBUDHp7Aj/AZLuRIv4DA4nwE1o7rc
Pj02C9sDDpfwY2kAeneb9VZw4VmONoEXEv56FAli+vc1+KQ6SIej9qTB6isDMtHNSaNqGebY8q4E
AjsME4XPaKJYYpejqHdHpDQ/yaMIcc0fuA6ICJEnUcBQ+3rOP4sRtW6wjwALbL1Qgjj0FstooBaK
ZKZDZQexOD8r/xHdQ/yCOvJ/m5GdC+cNhb9nJLjk0wuQrIJ+1tgPkRrF4BeCTfe/4XVGqT4gSTso
+zicFysDHmFBTmIwcpgJ6iN6F2D7cDqWh7DlbLNBIahV23Y2eYXSW4hdSU1ZPMBXFpJB0xBn9jRD
J1/+hC9RLNnAr9k8eqmArZh0HxaVLVVWjGnrUg4Yk6IVnEEKT7gquTzt7W2dZsRCj6ej6biOFsmg
UHl5gbu9/KlPaa1FrBYh4mUgh8P0F1wvFu18TaSZDUS6uP6h8fuSjSRv+W7D46z5zuqRJGNb5zqt
6Pu21T5eSY4iPw7NkzxbcKRua8ROrgZPHNy7pH+O9bmFQbKPqEyVfpjdLlC4GKDeCCibsgEmZU7C
S75ZOM7VX+8JiW1MevzHs6kmJv6U5OaDCLHeqRybNcuJWyQYoatbbtDQVGI5Tvvi2s4R3dlE3kY/
1S8J5P/eGB1PawaMMepHYbanazjtUdspMG1jZX8V7PNarOHyoH8niyXo9Z9zVdjFVF4CtTS+hlc7
muJ+tw/mVf7CDLaR0gQHHeHzrd1SrPTJel8AkoYEf0ZOnlUF3gYpq1zhum804HdGWR+uU98jfS3z
Uc5ape4SQmghnm50oXOd5sRNakNJ/IWd1GiIkQokiJJJpNbc4+yeHm9fMQHRldHD+FFBdrvsUjfP
zcSfancOG9Cybn/0z6903b/hEPAk5tXif0z8+b94D25CuDyL0mqvsWsMiyAW803KuvqPAVXeQAYw
6+K6QyiPOXrx4LxhUialWMyJTdZEFdA+0iYTGK18oqmHD8Fp8WNLTI5edmFXUIdba4sJ4mH/2n2Y
Cyx5xcoCyQPkY2PaxQfez+TCW2jgNiuSECLqrBa1zsVyot1owMnLVgaf0qTxE+pwNa1yJCxRNn9Z
cmKxmlTEq15E4FlXfJebIrZ7A2Mfkyl0vr8ikDfmMKCXtOb8yeHN2vpdYS1NB5m9qHQN+PY8nzyC
o3gmxf3b041xoTRPa/5Y2dcPVy+1XclvgK7Ir4fSrTML1Sb6f6DDyEVgn1uStPH+dtRCCIxME11V
BmenMJ0Oao2mOdwBIiIo3qEa+FiZJdQBJp5bmUP7V5Lkf7XQzsR6OJx5KwN6OPZ5QENArSrlGDbn
Qhs6sqcu/I5Va7a1jW+GCpAjseK2T6dHaKzqsekziWo4K/jq3Y1gUfUeYtI12dVrH7Ubf7qmAtXp
GhR5zhbBtYTGe3E33lO3TKAB3W+pAjnzES8sJEC0fDPb/8klFnVLeVe+ZqsyvFfYKyS97GKqjXJ4
H2mByx8xEVBBDmWPNo5SLsCKva2d2yYUSbRFQmmBNIlZ0fof90t86GAFIIAGerCu/GUKCivNxp4t
7BVUM2bDJsQgPMTk8EaJVc8pUiPCzhTqeoIIh5SuSfKMAd5MjY7zNXc8AzB+vwpAaiYuqDcOUfZb
+KJC4XdvUNx9e8K1s/3gt+neLj75nFud5rSHRWSUSWb8iZX96SyMG/FNbNsNs76PLvQdiyj0AL8G
RzTpnf5mlDi9VNO1JXIYs79tnwpMomC8aErtMimDQGBkbiwpOMoLDcQ4v976vN6CnfxPwYHg+X7D
TcPl/VK/hN4g3XWI38qLtdyKLhZ3zNH6YaH54BYmPnaGfLCz3MJr1SWbwVQ91Y1DL2WAoSPbBE+h
YxMtYh4JiFv/MzuFRt1RNWUukluEBTaox1OCAqLHU+Kbmgmq9iTkolOBGGypzyVwBLtfCcuQKvHe
1mwvcXTMhNlgPGd8ohQ5Jg9AEFiSxaH+04Qrk7tKB2+iInCLkoEkG4RgfJq/y2obGlpYGViCrDgv
ZEFfInf6bjTeloK5g92Lfiqf+61xjU1Kw9zEnUR2PX5Lw3ZNJ4lOYbfENY09Ij6UQ7SJe8rtDyyQ
mAkq+0UwQuyLJERqYgOkVo7CCRbMDRmJVi9YZAP1SXTjmHlpLqTcovU7R8V2rgL4BUEJA9JJEvWc
tX01uysyfb3pTmUoVeFFHAvKYu/GpeJm7pHvJa5xkztwqX4BUP7UW+LNC+v86wxkeenMF4BsREdi
OQanEQAvrKLgdFJui0NgAjUbSqcrQ5v/XmmLCexWu2JKi8ZvJHpqPlOtBgKtYEr+YrPe7+outaFX
YFzT4WJWijYQDnXQm6AZ+7TY8i25/jJdCMr15keiZ3agFIL5Tow/55/cunwLfW6jUrdxJ2jS9pgp
xTR827GEbika9z2MdoXoLk5iXT8Ehg3akT5IzD+ylxELunq5RAod/epoy4pweRiLbn8bQ/TwYEzi
qAyqe+Olp0Sn9UlrUcgkdyZNS3xqDbuYnegU/bwFw0OYDOOk+No/k0jGDoQhvdd3eJ9bq8RzE5Lc
qKm8pdTxnFrai55Nls+iwg144izrpProofct6NPIgHJLdWVmRA7x2y0BAj8OYPNquSU/oHy5k91K
FSQScWY2M+mlyQh4LGgL+smCZK5+bMPUXYaxmwR3VWeeK8UKmkSE42L3r089KYrXcMvIdHa0bbKY
5DXf3SQfIOEM/NsCriX/F2DhanB26ss+81SgNyPQVOVnEdcuU+DWdLa/4n0nDIKrBuTAJuFZ+pTq
ViTqrJtwMXRRf69t2C34CuEl8gNBX2KRQAmbmOkrdKfE++TfFmwVcLPkZ1R5T8iHhppD2ASQx8Xb
uBFIcmGq0lnf75jWkogVVnic1xzdDlU7nv4mKMoJEZuzThIieM+nI8Hlw0CZFOkrqsklamrWrTiT
Xw7a/fzNzVV+2WznSrBzRDxE1eJ5jwNLJbzDwmY8mPwyp/GQVO6BEpVvpZq9o6VEddmfypw9+kSZ
VaJsAEKxJ3V4pQLKCZGwdIXGUrWlQ7dWho6u6DNWIj57ezW+7t7ehBfOsy2Ble0ebXIPSGLo+f0s
nJng7DYksmqksd8tt495PrwN4OhrI7Dxjuox50fDf7nbrmYqr2GpxgnqiOI4YseUaVWhVNcJUV/h
LmwXzq0lMFAhWJsKp0rDI5fxUip48ZLI6g6glYu3N0WG4hU85lHraVasAnslZthHXT4V/ymdlTmy
o9u18KaLkMldr6hJslRdLa7vlRiQf3jgdBAI+SeA3VP3xoUcUx4VRRW9tZDEstdo5y4ht/dGU1gW
Q3hSO1UpQHZjXv3VaavESCvxKap10WUBjeSjwH3A+r2gNs0KjGRY7Pjykr27tNlRBHXJtElo8tfj
H1RyAeZg9Lyaj/ximNgZOLXVZK4Aey7B+9p3NjinFLXI/lwpA67+BzJ1pesWgE7mtFkmdJn9F6wZ
461bzVh1B/AvHz4weGxm1SM178Dh9J1DdvAVBy9wlgMwwPOSoXfBGKuK0COTCfHwY3MJHUj/bkNU
2S2F0iw1wgHofe4RuxzHZCbwLZfb/ujj5gQ6RyJIRIKdZnEMMQlW+VbCUmAFkYAzxLGZzYApORL/
kzYhpsz0VvL2OxAhVuOtQ/d335GyHDtdrRl/HP4RE3wEYBadGcsNMnAeOQ9zo2EC1M3uYgyF29sK
x2mKk9mqOTxkOMNeh2CCWNxRLhNxPIGzEeOOcGccvbS+FE4B1XTZXFSntMqj3dKK1xnKizohcdVC
zQpKrkm+jG1nJ/zwsRH4oEcOprCilNansFmHBxpaMwbIUDXYfNTho2ehL9IRHTDQetvfxHTjOMfF
tVC8MT1aRWez8Ehmy37FnaI8Hv1Ga02dOfF4T3iIHPaHe781j9lnq34BAWU0BwNtBhQati1IPKd8
a2D5HKoBJQreJJAvM/wFPSd7u6mgFMBgfltPfk6zGX8yMGm40sSvkza29Z9ZpzlqDQfjjbdA1PUL
n7FdwTxYFqoqZTyyzofiwbh2JmB9ulMNzn9pUM72FZ/88ciTMSHTN/23GYT2Qk+NTznkl0peTDJa
tiFAR4B5ZZjeOfBaOZKRqoQs8HvJDOPPZUt/ZIpecN583gud9YBup6tlmL+GlyNIIvUxJV5bpg2c
QC4j+5keIw9y1hdOcp1/ZDZMwvnNPgN7oCJyubm1tADFf3Uva2LwqYcLZZugmypJfjwQe4C6ct3S
7lprSvc2KVpcYPojoVv+rCEC4g2C8dd4KrEBfmf4994n8t6FNZ4+RxdvOdZTEosryYfACKFjfod7
emTB1eqiy2C53NmqkAvFICfLBEwyLiSXqF8jf9/YfdQfQiNK/mffYhCb4TEPT/D0dVObUC85/X4c
mytvEFBsk8d/xpCG0xaWCJgFuFfxCXShOF+MfvcM7ZFnRF4I85aLg5e8MGhkRsqHOgg9uY8jjCnF
cOlRU8bcr/jeg1igbq6t3FfaVdPQHGwUw9z5T5XA2RYW+p9mJ1kh6oAduIyjK+yvr1hv6gjcU3Im
Bg1p9F5GSIYxNVxXUyJqcdinHcga1AtrwyZCx4ZsiXwQHsMWT/MUSYbUUMLTPP9EbtNAGyTC+sa2
QUCGZlDBPFSFeK6C5HP+rbHjruAJzVFUBlHk3sHUDO18IO6LcNWcFYM8AtFveSfZDrlFvSqGFxKZ
cz50T5ytDXo7QY+d5/so4Id81R40VECPskYF93e+veFNMh00Srti1p2mX6xk0SSF/lERRSNqo6h5
wHOueMNLoRBK3Gspw3jgPeTlawrc3kgu06gTXuFtOjVe+VsCyHxByd1i64RL3fU2iqNFn25h50h0
RokfIp4C0l6vOSi6tUmVEX3VAJBmDUfgtwjU9aMQCyN3gDanntBdFTjJgj30OJowKPnK+/djo4JE
nfEfuWdlTjZzi/1Ht1l8ya9s00Wzpw2S1yHlr8cY5AwuN7g+dhbZUtZND6laaNZIRZjSA6C6CoXO
5C3qUL/doFwnHm3aW1kwHDNNYfk6Fn/WOEup7JPv1YW5wavi5+iCQ0YCO/svY8HXdVALPC8uB56E
4u3iAEvJnd9c9hqKP7h0zFx3XDCSPlmx8I5LtLy+i5PlUFTjbK9TfzB4AQ030AvjEhLgPSEoXOs4
9Gs5iYQZUfoTL0+t2wqq6xAdvqHL42xeakO4v29YVOzVLidBKCKWBgWUKSlPkgZMDP9O1j8gXBrb
AvtbMF9YrUEU9Vn7aS9yYv+I7Rwq+oRQiFS7mHKEeMNafsSHsJ0gfT0nwtzZVc/fp846sUpO56r5
WgRZOjRKcNPW9GFn/zFTFnOADqV9PQDcv3HwQqiaSyR1MfII9KwwR5Z7cp10aoOfzuKBR+0AR5sX
U/qIGvU70v4YXMBredjz4HucRapCecgQgLC9H5dxJgb7jLB2nLESnS8ZacRZhavDDhI88cIGNEYd
IuimP1h7k6W9ekl7BQSrVeq/hWSZ7dvgfRVmxJrcGJwS2sxKZRxUIprYL+nUtn6AOCec+9HVgCwt
rQJo1KQZ5OQdgqwi6NC1fUXXHC475DWpktn42LaKaHdRlJN6dK5smQsUiIjn2q25r9WaoyIoJY+T
MXnNNS0dU4Lby1Psm/L76fbAwgWlqOC7gSvlph8A5upwMO2vqvy25XIa7jM2q4Y3jwOIXytgRSiZ
gKpjFLAoodyh4Rc8CtVlG74drr+auYB4jH0BQe4akq/rcO80ltCD+u8BETQYyspYbUaYxKE2DswY
d/8Mswtlhf1kuk6G4TlhAC24JyVXE5t1FFqRBY71m/oDf+uD3luRWWCrUVVe+byjE+yKpBka5GAp
RFkj3j1wUYEHBNMwdRZCJKWfmsDCrAbP11deNBhVhROpWZx1G3b+tOgiqApBM5OYBLgiD+IhQk5b
VwmJAVbjE/wHwLIhyx0O4rpqac6FiGplGgweRXaB/+FC9t4bGxRHqLUwuRoovTWEeD9jqw2Bd+xc
JLqC17SiK5nlETK2/Tm2GnJIPi00kVzmWJFqFNkiCodbN+rcJX6AxxGcJvWtmHLQGKWb0pH2+0GC
dJxyOkO+FSIvzpEiPfdLy5zz5ogQZ9QZo8ay40qgX8VH+P1ydY8DIqpz5nVBBcnKck3m0U8LVtHI
LBG8dMMX1c0sIq8CMJADMf5xq6to3mG+8K5y80O67McD9kAQXcckJh59T+XKk+KJ207fqENSkqVO
a0EH6/P99GFGFa+1sdlXMy5Z+oE5XzNF8mWC57o6PMob5hyhilCqkPKCABc3YgR24irCOWPZbyzg
u47wjWIgUl6HX6veXPP7mb3wOGEB6UAQ8EDsF9pOzdh56xnVmw+CEumUXC/sYEUuWQaO41uZMw+Z
lyZTG6JsMMj6AGWwzQ/1vYgSKpAXZJZOAHW7Gvhl+MiEVVshFR0emWKdw0+kDRp2DzB4ngAUWnST
lqSS5TNOgBd0Fp91z98RKDfG82Tm0GpZiUv3gAF6+aKXgqJrnu7X2e2Aldj1hndcdugK/4LmPQ9i
i6CSBH4PV8CKTaz8d+bL/CBXYr/xvI+ovXx2nAIg69TJXTw3YT68ogvdZGELNXeG3c+5M+L+D8Z2
QKYZAS6yn8f0ODIOYXm1+KuijU4r+5S/bqSIatZNB9rfQBdo3I8wfLSnMwoo7TyX7nO6956db8f2
fRnIvH+vQFKpV5iMPNNeNa1q9Opl9dlAClFn3Cs2CATG2hokZzkIDxvcl1TwEZcuOF+Wx5qRzLUT
DzVujgEmNBV9b5w/KBsm2XMaUgUPUcBlbKJYw+NEeQMUmYsJx/uSvL1cST1ug+kxXdy3ezPbQNsO
QZaOi5445kznM6rM88l3Er1W+YU4utOG/fquK8f2bB0UnvDSCb6BlOe35aH8aAU8/X2Lewa8sSqs
G57WGVCnVw9dT4Ii8+HF91YyEEZ1Wz0Tu7rKLv9ZNx2kYnt7oQZ/nCJuc97J6SPj7AAhML8m9kcU
59p8hMkJWMHhHND7R693dgcLgHD9kdQ+XiZO+NTfearRkQ3xN05yvUHzL14R9VqKYi9zBF1A/PnB
G2FGK/loDIIMMs/m8OQvjGvB6IsQ9xROjcqauwmF1bAdkt+z9aqt9Y74+IyMS3D2Q56hX1olMk9u
AYGcVBVRd8ZJVI+Bb+YfwE4nyxJOAk8nF4k0GrdhedLVZIW3MohvcdKjpd5NG+wpZA6LMZL2I8tK
g/RCMj7BSOKVeNa4eAqerZSPR1HsjSud+za0+qlEcYynFN3EcwiGyCO/nkFdcE39Cqmr+a7mMAiC
mIB+nILI7adCZSSy55xyTitCjc5puVEex8ZwUrOQrAV16mp5wNr6Q5uUbdNngU6MQP9xM8W81HcP
fDluGugW2ivsbP0nHCdDw5gpZ8sj/wtiO61DeysFkHW2ptZE7N8lwO1MoLkhgAeVFJdAmBpx3oEo
XJBDhR1nyiSUFL1nXGEnl/bQn5j432q8QbYcmx/jH9uGWqFBbXIYvPW0oe1wu/eY9CxyeGJhSnBh
6nG30qjyfhP/pkezYd/xMEbdF/H9LMFIzQmUKZ8FOrrqyMYxl9cSdGi+PCu8G34ZwA0j9BpVS8DJ
1nWai0WNIWzbkj3z5GRqyeRqLwgfxkxgFzStISNIu0bhctduEhw80intsRqCXR8F+SyVW8f/d90T
n9fxmiu9rj3LUyS0OgKjtq3s+CIRGguiuH+6Fl0OrnLsGhPbIaxgSkcdFgEH5DNCe+H5XMfA97N7
ofroZU2LouPVxieWNvuKWc6vJ8jhMeGAg0qRSaal4/yV9qlAqQXfnf8zq8IHSdH3bvfnnWsKpWLj
254EE0ITy3u1x5HRBMOY0flt0pvkhcm/QFbh+89GCawQagxtR3hYpiJ/pQHvn+6iOKT5tWa2rqWo
5RfKO7NOSSMEZPw3t179WaVPHIaTVRFrM/Bdd9/LH+7z1ElinfDv3MyLM7YAJY2pMwOvGnysh3XK
0bYLQ9w80da79VidxjhEZFUhm1fLA3BtldnWWvOHUVICz535ia2OLGokutQtcEKP87VvCfalONsx
Dad8m7yOCInPEwb4DkFo85bOhyNUUSRrxj0/eVcH335bF/b99I6kLVpuIj0lwiLT9AEqsV/Fe/wX
Yi/F/wiYaCn01/L7D99kSgVbC8gBp7LD77rX8MXZTh/4BhQFQytW8ES6wRa2xR1SDyXgfOfkGbDr
Byqi2MonbI3OZ/vPKU67uIDhIKfO6u8DdDn19E6I9nR6YrjrGbubtf+hPiHzX/TGUDujQ1YBflH0
y2KBsm6/a791PcYGrbvvyraJf6inK1oPRTfgzdCOa75eMysq2Rtxy6j0BR8WOhEo4E4ZXZIZzHhi
UYC95FBzrPjOOjRh0GWkn3Cjqlz/nZeb6Fyi++9+SiZu5VNHLGzbNSmdhSmvlQtEus2xHGHzQkMB
UN9q5//a0SgFhAWBGKCA2xeMeiqUGlJ01ec/CFsedU3g7nRgDQvImUl3/BEar3pMc+3FwtEPUA6E
FQ768AahT8K8JhWykJg2ntb2K7IZLGnPbwVmm2p8t4+I/StoL2Onf+z+Wulx+GBmTljbfRYTq2jZ
UEJhmkw9AwgE5lNNzKUeYFgAcXdVp1pdCJAwLI9hBHUJY8OTPMJfUGBg4FwON9tvuikB8ANM5Sqs
fIS88juM8MKy6te6R55jd57EdS9xbKnyZ9OBD4IvKhUlmuEHjbDAj3wZnjykAWpR89r3hAxoYjKV
QqXRJ/6/TLVmdV42nkZDxrK5xq7wc/e0hi1uXQ/KwROXE+b56htjW3Of3LC0Ebn1LpYROrPkaCYm
IlEd6AgAnutq5E+3lq3bgYJoCjYAwv1KkVsILuIrr0LiqqQk7JTTIEaEJ80GTwqGS+VlOlZHNo9f
ZYXNGUN8z8PG23O5l8tY2iU2xPr8J7QZPB453gR8rdYuAItE20lJSm4F5m2XX2QCEWj97mlrUGsa
jy0Ew7TsPAVvEt56cGRGv2p6Su+EMAdwBG1aSmk60DW2LgwkMKafoJTzOrQBXW0MQgSmhjGzBpMS
y66b7oJmWECV3w/9ttRb+RfAHV2EpUg44kYN40MJ9JL137sQC/81Pgw5qkvz2/PWqT8A2wpj4VMj
nSW6CZdvE1Q9JHSwlEEU5GGrBRq4pRSibPZ9adc4eWO95JjwAnOxUZEo9l178U/wHs8lAtEHDcGq
P/Dhx427lW3cN8EzzqPL0FwssQXGzw/h2x1uyWCM5FSGOl4Ha751y9pKkdUiOXDyoQSTgVbW+WJm
34Zkhf9nygntfdHuA8a9VXG8YmCaU0syH0FRZEu8vlauurpo+hDW3Uv22w1kaUGUQOrISGtPpWtF
xW0qanvsVU3I9xDTHrlUkVgB4/xL+CbFPdWsb4x7xZMXbToQxJ9vPSZLQfhbWlTw1kBs0TFGc9+U
sqo/O9UopfeIMlcIHNx2j5OYsMUY4X5IfhNkqWCAwiN+VfL//+LhkgxEv3mwgOZUnGjyE9IZV4t5
wZVup2AwgBhBgDUN0XIw7F15li3Kd0+ku2SqxQwJguZPI9YaVIIuIOcEJ3tsPMMxuF78lgzTbMdY
elePfQbH1BEaJPUMM2/C+UKA4Jpxj6CyrrkPe2fV8K1rUb2IKcduC3lBdkIVLrsKZ27qaXly8dWJ
omoUTiR26F+6lLLNrylvEyphwvn5jkygxnU6Z/HlZuV7GKzWXdT887xALE2VREoIT73tP9zxyDvG
baJbS5L1K54n84NWse3fKpNkw7YBolugGSTMoDOX2Jnkzs8rNOnOGHgD7Prh06xUq6UiV+jOMvGq
0yXv/73gD+Ab8h5ngUZ3LiAKiLVX07uuHWDfr3g1hpY34cz/FSsx8I2iIi9g0I1IcKCE5u8eQfZp
vFZJcuxbEl4xEzaGN6xWu4OddL2dZEu7ZIAy7LNwMQXYTQNqhEt/Vn+tRywa8+2PQhzgdVJgzZlU
P4P4Ww8vecS0t9IfWB655zSDIqtNLh58Q18OO9zVmLomgf/WkDOb4PElHbLtHyJeeF7kfAS2u6Oa
UwroSKVaTmnkZCw2mbcaa1mAtVsxDlNJv5ovRc7pBwpz6sS3Tbi58uNhJx1cumoysqEtWbcSbtwL
SFUJ+WmeMM+t4pxS26U2ry9xH661v6tG6h+IWFgH93mRhWnJzJ/TBGnb+CMGHB63pOTXVgmlf4Il
HD6ismZVOW/fEuE1c76w5ybuQyJ4SflGo/mbM661WPTMxEzcFT79Ki7xOSvY+tEKi09PZU7yJgF2
NAK8YgA2wEf7dKKC2JcDjVgxR7d80neVkQiIk1SkKCQI7IrxFtRBLKEs2DbBuVI/MSTiLLVUUGKq
RsfV6e37YdeC+sK0lDvL2S9xcXd9TsMh3X8rSvv2CX1x9f9BMNnRyUWWBb49qWokGfZsMEcNUBTj
XGS7uSZJQjK6+LMWwEBZq5oRC3jOpqbxeQe8zXLddjXNQGc7ruSo8yOAlRJo2nU/ObqrZLJbLnS0
MfvUv2CKtLYgqzJlCb94Oew1brCH7CmuDIeA8bxofKZettyP9Q8nK/cksEU+nK5WcejXBrGV+wci
fEIj7BSrmZzQ+Kyrqdxo566SK9pJkn7l8HjqZn0K6Sc0+Snp7wtwGidAjDEsMqGGGMmZEgVgLDdF
RHM29yvxpmoubi4EB68hWUJG93FUpr5fjnwnCgsj13oLuQ2d+awJ3adbXn9gh7ii4Y498EWQKm0Q
UYAEKBP6K9sgaXEiRt7A7d6xWbKotyOLLHK1n2mWBPXsV3V4aU/8Eug0zJb2eq5bTM5jyMtS5o0E
TOPEQNSvNlxRn8tJgt0rYvv0qT+mvOak3+jBd3LLXCBKdM6Mtz32Hah4XRizM46EjBDHsPxBNxz4
emYYA20RPUyIdjdRd3+kS08ZXIz4D7iZpzNMpI+6urVXdLhsAp5HfQpgpthJ5ywSZK/XiqBVix63
8YM+98yTjt6g29Ol7hnB149I+APVvg0Uj2JbIXDUVGixvdQosKJJPmT4gs6HHFh3AKxixIHIujhy
ivI7FsenTH5XR2QOT7J4z4puHD+lFWEZcCEW8hzEdN6NXG4grJkb2i9p+LgJzF3b7MR8iUO89ffc
nrKG6GjdFFLRxU/kiVP4QSA4uQAIe7qEPBrwYo1UbVLn/2gefKu6ZHy8I8ny/TNO9+sUMFI6T5uS
4jCjGkOBvT5BrSqfV6jvRcoSCRzYPTEi7MVHbPd+bejxyJd27RCIMoPP2ZTeEnQg9W9vRJjwzvRj
puqleUnSB+h50rQvcBr0qCF3ccSZWQCeoLes6tqs6W0x7SdmXTnJVEXrHNGBuyp6skjLdzcNKX2u
dmkctF79dchJsiioRCvmQha6AKZMnauOoWGkjTMymLyP1l3Ki/xl0VSEN2g+WhWfeT0bEAi4eK3h
dfDTk8d83YaOqmrYG7WXnJiLmY4WAc0aJ7q3D+QNs4Sn17onnmMzgAPDbDIiMVi5kEzd48YRPK07
pV0dh2N3FCWkuPwkWVxecpnhTJV4IxO8uCYKqaEJlWwTVb3rsxsM2NN6HjtgPjvvn27p7kJN6IKa
LuQDhmxxWL9xvW02lNCvnpycpSpCMzEtsigMBeHtXJrF6pt1wMOtUS8caueKGm/kuRsQNqXQ4Tu7
AthktOSTVQihBHYn1KbITZ2ZCCMNTSYJ210RXI7YoWjLk0u2/QQHK3xeqVc/fjvq6hYsoqx8BllU
YHeKAeG6ipXqotsszHgPwcW35yN7hrpoYQrvxZ+OLG3wvbKhcxotxOP5AUZaHDysFaLiCdN07opF
WnvGhDnGTeKgXb3+0WKfa8gZiuhBdPTcqCJgYVnlZoDUP53rB/nwuyanIlkLgXjZEviKlhiFJXrJ
IfsHabQDfJ1AvJMywoBvRS2wNkc5GEzRYkoA0dzjO6jbeZ4o+O43r2TJSRxrpN41ev4Qy1HmSDvm
00zoS84oS8tYRv13Kt8LYFujuBPJR6Z2SftR4WXLZUPa3B+8HgDCyUaWljqvhWQe0gHQTTO/740/
B8uNTfsGF2gwfY0i6/cR5DKopp8C0idl4UeyoR0VhP7Bc29nNgC9vcIR3BKB2auAjxnImjb4EzaP
0kchzeI5s7g1tBxNpKYlNIOUhPkUK9lL3Qb3RaDCRG4O1KALNYJoB1E7BL0MYy9fC3DZLGX4Yilm
cAH80/RxkhIL8USTZZywZcAaHOdr5gs0nD1erYq4wheV5ApP6WhwxRDX3POSDupudL2J7HcUKpMu
72s0fDlMhgewfiLMtFIVY56e/8Rj2wE9sZzfHfqsFHLlgHTqCpGGHxE6+h+wHAkIC2K2xgJTvBlc
ZKal4ZGkGA3jYytp0HmfG+lRkLR9kkv1iwsDrFD2wzuyUyBav+Pk6JbG295Tpi0addWQgLF5rrmX
XLcyaR6sFVOraDgMx/6HZf/fEJYIi367BCSCIECFaVIGx7K5IR4UlBNhCLCoZeoTl6b0+RVz8phW
LRfylhmDqxedxshLfHJhtcJ1RqY38yk1h30jf2+FxhfVpvlwo8QS4UrWs0uj/BWbEuak3HORh6od
DJ0bxMeiWVICm9jip4l5V2UVUMouOarM7vKxPQ1eH9itkX3LgNVsuwNhst8+N2YlP6+CHIPqL1C1
Dun7OgyArI17dSyACmK9CrVqA5edK1SRQgDySdknfE/7STnz9jYXJPj8FPNnHBpOe4CJOZIbYfi6
BiPRqtTi0k4/evyibYH/oHMaJXzNX0urhDPAzjQP2OQ1wxGTycPyaemGvz28EHtZwDHkwmoRe6Sf
Bpp4DpdmV0nbup+RXiSjijzwWs+XV/mskGUC0NqLjQ7F1zM6mNLIEMKX3DsJc1WE7KTVTdOYuRel
mf+mmqDH56KcAKBZ+05FYvnPJzTmvkn5wHlRuAKC+fUca0xz2NzbL93LsOHG5jAnAwAKAyCz9Y4X
/hmcXnCL74rRk7LkQtOyrSnWmhPE+je9fx7GnY63bCEp6h+po63JnnalUjMZfrUNYfxtljUaOmPz
Y6SFT4L/le6VJDXPFI/kri1nS2GE1VI0gCKuHeTxM4oe202TWKhg+krUhW76O1K+W9tTOM9zpFdn
kf/lNIbydiiaYFqWn1V7jHP8DzDgHM9P/JRsr7eYg5HqTteKP5XKxqGhlUhvAVuVJlQsOyle6RpL
IiCRrGGSyFxwL9ExJ5Sidmnt7BwEyR4euFU4mSww9atK+cKNoT06zKYiOoe7aO+0WZMsDCNoA+DU
9pUNjRfFptKum3z+7JerVfwYoUXiC78r4sVOTzloX1aJO8FkyqtVt3rue0u5CLDtiI8cSl3eE3ER
wfxG3wgUwpzuKv9b3VF1TCHP1jDDE6YRJxFa7WGHzaFoXb98UHHBp9oWOeqbsyiJVO42amrjHcXq
wNYkzP91j5nFVOWjnHEDHNxYjxxG9C7vKR6A8BPlUJDJ88s7Ckl8Ey38bo2UdCH29uEwIHk/Gztb
ScoKHtl5KGYpV38lsD0hOmOuQQIUarn8aJWQakM19YXv75xRVUTZQiRzgp7jBVB+RA92RUbQCumb
F5PWcovOxTG1A+WK62JpwDOsAwMbFyTbVR/09OjpeHZ+5H0CKY5A7bC9kdzR9igXYWsVkA+upeII
/8D23QBRxCbAXEYkwksFyiGkJcFZ20Y3PNpZB//iJKF39b7lqQ3CaSppq//cJBcIALv8vZFaN6pr
uxYueJ7A8XcnRHPuYdJ6kkzTzWUACLjrDwKWQNtl6eR7iV+yUqSwLf8FwxBzMpqaQ00tu/pxvOof
9qOdeg2z61TEA5mLQE4pgFjoT+FSBQyJ1GufzWfklEx3QEc9g+qRdq9eGWadI9Ms6hscs8O2pUFf
I4fK17Ork7aZ1Tu7Rexsv27SCvNBup1Mc7tHhjqqAj4HoiFn9O6xRnr9w8O3GxLXuaxh4QjYf4vr
a4NbI2R3yORl3qAh0oUvXHVJkRpiIlvUu0zcqZmQo95RnIXCz+obYyypjA88Qcl0xmn+Z8TLUsWM
xZiKvOpp6YKG0N+nO8qv9tWJsEi35Jzyt/aERTUxTf3ckqRaZhD37/qx7ylEeaAn0ZBCkKLTROy0
URX1Tyb4my2L4bodp2lE/Mx/FVrXS0/SLFC8z/eS+DS2PH2IcxTsEKRoNaEctEMBUC+7sR/lB2W8
1KgrPbshY50V/lugtSpT8hPLnMB3zSnDki0Eq8mQOQ/mTvU03alykkJnVWliL0gAzuHZgIQhGihO
bWEPBSaZrn5yjMkRkI015gBEURvPYZXRG3pMdiFm/Xe2hMiPcb/OtAg/kYCSw+gCMRYQzi4PcrdB
e05dGOWfK6VRSjk1zpJokjZFSJuY0Pqhgk2p18NyOpmMMg33CAXfDf/YLXWrDEnHR0cjrheyLkYT
lmem+R3u4vuBP7hPeItzrO5+rAh8DyU3TnlLRF3zHg4QjTxlPmQRTsW0YaxzlkPS8HqrhwLA3Bof
kKlDf3mVw//X21MMF19SNjxaEIfHybrTh7c603EhFZfKprFqYPeKhSPHonAVlf9A0NF5BYBkpZX5
fraSoDvNSgQs9fppDwsrkaPZSbzjr492c8wzXWdhs1ftA/B3h9YiBVGUqz6PiAmaTkfANF84ydXf
EOuBFP0yRY/oUO97i/s42SFlFW6RCjBhq/PHtUEu3oTnjvKp8OrPwnXqugBKSesbA/vUPExfpW6E
qjcd2wrK6ThnLN4cf2S77H+yNMmHhQSNGd4jHShGbu3ol3DLFort8NTOB05HZlk6zkIMYzgoB19+
uxSfBcPlFItfrQEDK8dztdIMh5nGNEVGu4Bax1dwXCegmTnCGi2Dz5ZIfMw/ljkuhOYk2Zta6lvH
yw6aGCrQFiOGZW/5FKW6l1+rpkufvisjJgysTXpq6t+oKUjGmqCMy7lrjAmAN/w8brsP8pmMcKwC
uCpBkgBoWHSXpVW7zqSZy/tKbLvGAhC/RqUXEjzDl7BMVdYpiLrqCZ3XtHfzfD5+yEYEcLWBaZj7
TZdn0kIuQDKATDQ3NKBB4OvstM3SyWxfCcaFPHkMWm7hyjHVETIPBmX8N9NOkYM4MwlOOh45wHXY
dw0frQOygbi3g6TNpLCXvmygtPGefHlrxbOFdDlOTm7qPTBnOazryeidryCOv3D6wzvBLzPXaJma
JcEBhZqIj2WmM4lH4TeG4yHMjmcGdugFHkjh3JiPNsjp6iOMBpN6zaShiq9wjpYdOaibCo5EYc57
hhwsgFjs8O8FbGI/vJucNthJ1tST8+f1iMbzvocEpBjuzdvrLorBtIDQs1MnoMsvdC2i7hKXGx/Y
QPRUDS7MD7VONidUGaaIYg1oYOQDLPQTHPrffQxQJMvRfAa9brFovaL0Bw+Qkt3s8KvO5H/IxZZx
o2z6eX1Qo3E/Gu/Ki304SxFAzSs0S4g+/e5KC0hZHl1VYZuKxgCuo+qcnTEod7bhkk2aUzMZda9e
gvnYkYK9kaExWIOeJ5DoB5wfPKIWNDWAkCQff3EuLXGHUzumnVgCSageDD3ZyFWcuwU4fVLNSc9r
Ovz3DWeQWFVNWdSf3xVd4DdgvldIHVUIyOqf63tpk9rRH2ov//Yht7czy9xppmPn2EtootgBh8+G
68Llel144OUpufE73jCxRBhFvfT5+9NVqcFaGxK4ch5in9BIU95YxRbQqhHFUNTCuP+F2M6xEEhe
LcTOQiGfwxHNrnDstVtSO1QJFhsNz+CJcaB49nBvqrkdSXbCSULp8OhX8MDoHPheZDXOuVxo4tLm
zmn5306H4QKuZSTdhv0lrBQ5Pqvu3VBD7eqeT1Xk7Y+pOhs9BjSzv/wI71vMXiDxJ9ZFCDmKBDzB
gBjog14yIg/waqi8rMOX6PR/B1XrHTN4Zcg6pNSqGqtsm4OavHy5Ji4wcN/XFuNYqRQvhoCAlE4R
knHROZGdAfga5ZoITUic6HVdYR6m9dIBvuwMJGpnIQOl29gTZV3/l7i7ogq1MmTxNcNGuWcbpfit
i3BsfXkLpvHXMv801GuwPBtAWeasELUncfzm5gmXwNPsrTXXSEWqPgQpdr1Xm+mcEgcCnz9/Y4nz
K1jf4i21Ul0qAliwv3+30E8UE6WPnEQ5Z7kTflrVisn2dkJjbyv36Zv0xNXgRGCHTWQ8k1Jxyh83
NcNvwxn+ZwjIvNTjo6sjcBDsUjRfudeQjme8qWs1ny6ZGson0Ver+vu6EE00yFzOMFNWoRRdDSLQ
jCmm/OrSsNfztthbG+PrTKXTXBwu3WIMod0UfOLEd01yDGYVzzTer6+v8xWQf7oeWnJ7v+9mzazY
Ec94+cFhtTrjaW442sQ3ddUc0+3z54twwzOegRSeHFn+tFUq/Ax7wexBs5VOrPx4jFbBViK2VAuT
kZ0QkpiYi5IWwyHbMeI8OTf+HnZvmZNqhrj3hSSwV2stCswKC4emQbpzSa2ZD03VfYPnOaH7gtxn
RyUyxTvSvongUQsh/dneUQOVZd4R10j8RlQJQrmXRO9ojvI3Sg5H1ZKStK5zhjw87BVXmSeBR48S
cYub2g+WNqg/+Ue1Ir0GU20TpBKGcQ4+WDLt2c4ObNYCTi7vizn5Wdv3KlIEzKiSdr8Abxt9yC32
zoEcXZdct4PnryRUl/1KaSPkntS9f4rVxtlrPZdFOyOA8XCYsscizek+f5H/K3Q472udK+RDXQfI
iZecWiQTwwhdaN48+uviF3q0UJJXasA1dB1oH8qjwKD5+RAuaYRmoR5wLrulvgYdYEvQrd1jeriW
bRZIja1N3hX5SYABSbddY6Mi8Tkj8kEhl7iDZBWeYnKGVHBtc031HTD6pE+CdniYjltXTKJ5fzin
ljwAlm/JfU5UHkfVQ1YNx/yve0C3ai+MfRX30GdUYiwXW0FESQrx+kKgMTJVn/XL4hD0qhLY/PM8
Cc61zw14HK7REr/OtFcrDJTLAVEF+CGksZnQbQAJPGE5C/dA+Ojv9nkaptKnvVC/iBic7IJtNygu
GPscUzJRs9dEImwzgWJcforjPJD9gnSCZlWIfNYIc76ArzgQhEvsFzJWgVtYr2H44XlMmNQHsLUL
RmTVGKkNX7WukG+ut05YXx5QAa9bKtNIdfUHL3CpEX30xjka2KMpZ8MUZX829nVf+BadBcF1N6np
De7gU3/Z/mTXZW0qVST20UOFfUi6oBJHf8gv1fBF6q90H36VReLXum/d+Z2/9o7WVDl/tKNavaTc
yMnmvVyR3qE0Bk/whsX4Bzop0pPjBfeNLm+IEHyjd4OyYxhAHvA4eNh+b5GvqOOOIg4O63KJ8uo3
LyMPy/lWLSU4ZU72sO3BIYvqMoUimnyftn6cze2Qgs6NrLCouNyszOrQbedWQRceCoKVaNb8N3hf
mY9IjFFN+g6XTS/MRQZmOBPnrDKuvE5WQrmCmMOol+Mjm9FAvvAGpYP13wqtyoTI/ISSlxCi18ZO
4xbqZ2eRSGwu95x5IAIle9pgX3t91S3DC9exGR1Axo1pDlKCnG3VPGBer8MBnqardjphsmWiwfqq
4C+w11qfujABYc4F5fh8FSn2zasS92UYAE7lzF8rfPXhRy3lU16TpLuLFkzGOUigXH7EqK8K45s0
0MMvVZYRbW7H164zOU5eP0ZuCXtzXcy2NHJZwo/fC4NShv9duNbPa1hSz/mxKlT5IiwWNlYIpbfM
lTiFe/7Yd9Kf6TQ4PDUbIxsYuX7ocn3fa/j1v77/IeoxzWRU5fWBb/9ZxolVeCdFzjsp/zivFp1p
5n5BFBahnAFpuJsaAB1IWKK431QsrzdwmQh/5kUUehupGsFJg4rOBVpjYlemyAI4bFKMwLAWPq0M
sn/A35dFR0OEpDluxsftWh0N5Q2ZkZAtg7y9P1fCfidl8XN2N3ygD891xaHTN6O6mFnHOZyvydde
Sp1OjOOiL6f9TDPhX5QTnHx6bMqpy5FhJHJmSugvtKynlauhU13sjsaD2Sh9ER8f9B9mwFXNdeB1
qN9XVyWtJhXnM4rfw/8woFctoLD05Co1fsBeCisG1xWd8H+FBn76AGSOFPwMkneW0ztnF1wJfFeg
svFkwNvVNAXfIEQs10j2fdlagfme7NXS149lsD/iExp/lftRXXAzu/klfrx6rmMhPRrtBeVYEtCx
p7H5VDqYPiJp22P7QjZ54CEaqqGZhN18PCRy/0QszSsDgQmiZ3hX49c58fEQl58Qed89HhxkIqiX
tclo0De7SzDg95T4BpO+r1dL/S1SbJkFrUXJw4US/A06m0kkbESqDIu1pnvxOFH/6iOuJGpThSZ1
tUXvjJ/yYce7oomcWDx7m8IUHjQ53Qm8jf8Cw6LBvRqt+3pMUAmZe3CXvCho6hcmdG27R2NEXe0h
K3u+xbltReYenZyrvlPLikYgJsUhVtLl9+NMGnF8GwODFFQpc8EEJjRwTU4j+bKkfHo7a+t+pNhP
jKfc/NwjOWtuurpB/zl/rJp1K2JbzLlNK5F4fKXyDklPltT6CjPPF0jvLcwZ5HGKrEQexl+I/jvU
Kp4Ji3Rp9qdcHYWUW813uZ7ghSvjsaAoP2YNIxsXtRTAgJT+HUZoGNiNxxabQWenmV83Hy9e3CY4
iozTQt5jT1jUmdOcpgMOm30E7Ucrp18ERoFqg9tgFu+uFDIo3nsPClonDxArC3TtEeRIJdhocoYF
tE3zTvuqNIGdKfDlURTxDce2vFLU8bvUE2ZcHYDFb9UiDxM8IkEVEt3uRcVJ80Ww9TPqIUSMOzJT
QEdamifv3wKQuK58839kjlLnU5YntGV8dQ7UH+n1PYnc9Hjv5L1dwX1Bi59Ekry6l+LhNDr+2Ocr
avVrCO2HfK9XgEqTXFz6T1sk0qz/4P1LDKfG0tSgGkjIKzjJ4N5YpX1XbQOLPWUiu12BVUHeMzzw
924mPepmcAat8IdvHHaURnPkrEPYg0iBdYLgByy6X29PjLYH1pcbR4q8ieQEzohTjCqMAekuqRfL
vAcI6DmBWjEScOkjH6NebnMcpykFlhON+lTEc23jcdhBjvqssk0bMLMZt5dg2Z65NRZ5yEtJb797
FoEvxDZTYHTyUSu+yipJhEjqpp83zIBDeY6hK4wZtp54fSvcIX0vuCb0bbuCL2RxR8Lw5G+LQ8g2
ppEMJpehLOOEGw2FI6TJJUBEevwxtpCWjTL0kEKe39tX0Ic1yv4b1NJ/d7PQWdQV1JKqE83pl4Pw
TeDabHC4jIhCnznmYl4EOJJ1gFfKIo4AernlTSS45CEJPW6Xsmzg7RnmYV6omv2uERmK8+HYOA4f
M2KYOPjdLrnQCzvytsu/31clpfbDcvsczvXU4D9P6QJ3EFRUj6wdSuJI9C3VUfWWkLQIuMmv+nrl
5D+aCl/IAe2DI9ZuwxlGyITDfuWOUWxFVq19PBdEqbqm+s6Jfb2mpoVowfMIFfW3TGsciaE9gxnn
p45i3iDqqINxLXzE6/PSf5Pjh4Rh3MVVbsy5RjBT8am82+/mPGXe86zlV3+hyAeypJXSKKlukS2C
TMo/gRIR0d3xozdTTIoM+fJgWxrwUgdrURo7lG8dl/z8lCXVcdqJysIsz+ZoU1adrOnSrE+GC+Rd
QuCypZRG6B5HHMEkV4JeJp3fnnMltAS3q/FSqgYTbzRPbrJQ7EAms9/dfWJ4n8WY1eqO8TBkNX3d
SorzgvCaZ3YaZ8m9xcKxnaBrmhh9Hoi8lzoaKNq0TKZfYNAv4ucfJHjs+BWvUnYUcIJetTx3Md+n
N5n+0gMFOn57oulh/YxjNhHvjzbQniKz/rV1N+kYlcW8qG2jfKaKC3oL6fd780LZiPcPCXy/9aVE
W0bpyz/DoQOqMWDmTgOCd26IVi/eUtHYa9cTIqNwMr8C2oYdshsJgHVVN6abKk/qcmtnMXAKS9z+
xPbSUJ6J5OBKtemWDlUPt4LgsTbfOLMUKX68BXHghWHh0wQLypK9RQ8b7onpKvVcduto0SRhUkij
dwft8JF4thxsL/vdN1y0IEuGkdzhILiW3qzVTzgYPmu2L0uJw3YH7G9h1TZCAvQfrPY6dECUJ/QP
GQN7cn75dC/ydZgrB+dB/bvdXVxERHMkn6lEj+XLmPhyiNwEWy3O7r3DCaTBFDMTuAvIN9zVVK9f
tTDfOCsRJVbg53JiCdAvS7Y48XZbart3UACzyADXrlntsjsTzP5hN2i6HdUzAwmCzC/EpKP3tZWu
UN7SJzswggQC1FUOSLQtoo/ZFMVCYFMyJFOrz1zjnIhxk9LJIe/TfLVOT/HzndsYilQC7grtyc61
InMbvNCNTnHKhvQNCYc329zb2OoJ5Qa/N57KEZOsK66hfKXL7LCB6itAfJy8awlgVFSCCZMDGvi7
R8Ih7MhnoX1YikKnrRGTKhwnHjM8RQmkz3kpUbzlu2DjbMgNRaW3oOnGUL4OejFyd5FtRtFa/Eox
pkDmoPS/IslRiyBdvIzPWZOuL01a33VUZkmzBo/aHftkD1TSsUXfizBX8witqSQCl+Z3cHYDA77y
pFGugMKb6b4IP5Hkw273HaYLeJhiy/pc+FdbWlIvumz0qGl2Q4VDOPPbnE/HoRdtSjuIFa3gWyPt
OtbltMbJhaQHFPCsJrtnIwxO1oVl08wMQJc/mGvx3TDmuo2Dst7yL+m0Iib5GKDPg68SMsZUQExD
WjEIXt6jdutpgheHsJH9nLJOW7ygVP/opWwrphvo9jaERVE+E20h8qONr+EegmE/LtRjwPSZRsRb
CujYdj4KnRaJcmuLdIoB9OKrXpHVDEPBvI1ftV76fsbG5deEOYuWUQStu+UtbA6P5U8+ysq4ugXY
XnHZNdiewnVFWfMZnuTajRk4+l9IUi9Di9oSNw16DOtzT9qDpr1EuLONEPGWCfQU3TSqLvvdNlKd
8xq4tvTILVJQme7ZbojI5VUjxBYR0lYci4pv9wm+HfT83daMAbZeaECZq76jZhDuMfNbJ0Xi5vBN
cvMY534yQ9VHbhbhMYVTryfTI4srF3VhCucSVO5WezMlannSvkZEHNSbfXD+HfLWCkSHGD1QKYzO
S97Sn+pkG+TWQ0XF7kqUl0V5aLprr4PeLWLG75F5WqaYtHOPLjNFv3qkpVFfvlzwuTe3UpLbQNMA
tS1XJZYH7vhVF+1RRPdfoLvJ71XxPfncobBiOK4/u3OH94t00G+eYw5B2SqKOnXBBZDq1EUj+s/L
CtcX2Y7h3tUJU85h08p51N2NyRlwoxHlKPVAN6ul9aRrG3p4OYrDcJMDsoDRCebQwLZ/iuHceY0o
6NITPJw7+88MC77cfkA+6GX+zpxqDRZ57JkvXtZhP+M9iwoKRoWjzKv6VHZFgHZlLAEsTUp5/I2p
J1ubPdPF8EbsrYkzcNvfyAaRTVwFPlUyobQpp3cyKTZAD1m1FW91+TC+mInauyOVtyo5ciQxqG5f
qnJZeqThrsJ91D++c2NDSfoytxMZFDjaKpmegsG61nV2f/Nn8xPYom/vtcF+2a+iqexVUgwq1iQr
Fb7+r2LWxGI8UjYl6rN5fyepB1LcRsAt3HVd5JTA3r4MnEgAIe7Fy4wRjh2arvnOeZGFUvHYpI18
Ilmy9VHtCRbuKrIMnck9wossCMGH6Teu9OLv/GxKw91c353SHNERhkqe9LiNZieHRUTrMLr9aXcu
4mToLgBHLgZ5jxkLqeC/3NBt9a2HOb9Jhx2bzd3ymrXg33KK7RnU79difOvrEKemR2wQ1rr7IJvB
VlgH93JSTI+6Re+phD2UX9hKPvLG+fGxhCNuJsmAQGBoudCYoWsz+Vmh/D38P/m7SnGXYZ5YjZnq
km02zINMxdqZChsEbolv/FYr/VhNW92nHPswooGFRx1TPF7wBI44G7xBg2YwG+Ze3NWAPF1ewcTf
u7shyPHq/P0kZCLR91wu02WLGI8F2NyxhMAlR9wZWh+olLx6Cv3L5LSl0nx2t2Y/4aIV8wy4pPmO
k9WhbLNIgxdCMMKzBUm8WItmhQc7XGq5TNtlz1Ygw/gSV1M2WOWCkXFCHtza5rY+goxF7zQt6Frw
lnZLXFFMDvvkbyIduSFuWENXkpSCP5K2OcOBCTwwgiiBZaW9VTuq1KVqKK4r4qE8VxD1wE7YLp7U
4O210f/jR2+yXoQRgdcPbCTyTIhtyeq/bEGGen2QDXbscbZngeqZS1aW1OPFjocsj1zI28vi3Ugj
lV2NNHgs8EzDRyGoklmzq5Elk/Qe3hZqWb+XLtwMq9zgri7k7DaT986VHFg0n5MbLP5Te5VQJh3b
XKjZ7vhajvm+0nmT1CnkSkg8A8BW0uC+fPhYjtO415QMFwtRfLg08HHYXarYgT88CqP8ZSPk8ehB
cjjiv6keoeivi46z9r12f6uUXRjo1bylumc0SdxsxsJ5ZSlT2oASw54Po4EQqw24X84DYkXIsQfX
hkFwvF1K1z3b5jhkuQ+f1+gf0UX1CqRLa4YSm04pUzsuadwY+Yly3rk/ULcJCKQZI7Y7P6LncawK
yxpZ5a2S8fMvSYEn+y8uqBJHN88Gizh9zd4VoquXwqz+2gs02cATeRwzhuKcJ+vErGoY3/4pFp4b
oO+4OOefcqsaYitGIJ30SP59nf8TryPLvyNh5dfFcyVZnKYxq3jGBii1kO5hBfj9BhZVfW2mkC0w
9vM9jrCivQuHIfjTsY+ff948Y1iWYpUWEU70dkxsS4forJMLjde3oFjDwAEUPR771F9+bg2ZJyMh
mNZM1tzdHQQf9PeMWb0zKuY2CGPvPcrneYDmeBb6hQoqHX/fXAIhyjqwfn83xWP3DvtQeLroQAhQ
nlWgl/LhRBzmQW19suQixGKophfx/WlA2yRLd5aR+SWk0vHhyxinLJHzjl3NUrrZb643h065MLRe
YYP7Gy6XVoARwU1E6CN68cDWiVetpJt5fd/TKQ++RMTFCNz/eb+BxvAweLoPybHzOh9bu4Ss5M/c
nyiNLdSpQ/krKm89YEm8QlcvxmuIshbRTKNalWP18VpNM6UT0Pr3Xy0s/8YehNp0YAr18yV/bbZU
AO677h2O/hOvpq2B+yNlnaLBz2aZzUo2ptE5N8PhHNRhXbZyfN16qsdWImomgYt0EUring4VeHap
M8+nQ0Brt5L4WJTfNKwjbhTk2hXQ+Rbe7jsJjbLMk3DCYg7KftRh+4En1SHvNt2UE1u91fTa7RhO
O2TwzRYQJamACAuGLIhEPZt1NoclRY56MCuSdw/N9UrcOEBjc9nS94kVgDzCmCSROp8jKNniB7RZ
XF7CRYxKrshKGYlFTkS+nyth+LQri39Ey2NKaTr0PjPqp6ShNkpL8pcmfGKiir+2Fj24TbfzF5VI
JY+VNWMQBOkhQC8XsM+DMv3uXS4RR7gHp357VEUqH8SlWDQUxbcE1b6fM4ab4FIrsIq+wVP5lsCC
U28jYJdPcuLcg+ZwJ0ncl8YyVEjS4asypcWGyPDpSJXlvIixIi4phkkqfLknMKQc0JeEWWIZk9SE
TcpVhdiD/W2nrBIVxwLrdg0fEsYAGjqKHVMu6WjBUfia4ajIFahniVzR7KHMuw+DQM4CYS2whmVG
cOjKKEem5N/3lCVBy761J5/eLS/C/O5YCwbaTzoaN0BpKw1zqA/rK210opA8q7QnY6WbLHh6mVV9
0RUoDEKHKtSo/jgP8lXwCj4oapPKNQT5fwf01i4EPLC/dRs30CsbgE4CqjjaBCW8viuCdcUOpFvC
95r6oS1SqMUfPDX93sCDthIlTuRI6mV+wN7+/rATYgbKf1zSHU3Nd24WNPjg6a7/aQoAcWGcJDyu
4QYZd9traiyReSUfO74DXGruuP3qLB6yxZGkaJSQGjqARJP9iD/qw1hrs+al8G/8m3UVdAjxIaH3
GkcIX60TbvPQt6fk/FN9y05s3WKaefK3yzwZQiW69wss9++x+1ICwfQJvV6P/ma21T+YZEJ0ZChn
jrw+4Yn4ih8IBwntet/XTK4p0duhEOtqF5ZxGfS4IgIX+nMRw0GUhnhso6Pv8rmewkzzbKXJoOFw
wOFSzC9VCbUllcEqxL8lk5aNbBtShlT4LuNK40HdGa8s8C2MaeVbDRQTCTs2SUSBVBTofCuoI2qv
/1Vej7uf5KlM0oUICQ5aytMbCc2OReJ3CkEp0xqqSaRdCdI+pRKVMSwAwbU4Xgi2ssgh4CKzRmcJ
GPFTfBoLb9JlwNHKT/GyPRVl0HlTxKOEMchYCeIw0mO40tvYghFwbp8pkSCzAInOQVDECtfuqqgN
pkqcZdtPBG/51puNiQsFSmrQF82xwmuIGCvQyvgZ65Y4/4lIbDPrJ3m0QfbMUqJwjWLiPaVEvD3Y
K0WxaYk5/OYbUo8h5okCxvAwItPc5lQAOlOsQZc8FQ9O3IL48jNAdiYwPuyaFizXI2D8o5fiXBkI
ov71MZLc4+ohP22vpZMzkCbtZCpg+ESUhMvdr67E8zdhJw73yfEm+vzdbIj1lRSfkpXlN7VhXv/a
3BzbjJ7EDIAz4Ou3e5IRM3G1Daidx01VmqHOZLzPnvCDzjiS3kKq7rZM8LmuKgDN9Q5NNQYmqmNe
H8iSbvQ6Na+mcd+SdlsgL9Hosa/EFFsHrbloHP6ql4PwkfiUbURzVNlebfhd9mtuRA8LuJU0nmsc
7PwCfA/Yeb2xVjJ4F+hcz3d1yVY0wBWGjMUMUEDvO7/UgR1E+Sqcm1GSTi4XSRZmfcyWS98kfUxS
jUxQxLyeJuPPDX/XnZBsE0/STY8TMXHG9sI3tbKSih3PVe4HGiwB+djHF6IKWJWVYSA/Z3zaY+oz
TlkevYfOufmKGtuxZf+X7myYRYYG/GorPi9i92jmdsKdMSPdIfrSebJYFRfHTDY9mB/0Ci0yLr13
W8bPavnyUtP2vkOXXP0ztwXwgE/ZFM+oUlAVEOlF2/w0Rm9oBMzeVG+ZZd/UgoDyma1VPH6n/kgL
5w5/ZnFMfNjo8kzToqKbvRJl0qPKurD7jzSbI6IWJp1fVmz/8OAfVpIaYxse8SriXDk56t8xb0SZ
UAeFTtDYBTz7hBUi0X6nCAs8mHR04QkwPahWCDHp4s/dpZfn6Ws3bS32NEs7ewTofJTC8+ugJss+
1j1UNj+J+cre1Mv+EFtlikQS57UHuDdlJl4U4SlsIVb4oPBj/TwFOSVvpp+9wZNyV9vpuMJmJKur
F0P+q4T/jWHvIGzEyPbXjEWagZPzNBaSQSUUgXoDZJmA4h1D53GOH2TthyfnCj+Z9uLrULkTHdie
+HUS+MEWV2m0cCIHMqFQtX8BGcTuweNhAusC8x7hIIpzHmA+i2YnmGTp67nhZeOdBRM5pnvlyvsK
U/K4xTVcZrUQCdMtG22UqiuEjXHvXeK2P/+0nTrm8kAPcP1zfmhC9GqKmpogsittIQ3Wb/RgWWeH
8VdNa3CLjSJOyXBuV9peVmxPLPF8wmJyC+6H9GSQEwOq5DFJIZv00ylCt7TUuSM6yabwt1duXsmI
aiidVQWncuYaHmspFhGcX1Y3KHaXM1oy2a2fklygx4SlvqHdjrz/OYoG+yFv6vCZFX3pGssM1QGc
dFoHwJsFChq/UFRs7P791XB/f9cduN5Dq75LMs6IKt0YxRE1JKQuLuFlYJm1C7xE6NlDt4f3wZ42
M4WJQ2ay9xq3k7rASvm9Gkb6DiUmg/8lUdfLLcGnZYJi7v3WJwEXYiA5ntKA2cBs9Jl8qM8/f/ua
pkAMhpqcnsexZ2PqlXPC3dOD6qu2CTi7xq04xSrBPavsceFW/obnbHQRzPMtv2YJEXacXQpv2DnW
EzPyLvciecDokRLCSFP2UX3g039RO73QG3fLeap6obzzM1amY5VLHUmETsJkE4XVG1OunUdR7bSg
rDf6HMil9nRXM9J+pmF6HuvIrRy43JMHwv38w/1NeriTmro4qFT1OUm7bWgJx6u9UTInT0HKjvSh
/EpTXBNDkqse4GQkODCQb1MZ5YPkUGrN7dQKMLYKzRuFvFawuj3zGUax3ed1xhnrE7n0HuACsy/Z
LB6uzLUmxMTTXSjm23mhTNcS2MTdVh/ghVINJjSddpoAnIdN61BTX2ZnozHpeNRfIxaAzBRZlwln
aW3qLPVEI6Y+4yy6YzclolPbZqtL6Qw0nomo6ii4CSe2lEkH9eZsKHRkzW6dOV9Y0CX6iTylLlpd
4UITgiP5pcECUvSuoKiSugCr1EAikd9coNHVHihnosRxaKWoLelZxEZQfv+y7StSBcr4k0fksxYR
ASRpreXPVqM/5YZx8IWJevEV2EnUTYX1VxOzCr4CVZYwL42DboZ2CJC0qRsgjs+nY1tNiU0P+pLv
Ww5qi7NtVIoIM/BH50Y+alZwsDfsk8zMS2x+VeiJjCLMSE5q1sxATKzHSXVK8D7tQPbpf5kciKbb
eWwEOZqfYxYYXu0ngB3YOvgttfQOODUbuFS6Dnqa89caXEXoHsQtkpW0k5d1jbRLTEqa8jC53Ky/
EFqrTJpCo5TbI8dJD0xPN2sqLdM4cx/mnhe3DLLSYmvo+0QuB7P0VqmdOrn3T4/79FJ7Zbp16oEV
vM2WrWKXkzIcfv6CQZcbHhvZkdOq7p7HYKi8MqtqAjNaZvRt0grE4/KwC1Il9vNcrCgGTYwQ2CVi
5oGvh1NAb5VLsneZXA3bYYhf6cFzzVTaA5nJShqgRm4ciAAN8Izoh/d7qbeW6XgwVOe4DzAl/Ov7
vfsd+EE1Ek52QAhvV19xrxsLf77L0upZbIhqjxxxfl3scGDefVZSHmd3iE+YkEBJcymgsm+TJXb7
eD2t6SXl/BCjQCVgObbEOCM9GQX42CUhNvXICq57AbdG3xGMZw/P1xhJ1z7C1SS3FJshMolYhKnk
i19l6s7wknBIWMB9iLrWlaCwYB0e+I9EjwA75js4v+7sDbyFONLlLymFrFRPjbXsDy1CfM6+TRix
IPwunnBCNxmZDMYOcmPl+P4IDauSA7fPEpeyW314XNQK1SI3GUN7Y/CERASQi+hL75q93l0ep1oj
EUPVWTs8zruczmutuDvEWmZF9DElNwXyJ0pt6VT4moj8K732TuCa+YE3E+r3C+dQAkftX57RARSJ
xPq7pgKWFkUKQD9fFIqbaPw2ZjSatg==
`protect end_protected
