`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
HOoJoKm4NeLYttCHiPxtA116STh074SBQrVHMoa26g5USSyJPJSs/mf9AOpS6Z2SUUFR8Eawd0Lx
2TCHJJvljw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cE6yQafeZkHY5MshBJdAzjhvBIi2YDGA4EW9R+BU6ymxnmdW8wfTdRsyU6u86QK3CSd7FOkrly9g
vMYQxDOCkmBtSdvpzaBeOFdb/N+EV0mt9Z5962H+0ALi9WBFhBlaoqgsK4ypJrmx0Ea8abzHYRGs
jkAH/0+IVtITWOpTZP0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qAhDlk961K4KzlUNR3aaYToYQbOh+c1woK0PFmcC/cnY6uwt0Gezie3pKGFsVyzqeJ8fb0uf4/iz
TDuohF+/gl9BtR9Zd4i35Xj3LwtiHPqpBjwE/PzXuuNodCMs3QYOn9jsP4PLfSN9PtFJVi3Z0QmE
B6sRIUmzBM+edV4R11WHf25WFBL5LupMxoghxgXU2PSLATmQPrrQ4Gm8PPPL0AyIbIOKMV/75pdR
XJBTxvDr0tJXid7Z8ff/ckLKyaUinfOxGBWTE7Mg6h+V2argBFyfF3HuA3R88d9sXYhBlulZVx/4
VxYp6GFzX/svU5RnIdJPnVCxkTx6MV+Z3r/MKg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YXaotPHw4S+AEZatXZK3X8xqSybo1ocvEDi+ZybfF+uq2HScWau6X97qED6VcrgNiRjp45cQDiSM
/XkQjQYraPT8G0vUJtUrCEZhljz7FKLxnPudE43ptH51B0tiroVM2BH/KQhxcoTdqaa4qAQu4msB
q0UjBd95vUXhGOGopEg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nopy6Hrv6tmq6MinTKIG+45BwSwBIWu61Bez8tBobtM3CW38KtKp6cwu0Np8dYKebgFbuVRBgTFT
kJDX9u1Lv2b3nLb0lokBZZTwnFKwKcbouMVNpmlA1oDkUOQOkee+fPq5zpcjEVDEu5uF27ABUx3a
oszqHjAghRIcVQPgJsM91S4rfC8TmK0He04Em7sjnywtp6Ykv/2sHFU4xwzTIUpjW+251034SmiZ
n9OPsQSHl2ylKr4vufbHcxV7zbymLmSb7pfv1lqa3hL4PvrfwHEt3E0H5TY2Rs5hbj9JzB8DwuCf
mi1z3s5/DnKCx4rnpzBIvtMyrdeHUheKp8xFXg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
omtUE89IMO5TczsShD89OT435eQDFnXVCDCD9xXarc1uRWi4zC2tUiosk9WyjYHo/LFxEDxr850U
9zB0I/ppMyuZL/X90g07fQ32SDf4hTA6fHC9VxDPoL2v0EpLhi/vmZi3RBpCDkHgllIHeeLX/dQi
H9W8UddnnfKqa7JUayCROmupurXnfjut85dexXltQUJ2ajeuCCy+4ZXjJPlstY88NdAIjd9Qnorm
/ZCMnpqo1wDYZuJ+EK++owX+0aPceDj5sFrtTQ58NCcm+UE8iimpRsQOSHgBrZBmPRujJYqkeJSp
GMd6cJ3QW3bydhbF4Gx1Fg9oZ5V3rJrKnNXyFs8Yx0WJ1aDBGX7qayTZcDVNWBlqzdXKuhwnyFIu
nAqQlLQCyHCjlklpMKSxNYCZowPKtwVlzSYitkFxSspMN3Msf+77XODy1tjlf42CygcW4u2XpMRc
9eJrn7sWbrcGnEgrQCJyzw2tdgFN2XetV6RrltPEuoWOcq2bdhbIfS2qyvwRxpKjDAkdUYmRXC0k
ktNCYhglLDG3xdBUzsARFjCxqlp53xpcuzKswmbHq+3bxpIFWX1zlTuPUCiISmLtV1hbSF+mcqcr
agQ5eZYRTTPcNyKNmEUYkyfa8jPBaaeiDkiJi9ulrdxrIOMnQ0YsMVhalMeHrwDmNPWANHi81f/7
9WezGHW++aaeSN+iWnIDTArUx6RPxtGROU1anNFb6LDf7My60FbTdi5WGhvHPA+lsrshCbuu3Mdn
LkXEjeYIPST5537az6WxivgHozS4V690dlbx+NToRoB30mP5QXBxHJ2coCXellp7VxSpeaaJlShF
gPpX3DpKWrleDw4q/FBG1hkyUkusUcTSsaKmleUaBOkAg5sf13Vpaf62+Hz5DvrnO7WIq/7jS5t0
G2XGvs3QcpEPQyBCeFsrXjG2694QFY+shu/tLjN3C53ejDo+R4P6s2Cby/pg+nWePnf+satuCuzz
+c4dSW/rqWHH+ordw+0fb0TTXnkacH+AeStnn771n20GWfwlQHd6jvwKx8W07Jeism6durHy1+OY
w0QlWSGECE7Ztp+wdcPhKhNuBO/xoo735xJhZrWWyb1NyltxQR+ognChvtD/pK7v7S4PzZyrbQSN
4JpdTpkgszCn8ZIZlYTN07fhq65F23DPISZM43DxFBFJyXViSWpVuGGOHWs1Psv7VyweJvYaQ9qt
vmujlqUmKceVAIjUIiIuS6y4OXQD/khlfkMFIG1R2ixp2ZupZ1ihesR5zin2IQ5vNg3dIaCo1CLi
g8YfgfiEW0h8Ccg8+TPCcFT9ynjXhhoE5kh1gNW83RAJVy1P/lwORzYbrv+5pB63ogF60BxQ9l83
x6Xhy8B3hVrmTJQ0A/QsbFFTuATwKWw7Kmzd8Ii3n8JCD9bLPxkhd2YnCptk27PRg/nS3yQ5sl7y
g7Ou/o9w6yTpSEe5o9RbWcC14w31+6P7cux/uMVREbkdexWN3Ihxz/WCw3cvnGmiG+9DhXIoaIar
vuXbZGZk1jNBbhtgX5MiR2Jtj9wVGPuZ5zrB11oCRcQn8q5c/2aCbs+Kgr4S4hM3gFTny7sdyhRz
7ZsjbK8UaQ2+19a0IMKzTojA4b5PuC4hS1Gv0RZWzOFgauCXpG+0XIZ47bK7HiKXZwiI31fhF3ay
762TJK9iVdZkQm5arqEgyk/L57M5cN6E9qBybp++NBozKIjyCE1XcQ8Er19Cw4lCJlOkLwqVOs9S
iyrFbZKnmS4JtSXobXPVTHTsQYNRMguko6m1bNs5/xZAQlEy4V7kRqQwP2bKFDsBLuymawBkUL11
1y44xgkgFgL6VDdj4iHoPZ27YtWI5Oawuk56eZsZ8H25wgUm72EGIF6+Flpkx7PZfT6pycjMmiyV
TH9nxyL6qI4vdNvr2GxaJoreANx3iMR6BiCN2WGzYe36zSbhLVuTStZ4FkbGOBYo/wci7KuR5KCo
/VOZMzr5y6EWt48n8eeedWDEQXriDmQBVVNIskXUpHtYUQIlwW/9QqnidkbI9Ozb0X4YrIlrsIAG
+ujzsinTXZD4sq4gb8o9qldNcFiO581QoIn1Ksi7ybQz5jJO2TNR/60MWi41I9OOLt7z54BmbUc+
yO7g6J0vhOfonS/+vlIGv6e+IzmR9n9HkT0zon3GQJEIAndRHSPmSpqjNCZihOOId9GNRFE6zvwL
b4Z/Fq3Gc+pKeIM1U125vx8cHcP9GZulzZQwoouNuz2mc9j9q0YiYd92uctb65KFD2mG8xJkphu6
yGz7pnfexSf/nuaUtR9psBn4OmTIudZa5LJt4tYGHeaeywsDJ/hWj1WQvD2mO5rUbzC+wKIt23fe
gonPPAwtfJeK62jqLazbu/lL/O/xGP/l5PNawyVfxI4OG73nbN+gmh83ycp6mxJNXkTcdzhLLIJb
e4mZFDPZHqBHxkWedzFVgcYqfQCOOxxBxHeoQSVW3sxMT3Si931D+YTNt2MuUBgE5pc8yr/NxD0c
cz5acrIv48kkFhVZ/7HxZhDaRebx5u4kC6ZN4Dto0ojm44G4CizKLPTW+j0vBeyErx2iuTuhGPbk
Dt/zL69C5ZpwcyLJ/5QxBzXe+PBONK8x8Y5oitA3PFuSOlcnztCh582hkegwGVrtB8ZEnrr5pQu9
JWWNdyva5XyQUMnVGxtYKlESOFLWA1D1WuVVLJ6hNinEL+5wOIuTC+34/l1++qe69+fhhq5zVG9w
cp+HkhEx3rTczJ6T2A1QfSII7EUNmQB295ldNZoRhl6nIPhaKLdy9b9W5UKENF+XmoeUbNO0jyTM
A4iZJLoDtJkjM074NJHgNFKSuR+5IbW9Agf/xs/1ec1E8P0TWYydU5l4iCLUHLw3QbX61Lq445U7
XTOHyji8DdHUdTjPVL57G8pYrEHSd81QwEg1LSy/Jiej0cyXflmGiIJBKpnKUY2KEY0jpu+FEpNx
LggHliXKftJYMGP8fvNSGQdux7fd9ppQNIUtEeqf7eY3ivLUQQX2CyR4tG9X82U/uHMWt2xasxDm
bXIR3uImr4omlYH21h3B+SNHfL67jyVh7OexhH7uC5W6SsNPsQ6X6gycHo5Ur8gBmgMyrelHKQc8
XgNq3BrelLddp7K4JWwkCck4aD8QTig7vxzlMA4MAgPJk+3iex7xPf6l0KOSBBaY7l8tHqnL+lb0
zDzphytr3NMYg7mqZ5ras/VcbhMYCaproWg1umc/TcCJXOZYZukumZ6SyMm2bODT3VT3tN7v9HpG
+nx+nh7HXeUhPmG5F9P47KUYn3eBMzDY+W4bZfxD05/W9ZsaJBC6cIG2SZmjgTM0nzFCwrjRawaw
6r72rADTvm6u6cgxsSR+T2boL8PWOoRWUm/LRQDb1bgRJvF/l2i6ZxHmPERMJ2nI1fg+6E6fZDdk
tTtnZCgrrpEnwaRP1we/gmnSLy3DRv860bd9bYZdSsr9a8I2AlWrwDzsDoZ4ZDIL6+Ts8dztv/st
dtE7Ngr1uJ4AK2p+JaLcoKKP7S+ygZtkJpN3OgJmfSFcB0dX+WKiAUemogUnNdrJ91BQU3898Wy+
dEV/Bp2WNrXLHLpoLNLikGXZ03mItVDnLoOvD5IVQPTj+aBMkObQoE3m1fN8FsZwXUGJxodRfGoG
yCqZF4bTambsynJjUXfx60Y+nTN/WuN6Xat2knuw9ekarDMGr+UIk+T3birRqH6CiXjIM2Hcy0l2
a1oWNBAs1jpPOQy5My1gsTA0yOcFmJrZE1PhIJRwb0ib8XiwYCg9by1dJunz4bryS6vd46VFjCvK
z6o3o9M3mCm/ylZc0FjUOPV0m0VDk0O6vYkTjxRrTF0Z2HQyoFr5tYCHMaEgeoHf538Dppm1PcUb
IJGlRu/C8fuYQ+a9npUICzhoSI8NO//iNDkXGVaJl+e7pSfF571kT+m0HDOjIU7Tm2175aNYP0yz
cXS6fTge2vbQAXIbIlbSLJLLVhPvVhxutp26r2s9ZP/3p/MH4bEyShAGQkyvxkyQgmOPQKYkVmGg
uCbDfI1m/5IWUznZVGw51cQGg6C4SaaaH+80XE3fdplr5oBuwIgUqTbShiZihIH2lkp4Cm/CPeZw
6TuoNfDjDfur2Aam1KSFAuKH/4GekzDl2fIPQyS1U/mdUbzZZY1+1uiNZSrUIA65k5VpME7tJ4qK
dX9y4eBq/MsqzHR3nb925mUDu/hP8gsN8yZ5Pg26QWe6gNoTMd9oEs/PWdarir9Z8hg6BcikIp/y
Pj3ec2ajKwRzuFlk5HXSYMQnCAsfBsCdx7Q8+jApNDvk6acZB6Mc6UcT3m7OURcPHaC8a448VMEi
s92oNPWiPO+4nn+R/T4kNNjDpANQ+dhTm2VZTC8iYuFYKCAbMr1lwam8NNwuDhpPDJFrDbEB2U3y
rSdeixdOmMBxsTMuOuL+hVDXbjK8BEzb6vqPSHrCvuuZ6QFDo9C+txDvhCUxvA5DREqpFu10XA9y
AqqWsw810GGbmIHnvmd0hq8C8NYdfFIfroK4mwIQpB5PkjgkEL+ecmC5EgIs0n1n09bpHzvBvU5J
RlJhTa2JsjHlqjiPU/Q7/XmpzOKUCW+0nlA9C19G0w8mcprq0oOK9ZBOAsFxu/EivGsoyy2Ki4th
IY3uUnF+fqcMCpYzDgCMIL0efICMMn4ldcgG5/jgfvqBlXgqZcdYfu83TaoPbCybm4yQRY5TqgNW
Egn7YlS0rWfZlaJk5SefDknXzOd5Oc7w12Rt5ZRkdzqrsuf+pFFcQqXplBENUhvC50f/XBX86x9n
FpHxHkZGJ0KDXGRA1sd4oUyZ1KIfgkhtNphy+mcPyzUSxMpO4RCsR2Pp+TCZnVS/Z8Lg+3XKVTiG
/4gFWTER443dhRRjK+ySEy1vn539NNmBqFNzIo8GUsMwuXnB0VHsFsOXaPh5XAZn92b3a1IJtwv+
33gjvCf9nefj9z3n8O+EYMEEgcugiBv51N6XJ7fOnfi+Hufx7Elqpscb/Gzp3OQ3nUeJQIGYXsId
yLom+ygF6APABXCtu92PkQ2yLuQURK4XNsEP7QyzRfiyO1999r/dUlRcUBal234xtojF1BKVF/a2
SAEwe7l+AyH7bqghDuU8osrYBylApZIc1QD+bvdYP2siUmlliwF3p77KzOEIKw1tOm/xxTCjzJgZ
FHfFpeug2JcS5TIoJ4M6dHz7okBvYTabDrbMdjjurIWaovGGgz2YZ9m3hVdDxb2tRMqpbbuquP1U
Xxq2tLbP5HrpTkfywvGhI9r+13xKxI1z74ZLylbOyE0lnU3VR/buT0hEhVugndVYfLPUkivTMIKc
vLpoWMpgxNpWd3+h2mh5wg3np3teZ8A7cXiEmYxptQWn9pePm/hPiJYlmd3/eeBHq5550p4F/0n8
YRA9iXROzHRk5h/szxJoIwOwBKajW3GNsd/ZtAOqzEunL06L5vazc+w4fiXVnnlol0TXh7khEP+V
92q+8+4mTR8W8MpL5Kpts63VLbAPMKrWQRHyx2eD02wcenCff2CmCuozjlNndIMW8BhPlghmIsdS
M9I8MJMXYFgi8xOkUt0Ruum5+R8XxteiNAKa3qkb6SSpC51xys5Oa3w213IK2W3sNB31FbUZFp7a
hfBNGwV5kwM6TWOoCMEzV+XKMN57sIHNmzj7lyO2ZGqWFURd0E4Wia1rZAqH7mZqTNGhDj5sF+O+
bZzR0D8ADw1O4mHhAQ9sYZg8ycAMDI5T96jJFXqqJneLig+YhtNoDRk+Do1h/vjOxxBGxztiMVaw
SAT+wFQWWyABrwQGHL4ISgjXf5klzMy5ThIqj6AYLac1bBvakb1zyA5gaBCJjY7s9jkFlOszDkNn
9s5FIW2pEakRg+PwI+SoCqvm7w4Kar+Uc+ImJhLlvc76Sxx4BjDFK6f5AqZ78ifNulSF7dhv4/VO
MjATkARhC1muE5jxBGwh+NGObkUzz1tD8LDMWVgmTh0SJII/2fqmRh2967HhODIHcIgThUnRwNRK
bQz65p6LrNxd/VH/917yz0NTQqwV3uJ4ak8uoc9jOGdtqli9LZwWWLBMiMC6bpBJjpVDWzJwIFJm
TKShzamDzerXMLja0YhYATNtEScSfB9ULWc1Ml73sFeHJDBepbTpvOVAW1kYNRvpjka8ktj57Ovt
uqZqTfYS5LPm42PsRqpkbiy+aVGDTXqgH0t311hpkKgktIgQQZwZP2y6AUwnQA+1w8nvifzJtdiF
SXP9kZiPOPzRsRMgO1q/9BUgq7e73bRdl7/X0e03xGQbKEaRuWV1Q/imsC4IIJ/I8j2FMHgVmmbW
lFLbdQfuohrO1tL1Yc9HZeJGB8oTl4NjB7LZS8bsg/lBlqo06G8EyE0rAt5aXpj78QFr3M0J1T1j
8tDT7WxNjxmGKbbl3bh41H0jIMJVu13NT4Sm+8itq11dzpS1Emg+sq+OznqEJFOZSAGHL5rfD7ov
J1x9d5RToa9wbIiwi6lj6aNd7n8efZ2tU/iwQ6q8xApy6ShemgaonuAWm23J7cqp7cnme3deWgYr
+LHbVEKSZ9ZRMQ3rGfUd4fSZQclOFJj8CJVIIqDriTSEciNBDGSqLdkcfTJtZs780bcUU/taIog+
zQ8HiJ5b9V4KcntSfXISjzaPiKVeirSJu4nkKcNBejSJ3drN6b5mrOqdeEep644qVc9fISY3ZHcR
cvm/I9+ZzH/0XNaQJPb4KsEs7w4N/EJCItaI1vI7ZAu82mMCkjVNYksMnFX9kSkmIq2VeWtQjWei
o9tXSSI+q6XcPko356BopBPqjMbHDnHLB2HClDZXQdUxC02ji6gInjApFdol+o/pDPyjhE2pSKRF
9ayW+PX5TpnLIG/WtsubU0/Uz79/73nMK4UpXESdHjHhcozPH2KKNMJ2mgy4nyAYleRs4Hbmt4aP
v0iXX2VUmNgVAE+HM/3nAAnkwQ4r3XftqMpNB8klfqlfbNOp1b/DoBtxeWF21GLVk8c/GEQiON0P
tJxCRXC31/wXXXP7p3z0LPng8Z7MNUOceHwu4zBze/au/Nb7iGDtaDq3G9q0G9E5jhBWTd7TZo7/
dFt4f7dBU5/2vpIalku5LvKMes1g+XZD+wKPBWXLw2eKX7UnwFL9Cs+tJlI/fVRP4jbr3DOcH14/
Gvd56ajZ72mz9f5NjFVw6RtGNfC1/TPXx9Wy6Iq96QETewE4rRw6pnxdyX7fgXifGNCBvp++8Uyo
vz/RVmByTpeNfB33gg6Uii2TwvCfYczb4hnxfUD8hAP+I98fv/N0l/DDasrYs1j7pd49OElleI1Y
uXdjr3Qk7rtCAie1T1Wlpqh+Jc/IrKOmDPY4CslWtXeVLZ1Z87/d4X32fpqx09+LUVUgrz04TQWw
e/g0pQVoLhLT7SA8duxnXNTCVZ5OqYPV1BKb5Wuq0BJA/GffiawATPZHHMYS5dQbkv7NOe5e04Sy
C+2SnZZ03cB8yXd9NzGZdp+rz62JejQQJeODTDUJuAtgckUsJ9A2ccUuoRaJoM03xX187rkqhzUg
UQA+jbgBDJtzfl2uoP9G+EClvkuPaseRxJypduj0MIEasyVkmuDhk/Xlm//Ql7q6ul0vDP7kJmEC
7DyKk/bkCqFWUOfAtITXJPpE75/t6qb7BiRRz11U0epbSQ1kLTuvyZ9tSBZwUepsCq6xLx16cS3n
qH0EWp0+oqNjiUZNuFv++OfZYYLIiQToiQSW5993ikny4gqxswRca/FmL8tsFUeO8Q1VENdBJQU2
Be1PdxzbdP18n7uhW6wkv2Ke0Pp2k8yunLabH2JvfWOWgRwvdTS5j18P6p6CyRYC8MtO3T5AyZ5f
2fC9H+kwBIay3RnN3YGNo/8SnGJLOZehqtFvneYOq2Yr4Xfn7kYZLclmYD/H8NbaM7kDjYG2h2gQ
fkExAKqzJ0kv1btSOvLvBx8ohhztLUbEzRMSmMw3XITo+fWSZeIsgx6DWh3DnnrLKlKWjDyM9Sx7
6m01503xlkhjiaM8o596eOSR32bK4zBo547lWHlZWm2x57zxV9jyBWpiR+y6K+SHf2w+j+xjidF/
PlKcS+RbbyRv+KkbRm941jV8BrtyYWEVturOkl87h4ufkNjYXu5SsbOLb69Me5QRp3JE2GS9yCmJ
evq4M/osQyEmn2tibNpjDW4o6/KlG1/gYOirGcEqTKdGTWL1tcWDZ0snChfsr/k1/quNCevPA//5
RKYi8IHFQPv2sUFvHTqfXGdUm3oPZlyG3xCDloXoqEYCl+uZ6r2PQem0TVoYLWhjhQSQdrdGKuPs
rUx8WoXZAm+K6eFGvBaxU/H1ke19oJ+pwRNIneDfNx9QIvGfkMi5TBrVQ3Nsb4C2VYVxKCCUIC0V
P575vnzvWjJ+2eDctjYMxE/8pmTcomZlf3BWRVJDl6a/jH+BpE1s0ul421BTKJwzrYz9yej0+uxs
Lv1xMOppwObkSuPVrolN93ZaX4Jg0JHQFD7MI6TYOqvtdFznO8LjrNmnemtP+JegA2yS+hU3CpQj
xcBoDBBsRtmjnD+wfPoPTu3rBwRu1knx97wIpZ1cyuaCEbOPAkv9Uczrq/weWnqxvQOtfRJoOG//
IE8XnsnDSQNWv5DvlEYQvQoKiSau4s48l3vZNHE39XJs9GUgMe3rHATtHE3smzj1bDjlQhyQs280
8u6O9ZWLQsJE+wZc/FUVElNMs7CQwLNzbG7Z6qKcPqwzxiCePwNrRryMdTMNBy7lU9FVUhl0UMdD
iqXHbTzdeR7x3u4kQiCp8BOMLz0ASWygIy0sHrILrw4kMq2xNwYo9tiEfQQxT0eqZUuaMr88tUYI
9sAFjgoBOrKQirJTUjvsj0DfLmoQynN8CD9a53n+WH1+oMd47DgvLI/Zv2ytHfYaERMgT3G/SZw7
NnmuBgqt7KBwwJVKTKSt1bQ86MJ9ExKaPU8S48eaae+4QvmEnE0/E0ZkzU4hyxKXV4TV/XIyjnxB
EDzBZTEqUmg1GzPlmp6Wg/IpVwDSg6nrv4TD8mGDxaullXIoHs9OnV5mVu/ngXYTkOmGtTMo1ncp
4i7dfUUUMs6XN0+T7b8+Cxay4JxtZV81JcOnWTryubdSBUc30MIMbmTkQcdaIxwGY7+2O8phgZBq
3RupyjDLo65GtMGczex3ce8FYpzDegZJ2HsfMbKFXLRdSf+j0om4bR9jIxghXG/0vJRocFW/Egjy
SjOp61m0CTonSFfdZRYLtrPgFZTKZjGRbcwzdUxy7GYVBtDJo4950F+9BdyETPXd5c51TojU5Mp4
uErHiNLQECPYO16NIbEik3wrqb1Jr30LueeowG7aZXQgJJ1AsCWC/iok4z49p9FIE4kY2VyxngeG
xBYPBUjggo9OS4x9eEe1zLVmTfwvElouis5vnGHaM9UXyykET9fq2b1nSO8gvRxzLNW03F2wxkxR
X9KbUCFAIG3xVfjiIg1mBJ5ol5CnR3+zwftfg1p+NzCz1/Bo2ySZhJS5y3wqU0TbOIVm7rET2rtH
/1TlK2uy3h/qhdvPlT4+mJy9CvqGxELvme8p9Fgufk3t4NhQRxH5jQzFL2aAiNGlmSaiDAISxHx1
BbQ7UodmP8mq0ufEtDSgtH4CUNWipIccupN2Y3VdzD/gD6u88aeajtyoxjTEU0aU6jRnixpAWd7+
1WL+Kclba3NVb3ZvUcmtXF9zM5dP4nKUfPlPQXng5sDQmCWVhNRh19hFfwn+b2UvBlkJr0SMQE7l
HtgkBWgcuxkTSt0vIZc2fVfviGIy85P74VOCoYedl8JdYHFEVSYlr4ngC2dP4+BPpCq/UuY7QHnc
11PK6eA9qE4NumahfG1dYWUB45Z7dnOK/H0enxRdafHaVxf3hKWfrMUcvVM1jANnNVURmOeTDqqS
4JOTLL+2WHke8cO0obmZ80Ehb241pSXzTbZI1cSlUwJ7dFWSmPyHDU53fcoQGENjC/sqkxaxG0+5
lX/AqEhqrO8sw44nL5FmvnMf/mAiNb7nnL94XAai4xQ8fKbXBvN9gHX3Lj+aec4xE0JD6JdwwgNb
Oo1sy/rCy4omKASbbc2iyDDsoFt5F+g+dBGkmnEFBCMS6Eye8PHFKA8MaIaeg+tfmORy4luwEdV/
ObrJdp8WCS5dvpsaQ3ZcoQoHAP4HKl2Y5zrKMHdlFU6cy8BxDI0OdBumHCZOKq200k6ak5sqJUtS
9Jchf87q37y3q2N47NGCMLfxCw9SCh8yRTn4Hw3bz18EnqKVJYHe+jb7yfggDzQA3Blh5YKED/aS
zQwM/Geyg20ZKZPx9zJAdEJdYAuulaZPgIuuVbiBDPCzAdbd+mjUsB7y9mbcifYfz0lMt1uIYjFH
S78eSapNZMIyzfzafpCWaIzGkrs32yo9JS99fqjmeoELUFc5moKLg9eyGH9KOwij4GZ11lWRD3Yd
s46eVFrFHesmJH1bXgzA4skz46t2Brde2CXn6MVVcuajj/qQub68HIlGoqFNDhEc91m6FUPYQNSS
h8SG8UXl8Eo43dp58ow7LQO8Nb7G6TOmftHKeWThz3vbBDPU1JJ6/kYDOcnOla+0JpOxJZqL4hrG
/8Ir856Kog+DvcT0QjXWT2FiriQtGun2crrzW890D+JiK1O8bAAfH9+5XHFF/2VDzZQ974u4wb2g
c8fNSgVDPSOVCXLiqmFa52U5vMNYf0if59pgMjZKDfiPR7SqrQ0ca+28WDeFzpSaQY9FJNHSbECg
0uydY0b7tyUGINCr6NTHTayzNgkMOGUyNA7SgQh62sxse0kYptJ0/HpMpkXZaxXEIZ6afCjjmJu3
1xbR66RvIGVfyuITuElHUwT073l/Jc6AX+Tb4ruvEuYZTjiFcv8GbrKmyvTTODmkelz+Hrpkic5f
AMZg0H72v40CPewhqoqItSHniGgmpOZBiy8kiAEwFmohceL6u62qBUSfvp2eFg8AuGRh4rrtjtTn
Pdu0vggMLg62o1SYSHDW4fO3jLChbCXx6feKS+gvSnrZCCmSZTUduIOQ7p4DhH6kK9mCxKfI4qRz
3OSBaD+6etgeY9YCHWk6i6p8DSEk6altVlQe9S5fpswFHxGg6/UWMpHXsgY4MnMTTlJZRXEYoOzw
vvpTgNwpLwl+RgNpWHma7ebRUn7fTLwxy6+nnB+EwyIJDft9++UfJBvyHBa9JSvOI1iSPMfrYEO7
Cmkdf3/PlMqsgTc1hp6ltXnIBy4tRF0nua7TZM4MtOEQ1VmhZljAHsjPHmC+Hd0jLZJ0XFWeSK4K
ODhXwFOwrb6pw0xAYsJK2pyo/iydxjpwGg6skBkQHSl2eVPaFo+Kbry04B5ilnsKXP/C6FLWboIO
vwq2Bc9qytpu4v68NZ5N+KffDoqYuc+wJ0ZVNSMX5YJSb5QULA+szqOxjccVJrlnCGjkf7eqGQyU
zHTVuDqQO0n04ropocHQ2Uy2jD9E+0M0at1C/wBJSP50M8gBtfHJPudn+aHxLdg7CiplNdK0P06r
79wUEN3bVpcLcqV56w3FNOjhmjJEGjpPXu8Tb92yudy5+B5U1KUpC0mf1ZZjhMEkYhJ5BI1HNZJy
5qoUUrGJQqToneTLwF2nP6uwsdAhOu8utKijoX3mgpOfc9BQYsp5bT0udA6H3JXoNdDS1edefrYZ
/NYCrfuWZG6Bcdjko0PWWSDlcWOlHnO316IDrn330u+q4TBoyX8lY77A+R0ujZkchcEUbkgtm5rA
8HcaToupzvoX3LIUJSA9hFVE17UQSGIAoggsTYqJxgwYlvspI1x8h5i/hELSK79oqzS9TCqwhw6Z
DnOHT0AdKZWrWZO6n0z2YM560OB+iWmrcLosi0pZ6/+y5sC84k35DjO9073Ev08uwKiXUX5crs3W
3owg2qNd5vClWcucP8JROrXvVq0j6sK9k+0SoMR2vJJp+XaOzkAetT4ZsHm4jzgXRB21tffjHiu7
yQP5SbK65Y3YZX+mJPNz1yZ06yV1C6+u9PCJGs/9PPQmPOYxFeVOoEXxcc18oAREQPeLGjUPq3fw
zE7rhkWCYMSazdFrzUE1eyyGEFgQGtdOCiuvInFcVTYH2+wN7SUtNpoFQqaC+QKzuPZvqP5Mcc+m
TnKsJHVtWhcp0HQsJkKwoGZxzdhgWTmJWdPh6iC4964gsvd6q5iie4gT4fMSJMmG8fXqKtTheV8x
8fSkkOwbExvVjHvBePEMxJuEMQZmMuxiiZQOoGSpJxDXYHblb4xgApWIFhbypGQVXQAd3fHEDXnm
BS6j2dBI3BaoTU0dspSipVnscte1ibJ5e+YIUkxCCTU9DLSN5eclpym0r3gb68zSxZITB/9GeJhZ
7DxNd0fRpmvvL59KDczongUi9uqCGeqA3AHQ/EEd1PF3wnawaW3LmBNWdqeFw01rOTM5XpNyDRAi
vELfpbjqIhhPB3nTbaKoxljoCOaObAfq5fM9uuFgrGewDtTAwQq9OuTVrG7HjPnern9KAo33Khc7
3GXN3MCcugHuJeF6JaVYLT9kP4VsYxoSvKDvLpSwGvzgXTVUA8UmHkKyby04YWclpp588OJtlTl7
2ymiih3rp+yKDsbDU9fxEaN+heWfUtHZgjKSPbHJBOH1UF8yvd4CuCy6wKW4v9k9BefUYEmDhN19
H/aypHT/5z/9cFpCMsdBwhnk+LBXLtQmVUqaclI4MByE+Kza9EWa+R+PaV2kf+DdkIMjV/XoE2/j
OFjd32uREMLmDtOzmM8enIb/0O1EdZzA/dyBTlcAIxRnkiVuttPfuznkyXrmCoC8U+p8TQI729d0
GlPLPOOBjyI3cJPY8Mie8C26VaCy8t9IVyQCuAnoW3mL/b+qZ/kpNgKXn9uurAoN13GBuTpwWHeI
GxbNv0sjAIGwAZmO83yDRuEVNYyco1na/QzpqLITCx+cVMk6oJX4UdffKIEyUlGvrsb1wD/uiWOe
j2mUjVMNURIENCHKiijgNrn0UWJvzCXIB9Yi8Z6VwA4WjialR28GaYLdXROx5sb83E+ntIR7vjcP
qtdu2NNN7tGSkMh0hD6mTWyymKhu9+FPyDtepR/lRcdDBWYr+LxYnn9LIuFTIDK2BVy7CxGZXDYH
TUPTrEmGJpEzDElJ80lTmxeWgiAICgeAPKCeHwajj+sfZhtqtL0R3nLBLp1OAeAU/zMLL1jdYhPo
c33/ZbeJfNjHdTN3vsbT0PAGf0K/ZmdSOV88gZvy4/AAZao1gJBhvTKqftimXsob2/7teKeXCCRw
mdtDKrqTti2aVYITmBmzw8Rj4f3cBnBwddXPyhu4rG1gEWOXxPZdHJKqUMMu2MkXDILuIDCtigSI
UXre+RnO3xn4mP46BRPgpexcycE9TdISy5BHEv0ee8BFyDl8F7YZpzM91vA6MPQ7uurHNKrLGaTf
cC6Lb7HM/DDRWXg76ePw3FjwxnxEUpWj7l9X7Ra8NZIj1JwiiahJP1UTJ2i3sT6Vtkmu90oKgCJu
69LB9YFCR7RQi+7CLtiRS7PnkjIZ8XwOOmZgqNhKdeN/s5LRyHYdVzoiH6SdeuHpW2bMssuzlR+M
Y1I18FtAiBclcAy+hajZ0kgLW/3T4jbHEkNSFk7zMbsSbFikaZpFSxXcODaah3LTQDgRerGd2VGi
2M2HWurnfIwrmbi37Zbhdqhkos1aPm68U9y1pI3ojto0CC/YqaF5JsJHYYs5e6BUbMal3Vw6CNqA
NTAOSyKtAYwyO5t4NV/gSUjSxKz7rtqePuc6IcJY2zICYi+nnSPY2Kums4ExM3IVqKkij6ZKNb4O
4pt+fqC5X/IxAjEkGKUTPpPFMNX2SealiTzsga0Nn8PRZx3//C041En1DAgwftF9OCPX9zOerNtZ
VOfjqE8Ms9m96BYnslRYc4cSAC1pVjV1f19FSIW72tacbqU3QhgGAPfQoRB165L/+fNlhuSc3MBY
2xJyMOIcIivBbmYHiC4bLJeFmEVhW8y6lQQ4522rGSdrcKX/E9YBAfo+bcdhHjDuG4n/6qxQ7wRI
IEvguHzuvzHWPCeHcSkkxcOSrESMW1ibTLPeI3HHPv6oNZk184WZ1Ds/mA7A7BPsYKihNVgEQpp5
hMmsYZphgTioa6SSC2rjdmj7upigzycJnqR/ijokHyf4CI5AU15ZO9nCU4hMrxzk5b2+Zb1Tf89r
FwPN10CHu60mfjaYkIeMcJNu/R6FWEjzEw00nC/4KTKuSJesxdcOY4qiEV7fDqaSl92ka2RrMY8Z
S/i5QoCIo6XvWn4YGWGf7+rXCGe/MO0A5c8lr65jfcEKrjEcS2eTvcJTI2xyorRmfs94zQKaR4dW
nISWW7wK2mxgKbtRsMzwfQ3VKcyGKc3n9cc4GDqNXmB1BwLCnjkTle03XBZ6WPpGpOL7KsVcPpv4
PAAnF62u5jGVTvODlqY83kadWCa80+pBULzr/jLF9odyyNAbJtacp5oEEMrY8vczEOa5V7E6FX+a
qY3bIytcgRfj2sugoDZqYU/LrUO3tB1y8Rpa8hup/Qo4SXrAc8RRskvehoVcV8n7ozZ8CBTLuDGZ
jzsxkrK9u1E+u1EK9ohxWBPjibgwan/eqxRfoCbY4HXAnwhLTysrbDYf+M8JJBoL3sb9SUwCToSj
hk4v1hocOAKDKMpkgByn6Y17qzErWvgvVfZaUbRWVSzg29FChJ5bKI2g/FxtNUZfaSzx4U3ybcZF
TAEkbOLMqkq8Ri4+jWDcSxis+rZdXZWe9i+MvpMZO3NjlQcJf2D7jIoOCYAca0ytrlxXsgL3F3Dm
C3YBHqewyRhvyl6n88t/T43VejOoL7e4+q+o18bHGwPwMJ3zIABnn9zPMVXLEkEYEjBdgayGfdzf
O/WCWTgBhcQytjj9/9qRvq25ZmPZggOcKYOShMwUD6PvP6SVSV7f6jwTTCzCZpQvHfwlzqCjNLdP
27K+DqkDSZceUKdu8cOfWqMgNw86e7l99I01nJq1M2zz3dPtlf8QQU9j4fZo3ncgPgXnO4N5VB9q
fVh9Ex8AAtXL/hAwMDZnH/WlMT6AKgHJX+IOvTTWZmm98PPPYkpcg3gBFA31ngaV9l6iHR/RMO0W
X+8awjgIg8d6OZVXoDtdt0R8Ix1BkxXbTtvkiLqafrbptQPJ/OycdbdxRd8akNh65eD+BFAnFmtZ
77FPeTwbwpY4wweb8HisrLfL3SMJEuAHPwkZb7ZsjKATMDZEXu6WJuw69TRaPLebSj7aGOjfy2mj
l+G9W1I0gzzl4X5CapQhs1QzeDmnFevVZeOjsj+QtfOhygOkpswotH29oWQ0gK7b2SizkJcPKWws
YFgo/MQAnBZw11gFRZSRtvoOJ0sjT8ojP0REH9cRiTFQk9q67Ktmj1ty7rLvvGr8GFbUHqZyrNSY
p2vVT6qGxnhNjnKoLdH1zbOtRAyRbOv2+NpeCFLQriSrFgTE9I0xPuz8CfRpGlcegxFl0zYE5ch5
M9W0vayTjCPuLvUGUmP/WYupIC1dKrQDs1ZBwIuj6/lYdcTrGY2cV/NoIrwhIzupR9Bdu575CLmo
I86VqBrMcTTY465FQ3W9bt0gDBOFTiRy2PltypNf09m8n8j97XHCa38/b4bjYwQ73/ZuoQ7h5kPn
gauKVs4G+uOu+3UZRDALrYPVC6hEWbGM603jxjabUARg6yXqJ8VOdVuv1d6A6M3xiFwN+8qcVLVO
xoEc17ERKdxf+iY2AxYOTqKySl/zE1d5FPqcfggvCR0igU3F6FPGls8vjw6sHSioRVvlrRuKewRB
SxGwDBZviFIIZTSx4n38LdSg2rjc/uRYrVEHpAr166vv4ZEQEz5S2K42t39CecuEVOcpLkeJNuTE
vDGpGIQyPBUycNpLIfxoAHPLgEkZhsqKd2lLxHDnmrzG6pkgipTzUq1AuQfVBkDVYu4HKTtW8VAd
dbpUMB05gcYI5xMXsBsFzI1rzxTLS5SO6fa5mysG9W9aCZ+S89o+kJM6m7k/K9yfT+3vexyudmT4
huhNZTygHz8Gvv04MTDEBb1O69AMeauFfxINceb29685ETtskbxtwm7EIY5gkeQy0Y/8vyM/O0m5
vmcaf/CCUD0naxtpmKSmzSHjI86z+rCPG9D6PBoUFU9hpCxO8LgluljSV437/remU6Q25xj8jtus
NHncje5d/dAfyrZ1LqYEswI7FKklAWM0dXZyRiR2X8Rdya69Q+E1NldHNq5sdEKkuFShfgVVEfux
3aaW8AhivgS39tQZRGhY8iy3RxE1F9ls70Bdtbfx9o23deILNdATwTD5uSReir3webperUxE8A6t
hJuUWv8ZjshJKhjJKJrACz6mAeHb4pgIQRSGHxx+ajVuRaugwScT6fRM2GgLk3vNg2CY78nqzbCc
h4abtgzg+IaO9F5aAWwIBk3UWEXsujUyGq8UBgA3TnLQUr0koJHMBcxFnZqciRNi4TtPWBZ5ZeEc
RtX/LDa1ilesv17rmP/QSownj63HTcecoOpaFKCXQff2Xb8FAJeneIgIj15FcOMaOrQQC0Hkr0Fq
JdPUb/gFTKD2RCYISaXllxlyM8QPq/UMSOiwsbixYXmpMHVhOdKDnJ0igTdxfbJ4qxoAot0OsVD3
fr1+4QmWBSEelr30HRJ0dvx4583rfnAdw6J7JyNHh7OY4eEVQ3QR7hUH2gm4dkidZewBS2G/szVG
Y2YWWLJ6l3052x0zt7uO7HdnH1KaqRPSw8F/Y0sA6+JFQeItFX6pc9c5611KVsXhFJa9ebcIwori
jIlgCePwczv+mUfXTbThv+rFzwiClzDn0LEFwokeQEldclSO9vaqal6x0vck1V1zeaDFNIyhZ77K
lAaKsWO8szdtRis=
`protect end_protected
