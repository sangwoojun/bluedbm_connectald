/home/mingliu/NandController/src/ControllerTypes.bsv