`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Px69Gw+ZL1VDfZd/kkftYwmA5j1zVDFcBwubGWn/wPw3zz+3DcRreAPTP/2M0TSi8aXL0bWrDd4O
qG8l2fA0Rg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WTrhrh8qEI6Y3jEm6xadY9aq5OiyBPNYdBnqtmM5eUSDddG6hIRf2g9VunObrK8pnMJcEhqLzg6e
ZxMXaLy5zEbQXzmZMPJUaQgGIrHyqg/gsPS4VO+3ohWGrYpoFeRvzsHybVZEFKppByAyi8HPKvwz
Xjfvhh9705E2ZHog/ro=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qhk2qE/SyaRmP3Qja84PQG0cmwDjRWo/xZSvMPJO/wDyrzf+/pa9dc4o4VkAhyKGike2YkISJStC
2vDTfTxEOT2SS1DbN90DtAZ2nhK9LO6jjf+IR/TMasTSLY4iEt7zJOYcuwDDKPCgzczViHfYVT1p
cv9rSlUglR/3IIbv3Fhuzjb4+lhUyjeJxdFo6/QxAypwQzbP/8CIGP/JVWFPjIWLxTRDqrXlXeqW
iT1NbRiw6R0DKtaTLCyl/ddVl0qCxkyz8mjPvgU7cakxZKMiTsBy+RH6SDlpfj7MT9ehvYV34C5f
RPc6gsmeVo3pXLCiMlWm9Oah3gDkLj+OkDOg5A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k573soHMbF7jjkhzbbPzh8NfmQTN0/zgOa1MdZG4C+55R4BX1zpWgQMZFzNyxNNhsZMYiisI5xZE
Z2WVWD0yn5OKFAQ6PgHCVaPEmh1ZoykNwI4WglAAqi44z3Ck1F20y9GisekdcDXCguBNlRk2pzqv
FwvPemcLPWhw5rOZjPI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R6nMS0fmmT/5SksjExLksbtdL2PDC0VYps/LGB3/EgNYK8BLFTTJtvdhxKqT047hn9jqhQ1v7HnX
bLRBAvmBMNU+djm18VMK6M4wJYtshLl+UTdvGlevX9Y1NqmiyBWEeZHMLLgxQwAY9bmXoGeiERxH
welz+7B/hSeO5bCegfdMgRjeWFZ/1sulQsiwD8pJfl2LBwM3pVO5coNN6sSzWh5VuHT26FiOIw0E
7fl/8p8xLrRVHPnojkgGN4MP9ILJOdUCuUhKQfWfmiGdecrcVtCgDseLjg2HHBsWeUfVBDROwQZu
3yIKzPtTE6d2IGt9NUtzPXhbQnWaMWgWDfY+IA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 41056)
`protect data_block
/332lgOm8PyC0hcatsylrEs3i62n+CrmtdUnCcR9Xd4V2FYIa4S9wm9oMHWJ8crOwuVTUcivG3zm
AArRRLIkoF4GgEfU0ZpHpJNfhj0uLZ1Br0forAgetdkgLQxSOisdh1+NsjPBmppFvLaP7RSaztMA
n0EiP5HdDdBY/ZQ+9W2Ma4ZWsmwvgmrQvcUoBvzr4+eSxSMJERbKD4jsw9qi++ptKhUpMnDnJfzF
gsoUFZ2lDp8bHCL/wyTvJe0Q8M1ZmGxgg7uRj7gVV5/c6MaZqCwjOR44HiqCfiNMezDrqezD/UBi
X+YdD7wp6DggcG9kiAtOxvxEkEHDxGXjEzrPmiKkHF+ai+NJH/A/RdabOhcVKBCDURgfxP0Y5aEB
t+/WlGivT7vJX6lEKwkKVH1Hp9uh2JTR/Mb8mWMa6LqyZm4H9yKfFDzyel1MTqwtIXW2o6dDonhD
Zg17f9xQYJ2DPYXKX7qnlyxSf3OQb1ltDEv6mKDKahGw6qeZdHrP9V9G8Uyq3itq9cWS1xkWcOT0
je03vW0MrYVP8KM7AmG2h1j8ACNNWCP8lV2HWBT2Qbrtr0LHmHfR0hlGHPH9zBQpxdE/vWSwFy6W
AGleDxPZ0ITBsTDbLHBvuH/MVlGOLnclPcbuK5q10oia9k64mGMc3uT8PGVO1I4msDf6KspTLB3M
ZcX4OJz3pQjJroO1wv0UobMoGaHuSjwbOCnUThAJaWTNApN58YHoa2GKnomGMXKUmePsdwYmyFXp
BX2A75nNNPf0+4lFDfzAsAzZiGpS+r2/JW8EQeqHEcn1dV3lY9yTuXCjw6p2Ib1QUNq7119SrOQF
3M+NJrrFstFD4Dsoj4VGEgS6TV80JoJeHFXniZKMl3E1mFmNFUcsWit9/VoxoqCcZsRoVXnHTV2p
YyQMysUbJSQKp4MMT49Peu3+98bjm3Kgl/7HOUsTLeibQCSf1J8Ud1DYU5ijoy7XNO482+J4qrwS
9CZJ80U3N3FWVBcGBJR3Vd+KuJ3P99Ese21vOm+2AqaEw3IGbIebonJaRNFEVHXlryQmiLR+zIG9
b3pDqp9WAxGogZUkwR4pJ9daTGQUv+tS37oaM+2Nivt+S1pRjEw/0bWqrTB8jkv+pilPT3dLpJfs
r6XvJ4HIA75JJ+LqZDOt20FAdb4xNP9oc/SDlr3aLkUwCCs2kl+0a6dofIXqnRiLdiNQPXq5bgVo
YEJU1A65vSwjgrvX7vm+H6U21jhdSBovm7wQ1vBHyPqrU4NTv12XBTH8RaE+lrR8UDcmI9QZQzPM
pj/wU0admXxO+cVqcOLucLaiKPJHZen7sZxGBlTfRF6/ME/0U7yRb/DeJcpFWft0jcfvnMySw/2C
zlhkIGb8CJ/xcOPv8ZEx52nGGrLC5VDteSoTtMCzS1G5DgUOVHLQOHpaEbHBSvrnVS9Scc5RNiil
ZJWy1EyZTwCgRndN1++q55e3cmfqmkzyiOqT6zhC3/lQau/Q8eENf2qjX7Lf/bq4fWOTQCUgJKH+
ddh0YTa6JFVOWOcfC1V9kAOzhGkLV6a5snGzo8/s/PEc9H7/mekKftMCbqwEFGnVRS0+givh4ZKm
ZWMVc17yL++3aC1+OSPzmZKiv6wFNzGxFUlCkwoD58OautNDKiuCKCvBeVIcGdM8v+3qO8Oqjjqw
J1rsgVZzCAvLKg+reC0z82INlDUPQN3bRIYjg4uS4aToWzSUNidRpNYl4GINAHdStO4sm/efPBYo
dSQ0wUMaAEF/IaHhbmFWMgXRSxnnpwMSMrf0yGKcZlVimxlksFZXkd7QH8vZbQNPHjaBtxzj1z+R
pWjuRgs9ehbs52YWnzZj0J3IAGE7M38SV5lci7IQ9x7Xr1jzcH/NR0Bb3oZcUtt1SanR/t45fCx5
tKRLomuyJHVEn9eWufN/1MjVltvXiTJ/aiSv7bAUR+CAv3vHe5+GQliZv9HWJwcVHjbwJ9VUCGUt
omXHUDPOBPaFoPpwgPRHKogS8/7dy/XxovQP/NQ5y9iXlI7ppWhTVY4tQf5/n3jaOYWAQTocb7ma
RFq2Cy7HDzfmJXd+EmFrden00ewcES/6mT04q/Rcj/Urg48cEqnobt4fODkyy4IVcfQm2PYs6hYS
373cRfzQmDztAmXrUMJWE+o9h4D9iZeFuQk2b76V8ShMCf177ANdzbjav7tkbV4coBfhPG8aIoJ3
629rk6UVFnFhM8CGr5TB4RCZOp1nltwINzrIiIAjqrbtUoD15pQ5+bqkoVud8/1MF5vo5M8GGScs
usR6+MAU+UXHF5XJUD3ldjN935wvhfqXkxK9c4NATV7HSF9AfrtIy4DohYZoV9FzUhNthFodjIW/
k+6yWn5tmZMXiyznpE/yz9KkPtsG/Wm0AbVjvTsYPS6ENxRTn6hQzcuHCCMAdzQuqG8Ud1FPp8fo
AWk7Q8DkZkBqP65Gk6VuN/f1y2+PIh68wSN9gsh/62RyOkgD/+2rTeDjQ2nERGVQknkFZRZiOBQT
NPXKt/xxEPuHFxuiGkfhBAvvSVuWtl6ayGRJbkH9Qh4xP/XJiRtKn/Jq+D9BUY0eQ4c5qkm6UG33
FP/YKVVE0GXO4KUrlTi4ImoZY0scM4goXMUmLqVV2MN3ScplKTmz4PDONk7kT/VZAr/4nmbXIB5P
bjKFtuV3wA3gUw6q9LhgCWONzGFtLvPTyo3NHDcbCbXfTlUegfOCiKrRuxxkFusefXKssturn4KJ
Dc+6wja0bl/ywvr/GdoVwXY9Y4VERJIU6l5FnYfaMJqTmo+eHcV4zVltzJEFW7RbCIrnXxGn2bT2
KOTvpAbcCE8FfcUtOCE13lc44X/gj5a4CATTXDxtXJf3xwbX6U+m/tCXV6IAqwWbFk85WNhWxSBw
lF/2Z+uojOFwLVm0kSp82RWZdDjbTsUs+OGM5poAsyrV6DhsMPb2aSjh65CMcp27AQJzx24y7hkJ
Xwx1zuH3KUxFXHswLqFbZNT4nuQ6WMgyEwGRncd73JELd7pYSS89PN/BtBnyZKi+TtTQuKi22n80
Cl80dS5Li1tFeJkxacI0L4wcpP8o8ORrkzuIWyYbCkOp5GyOWJ87be4EhO+4Gv+wplegFr2gj6Md
hZyl2UQCRoMPgo6e9TaC6yg5q7/6vT1V5QSqz9NeXKhbXoWylatyj7qfSnGlCbFE6hYYK+pDpd66
tIcmwytZn2fItBnTE1dpcip01bBZiJcsYnJcWd5anoy5W2plm+gxUCYfz4Elu8d1QiG7NZgX92kp
l4kEF9vt7gLP+Pjn1qUOXBKerhX516xcd+URIpjx/wwnfSukmVK4FOea3gfG8WPpSTFxW8zFaGzj
/laUMungKw1GiiBC44I8J8Pex0c7RqvFZjYlltiaaP3URvvnLPeRxRgHIy6nJc7tfFgSXGHCwbPU
NH2UoxhbR2IuH0yeibBewAuTkv0+kNGVDaOoaf5vUvXy9t6H1t6V0bQYXSfjDITqrDFBWzUmSct6
qyLJdmvYuTXOR+DTYYfVSKpSjjk41aXoi6jIt4353/tsz3nZylD6pgsSSsM8sGq3IDV9n70Qpc/E
vP1O6M0TBRONX+7QJsP+4dDb2GRlnnhpoO4HUvsPErz+fWEf4Y/yKIuk1BbCugohPhNdhM8n/h+5
QUJm6El4KqsH0QhZyX93xFMz7GCuixaKBvdxhio8nKrEe6nvtWfMDWqqGTgyQMtVgL339Y6zFwpb
nCJBhDxprnCAsUuQRUIGeOrc1YM7kqWT7LD1aCezPS+fUw+Eo4wg+tvAohmZBMS5MF4PhxBdCLvl
UGP/u7CWRZNWgOxpQPTfabKeWDOMSlhCC4MvzqLR0NdtW8Qdo8L9poY3nFo0pirmR3owmAnV9MtC
SN1EWR9cqv+GDaI3peY0PWFxGBEyTXXvy3PVyu5ayEW121TJfPQjvFaGTXBnYFtrTZxCncHsz768
VjAKhoeyP3FJOgL4R+tFIJSrwbLzHd1YyXSBb5xPd45ZkxHeHmjkIvqNEvGz5DlVkJR2+vC6SSnS
Ox9ub1IEe0uKjNZARzXA+2a4bZek6Fo9RYJYtNTkwg8Zw2tuMUQQ2M7iTl95XGY2M8YsAAc5BCLV
x2PdyjMcUzSkvDH+qnaJNVTZFh2w9r74hFH2qn0dOxaGehQ3XdtDXiY/wtdBmAndZq8dpzKlPjVb
zK79WZJsh4YHB8bsyBBa+l9Lk4e0XyAUu0Ww6t8lHUdN7ZZySGGMPWibAlnPtpawLB7nKjW9LOYX
lASWaoiVS73CdlYfw7QQwrIfgp+lEcUBb/habTxTW8wl6WCJYlGPcwUXmP1z5kBUvcRMVSn0hf1S
ULrhhDrJZUcmXS/kEJUREp/TtJv36BPVmH4qCRgPeS7ni/9H3XJTaHZtdiZrbbZ96vjRb7/OMxVj
EsBxgncDfBUeBTCdyVWhwTRnWS0ecaCPkpvfCEpYJIUeYeP/bc1TNozAG3+e4TVYJPkVaFFWqr/N
ag26bswra4YtltWuRrgSqFaGHItNT+XLVnfoEQuLQAfFA9xPrPUMDxIz+NidGFHVRl9deXi8BT4o
z3N21CM1CN7xZnaj3tgpcs82y4B496NHEA9ZJ9Foj+cBVCbzjQdI9gqxTLYD22OcCwcqQTpf1I3p
vuxRL6lcjSi4U7ShusRU0zyr2cSeLhqFsnJ+4Sh1XzkMI5m9jOFzrC3L3JRACBjupD6epproWTQa
JFnlEI9XquUgnYlJQa57KPaZ+VEvS+NXrJ88OoUKfJLSI84ZKI2yZZiGzq+jNVCnJ6fE5+Tn523k
me01N/9ucEz8fJZQPkEn2VwsB6XEfNglmOi0I5OyXwZlY7Z2/MK5aUiUv/fPjcMH9qFIccfwEqUI
xhAqPyb6rRPFUplbDIGUi2obFalQ+NrQhnFBg9Us5Ov0AsIVXWoOuAYw38+pXcPj5LqoydmB7AOn
oeLOVo4M1PxX69fDTNXs5AxUkAmTjGIozoRJQKlneITkI8k6TKceak1E5CySG7K2KgQAMm7ZvFGY
sWav5dLWR7WwjsWbGDk6+xmqHUl+gkFzHZU03AYnO5DHA1ZjYZe3eahbTVfHTp29jxn5M/BitrHv
+qcFRp8dLQwBRqOAJK9cJn+4a2KJO3hdf0SrDO1aORk0gWOzA7PUvbbIRnI0njWvlgkIwpi+743X
44Zaag8qev2d2X+BMQ1UztMkLcw65OKamFGOa5/y88x5sONwWuNMtyDqvywmcJxDnw2QE8GZjJsC
UvvY2MHHYP+eKRlClepypC05Imn1jCrYPLzGudAhZW1HnHKrecBlZ/j2T2+izgmtj+FRWM5WCBzY
Ok5kOrZ8Ojh4/ejiR8CwRzmQUZLXHiAnXNqTn47UahA9QfMFuARtKd2hAZecQGzI5B9zLycr0G6Y
vaHLSK+6nrnca1gxfTkscZ6c9V7FOrfDIvrUk52WXlwrIzR+VFWDotY8EuT0nkLdXHuM01WbknQf
PlFPz6aWSkEWoV92jhblqn3jDpNaaDYyPg1+bjQvHBiplnqjo71fewlL+gJPQk7mjJ2OwhJhaHsZ
f3paVKumf4My1IPYtqp2fUmYip6KCS2Ci+Drz880RGKAgnXntu5KN3FflszWzUw/Ew41vRdQ9dEc
3tw5hWCoctpcGZyFBvr/dbjF+hULv85CgAezxTbGvWeR07gOxnqBwgIk+49pZrhT7iaCSy99Ft0X
4l5eksKkH5XuuKctwYT5l/8e9YxsNeaaoSl6g5pZVGPCzrM3VfuBWVGPjoHbUZfDO5vrg2NO0mOr
0rcgucwDj9SOOQ1Y2HkpC3nZa1n94SBf28ROflrDzb32TLEfqL8LC+b1MpJuUjCLyAGVhPMsl/vj
8qRks/57yLEfSU+kPglEhlGrcADllII1B8y47tMIvfUs6LXhpbkOTUfaBKsj8OzxMD3+QjxU+hx/
tZGiEO1ZD8zLgJsiaLUr4CMV8vEhLdec+9BYc1lHDmqGYM2Y70MHgI/b93aFqR/f/1Q5pR50ETFW
sImhIdwmlHJfmTPchn3bQw0HrObLEUaEuUJomD33sp4rWmzHKfjG8iSdBNm/qfYGTCJ6z92SOsWR
tehNMj5odPFZCNvjpR8vc0B1bphQQyZ3XBq9ZxjJtab/1WI1y//H1fY4KG/jAQDgB9T3mAOMeNIe
My/e4pkiSVCV9ZpM/kfYRwULJI4sozYcf4cJnMR7YJeyVozaK1wVkpg0spJFQyoedT9Arhy6kflg
9zrrkq5Z3IOBGoW/HqbcjQjEP1ZHntzch8yR6hDy/1SU7AE/2V+7JItCky8oCQ8zlWHY4KDQk/q+
JTEAOF2g/HrnBNXAaZ5vg3VJOktdp58m2Q8bowHzk8PRWWN8beywEs70fkfti2LGIiwfNt6DfTO5
qIMYL6R+tAKBfiF4Hj98hqUWtPyGQQT5DUI3YK8chAjIluyQ39vyfUL8QoJ8DT4dcdvyOScVAkRp
6FVTQjF1VkzlFXFNmEhq1CdIUl6F9sNKLjwUD2KTEplexBsJMVtkow93pcYwkQ7UdRc9KtqxePA9
cNyEwLYMfnE5ZYnRCRUszKlkIoHIv78Sch8+TolFk29Ljx0UUXeXQZbyO7nmbjDGn70oOn22lW2X
KDFRcNb8/crEKwDmHzik1xtD9dMkKMzaeV3GMqQLUL7lPyB/xKDPZS/AYTOI9zwjQrLwS7ro8uu4
8QsOPHPxX9o6Dcprr6uaIl3qS4cn9gQK7IXQWrkxx9EcZAxcoblICUlRUgx5vfAJ8KG9wM8TorvD
SxYDC7kfpFyo+IhZ2Xq2W1Iqh+dSMc1Apt/l2ecmNS94HpknP0Db8Uh84f9oHwMFOZ+td/UgNGZG
o3EGs5E4dQQM1Pzj4LrwfrGsG4BQCxRc/VzHN6rInVYQukFdrHlzf7RIoCbelb/5R6yNLCNbeOg9
TidlnaQzbnT6VBVcKddNW0hDYXtwKtybn51hw3b7YCRpbeoqm5m6RsiYxnOz7VOBzbd8FBZ8E+b7
JXHXz3hHjUek8pEaMNe9ukWjaEwt2M4lOyCqX03Fo3muW7ipO5eW9MHuBATXxF/Zyqpn7eA0F9mn
5NJwlHJLxE1VO5o2cRw2b4TgNSAYwpWjJdY1WHmWq5QRVN2MVWbpgerhlDMfcd7jWSPxh8MA6Di7
1h/CLwHclySkNtvGzjewbaikeYmIsB9d4H+ddN9v5u5Be/yDjkJyRehFcdpt3ARW7YruwJJabbG6
UnqYcv5qPdeI9EpVcCztq6ypjQ4hBOtwxAeWSEmGXKCzbsyGP7tYJhiCbTsqyQH0DhR3pOV/fia5
XoAw5QbUb6iGFnUBKB+lTZ/4hKudv2IBL9+VRDSWwwRjsVzJoYpn9PQMPtW5DH5i1AKPCDPXlnY5
ZCMJXfrD1SRqZ2R4IqJ5t33aYIFDWaxdaFNA+vzNclIQH5VrmqFNBcEj/Pzn/8XCiP/CclVMZTJj
h0AKDRXnqGRIDO1hFZd8y5tkGSttsBze1SCPdN2uy+Linh0b9UgrvKvpSB6ldrS0Tr+ZP9d23s0b
RfMizq4pRTvtTTcKM4t41KJ7TU0L2Vux0+vgzHwn0OEyUJV+RRxpYMdn7o8CeaifiHl8StZfvqyg
X6fvQMROJsBAXlxWiLka9szKAFf24Z8W9ZMSDAdPnfkHXFPn6XBEkC+7UcEWzpyuHyDTAO6Y5bap
b6SmAfRZPPhA4k5wi36aPjbgiiBo1Jh59BjnVmCtiWKUbdMAYXRNprnvvKGCcspscaekE7CCuVVn
tMEEy34GvSXMoxUQAuWffRtwP8vbVUGExWfnnarenALkphZbfN+wrocbh9IePy36d5qJmya+ZtAj
2BKYzFJ3ADgi/PL0DFp2BMzRRow9hPWenNSZh+MvJx+sY0oxUtTRS/f1itkAx5fdwXbYC+92dyle
nY3CEE4ljDxdlulf/5UHCTtrbFGgcawKd6AXsdel/XoyTltLMwwK3msOjd6+MxXAjEE085Zc+j3K
qJUuQjrCubVTl11lp+P07pt8gJ6sK7Gnh2OJNh1wA5OHk4Ku5ELXaKFU8/LPElJpS5rNe5WpaEkG
RpHH6rqR86HnnFysgNqyAyPSpODBwjmzzj/faF5xeV1uWNE7O8wS4YK4xSEQTbcwYz2bQZqAtoLw
3/evJY3Q9le0IZ48Z96PYKWbyWnnGU3kBM58v3zptE/8ajFeiWZ5FWloZmFMfkbiv9WbOZrRA7dP
j/aDDqpfXSx2zjCWktKzeeGXV4+25kA/nytmGtQrKjGs09gVGUi6SY0ieNyPKSnKvGHXcQVx13v4
n+yK+QmKqRm7K257lU+o3ygu4FA7KdR82mRwdu80Z8MTa6C0DQA7M7VXH9nMVS82B0sNFEYAsQFC
uyD/nn/0tgFN8M+751FHudqwuLfXALJcBEci6SLrZXBE0Q9sK4n5TCIi/sn9ZCZg7mAOpnHyz3Jh
dF/h6uMP2DYnCDBht/+jOKd9WZpZ8J6oU/ZdCuVVJ6n1Ow3ESjwHDoItGLfK+UeLYcNL+iwqaNcB
coWh5mU2rfD34PsFNSHUc1HLC09GIPImLxa0VuuJR1WdR6IfQU/ACRazYLdEOwvUwq2/61cRSw0I
0vzRpQyiUnmyZlO7Z3KPjVbapGuSCMmZ7lwlcrLd+vHklbTmwKJMa07oFlTIJ18fa+FsJKEi5kI+
ak/EwD3FXWBJXlabRSgBzMXQdETltbOrYYoPVI/ZmN3g1F1audHfYMaj/VmqOs6vpy2i3Sjmmbt2
KK0SR+Zw4hPqyzQxiYxy6pLQKTMbBw7phKD2mXHG+T7ejwnuFtOMpVGOyy88nyIJtXZKIndhfMC+
kDRFl0MEQhb5tW0LHPgozXCn/ActmKwnBs2toOgIiYS4apA3ytFe0m83Fx+HMa3+Z13VNFAgqh61
A+HrP+7rjqwNnEDR76tYdQg2kynJ7RBmuSDqfMA1D/0AambNpPEBFpw98VnnuVLPZEYiOOsduNtC
tw8Gof8dOPJLspXsvajYy0mZOfbr9iVu3CHobPIBZzI8kQBATLt5PWZ3Ur4ae8XwQETd3Xfm0Yh7
pNmD6lnplfSg26WIooDCn5SNxz2D4OKFBqqX2OP1BoKj3nlimg1n74kUq7DmDuPp6vDi/2u84+rP
KyOzcZ47ANNlBkr/kZdh9VJlWAG9TZMCG+YeoAUdOTCBPgyyDhslUfwQMncJz/ybuRhwVbyW/w3Z
BLXAeve4jLVag3+AoMowCeTYHdnv9nR8fQ8+5qXeYdJU4y7OqgS+g/ec59Mc4hC4HCpAwI+P8xYj
Lmx7YaB1DYrcTvFoe7HxAGUtQcb+MZfkgUTKbFCHNU+YAaq3kqIuwRdso8GS1lkufio+zpth/E9R
0nAQQunO9Kvs71Qi1xnGCOiWZkUTlqDm8xTqYoSre8KhlujRCEh9IImJHzhP0XzD9zxZLtyH7bWP
wspqAz9obk2OEQ6rKFnno6TRGpdcoVzadDCebz8zyPXTF6eLJ/sxy/WIDrtsMDSCxlPZaDC9AM3s
jsb/PsF4csHN7yrq6WF1fb7BrwyfSrkMsXOJuKyGzE3ECO2hPTJbMJ26fJoly3DUZQV+EAmlQIK3
rfK1+Ytdsj0SFK7vsvub6iw1zgVHZGzwFGwP05nce9ZPGdR2Hof+sUxyh6cuZGxUjd005GYctHn6
0gSJIPXpWALXK+rcgSeBfSxQa43HJ61Ip9Y2ntDkDguxvJbbv+G3aaP5shncVRd3pInve6xxrhYu
+B+ukOhtmkRc/1eHirI1CibeFW8lzsaqdvdPLDLbfYS4C8uZAFUPwVo+3K8xh6N4faAMLukhLdUh
jdiOUg433zx34b0LMpxpax9dE324BC87OrviTre6L6oNZoIIIzCL4PNJaxkKTOYDSo8v3w6dsy2v
KWCp0jMQXacq8gXfOU/HWcCaBhbaYd5dXGaaAvP9SU8qmga8/5rMRLOarAR8ro+ohMLuktZ/8sXI
Pu2ILfdq0+pgTQRozmRFv2t03pVNzvweD8vSQyVptvVdOHEWfuVvzmJjGZTvOiP0Zz1ZSu7drpSE
6009mYSSZfl45uxQFxXAT3H6h3tAC3RStpMXiayWflJ4tQQ2q5qI5w14uiAlaEKaGjOiHj15WOuK
zgG8g2ZegZaJbEX/dT55NMv1ONZrtVVfiTIG9fRV6nidhmbd2n656RtP/MujnNhssELrkRCnSn7P
Uc9SVQiI2IPBnffsMtv6L3HIFnDXONBWp/DCGtKnviIfVDMuHAWFI/Sy0Msp+p3fau51uj4F70GK
059klg0orhiPRcUaRVnrCeEMerpzgWzQB8PilcF3tN+ZhIUS4GT6zCuzHk3/c3raBVWD5x3RaXL5
Rv2XX/WU7jLDEghTH/Sx7pRDBEiGBGN6g/GaTBylc62vim4ZgpL2Sri0QD4gY/o7I2asvW8xU7yT
KanvShhCR32c0hkGdAAHQ7U3NrYwh4W8osyT+vp6AUfsRnkbb5xnU7/xgzh8GcSPRiRkPsMfHbIy
w9C9x4WJggjVeDjC19zB47RJgQBpyBxIlGbRH95eNIGWcjxsUu9WtF1wRLM9H3hstUFH+XFkOY99
EfP4TlZAN1dwP00qk6ZjCdAeTo8YWBzuBMsryDQLGnvEXBwkc/exsUD8xcsvMs6Bar3O3SR6SC1h
46Vcv8flE15fPC2WTnBksZyLwgPdINSzIXKD53eY1T65YsFk3gdaEkFbLKvGEGFqZTK95GJDFr3H
j4c8R2i+MatNRGDphkm+V6PDsOX0uhEEOpEZh9fWQspxL/epiCQTvXZAM7dugdybX/UllmJGLdn6
7KnSKXlAQ8RRXsiee1pmduJfgkZGhTU83Kaxzi6f/p6wPiafDuHFMRPfl2QzoQm/WEe+bR31dSje
3W5Qw5zzH7+3wukyJiNczPOu7vfXgcJNwNonGqLQDWBjIhJq60/TAvSNaC9kf2JsDqNP8vssl6PI
0zCfDjGpOecXnWUJSzeEHqkmPAPgHucUxexQQxrSMqvehlpKEvoUthbc+/VR1EF3gZL5w4de6Qc+
btIfRD9Em21wzhw25Pwqikx/YlpCau5X2sSgSZ5fcXKRM/3F/6H1O23+UO5fiBF95ttQ4u39B3Wb
XQe6Kmfu0QvM+kQKBd8i6l92y+ZUIGsYw9TZ3s3FDR3VPf+ogiZtwcF0mhMW/owaeBL3aCqXUT3p
YfJiJQmMYdOWxcOS7HSq1P3HTcMcojrulx4ML4iOC2v+myhLN/OLkoSwovH6Y5li6w9yycQgBuiA
+T3l2Lzo15rTnFlkm5kpZWtgiKq2aEts4OBZVmOdwCbShCX42eeFpURvLthQ32tAVm0Sbi0SOvFs
F2HVU3vQ/OLgc6TcTkn76HDXRam97OANfeus5akg/TWmIosrkr2M7rKnTpSjBjyYyiuCDQmj6ZZs
4nxxW+H5oGwvjVI/O9WxjK21Yvy1+sjbMPkZQ7j/WM5qcLzj9lOqwX0FiWrLs0YI90L4dmCuMjKC
sLCPG2vt5mi0kJBBLY7+Q53DTDitX17HA13++ZLcaHtcZ9nIYMRf60Py9EDh5USjs2hKn+pKb40a
hLN94+6guVTilsQVFR/yZCLAzdyIV5UzBrs6Ixn5VCblsU6apq+CQTsw6uB0KP6WrC2qoOXJn+ey
iZlwe3nP3yx/4E2NB5BPx+oXDeN2Vp6wGvlW+mYBy3Nl64bRHvWXdKJwybvwNjcsY+V2fAX6IRde
EPMl4HsMZ/gMk8TqguKC5oXAs7DRfe20Y/6VlZfUGpDjluexf2hlqNNehnGli+b0V0Jt12DUdz56
4478BqeUv2XutcMwHvNNcaTboaRJ+u9Xireoq1o0eJXONEJAL0fEKoFiA4WkUyFJF1WWRLB4IEVs
A6GvqZSvcZvrTOnlzKylH+jhfj5w9fQ9GKSbdjt0mG+JZSpHaCssxD6CgYPT6h3iz9RHr6vCHdS4
5Ni4S7yWMdbtdOIJauZksIwaV3BWoLwtgn9dY6pg89FmpCNQzgjlGjCLuWgci+qq3QTYfTt/froi
r4ySSCa4k4VysV0uMwt4nUtYbSN+6Cz7jHmSdBRAadfYrxZiXWe8A3e+RKLEKvRamMRl8OTftXZ7
Gze2QuxeOUABT5imvCZo56fe4vYveZFPkYod+liqLohngURzBt3T+fgVGOYLDY4tw9yJ63upRjw0
UBVEeuu9WwiapPVwkRERhrVif3fLJ8C5klArlp4ydc+0hoBDnhicwJhFJWkbwqDg3cZuA1S5P5+w
wJUBuJ2P9vpEA3svAK7ArOeoUwS4z/nbl/tNMAriidX5H7IAzRQ5iKEslcXcWQI29TulU0LGwOsb
rj847YU3BoIPFsg2N4N4fWpGwZj1jMSmm8Nxtdv5k9Zusioz/gQGdeP5hGwP0vWHOpmhLPz4lY6B
TADJdFXbm1WmdupmWv1s4yfKltPCIu40WWeSRaSZ+20Lh1+L+yxF1l4uf0xovAo/+nmO/8C65DqK
kNEhiKR2wZ9XlxrOfZankfUwP+2f167aza8Eu+Fq46QhvFwIFfd3AH+cREFsYOJEDxwF6txcyS1S
ZKw07fMbVVbqLjdHCEeOn8+f3zPz7q7oiQEyjgCdcLX95w6joOanIuMMaYUQVqw7zFMH9lRjQOhp
RqMTB73hgHQQMMYodMSopfaaHao0TzPBzKyoiH0u0qOdaUke9vfEMbyrT7RnX0yh2de/cJXV13Mq
8T4MP9wLUohPQTZljDn2Ox4pN/8ut8urUBdiBxlXtpmApoH6tovME7r8K6DXiHqvh4MlJhU0m4zx
ET40cOVWMHnOo6D4GLTVgNYZ3WenfYKXMHCz+dqYHv3ETPCnYF7J/7klBLgUGNGYBJot2hJCgv8H
gU0jMAZQUxao+CKpOOs+Ync4i7BUSzBkNPhiCK7uEKHqX9QO7Luaue4yMu3i1e4sJU+gFRjxJozh
mrW3owtqUcQWW5ZhHKcZHLglfuS+KuE00f2n/nuVsuQg5r+lE3KOudBwdagvYX4hIyFsJTT8i6se
32rV+MGSgHTT83o8tTRiulLJmDKj3tcCUwZtYyAGWAxomMBN5yP0wRu4LUHLwWUXDHX7Vy2YReUe
bbN4zLDs1mHsmPp4BHE2kDwPCw+DCwGS5V0+vOQld3ehJI3wktgKvyH95WlQJrdkFliev5P62PNM
xQpFflXc+iyv3sHym/8+2sxFQa5YmbJc1+B9/Wnt7Q5KVmMt+llp9yhPfI3wvC2oicMRGdLstuxk
YGM+47OFJ3iToY7+XF6erRjZQNNk9dT7yhftulEDrrO76m4vlz4KtYhbSxnvh4tzpaqNFiw6GKx4
mkNdWQK+AZKWxvpCahKnq8y4bArJ4Nn4QakXiz33Q6ZHhCMwPMsus6gTI3dWhjC285SbJ8xr9N+9
FbaEfiTLoAS0Y3rR9PgLLruHsut43PXkXVFvPGmuIcrUf0xSYFIHrjfwaHhg4Yqq2mXoq4y2iq3Y
NNGbu0FPnlLjA9anVYGdn2SC439g1HXmLtSU2pqHLFMIu+PWOq3wU8WmzwQ4cVo0zYeicfX3CjT5
2Op2RPG9Ukdn4RKfQ+C35okkFF0abe4b/ZL/ihCm1LLivw40Z/8Y7XhJxVytcEU0donnDDpwEaAi
jgWZJKAStpG/Rqdc/gAfnSpiH+6YUP1oEZvYltoNex9FXPmg2nHW1szdZQQkjMV5CgXCALaPxCVg
XHwdIKB98JPpZ7LeHVG8VRXN4QhWZdaR9hn2sr+dGgkkDKFlJD301ITh/GShnPxeCcBwMZzYF8jE
LtfoXqdMqx+P526Kks2/ga4o4oKO+PIeDCZDLydTEpj57qNDxHMuyLQ7ku0th2ib6VePdsxmW5DT
WYEtVc+H4zjlEmCaUhKe0tFcgLG23i98oUsOWyjePkOus+3XKu1+rEJyp4ZZWLV6B/DroLn60myb
ySNao2iJV7GRIEIRzh6pv+cz+6ZYN9AUm5Uu6x77Sg1nWE7iV/YRsNRGsq+lm4Cx9EmrqzMhxNY4
VF2tUxZ/DUhymjhzyu23zq/MPK3q3+u89dSkDBG08aX04MsRdBwdZNM8hFEeQD4FL1g+mBYE9Q2N
P5NS7MO9kZNoRlEAkdFcVWglQEOECahHEQYk/5D2P52raVRNk6+B4MdOzvDybVj++nryp4qXrz7Z
N2fUTHCw7SIDxr44sk6rHLTdAhzmBHW+/+IEfmkiwrDaX0ue9z+gz3evxMl/IZXIFTdVoGJuq5og
OacMfdEK/61AOD2tyj5om+JQaNlf2bcaMK6ftSQSIWQQnK0NeSGzhdmmzcATpUw5SHGNuRizv2E2
wXrkA6axx08Kv+GK4POhFRvH6Lw15xh/VdEstYRc0jtiZh1fhGbfsequb8uEoo1H0sWUf8taSrPK
zEntYOZQ/UMRooKXDFT9KW1l7XJuRqoJiKfWw7lBUmFv1NxjEWhMKcG6P4jD5OITAdMZpFwWIwkS
aYfVucr6CQA0dvWRjR7I/WSK4vWVZfP03cJ3T9tiXCjkk2QW9LBvOkmt1NZmqk8m0p7ymbiv+QCW
2O9wlliBEA2iGbcgOfaAW8t1zmxpiJEu5EhgdrsTm4qUfQNxlA/XLyjNE4XEmoivKwMvlEqCklUI
/xZzi3cHjQwPomUgSUANyl90y47LVOilO+kvEddDbIn35g3MUBltGSErAXRW29vUGXCBE5r4DwyW
Lzx/e6QIrVD4Ys+RJi/7KtD9eoY7HV50Ez3WSKn3pMdM8PrPEc1DEr+YwDBqLm3lGD+6K0jjJP4h
gWY/iaB5iIOO4bezaN1ClYO7Diyz2qF8KP0qdkPbza3GXYo1B48q2szCyFtE98WOLNaiGgeBkq4G
MDniicb7AUf6oUMW0hM7K1oP4mmHwccyroOn7DwvYmg+4mSHkHxCsbJ7mQvgfXl9j/r7LUo1Qqu0
qIJwFMB/DdJKx+DU8mhJ2kEqSKEJnPOYWY5VdtQzmWs/Q/sEP3o4kBAEMg9bHyxdLxq9HtL2nVhA
LnHSw9OL13PL86x4/gjMkjQ6ajhrazxtNcsQtH0SOKIulfXNQwDVpTYny0P+vwK/6+o4ThTIB4Er
nTmmP0ldeHHWK39N2dD4kX51SMCMtMtZSWZmWjAd0kqYC+XOF2BtvwKjdGiKJ5YEYQ1gnKyjvjgt
vfPtDXYPvxT8rWtoEjcOD78uazmHeIxU9wL57XOquzvZ2kj6pdm2DAkAP7fHT/jTV93SIimPPWSa
XAGWf/Armrz3RxApIn3vwirmVlWf2irelZOwkAkBavAzS/ic8/QA+V6qOCgI/mSJSTHXcwqEMBSj
j2oIrfdyBZc0D5hi82rv2D0EBJDJgzVbwVp0LsQynkedBrWPHKyz0d8duRqEbyx6pqhaqDf4STQ/
438KkVQ8U8D+YoIhSL37mtmUtS/+MpDPsphFO4wE6dwq7cigOHdHHkFsVa9Q6et4VRbweJB5yrEP
HKfG7jkALEZNzeZzfqyt/aGU2VKocfz4pxFKJBhfhXHu7I2rL7WZwscAR2HqPqJJvHDg9tVEJtap
ZxJSJtjPm9LNuCl/rr3GpyMlEyvGYqkN3xBdPOceMhpNJ5xIz6L4Zm18ZmwlUuz3gEbTlUp5v7GW
9K/TTBXx1wpZuXyAEIhQWwDD8twGgUwR3q/NkaRszsCRXmx7vaAFdzXM/zGZHf6yhNkfRzH3ZykQ
+kHRwTb9jHBsBZ1yN+nKnjMCWcygJEmDichdu3uHQ1yEbv4RmVv3usehPpdrWHEUmMRbWjXEohbC
qVu9l8iD4pk9DEGuiK5FmZjJ8Q+RWvWLFnkKsUC5JE8MJ/UwPsS43fn1muBo9ZBkK6BScRXBjNKL
aHHnqvTyclP2mW+9RNx7EBsrqDjdusgLzYYrKnrf30rMzFs6+scsyZ6syZjbg0qNwJoxU2v4iunv
cB9xSKBzo0TC0XOEgGbQ62w0J9FaxCqDBgvv10CU6umfOXYQY59r0BFyZXETU9Lg2GGHJn6a/GB0
hwSV58dvQ5+HiAjN5OBNlV8IwAal7R6bVLveBxs+LVW8BAZVVlrM2uCdZKmdqursLarFouHICJ0y
KfCvjQJX0mOe6+AQa3pyFCJ9aTN7R6PnSVUbb/2BEhXXAsiX+yw1Wdsieeeski7EQ0PoBBMQjro1
CLhxI87bYTTjlPp+zfsFcLL0WyiQCHo1/EGrrdO97NGoGf0JkAvWmwYOIABoTPpAYtx2uxRCqlWr
yshMItNyHoAwqR91KT+C28PDr9Chv+eACFxnzQ/O8y2fcbsSaneqwTpBDu1kXPAu6jzE/44B+JT+
qHXZkb09v8En0zfBnIw1Orc9ZCeM4cm6CYBq9V+1feHSELx/BPFzmKlEz74PUJNClFHAnDrPvlaf
jD4eEg0sg9PciopPZBFcv2ne330/uibzvkFlXTdXg0RfkfjJM5QokxtlPP3fQmj+dkNWmAuOop1b
mx5YIUwBEy83gU2EM6a5SCCB/1uJcNupFqsEKjCLwBp5euaEoKRMtiDh+C6fpjhFwa0zvB5E7Bey
qGEQRQ8P2RyycvW2S+4IipEQmCVHVhEs7+uB9TUxXDsBSlnrOVhIoHLsAFJ9Tn5AIS+DJCQrwIAF
VWfeGcP4e2pQ7bb6T344HfX5h9sCA5VZTCg7YJsIR9MJxv/WKumOHHGmlnjiUf5OcyVzw1pG/WZo
iFUDbbDX4Nkv9VNge5AIo0gzbZhiDv4W7eWi6vIwJr53MebDi2TPNQgB6a9Wy5sR4K2TFw7S8bq7
xtOczcnWuhGPpBpGBJz04JKyy/e+C4lggcqizFD9b/zJybU7A3OpezRqSnsYUDq1TgkZ9HuLjsUE
UuXspbc6MdQ/6T8rc+9b1bvgWE5EVmQtoa4qbCj4v0k+paIbAzNUOg7yu5f2vDHXToubkQoAEq+l
e1lRhl7eCw+TGURAt3IdzZtewwz5+CKNbP0T5MlB6g/4RIWETrxT+V/T9BY8npdzC62q83YnXb1H
rCZ0ZFEo0EJTZq6ZT66Qae+EmEdzRLciuUqestrs8L1ZhM4dAwXcxSJKassAe8/WWsX0Aa0kOQ2k
LNKXR8vVMjrAqjaeZwbZHe8Vc3aLnnVR5ShuO8TwllYtEvDEboOTM9ml5OAtMwyTDIoG6CpFV5Pe
qF0kqQWas5ml/i0Zbo3QL41HUvMLwqzQ7vSeKZ/HiMZbbALKWqbo8ZutFpuLc1jmMJMzvAliFSJ6
3392D5AlACBJ2DB/Cf+SoHQWTIf0CqCGG0S3dKBIlyqVUvgFc8/mWyPeNmLzyjNbVCDVSMG5KsF0
MlQ8q2S/AMkVZ7isDTDC0P88Lv7HpicOV9qn50uZaB9y3PW6eDn+ous7jM/nqlVJc6RKXxpDBSbd
ytxq98AMSR7k0Juj0zMhm1Wj00/v3we2rvaWyAyj0jgVtCCfbi60qrVC8PZT3fbaoxJJV1O2Kg0+
rQ/tvsf2llx0CAyqsRCzPt0dRhBl4A6MMC0Fs2LlxzhbNGIx18MWYvIhTrakzUxFQHJN4D5Ba4Zd
4U83EF6Y/TF+YOtROzdRI/uC37WAG9zECQ1RWDOC9TIIkbHnsy5r5r7T3PKgM9/l7rImsXpYkYat
E3OBIiqoKOgKREsp4SXKfW+5FdaYqbK3ecmEo79Z2IFCT7tqi37GWN42xFq0rCE+7lDV7BqrXsTv
XnbISRsPMWfLcaPc4Kjhadtry8t7/mV4wc+KJWFKm+cwX8pvF+BB8GzwVy1JDOHDArH3Zl9WS1Hd
IckSikVAFbnjnCS/leze9HuBpa31mtfGVHnZP8n9fcHaAvUrCIthUdZGFvV28+04xnzs/qqtcmy5
RrC5yRV4beQ4AbQCLOX42IWJVuXywTkU3S98/2ppi6mpjwpQ5NxYJ9Tfvo9Lq+5B66Ummog+NlXw
ZC19DwDaQXP5vvusxCuZYYp9hQuttP8cX4ufvgnUelDE87dRYry8HH6xfzGhB/azCrYnbFemKbPW
nTqWqPS+xFWBrI+iIdw4ky0rVIfAd5UexjpbEpIccXrgryYXYuthG1E1GZLuYT2CF0W46Myv2uOm
EZwWmXVaBark4p3xCuIQMRMIfP3mBK6wn2bshQkDKv4Uv/PcmGNBD0HKYAFVWYguFdLUzah0C/UC
Wch1SQpckg6TIvHWKpg0lOZzgMESraAAposzckxmTtQ+c31lI/MxEnhUQwx9JKrOtgI2pZJJ7hDp
Z9Addzh8eESmU8xD35orgiO/NwHmqrZX/ZzVN0IC+GO005K8OqSrZZ+Dbksoy5fW1uTko9LADsrN
beOWKe9Z4xQtYYq+CxtOfK5QBpeMWARmdZ5v5yR8yFGtSFmMIWw3hcJYO2U4tW0EFt82zp9qIu6W
Rm2GyfqFuVop6eYIiYOhSomZ3aezEIXV71JBJAwNT4/iIw0iR8jijs+t9Wumjc2XVKwpBTXVXORb
XDSAjFIBQNfqoqZ7u89RsS1r8eciJqY1eq+jbhfBk9uYU00gidsqDovtKBWKOF5DKrst1VljOUyf
q4WgesffyVQePJfck0YX1uM0hgXqPGAI7ymqJFVXn6g1tXLpvitELPcvHJhGZGJj5A1tbk2SBcmf
JiapohjUyLbmYMluEYjhdO3nPhi6uqK/fckwte+g5/zBGzyxNE7Rn7+osDPA2Za/vnTzELbQXHil
QZDFrIt5r8LmAvqOqrZs6NGkXUc6KXooxVwNmu57uhAzEydhiNUe57nwTTiu6jdbVSigxiavlSv4
VP+Szf9DW53u7Zd90uFMx57gEoHJkGsgk3RjsmBzvdUzDMjCLlWfCX9hgNDE9YvBJpmJMQP48Re4
fHj4MZ+nq9YNL0ZxTgBW3IaX1HjI3namePwBlCvuoxnKXZOegVPcZiyeQXhvvytXPbOx+G7sUcwi
sBp3xvx3h2HApM9bmOLUrCv7L3KMrmAfCFeRJqMgiHY3m7K1ZRqysqTm2l78LPcGkwIKctilCGsb
OIr697HPq2ThfFMkpgHowlHFOHcPuccs1sMPR2RYli0fGFZhbW1hkJbV5XiaFObMEvlw1UtrNPqQ
QE84T+fJ9j/tvq31mUtNivI6HON3Xfz/y8RMxMlYYU4k45yCpioAHkWt4jMstSiyjL2kO49LtOWr
paC9md3RyJR1l9ewM2s7N7dOOB7JHFsgH85JYz9ERZGigiCmI/mJqY8WQNByYbmJezJ1fnGQ/mfA
2ZGZsVZDcivKJDUs77Opky9Ywb4wI6VwX+W+5zApe5dA+6UsFJd8+7mNUrCeJu9mCq8Xq5eeSdoo
afvGM7U+6XjE7Qmbo2DYo8iimCtSMXlMZcvwJBHuFazarUZ6+nMJWKQ4iwjsKZ83fi3dYIFceeB1
HKwfd/eXuiSRJSnp68qq9rryKROTXgldPVG28zqTc5SghSSQb3253Qqj4wLCfEthlR4cUPGJZs8p
D1Gq01tEmG+vqmthg8ttrhJ/uLZZ2EEUsLB9huxt9ucniCen1xE2pFnFiRC8+tOg0GfRpmHtQi8X
aSIKxHiHH2Uqy5wLZYxkbG7tVCYSIrz9ziuq/8etjnmpmQyVi6dLrrNFjJtanqplLGWEYdcukKQY
Clm2lapy+CjcgdsfZWO2zZ76j0Co9Zt8OdfkJUrE7bEqAO2DyQOpeKB4R+pW5mqhixtV5X+M+Zxh
znXSFFJt0qxEJSE46MHKjgcbaO+YVdyGMKC00Od2z8o8sKgTgaT89n6+PTamS7/I8lulyLMk/k9h
+oiKhY9zw8aXAUQPBlinO7pyHKBwlbV2+SRP3ocOQ68FyyJJTOhzqDyGBxguzCMdfi19z1CdfXmT
JtjWQZQLTxGjmbNJq49wKU8yi4GhrKrf7RiYqdAhpBY2viD/rzBRPDUJ1tIOFpxrFVU3gmQ3jR9G
BWXceIJM6VVZImMMYuo3dy02Qq/r0e/Q/CkvEux4CGN7c+qMwiv36oYqLT9Ot4MikEqeKzwi8fLI
qK25IeMDiLPmevzl2Tohlbo/NGtaATgj0kzRIFgZvxW7A+a151Tf7QPJ8kyRIfKe69zCbyOc/W1b
ThKoLoeUfPTJBWTvnz/umCd23beGax5tXskO1V9dOvrazwFpVJh/1xBNhKfBRpncc/cvBXeXaIpo
e6cubz4NRqpcico/siukzEjcriiLNTjbq4DIW1geE3/d9uDMrNqtBeKjdeSmSnFBTlrWjumvkRwN
42NAEtH1OcyK76RmGFyml+XYwKv/IuMseTZZRaQ6IDs32V7IqV77CGt53cV96SFLpIvgqd/EjX3q
YfIyOud8mwwt+18ckDdac1JrSIW2s0LUj+xJqb+BVqNGB9Eg5reMXkw02bKatxRM8nfqJQTQ0oOi
vb2yVjBe4J2bLlnV9Qe0ALgCDB3Z4ZLtoarPJDrBvhcUaQ1/3krSgdSMvkVHULVhwHprGq4W6auL
Fk5pPa5l303eqjzR2OSmbhcnP3lBNbrULSXHJcg2Vp0fuVQDbWfKwteJfGA17J+K1iPiuuJTB7lH
v8ccjoEChOVm89JO2F2g5TBQNArwVcz0HsCTqtW3NW4NenO1xdwSBCoCBRQ6r9/I5+mxLt9sdCIw
aihuqLlegjMv1vCjWG1yXROxbJXTbxB6GrYIQ9I9BNpEJ/tPnmdVYqAAj/ZH9CVIEBkxOzYqJtyA
cwpMAq/7QA6jbRmGhtR6vzYsAhvWNtL80BaZ/ExGi8RzTZXwcDB/VR4Jgb1GIg0lbKAuLGl3YHgm
toEtabunwkwCdlQVlMyhP9j8u0SNYBtgxrxemL6u/D/8XMGZpoSYlDkVfGKGVOu1USb5uUs27Vnm
UOrOMy6kiORJZCrcQSoVx+YNWxOn4OUtRxLvbGL7CcgGt24UMkwuPhvhNZXhpgz62eAVPFJt96/U
xq3S0FWvYAcDp1nKga6O0G874hO3+bkAJ3Oc9qU1C/Tqs4gcQ+YEabhJGvpptJf7zMO2l8cQQmQw
wyFOmXzp8cSYbPBnXGjRTZWvhoRRMTUwrNkkwHC7kLCT613LV07J/xblv+6wAQ+kLyT07A2D8/QZ
Egb6j5BIy0EvBPYMs7jjRY0sMnLBrbRGbsZHhKgYwQg096NW5Ojet9RW7g29Obw+11MtKgx7/ohM
CXiznDTe/+pXGIey/Apcj9l+SdlVfPM4ab1A5LEAFleZDvRrZiIy6deWPrO2g/6ZbT8yx6cf3ccD
nKFlWUxhThasCm3qhl95DR/yHpdXo/+jKlt7AHfjY+ouYX55X2fYq2w9S8aEvyYjDJAp71qboG/P
XmiNvUbdsVMr5QdKLLdUnQXkHAhGAAFAEkCrJlNBh8AaR4tSCWPXtu94kAzONrob/1fzUoM01Ua2
HPZfo/oBvZ9/ZpM1lWYsBBVMXDfPXePC3PFMptFoiVhpUe5ziW3GVF/nq64McM9aC4hfKVy6if/m
OhSMlwK/4v84NGqpPadkvPpNrxflLwTy78SxN2Di97tx3S+l3ndx6LxO6hJMk37KAhFlz95j+3Uw
e6GHDSm0laDY6GqTACuoOUfsmBEYwarebQFf6Kesw+ClCkD7dwlXbUAHFo1+awmh9kf+ie/yrGXd
lwtSfeXQyCsSsoH7JZWCeNBDCBr7fUkIEk+TTV3KbCz5UuevhrbCaEWn7kLM+lIa/jyW9dLA+2C4
5Ot68CZNoj5n/Z3O22qBmxxW4dkZuRa2j0KiKRAB9XzqTXncs6llKNSOcbEAlpnK/Ge7TW5I1Ja5
x85azC+09Ef21G4J4zgVXZa9b9JcElKPF4bJsvPu1MnMPBpawfzQ3BbU7eJAgmLTvFBaNOFNX1Ma
In+IpKRSHMGJIVzhLuoy4ltNjuNK16bMRx2bQnHgcUVEstMkOUTedt9lr8bjEjJCpVDG1g+enAPY
SKPecGr3HRi+t0iYNC8Gis/G/aD+8LUCnjyKD/NeKzyIO7jifat828nQ4/JHOIgQ+mWbVCodLdMA
prCIRkkylIbtwEdLpLJ21196FB9AzfqCEgauKjpuSq2Pg3b6CCIUVE98YMu+tjeFkciNaV/Hsw/8
J+wO9I1fhMQ4zvzYSNi+UWNUP3E4eYE1WD3zQbSv/s0zOIyqVWKEGB0i8UXS7NVl+2v9TAxTiilS
TzHdTWvYV09TqOW7L/zhGFK+W/OAtJour7XgYl3gxWx3XMYGnZzK2u4lgmKpeF+tVoyUkE1PSgSb
G5NQlh0kZgQ2Au+ZEYCfDMEkBr7veJZFCwjdnF7YQf7iur1DG9mGdDlmIr5SltBZoRIqQKGs1GV8
CdmS74nWmGpHN1aDuFBFIe6M/hPKj6mt/yysGwh+kkCpZG3bokIcrtu8wWYVyidi4FvNK1FCclrk
aipQBHQUA0AA42QrMkcDJZ2JX4r775ZIeaNQE2f5no5Q4Y9LBQzkEAwvnMH6SiXbdPGlUif+Nh6e
exDgXZ6d6e5PriCwiAm573vIgUWWqYufo5oYgMKS5qVGP09fA4gVMGRN4e0GLXKm3ie8MtrgrCYG
B+5Dg51F8eXlbxzIVxo1WljmM6+fCVvCVV5RwIVcGjLkkIuZEmlH+Y1aqoHNvJbaVBJqBRfj7E66
JtnEtzYrCVwH924vLNexLryFn302JZ4BtKHPfwtZDygMUK9xe1PFpkuXI8cJ8PhElaPUlc+7oqyG
8jW8XOocyp6pJpx4SfbjML5xxBks/XeG3YBL/ZUUmGkJFUpQ7J9TnAaC3K1bb26c1ZV4EACLWcyw
kZ3aLDFLxiDE8akugl8gfW5R04XNNw1CCpkvJrfTdP5jcCzjOfDoW95J7zH9HTfhNYyKz19NMafo
yuCWAIAws6wA4e3ceq+vrbG0jqMAEI5TEP/RPcNqsVuli1EhGNdCMpNy68X4dhez8HS58qesFvSm
pGBkaxZ3IXHZmPSil0+wSSCNpzl4mfbsGqwQCzAI7M+MLTC3aVxZg31YgrxhC2e98HE9vtrpC4jn
HmNa2rmtC0/kKTOam4LI7IniAhRXiZ0y5uEanivYekmNl0hG98XROPJCjRUbRc5e3wbEBVq0qD14
veERhu/PqFc0sEY7oYpK/hT8BsFNYH/cJfG1MUP3Lgda0pgRB7NTKsEiTQGRuJTf/Zjixv/3DGWh
V0mkxdpGHS6FuWZbquZBE8ecg4sBoebwelJEzZVmgGNLF2yWbil408HNNad4+qBfkzfIx7Arnldp
MpEvwXO0wlIzUuFjx0+SBp4Une6XBOO1ZwwUMMzDkdnOwnEpZ0t48oO+yS+V5yAeWVtXrrtHATbO
Lx43sOAjm+Z8XxIuVcygPe/cx+oOnW25FcXq5JKyiCCOYQJIs0CqxtTx/m2TYY0eA+Dw2DDO9M3V
hyGiZBOMjCa6ducPAmG7Q8TumFePE25STsrpHFJm/azgGkZp9HgeKxXzZ/GbijTbf647gep6CvIw
FjyFq2V5oPlhkMikhTbKs59s3Z3zYYEMVmLacBS+7zV8GS0x3tz++tWgwouMmL+UafwY10MBKVTU
PvNPvvgJ8IulGyUbdI5E82XKvkwuVX3dPNLVLBdlElPAZEry2iEQN1qW06nH6L629oEMDbQVVtRJ
yfKTiE0LENTsm5gylNohyyWLA1/ra3X/j7boTg2G2xsya36pA69OhsqOmepNnSZQqzmgqZi2T4XK
undaJXU3BmJINXw4PUhTpC8dzpgpzFPk3gRkwOf3DFnK80KW1/5JO190UU8Cj6Laa/2Iw+ZjHONZ
vkdEMZnje6aL4VHqblXCG7qVZtrPDW1hIwkCIe5bvuYfy0llrgczm9a7VBwNfE8ocv63E3TEPDdz
wWCILE9N5pw3hcXHc5LCKOgSzYxjlLu1nl+XyIfbGxJseiedn+OOIuR5RXMtIbBU3BnaRx9tw7fd
ewD1rufRxwEmpZN81HsFPE7E3koUeuxIZdcWcpl4wgBgSKOe4z2V+0IcCYhKDlN1xTaomgPofnuG
Bw32OEaEeO5AU3ymjUd7rKnNvvhbzA4aFqEkumh6KKY8CJhvqaaPX5p9xCvPYRpfjyCwgwPU+eIj
oy26l5TI+ebB3UcacHdeV6T9/Tf9uFvB5U8LwYII1MLmjfvRgy6Ndqr0vI4dJe6atSXsyfr4h7sr
NvRvfX2WRKePyrMZec/20yyDSpca3aeyqmdeuGHM8Nwg+oB5ztbHykRrJBXmTdE9PCmPANBQLA1V
czMCyiIDG6E9RYsFP9ivVv2OKqvW4V56ctVGk3Yv0/cr0PmCKT2ECm0yhPicczmuUbxe7O17By4r
8y//BWHcil/u4mbw46R3cYE/MJY221EHKsuf3hJBMfWOmRWTIxhuFZcDV/YxsQWPjJx7qgXwnQa2
MVjsFIkSdyeZn+kv0VquDkHuZNuf12EktBLKQecRK1IvGUG8SG4ZKSx5pecylrGm3z5AL8ds+q+v
Zz9jgTdeU+SD0tmb68Zu11AqhRPiKC3Pi8lZUUQyoNIPNRZI/uZRPKatbPKBtb/P4DWn9J4+uONW
JP15QRQ/cWLDjHDwTE2c4866RO0z02+xkwpeoDS1TgJs8S6oILOU7bIPl8S3vzrfBy1DP3t9l12x
JFS5X01m6z3M9xZfIZWNRHBRv6AOyZEvHZFVbJusOrJ5JJvpDQZL7ZEJhb5gotCQmHRWtYrxFBdq
lE9EDbZt9ervh58bhpMd9VXbYgQq+BtzSF1ZaD721Uu2ZFwUDEjwMqiqtQrHsNhcW/+QHkQgJi6M
UcezQEgJN2WFYhO4Lz1NXeS8UJZp+bhRHQbzowzVrw9FWoCmEbolH1fir5m3XfdOWGhjwm3rcnvi
eWYSqL/h+tplTEmLHYq8f33SeAqoodIbEKuB4v2jlphGWluiD7Qbi+iTfLNDTRhk+i2LRf2I5ARI
mI9pzXJ9wtASSn9MdZz3Ff0sC1Ucgffi0x9z5plSm3SdK1rh6CPFk0HQ4GCOufDfz9JiREw5g+t3
/VS/PmuGP+oeJKujb2LvFtwq8YbrEsjEK4Vt2+0t6iJKdIumi08w62WmiD4GgwKPR5E+3qI5j1IU
alSvfodkGOWgiHJvqc2nJ9uHWWQV2g5Myqa4RYt2C78gS2pgGjAnqYAKDJPexlSKxwZSAeT7jf3t
P3Ov7NDWC/3cgpnZnOHxH0hhG+iZU4XISw3YCBJZhmryWo6ew1OaMuzWCe4TRz1aiO7RS0NVO7b1
qJcvKx+PcztwVYe0lwN9EQFpKByUtsUoDlICqBZp57YGEDi1MNu+b524gBsicbfCjG492U+zFRfh
OYEZcqHJmXsWWw3khPneOOc0ORjexvlJp750XmTD5yA8xHi/cnRbm0pe7lzBPdsSuHR0rpgTLr08
0ibMQXrhhjkBSb5Pa4a+dZdUds7wXlnMRmO4dtv5xUsvPXyuewjD8br5FZzETyarf5EK0zIS+jrC
8r3a6M8I2K7GB/IEY1SRsVB4gT8yM3ZtXeHkf8FU6eK83grF/EzMJsD64dvtXmfVxwR8fDbEgr5d
jKtP0qtmBiJG3+EoUU8h8YEJXxm2xfoErMTNSYD1oDUcOX4ykz5peMpR15ZQVYVsa6niqmK9o/JD
jaqBi4GBjWQzrDrzGs0AuB+QWiTWPF6LXDWtq6d7kULiznBv47kKppCvvpmfHDOJKJrSgikWEvIa
I05A7F3yPwrEn0RQIUvrsH+8128olBHw/1EA5MhHg3Te2suJ6/hiNqQWl5BoqqgGK9Y+NfQa8QkR
/KMNcZKkKG6gIkdCeozStw6OWcPRDPoc5pPyRhAI8X3M/5Jcx3IoL/LiQ36vVqJ2L4DW8L/cCN6K
GxxYjZl6mQzQVTBEajoSfTFOTuKRTGB2oHDjujFlo3GZacBaRkSSjVxcokQcIWtSTRhpBGrHssHe
rtRfBIQ+6ro5fyt0f1AaDTrwzrBgbaYfK/j5gE6NV2zdPvGh/4i95K+zAADI02lS9TkHoKwYwDlB
028h2seRjWdhe6KmYFiJmBUu62Qxx1JAfYG8mzvL7QYUud3Z5mF6ZYsVH48sEk0kch+g/W6Ixyrx
aCpl+KaBA3rq88oeLegRze8xOmeVLPIy4SHzgLiUItmG1ymjVC445eeewCg6AkVhlYL8pdmv4W3p
G/PohBpjtTTzXGeS6koZev/XbVmK0yaZQVs6fbOB04Ws5Abi9cu4R1GPgQ+rZLHGwy7zdjE3OFpb
L6ZHo8OUTtImYMCqvxlN808KCXUwGmAlvW+/B4axRe1fA4dDEHZO5eqbp+dwFY7g4dyQsrm9d+CI
4SzWDaluhBMLuWgvhusj1KsXlNWkxGzETfI4KTfnUYLvqZF9I7loxsrd0vNvMR45UmqXmCnZcoBK
gTXptFpXZMDI3k0KwG+4XRoZ7flENyjSDJucJX/Es37p8bkmDmzAo/FoZG1/C0fyd1lrb5C60ApO
Rq3jrXueg764mGwFucUknh1i/E9489uKVI4VpiCvJ28eLFD1CYlglDDy2IPhB41ynWXGnVi0lM4k
m5hsjYlghFDRNrm7JMmMNvpH4godvcCjEPAii2/l7Y7NbLNo7mql9GylFvGko7iKUrIIUZRkXRn6
kLVcPVCmwgp7mL3ymSruoCa1Ilq9UKOWk0+HFKCYdstvTLS8sOpL6WsiF1oe7EEsMxKtzZV2Ld3A
Q15OTctSlE88tWRnsGVY1xPKkeIS3NBTJB5ic0m0dz3DTb5HJ+nZT8Kk/wwKk5A8HNiMv8ta7n8z
dih8jFkRXFtEmSYmqY21AGYSCGUb655FMVhVlMV5EyPuCy7FvjG9eh8ZONGd75u7pJnjORVsz7pI
50DhN+gd0othyBpOtmsMixanFWLk50zlFXuZP8IGporXKKbL47a1dLVkYPvPLlqCbRlguBA3x2S/
EGLdjYsROWclg0QHxp5yS23+DZ3X/gkKrSb14elTTtj1y2oOic7dMpvbxL95aHoWwidzModrCR5T
DxfV1Z96/EQQ+ZdYl/fnQVxd1l91apGeaz00KcEYo7c0lwxZRChY3aSf1TcXUDaztdMhTDiUk9wl
4/2dpw1I+PqRnxJFeZTR1mvlks1W/BhVf9exXLCje02gXFnq37lHKVmL3E6qZtquq/WVLylyxY7h
SmO0UHRA9QUi0a9ob5INvClA8ewo6C5N9ft2C4LUpNMbMuXym0uMMsBcLJln7ZYUosz8mhTVtlpk
Kt5T/GVzadQnHo9X6g5RKwYxHRLCWQyS23SKGz7jNFTAUuiyF/0MHa/aqDTx4OoyLua107KhKoiA
V+e20eMaF3UZVaiM0tzY4lVKXs8oywL1p/HNAkMcwWLBLMo1q2/gnTXWd5gu72P+X1vrNZmTKh1o
hFEjlZJpGiiMHegHHs7WBT/Hbd/2eSzCaX+AdDcCbzrb9pQP/Ds8IbeRL/0dfkDnjLg7jSgZ543L
GsfDww15bIFGkb0T9JRNcgKzQHVa2+JhagBo6b6ApcXDNyKpr147uf2Ktk1jI3L6yR9jqWLpkL1s
Yi9uVJauN33wJloRFcXdv2cnSVTm1clnHsaR6L+1wNJHhzRWb9JUJOd1LDCxen+gb7KKc84m9mrW
8eWaMomLmQ0E12SPlZIT1iHWhZjC+GJ5FyOeLBL4++pBJH+N6OrSkJdvi66OAMjasKOvRsnDpwL8
Q0tDBfrwoO9CmkBjan256X0e+DztqkWOb3N0VVznrFYJIACHje5nWaK00VECwIOjgnA+6kaLzLmM
GbT3HkyylgurbQUck2v74OasQz5RgLhxmaXJgZzVVAO5PnVPJCgDRH2IgRLU2o9cxIhAd5BY2Raq
H1j0PWv8RiyfSU+QFL3bI+eUL6ltNosjwO2qHbIi3xUxl32OiQjQVbPrc0pP1CDF01DELdPn/6ii
X6xXCP1zae/+dy/ydeGKlzGdVdtOKkZHp9CyHQ2oKOMbbpnKBlbU6aUPaptCIOTuoOa9lvxAhzAD
0GlTETapBZbY9YN9tuXocGuF+YFAwv8gLM3JV6NfxfU0NVEyfbpzuQHYrw3v68weYIGvscqKHSsn
LiyZ60wC8HdtniXntWnPWF9YC4KE4qs8TcqYqX7jn9NRKNwI06aThXr3Ux8BkvzAiJC/NU3n8Mxh
fxa6RP3FdwZdcyiGBUTePxjIAxNu/8C5fLpNjOEon0zLvP/Hf9ALRtbrrhmUyUuqQkmgA0Mxh5nS
2pAaIulHgR9jMk7NQ+AJujdSC5FxblycY8IYbdG1J+F8gkvk/ktoZ18yap6Xa7ueYsEryrJiD0lx
j4tzwh4SqwQaS9L2R+0JHSZsoGkW59/qCtkqx57GeHN2plv3E6phqqotfIKMdvoDqj9mEGYyBf2m
SkuDPCOnbLeC6Od0FMY00BeNQfUHbCT+/crX+yXDrPUUFaAO/nu/rUARVTTQCSYJM8t4LMNX5aXX
QWvIzawxtPvHlbAfkoA0Wc/Wgcl5+RYmrmQUPD0zX1k5hLAejphnpYYQB4r9ouYwJsupE5QPc+CB
8ZL6iy8Q171MHWa/ssPSjf1FgDY8LFek0wuCq0WYR4kmDBJ9htNywrOUIROJxezuGVRzBGGuyVQ+
XWAKkUE65GrwumjPOkD92/5DDSiec+4tD1IDkg1EOjgZyCwxLgFtL9sKXzmvmqn/Fze6P7SakWND
btUPz4XwsuFTG4k8o1mmPWPwiu4nfkwxXCFoVTCScrJasac1LXpULBs9lbcbGZkLORKIHWUrfrVO
BKQb7OX1h7XIc1jagxwz+WPbUJ0p6oCjGf20DGFZrHHLLxA8/Y54Ohde4lCvMu6xamFaN/0bzvH8
gyxOTonL9R9LhRzq1siCsjqdXTkYiiFWS1Gc5I5gbYwBZYzOiaX23XK5lCWwz7zfZO3EihFc4UV1
q8T1IM8Gszv/BqFC9Thkqauz5R48Rv00yWSodeeZwq5vsMMDGff9wBKRvgyl5nHql265sA1oKwh6
B+wH8AVTTVlTGGBmj499m+PayTv35eEM2Jsql4Kpte0KUt3/1LHKpGzIFcDRXo0RT3ffS0d16aC8
4fonGh+Y9AvqZzvcZrxRMB657MgiGTKP4yyQY3UVd+5mkadocOhUYNKinP9xRdWisnsOPcluZkzU
u7kDSErGBOpIhM+EJGeuNmnFb/WuuDq8LKKvPTVgdOApK5fgJX4IKDRFQAU1fJ4POWZMIMKPgCzh
wgsJ6AZbQ5Hk1fNOdQ6oY0ncfQP3sVzFejP0Q3GUKA01V04sJCwKF5cLylUOBjxZ2LpXj1eGvueM
K4EPfdYQ9OPPzTdGwRL8S0/y8Ag83WPFGRqZe7m7X3Z6toH78fM6QgtmWvQahLGaiAahecoJF5vl
+T66CxJR80ip5t0CxtnrPJrnj5QqbHp5887aSGfc/fIbckorUd4l2Yoa9ChKaHvzFjBlM87CRvqj
olVnyHQytaOPkkFIrnVUYwIEEIuX04Sh6cyZGiPqVn3hSS8VUAcPEzicJawIfVwkURJll2Zb/w8u
dSibaMN8tJCfl4MrQM/Iwi7vsyJCvTtxoHjEGSW97MtU7z3jQ2yqKi+JDRO42R+ZeS0aQSJuLF9R
dcQi+hNzvU2uvzJSgqQOk4579hrIjFbd0OSsc/0k8+k6R1aHDB1piIQwRHPHsv88nISUclO1Usct
b/3xW8M2SPoejuepnHEpziZDQqqw2GIhmIxDPxXSerRgcfwtsOAWsJzKk2mxVZ+AWRREz7/er7a+
Crq28QPHnDKLxWNUrkEOVFIQy5UPrtt7PO+sany4TlOO1IWCvXUPwPf2PC2h9Jk5WHcp34FHZyQv
PIM1Ggp2T4wmKyQ1E5XvJt0+04ZV9pvWHJR8DzpTuHw18ZktkbvTfsXqZ8HqGwBlVi6Vn06OURmt
ghtxfcEyqdQH5dKrK6gGiSDxzU6Lq0XjMfrHEZUeIPWEFcJxJqGgxqtPZCUalWYjo+Gy7932oY56
g3fStFqp+2GPQtFxt+SwD4t5X/qxmrwGmxWt+i7xLWjST74dEoj56WRoJ0zUpYjWYgzXwqpczcIR
YlrsXQXa4OQzs/XRONeyCALEhxf+T306DFF9s7/N/stg51VC3EYnsl4mZxdwmYrNKYsalC/cme7D
BNjaU22bnU5itPU0ccFrVAwbAS9HGQ84P8eSdBDAUf12ZkgBFTDx7BWiH2hqJk4VZ3vq0e2/a9Tg
E3pLGXt1paxVF/+WF8SEdL07OLEVApP0uw7+kdxtvlrkrOstMr81DTBTgiua2tD0qceGPsKEi6O4
1bd+t/MZYOhop+PU09nOY25bztiFS+p+wZSCggp05ybpdVsiwhVG+cjcIxvhT2tDAdBg5CHBCbVN
Fv7SZPNspxe+4IVBKBwvz1mBzSCajClkiPVK21amIGQW0QjR5UkG4xQe/L5R6VH9g8ROy0HhcxU7
AbeMLUoFouk9UH+oriXKtAsCYskz/bX+JPTKXE8cqfjAMvhVXneoqZsXI05nc5qGA5AkI9wFyC9W
1eHFr9kcSngEStW9fsB1seIq5yOWPMv/2arDIv7M28g+ScA2z3Ew6U5dM031jQWQ5vABXcPML3jr
7hISVrGX0Rhj0kVq0sQRGSs6XWjrwjfWFliOa8MDUWGlFelED43jhSnjUPBeLwAILKnmF2e/iVX9
VBgQNRmw7jJTsyJYqcgHgRwnFGZ8rIcxiO6n2l0vhi1zMWC4UaiJdyGJDlAZlINRivJoBWTsg4Oz
7ua9KNeck/Zhxga8B/Tm+8kFJdQmEX5Ik2b9Oat1EnMwJzeCubTelA2xHM9avHxH8guf5xb14qwM
93tHoX66RLrF/dFqbq2kV6aru38aGvZnK+yMEqMKuuAYK79JlyIb6tzgHArcyjtIiWpqLP1AUdBO
si0oqPw+xDVZqldDco5Wa7ZX7HPft3LnmXLLGKfU/f1ZvUKLTqRwPiZOnEcFEdMg+wM+vihfHbIE
T3HxQ2ScCkaPIXprUp20WmmFK3jKCLRMFjciwH+yV4BXMkrR4jjnzM8wTyNZMDHijEotIOOPACZg
m4PyzQnlXtP1I6Kdi+TXYGZUP+ICwo/mDbmqNUMNRAdY7VI3HCXy8A7O9KjJ5EfIziJpFhUZT2qY
siTfq9cXVPERJiL4kKZlBDl+mPzbEuLzxz85yXZ5v4xQVFSxu5ncCq5GdsqtIOfhI9Dhbruv+kdm
DH20DDGwVzbDu6DjOKQ4Zk0RJ8wT1wwiCgnj8C1mPp/K94N4POyar44rXIhSDNjenjeB6Yv/NwfZ
89vR+xJke82ZUUmd3iE4PXsRk5PuYRcaGsvo8jfRx82tDvfOVOF66HOxLO/C4YpjnZ64doXSrceQ
tTBV/GkrIrYIWCEDtjpT1ITaLQaLb/1HqmVZdgoNrJ/A+dFEUrCUnhWpqWyBUYIzAkILYjMhOBJu
u1AGNsqHvbwAifUrsc3/RzgGqwKv0OPcuqtwI6Q4dhm7MBiQsQ8JemxFU2WgeX9ffnmAEOk/vfUp
B5tlUZm2+VK3NOZ581flAG2CADCjJz/yLhHginJVfFrH5bbW+vZoVFIKAKOvQ+TrJIWZsVCFo7o/
xJ3mPZAEN0Th28C9vUxQ5vKaoqdB97LO4u5CiRc+LT4UvgGPR4mnlvcrhEAljfDZKLVs1S0zJ+yC
FUYNJRDntjQOCoaxkn+EwFA4c6A6v1V0q/Vxz9TO8s553q0YsykzAQOu0l9UX4Ty0uhULK/nyr2t
SFNceEraYN7vnFVS52hgXyoEJvWtdM5MeJw0p7niBcn5Amv46obN+UVJ+5Hs5K64jGJKaPsGDNDW
V6JQZqvkjSHVKH1Zmj2n3+1zds9qQU7oTk3lCc/gCeRSdFTCc3xdB0n/KwsLAvRiwmjyCWG5Jeq7
RBbYPH2bjH5+VJGhjvbClxEis8ZX61Zm0Kge4ryhDtu8EwKrvvaBhzMxa7V6Me413oLp2LuNgad5
OmBe5veivOXmEZF/Tet00mwVmdQAWHLRictYnrNYRCvhUv3wxBIDn3cKQWw9qzOSbJB8V75I7zsS
8JBFtU+T68AHByo79xxLoDTcea23kVF+fAuczDVaO+H+xzS4YowVOTF0x4m7DVfsj/OphHW7XIzT
StNoyHPtmRZI0z33OL050SZV80GPATLe/ceYKtZbskHwwl12eaXwMjwFHe713Be8tiVn/BGE6VgP
JveAdFMU05y2fAEjxGKclKdtZQdwKwZxXy7D5+j0igGI3zIQawPqUqFnP0KZM8Dfcv6NIZVdwxIJ
MwCkr3Cm8U5eoTCgmbzaNOS/81VrC7OioQR8cB89ue0OaKiSxuTGePw+tlPZuDg/CijwwSrLuZSo
4dnUfR0iDJ3EIlpRjRMtOkmCeCnz6Yeqq+nFo/UAeR3hblVU9gXLjHIFhglyl7/TDpuvpDc8b/aW
r5G8eNnWpAW+Q3L/WS/zWh4dy6LVK+q9IfmPNzflxT30DkDB099Z8IyThEEM0M8hAJzj6JDXNoKj
u79+aHnn+nOLLp1dmekyd+lyPKe3RjotmZUWEaTMCEqNAaGDDQvqXR5ACR0racDt5g3iNKExUShl
JRVQo26qXFJ3SKtQwryWISNpBU7s6Wj9iaPB8J+lV99BQKbquelacWivar7u2uEYq/0SDLKlCUUK
gFbY8Lgfrw6xzfAr8+pxhEKJ6iXY/Cz+XpOGa2oyHJMlkNCdUhX15ZBK+5w3DnWG0DfqR0yQeRoQ
RqlToArfidcsxdNN9Gg+9qBR7PmkEPAujX/m5HTCLFlH6IwXFFCVLIsk9/cM27zo4Q6E1TkAnelG
EZj02gLzizhvUXRZdUzgtzcnArAnw2rliWj4jfU8MrOLZsjqDCNXEEcuokLM2ckvhM2k/0vLbBIr
odrrEukdpN9FyUj/UR2jyl8FwS/mblX9psiXncqqDG7kapfWuHSnL6hFKpz6FwlZMVo2ILITUX4P
JO+Sl4aDFcjBoqNPpCYOMsDL+Tmx1cAX3+Vg/wFTuKcnyZKFMSC9/g1Vy4YWB/mZHkDwZFF9bmdX
qhX4buDQ5iFEtCCgw59TIQUbijOQQEwjOgtfB8WbBnuDPJJIalz2jhJX+G4FXDA1vnZn1DDLgC6a
+YFjU5/igsmChMgZ2OAo8ULS9chTYnR6H89tQW0pXQN5pSKlJkcmBNzTWu9MyMK8mG2003+qLBeg
PuJT70vq0fOV804SSdVpdqukwKM1TlPLz5M7DvMtJgA9toJKE4a0ceo7sutPHy3oS4we1gu+0rN9
2N0ZN9oCIMqjnOnKwN1EYxFt2VUapikjDFjBOfhuy0JMB6SZCvL8wORygNLnISxgHjo3MBUJUWE1
0CA+lcbTugcb/AKuUMiTYmKUeHNNGg68+Ci9WUvp3rl3oKoyz8fs7dfAGKiAbTL2uAY9gg2SwJ+D
pz01S7+Da0whT1Va6orrK6gmVk8AiY8tPB6BOTwnxPrSRIXVNjXW27MEHeJIwXhyq77XmH8A8OVa
QAiyvtkNKr5XBLMkw6taMa+WecGr+uw1Q6D+sKlqLVMn04yjr+QnQ50l605hmShSrrxQ/IcTkXQp
PWR+2t9Ck1axTfMLEuiKXZ176fG8kDc9uSzbD5tf8cjcOySDCdUh7cwPRmErvkeJ90khfFMclFnY
IQXLOX8aorTnOjhDEoIeBOEFElVIf4U6CkRt6+qa6DwbCA1qzyfTlff7l+rM4jcb/cJK0CD44EAi
DcYSI1a6d0DxC7quwP22Y/hh2Bj6MyoNIXIn6iZvbGBDp2slRLs//Ia9HexkKj+tp6VwDME5K1DJ
ku+oO+mz92J7vuVZJj4F0LFi+Uci9+oPNCNwzw9F2fsLUSsam4X+Rp7u3sSXfNARLFmdQo+m0BFG
3AbCbMa+52rK64If+asAvhZIBKI0xAGNzGR3cxDtTBFin8kNy4QrEvGgP9vNPxZ83/tGDnnoMUPw
27DKcRBYi3VnUlzELHaSTVDrScDBJer8yEB8ikOUAIG8R7yTCGNdgqZV+kUzYUfqlidvPZWrO6Vm
GOATggjYO47N7L3U75P9mzMC/s+F0piCwz29f9Gv0H2GgL6r/GViR9/OZhs2TsYomR9c0Pvy94t4
SsArFCOl5G9HJ84dNvs9UogKmkF6tKPHI7UHnGLzbYVgM9hd/qRZdptfXzPomibBEtIfbxbtRSAp
l7JCZMZZMoy+yIy7QhfPk3gLzvbkG0RML0zjYspwVcZJqslCNV4T2Y2SmebwME8SJkOo9AkfeqMW
wdE20N2AhGxni408SNxGFqRZSb1NHyZvWX1qU2QV3A5xjQaDkIRaiph0UIATCoR9NenNpvOoNe5Q
aDoCsAH5Uuf/MaZ94SboouaU+akZSM0zauToFciDVeotk4rEiFC3fu8fio7JscSgxVf14T2VKQjL
Ym40xt4lohGk7bUZbhB8MkTrV+hNT/DJpEug95XmEYYTpI3kHGvKrfu82I+APKUbAhiYeqgIJZHR
xj5m2XkYxPd+S56sJuomHqV59wxb5dZf4e7DGt+7hKt/tVH771vaF696863R1ALPJRHQJyte+j22
e5DjbKzuUHMI+fEX6SGqWfF7OUn5Kxn56/KQvz7iVjoXgg/UhKNlObZoPLmam3nfdWG7Jxcsqr/6
CKWfUjUSxUwCpFyzT5MVJL1jFcQJ0vdA6j/mkjamnWHe/uPqYX3Vg51zY8Z9wjJx49kBEEZTE4b1
Z4hU0OQgxxarJuIbtWhAq6GWt7GbfhoAI4ln6qbVk6SEfrqTGXPFYeWXhlNc2+xIUqTq/tews+9o
lE+5jMYvlX2z562mcEDPCp9ik3fhgUsMylR3oqC2qm+b/QIFTAUZbPcjL9Lxcn0hhmEWfqt0fzV0
crj0dXXCoxNhDeKJve0IYfMAlkZkv9KNT0jMJSBoOKwyqxtXOGgSSpvQGjYYBviOYAAZJn9Afx2j
9bcvbQ8gCh6+9tOQSLmXLRdtNWXhMypr5T9ggmuqyX6kWALAHmB6zKthR8/4CAU78pEmwaHH90cn
Aax8shJSy7SasTYvIsr+X5AVFZoPmUWiS4gYxqRVsotL5EmI9x1MEc6LxMAv+wiObwZHAPDPXACs
1wEpQ7H3PF+U4upkPjfvqa2xzJ4K9VGKO58qt4ADqxHvGV2VTuCc3zRVAxD62+ZUFHtg7zCSVhrA
tAZqE0rJ8kYtd3jxYrwQvAXpVdtEqiJgWWmqe+FyhJWx1BByOyhKbMv6bsr9QwBkVXhhkyxZxikt
rfde7YTvBlfjT27ZmPJYURI5zrigFPtsDIY9wesfamH5s7+3b9QqbhAbfuTnWW9+hzW/yRYvasac
VdtZAYUQZTFSnkFamnfsKgg/6UqLCxSVvfrkf6f5OuVtO0JKyk4fmmqcRZPs9OGIgDw97mHrnlkt
biUht2aVrEkCHm7SCBfrxOwfXO3jlh2MMq0uGzy02uxDloZ6vMebiDiq6OSWu/sdywRmrN+Dhcvl
2V8uC1lIlQ51nbYSihbeB1yYGDKRiK8cOvsz9iy4gC3yMQlidPZAeJGTvlnn0j2f+DCWebJ6fVEH
IPkhcWhXQcOEiSVPEOwzE2+wBhmDkvoxx1wWZ9KUPAjYQXE7IdWMIff7+Avj+pSQrWBxkyOCS7on
czRc/aJr0spnsYy3vLOUXDA4gVKj0Tu4t4guKgn6u/TeLrxZRsM/jgXoxhFfIu23zF9RUDKZsdMh
iZ1StCrNAgJ2S1nz6VO7XWzFuBXFZQPKlufMcyuayr9nOQSDOp15Suz00wSddMXROUUfa6oonsgB
7+MWFAbF2gGQxa+4ZN/yl9c4PYVonGQj9vKEAGQYG1Wk7CTwKhZAwM99npo1SKwy1Ormp9KbDzgx
q37eHkZ4A8yFSRzBu+tv0BfP9buMQMH3QNsEjcw2A/pp2LeP9l/EpOkSqu8R1ANfNro8PN1dvwvh
iFDBtKq8wz0YuFiaE8GU84qU4vHQOTnXHn2Q3UUD61EqS2TCoMJhs5/K+pPlbxj688UI891HdMzf
mSQW4G+Q0IVhDRvR2U/AoUR/ZoTPjpoNt0X9CZ13NjLeg2hZSneDjIu5VXBXhyvZo+04MttCftYK
2buzMfBTlN5h7tdcJclUhs94ty1PeC6YsQmb1c0q2zom+hsGMPLQFMa5kFNnfJYzSQ3e36lUvN0H
8uj5uFC46lmY9SZ71Jryxdp1+oThhcFcvRIXzgkk1Rdd8bdc3ex8uhz1vCmBrKWmqIY/dVw8Goos
LjKDo2MdySNiEfCKxZTC3A6ewkncOCuOLDRmxB4MFxWBhT6dHYx1vlxt851Tlyq00e4AcV8+jLIf
CRD8BXlI9UB/yMOzRdNVeZ38zZ8C36EX9biLGkDxnDYH5Q9XeopgBfhIVMon03yXziAHWz1p+nk5
EBvmb5s3405VOQanmOhuZC1/BpX2Si1lvpdboZff8/dR04chkV4tzqC/R4c557TeGWxkZ3W5996J
kCeGON5+0VgQKAfmm9tN5mCaAZzBpaeVMsLorOCKy85PxJmRhDXLbD+a0i+Hrctr2NSOOjxAfAxA
NF9+lRNDkJNKNNy+9pNZBuY2LnV0eEvPM2vKWSD1rb/eNijsa84oq7DjdPWW5abvEb6r1vtJpJ3G
tzeL+9b+MOmY9nzA0uZR1FEr8Ik4VZcF6U2g8cfVEICi9dGCmzKfUv6EPuIW/AkTQ+ZRLYpUpRBx
m0U9nnBNjPQFauR5t9jWuSXGdPvxASVpRw6DWh/X11tfB4f6tLvb2J8FbwlhuvPBuAQcoOkVN839
MEIGkJF+wMvodMkyVy9YzqaGb7WuPQLPngtNinzAre/U5K9+XhEMmFxWI+0//GgTvzYlAdz6TXTV
HmfpIDfd37HYYWU82GLRsyyF/Tt/eHHJJVUfT4Cf12zoeLFtDm9gZ7T1GyT74lj8FZfhGVmLzLS4
5sTWjGVd52eFnjJHwr6Qt4btbC4gzR3vNZd34w79fRnaEJRNX303dduqhfAsAw/W9qXc8jB2Q7ju
sQDA5vO4kUKMrmDwhAU5RJJ6P2oTDv8FL7JPG4NAKBgfCpMDrUSztaNOELG66vdoEVLxEQHn+e3B
uKv2IKhw0iVQrpWktkK+QtxZP1Ejaih4RPakZEYIVsubrY+TvSS5W4FSji7W6jiQeewTWOXnWbBP
TRCIYJYjmuSv7IwWUCasHRI3dJxvzzIGVenuMeSW/UbiKyt98mTAdIrqoP/CFSkhjU7pUURcT7XT
R7m/eoh9Xj+VQTSQ/eCPIJj3WwThacfexGxCfxS6X0/JsfICpmo8wavBPFZcMUZCI8KCa5/StCVP
viFF8FMh8CXel6akX6mUyEn3DLwZ9Jw3KFcQ9QKFXPqEoPVbbtrn6T8Y5DIpEIxftigedReA+knt
Jlpy/0wej11Fi+TldRjN1/Vp3YThE294TJQSq+KWyotzzn8b8fk8FjpGuhxUqusCVgA155tLNyfY
MSSZc7ri1k4Et9gyo69iUN180Gr1pN/6xweZnLTx+HPxrzpUDP+CMYq69DJVl6UMBS3oPq1WUZpE
Id65kGnvtP5Ecy2hW+uiRCqsvKmxqhcQP+alqahA8QM5E+AVQQLK9f+EbfB7m+9bsRB9X/Jta7f9
AYOwgY9Vb/a9aQ7toMkzwvY2zt/qbMepM9bAMv47qVO14njkPlHwoRZKTtlHADOQ1A5u3FbdeFCu
Y9ah0LG1GJnSKAKwKVKHmmlZUl13rspRSTNwSHxw9PGm+x8Cppcp8ePcVVDPnI9aw0brh4Ot5TGF
+ykOIyAmf/HpqlEidt2Gtmo2RO7sbO9Pky9MAysAIIb1Dj5Hp8+F4cVd3jpUI8XOg9QeI+SSYyZN
vXQV/J4idqqyJNxUDPPSWW3NOeTNJEyGo3QsGAuoUYM8l9vrE6lZ3MyvPELw1cCLlhkafnR4LwHj
qK/nsRNQNF1ZHDN/WI6ZKlBqyF1vghifLiYyn11BRf03os64Eh3kS4hHMO5ynaVd/dGDP/8kUQA0
EKTCoN+f05rqC9ciKP+Pt5o89oK83bcfoC8oZVbUTdI7sIcz/UvuFshHt3D/ZU2BdD5T9AfCyayx
zf1kICHN9ucxTuuMq++7osvLSs6iiRsgecC3LUuy/7tvUQpB+wGR7zM4RIyIaHaSiteHSQ/wygcE
NsOsVGFlZXkjsVUax2J/csDXYgSycUoEMkCafIWb7lxlgyQlfR/3meyHBNyCwnful7mCCu8/xSRc
xpNnBT7KbmE869l5U9f5fV1O072RJmwAK15NV/1cXP+7c117M02dWgwDlgzKoTnC7Zk2sYvs3cac
wGskfjHOccdFuaAYhdiULTDKusAwMQGspDAonbRMkxaDQWktNLfFDzYb8tFqmCC+straft3UqyXI
jHmx09Tzvulk0h27TOAjj09fmKu3dO4horrGlt6McTZZprKkEzSuw71e7gxX5J14QeWNMwlMcdzs
kNpTVAH/xInGuq7N3CS7pNCjDnpWp/hVwbRuiSVCXAKEUjdl6n+olKeH6RaRck0Z9Mblr65Xsra4
4eFVYxgBo1fRClxOfC5sLN1L2YS1MwP8WfX3FG9V3CBlzxet4XuPv6+WQeU7f1dLYDkWutQs3nb4
orvFbxqVwnK2IagWQN6La66gXjYYvbzT5zC+KEJCaqFBP1owdrlJPeogw67bk0/fhL8MJHj3Iz/F
fGqx2ch7hGL1sgN97zk51JkyYnHQOnQ6QCMEStsfAEBNm1h692L7n9u+Eiapy5OK8an2ypLqMpBJ
BMFXPbTckMLVRCbSx50gPskd9ZnhxzKdqvuK6o65c1RUaCr/PMrtOfmMnsEBsiZDuxs2ADKS/G8w
1+RfUOVmm8ZWi7ipAi9lNYcuekBBYtx2Ao4rFPQKeoRTTQDFYoIxwEZzl9YU4eZREerm446cAy3J
0M4xDTXVyjeIoLkyzwgwurdZCBkhkILJImie/Q1CO7ePn4Kr9LP4D9NK/gK3WYO+/y+ynEYyzAV+
RrmJgxV3jUGY78KVW4FvZBP5/kliUHZwdG+F9Pvq1DdwjeYl/4uw8ceCunpcej2csDiGmQdXbl7d
8I8dgA9XtEnkk0PJn37EXBc0PuJdNPBTTeQKCirzc+JxVSodaicwNyFIiFTD3r6WMv7Hzt+7760z
WsqaabwtCc5AQ53bR+uT/Mes0EpBCjM8N56mqlmZwomnGFojb4SjzoXHOvF8+X119k+4NZgggQpb
pSgMJYvd0ijqgXxHfEb1kQAtazx+xzrUhF9zO26rdZsCOHDHvYL5WBRuMsVxeaaWLofp2ZRs6ztA
9zn4V2/DdRuH7HuV3KbVsefcODQNRNDvi2goiFl4RD9U4DjKVH8LC5JGFCUoV1q+7bRezeeLR6WS
Ae0Zd5CNUnpwTdRho5v9Q7n/s+jqE7agMRjDsVshz6H4Zn5091l35nOXxWyPQie0NP4E9MwG/Ybb
wGc6iAMSCP6PHUlTFk1R+dw1wE1FUMaF+6TzfvJvPBKrE9D8pPRPcDwgCmVBNTK2QLX8wi7sjpiZ
USPR8xYP+xL0OYMC1J814tz6vHkIprhYddi0XVEZYIOwbBIEvrigVQvsAdsAu0XXAbu7LFlrwr5P
oGfXmoHU8JWbu6kiHfKH4At0In2dd9M4Og1Ege2YBxxODBfJgXx+TBcZRWRiH6GfKoXAU4RHOrJY
yzCssrD4gnZ2cbZx1klgwznuugdrObcWna2qYUcZXDMiLR+wKRVFNpvvc0OGbNFUlmOUvUjRHsm0
oeHDMdUOszSv2Hj80uCSwY6ksb0rp74AqIGwPQ7rK5DAm4Cs7bgs1R8tSeWowkdhIWXLKAAQwpyn
RA76ukh4jqB7MMpa6xrMq6bDHyj1LAkT9sbOzzg+PAmT7oPGUgEC1w7+iuLEFk6lMSxXugYyHXAT
cZJ2p2/NONmd6itg9wbksOkQ5g981OZqk1CQAOP3LSv4NI5sxlkvEW39LzhzIVfWgeOLkuG4vYGH
Ph5ZUhAt7os7XC3y2ItWi2pT7gN+c1GOtYjj4LZxdv44Z2a7ooSn8QkIktD9U2qyfkplZGWnDHAG
yKPGK1x62hhUqYBmlKQ8gyw7eRfdFnVZnLSrhH7aS9Ns436E6UjnAKOR0T5XBN3/qYcyC5BqEJnp
h8gjMG37VkUpbRkWA6GgN09Sa+PhX6ynil3idEIMwzpm8/lhCMKjSOOs25adsh7B9DeC/YGO88h1
HFW9H2cirQqKEo5VCg3t6WIoY4/w/dNkmihB9IBHkApZPD32pK924N98R0BWQa+nHc6pDsnOUJn/
pSDySGr8cEIycKiqRS/WsyoEUK39PoYO+EBdQ42bjE7LPWcBy7jst2fYmGkIN1y5STogjw5yXYZl
LeVyRfOBqDnWT452tsc4QkrnboafjmJyXMBWdy1hef4GVfhR+bFKfOdyYOvus8oRPPPDjQg2Enh9
q4iHsIkDJlNDysNZ39YMQMNyCQUKitF2vC4U95YRyukjedaYG4VbDQA7m8PIGflO+51U1iSGugWo
6B7yk41XvhMegiazK0jEuEXV5QP5EZ+32N9oXXd6kYmPto1s1pcEoRD5r93Nj450IIJCzdVnWxKr
f2qDmZqT8Iji5YeYz1zVDFSzhyI2eT2Zyhjk98j4ycLMihlwOlIauzNI+NeMekxWmMeHAqhRhcu9
q2f6jdDIepZMEH5LDjyvp54M3srhHFr17naS4UyDZJ6do1Ft68dXqbsZa054GIHiZ/kZqI3qVfFU
X11QCfli54BdYzRk+byRDg1C27s560DKcRM61bONimY5FgVKHiUzbSQAV6B5gRANLXnjnfJYTO8z
vHx37UfZ6m1zpD98YXPIx8/yq+aIGd6KENjpAMe4agu2X7DtgHHhIK8WYy3ynmTOz/Mkb7Sd2lf+
oU8trUyA3jEAYdrWjMwIRYijii8iwiXXYdruO0DIsPepCJRpOb4PxlxG7ffpQMoQSMRrv9g4LFqD
slkAE4TUPBNMraT9uD47duXbSQhdDtObqb7TqWUherU/dL4wlQUqdTRx2/iLKhdjg6+oa/m1MPoe
bb5LSTcEL/D9dAj3nfg87xomYltstnr6JExfuPaHiug/8PHSbsgYcvgMOfD4kYn4L3ST01oPH/Jt
fWrl1c35k+aKyACqcy3cg1shng85TOUeJYahBbSha9Ar7uGvKiVyT9+T5HeEME08iYBDivVEGrdp
hecZUQZXFotXEjh0afoZaTzVEYbhAZvQ6T+EE2zo/Ti4m2CHhfCXh4SFK/PR7DuZitjdrEgaih/u
9E3elNbWr4Q31YiacLXxrFkFhNrpEM9YBOZ3ciXAtMHS72krMPz7qfQJPbs4FuCX+9hHfXZYx1zV
ku13uEScTOnzAdGofaiM1g2mvd61L355gIuQCbcZy3j+WlXsyZB4QyLLYGu4EY2Zy/qspFk5oMAx
IDYjwRNCM1YmGl198C8xdW6isZR9rni0IwaOV86YXyGrDOU2OuJjgwcFA8qfFHFth6a84JpQ9y1D
0GmNJPeOZCrzlkmNcLMzRGdWN9Lawq/MotdqjsEYXAaeo+gBDVS9icxYYvM3Y3/3SCZmEwVhuTrE
E/HxrQVg4onSGjQhmTHWny+B0VH+osSFyL5V1R/SDv5Q7UZKbphxmKaWYWgV4fWRitE8mwDZuNhY
QZAOy3QtvMXBovXI0Y3XShP33/MFQGy8SktwtRjeaPBeZ4RqOlS+7vUAGzPpDO+mAHI3LHw2ao7D
KlcIVw1V27KlfcjtWYck/2ni8FL0AMNLXsFbPR2zrNm6lnGIL1IxAIZvvQdEj0ls1TyljYvT2s15
4IjF8Tg/fIh/ApfztkYBmqtCuKEi6xSIHT22STdg/8AJFAin4imr1EtlMHf6rkEjZbBxbImFCTRP
U1zxs2v7SxcEb2oM6B3LRjbigBWQGnjMsIPTFkySKMBPt1Oo9/xORsqL0tZjK4FSAmKAXLYiHJ9v
1tKuDotyq3XCpIa2W1rCY6kRDP/TR06jdzaWVVtBYlmFPWTmQiqnnANYZnJ+lNmKISxD5ZC2udGW
QB8ahRSZ9qL8nRb+TfIkWpaZibSRDkljJdc33UR2P8LLUvfZFieQM5s6mP5UCTnyX10fOYrQBB/g
okddO4tJwDVkZXyVYLBIUj3uRS22Sp/Ho16/NEV5NS+mOvDR2b+9OLCJl+HmZmKYMTlIAJbJkA6g
N4I3knWez5HNKJoJk7SkGehSAZ33GX5qIwp5Xz9tefid6r2l+dVeatruijVM2UsxJEkObFoR97AK
lSZ8GW4kLKGaYfNQaWr1/Fy92ybfs1HobsfH+fZno107aBF3xHQsrSCwNIDyTaMkjN8Rc1LZMnca
hB2NVJi5pqUB96b3PZ0TVu2IkdpQKd+4WJqm0Cahy4oIzZQenuOnarB4LfivT5+rxzHT4KUF0r5v
Jmv78sctWg02dhp91AS1ptJhzgn0wlCqe2JQJOGQtrqCzNdmSygxdJ9/Ix7KadQwlj+2d9FCOFxi
4LAaTh3rs2D3vX+G4UMHgdujwJnUOl57WPiI0G5HQAXJMnk2mftIymIQXcJDaCVGavQCMFSsIJwT
R7OulXLmA6PnYmeqiyJogQ2Hnt/slqfksBZQECeoCbct2IBfSVoaIGD79jDLICMmIF514TSXbQ/w
xOv0ivhiILKx4n8nZL8avaMSdcAM2QhZLFlYJf+Odd4YLjxeeW9ebCesT8a2eZtm9N11mQYDWBQn
tKVQcHOgwmy+/FZEjs77K7+I7i6F+s13RUoqvbkw4vy/zhKrg45hYjYybI16slzOEyakBqwbQfcK
IHRky02nuamFNoyACW8/xs91nXH/X/W9eMqxDw5DJfb54OL+fdZ3Jt2IxKN3EPusjo3s0AREQ+Bx
YPa+y7REiWmeblIJukq7zmfDZCQka3cQJrUwaxgQcaY9WQwHWeOMctt6iZ8hcAUq29XZUW9S7NCL
tCfR+m3NKL/SKCIhnAYH3SLwJoSldUTysv4tdvfqAygjJcCq0TBrJ7Evj+4VOkx9+yKH1MnJdA3R
UMeTwcynpVr21EpPTOzrCT9DNgpPe9LJSI+LPlayKu4GHMSVa6CpTRGhxKFD6pwCpqPsIq4AfcQD
11hzLwRLLulN9t1P9vE5fZrZ5pWTpBcfdjDm5xyt/qp52uCE9bhdwMRWJGcBk8qK1JJ4rylCuz37
CZ7ANWg5EPVHypuLTACnQ8WU2vwjVeht9WL0t3jR/hzKagfhj7B/pHe2dkmiCE2CBfryGX/HTWv+
M0trrGGKv22zz2BJ7m6wftVkMag257S6ogNlLWZfoCToNwRuNd+PzVBkrBwq9kaoGkCCBg9U1Cyf
Pmst5StI3EDTe5BXoyuuilEQgNZuriJveL6ryPeFl/WM3g7FhewOzoucRbtYt50Kpc6YzsYwWr0J
dggoBJC1lChJ1ArVxzxzdRF2SEbAdzm4imG6WG6CzClqe9JzT0mcBFlT4P8+5zyMOlDXLcNylSLA
VVhlNQTzBVoiDwGt3NGFw48OVZCsZAfbWcIj0NpI+Z0aRaKa66XPzuBPz48RzaopFVGd8sci61ht
CCAUMwWsDqmZsc4Nur0FjSEpMuPE2QKMbhj3sKdvYLdFtASMTPhgQKf04US7HIN0Dl0AMh6PMxkB
pLlt6vJWQxo93PU/8ZU7E1XmU8ars7mjpUJdqFhh5l3f78EfuHJ6wALmF8EhyuipUt2CpMogb2yC
nKoIts9IrWbIDDtioZKmzmxOloBo/xjvXAEn0C419ZXZ2gdKOM3i2y7RPuN5R9/cN8YpD9ZttMK0
UnUNpwPzS/l7GFbfcRjMObaG0dC9Of6ugUq1Rpnhk+yxyyN0LdbmtWNTPeTwRQLp2Bb22h2zb8SP
iDB4yDhtX1h+9kobWrXrkZKsxNCpH29ak2lRR1wMmPIedFurUSBYv5+wb3YBdtJ0KHXNXESA7YqZ
x9JVpDlo0GV8Ur9/Ehy/C8HTEt2JtgS+QuLDb/QSHTSf9yhYm8E1MNOMdAV4svZsVNBRepKiMput
LA6wHv2EIPjXOZRkxCWQJLtNrWGhIlGdYljAhVP4ECdeszbx3O5nShFSYqpCmqCCBgP1ZxC1vIsw
qFcuPFcDNijkjm42XaToYMeWP6pE3/4gCAMStII7LY6HeP/aKiF4EAFNSChy3+BR9/E/48ZQGKvD
xQgN6P0NhbJRzRWsht35o2xt2aB8P6G8GYCjQ0iW4x/nQuMjxuSP5Rci4+YMPc7uWjobwQAn7uJV
/WTrgtn4qDoGoxOWoxN5PLJO1sTdcKQkaEH1grbB19X5D6NF1s/fJQnN0GCwsx+47zupp84YdR6x
zFwhgnh7pPms/FZ+5VzjsfOC+kkzW4jpbcFE76FKFdZM1lQ5sdGM7cpgoxt80cVBPd4cUR/bBem2
xy+gKx83EZLpgOWf0oliH3yU67q+AgfYq8QbG2X/xjlipz9BaNyc/50vMDiGEcCY9cXw8YU/UmoX
DSUfm1NL/LfFbRChXtVLyC7SRWw/1lVyMwsvWZ98yZNqmfxNS7+8842cft8tRresHKfnDr80nzZJ
OedSpzTVrgEktDTyKKg3PiVVIhl/EX3niHYnYurUgkIzGJAajPr0+m7yASN1fYBvJVjlRtjEW8xM
hmoreAT94STpCLd3dtuZ14mhCstx/9lokaZjlOSrBlCERiPf8JtwVryDvCn5eVwEgDPoHY/6I6kM
ZKrEq9toa1zDRKFrG58yD9exitRuS/eEA6XjNYQ4ypcx88BrDD+lYCDA/k76291AmPhWBLb90EON
oWhXsKWS06SQiKG43R89min5oVaDm1pToqa22gxpR+E3R3Y7h0oO/Fxg50hS/bztfnXbH8R3viPM
0X+V4QX3Mv7C7kIV57O3ct1AUBUhV1L/49w+bpOozDHgbhv10mBOEiRxOIbKOmNweee/W5FOWL+E
dP9BtPudB7A4fj2LJwtpQLMI3BRL5gTLUQUA7RuE2saUYnwR5GpPdw6CB02pecRz93XjcGfRh/wQ
ag+IIRaDs9kQmk9nYzKY1ZFeGKRdGPJ16jW7USNx2kM2Tx2vV0U4T0kitnyVWBA7RPGW9Ul+gfjM
tYjcRdEB4XDHCqtn8ZteIDIG64pRk/hDi+xxL/bza/OYu1rOl10czPOhhpuQTeeolTiIzP0xuLJW
FDLechqrG9pcLMthX6DoiHsQhGAY/uZbV8O3J0v492of4PQ2Lt7c9i3f0FAt+9SSrthlzjutS2BO
QH2z0/K+ewZTUp7F4dS6JJdptc4gQhoqsYGA3xhAFgpnVpp/cm5pNp6HxLxpsXcoqI9znXcwq8XC
7F63cIeZz8k0StVHMzESC+FpLFfGyVOCfL3dgePPoI/kjnEPVORRFpWlB06O2PVZqlVkr0d2WMxL
eDqX2rA0YdvPTA/zEQs0xbuJl8eoEB8taWpTEBOQoqeGHp17VJTU3PIabcdqH9mabxirVcnIpslP
X4s4gYK49ZPHEZ/t3vfV4uexJLmGcKMeCpLbgh0trgHkFVbWC4Vh8KsJat7M4VjUSeRTLc+G6Cpf
UsxA8Vg98ugkmEV215kXUIUqywuq9HwHgevUb6TcVsfQ8ivfBWZW7+fXalFEEw6sSk9O7rcZKJm/
xY8RSEOY9CpIT2tznu0YhK4+0NfTT68DSUTLDAINg+0XyRuCtMhAT3JtgU4GHPf6WTzS9UKEGsNd
55watSsIaFe4QZIRnpEtufFSBpiELaNzeD+5V8T8Q3RedQPFYkqMyCiOQm34Ijr7ovOQpLD+gCOG
TxFFL5LTfGN+awy7kzuqmzbrJR93L9KunclmtqqlUTU8tyv1lmRsZQjYWX4cUCY28KGv2gJgC/Fe
xpUwuCJTjUuqbYIV/ZnfEkkZqP9E8XtuUVlx6N0ZvSRAUZVp6i0ODAfcOJ0iCC61aNJ8ZOgsKnQp
mENTj5E+E0JUK+YuPp3Oyn0Rj6kXXxJzlKn36iCdrPg33EwZ7GwGjADxOFngest+sdZgbsyn+/XC
5Q2I9+hmAzHVhK7puGU/nENdKPvIF/vO97KK7hOaK9xheI3vLTf7NOtLey5dTV2JveERpp7t/whM
lK7LIyf+NQ3Aw+rPpDudOm6VB1SEB7aJw+wTCVbGbN1vBXElhJr5gvJxgrFwsUzzcGaesZ3KHt7j
+DWKB6PVimMEx8PlKW2wOs9bxgGJ6jxAnkUDT3jMuCKRaIqOM2GfC+J3WETG7FaqrmyKdxLRVfsA
hkfBaGPZXgO0fEcZL/6E0puOQTKqa+0Cj45vog/ey8I/b2oMW/5xMllBIHjBy17vY+UW3hMjNjeo
EndJsf9NqO+ghsdr8GbsoQb84Hfl3AEe5vHsvZL+2OinTcebkbOM+W4S75eXeaPqFQ0waymf67r6
zX5wRBA8h2EQe8/qpp/izDC4Ph6O3zifnvSn+QqcE2wEmrba5yJHBeLVbQDhdAilcPeCXGt+D9WZ
WH4TVBAgVb5XJpRBBuW7YGgXvVcfddTYmvZnfd+qDSF6Mlv2Qb6LLNbJVXeRtubSanChUX67QgLG
0+g1J2yAtMwt8x8jIesd+/8KbZjE7Ct36MtD6mjAm/2OLj6l6C4OQXa8v1D//8kVn+oL2cFBXt+H
fGl5K8+Ud397YSk38EFL3J/ELJhodD/f7PNUFQqk/GU00B3wOlghSRTpWKTdFjoHFM3l7krUmFyk
yJVZ3RjTUfRiaLrf9CuVgWMPmrjBb+K+7Ep80v1Iw4WnPpbAD+sRn5uGNTyp4Pe2tL+94BvTisYw
luuYijiMluz8whxah99muuO39zRqDC2ZIhMG2z4QTCuEXPB4lAsYCgNH5Y395+xOBMfija2OGs5g
dMtJ0TRmRv9vA28k3T2pOMKQzJDoNarwB4ClSu37ZZeNiTR2LS7ZQCg8/BCQy9vkZE/9FQTIq70c
Y4jIQDZLzTnE9dKGbHoCkvBo/vJXenAWxDlzwor3rOTV1cqC6pWRmAegdBEhFcqm89i2spXoQXiN
xPkUcAUOV+ObV6mGOCCqMa/oPNIQ4f+YjBGb7KZKBPGm5d4sUZqF0rVwZJZuEeQ209tS5FKFz5zU
KrcQWY8WoQKyRuIc3yjhg7ejO77aYaNjGRNK8hLBgtGv1qCdov/iRJDoM4L1jmdIkoi4cJ958C1i
3NrEo6iqJ3G67+fSJKbpuqnL4MivHJla0TWoQhVCuevAT4EglZ0R72ism2o0K8ok12iKGcRqlvYc
S3bSyCXRJQBkgmYpfjSn5ZGCqAPJVDDeAA0zLhtv48ao+Rc49RYHl+RtJj04JhglrUzBb351i1GA
r13XBKLTSek46bKutp70dUMdNXpMuOHUFM3ZfuEDlLqA5LCL6wn7JY3AXc90aruLOV5XAr376gNf
zZyYdKxFbhtz0fNkRsVittYzQNWAALDbxXv1kJqNLEiEkXD+qgNG3FBy31cJFTCyLGyeVfnLlIOm
rw0h/xZmRx/oxa61HQoGR/Nt2dO8b/bAP11U0/z+CfpNupA5DP37mNitR83ntRvAj8JfwxyVLzlu
rZL7tHCcDz9V+epDXMyByLL1HtGeL0j4IVRBrp+a0MH78y/JITOkxnB4/yYH/ZK9BzHII49pFkyi
fWph9uZTX5u0eqdalmyJOzepUmkXL/QyuMa0R7Ze8mHxfAUOr13THj6BCZW+l82oWU/QVPDmdjtG
4t+s3vFkxn18IazV1i3Cm3eJumExsK+xnbhsoy5fPUZx0siSFYFc28d3alDKoFFL+RjY7x7UbBQc
5Jbg266xNzLsZPTczNbHxMdr4S271eTRaBID41DwxjXptbGrE/t9/S9xVtdU+gv+nQ1ETmiqZVEb
bptXSbOwCxUWDdhDaHel+QDBwKcTWeC+oj6YQgW5QTxIqxWd0FbxDussK6jJQOtWHnkmuf9nu3z1
3aVfcZ9B9wkxaEXside8kdz/PGHVSd1RSihyLeRhz2nW9+++jDXXG6jw2+snDnVWfFVldLGzVN38
e5aHxMmRn+AYyaR+4TndnxP7jXyaXWLDZcxMICdHJUbDYAivSi/D78rn5/sUzEtqhb+3kTr9WNWI
o4jPEHjLaFxUaBR0AqzMuRqkirjqT9CATGCtS/TfTAyJq2d52I/TV9DQqMd33R+sSSGIc9fdzu3Q
eA1Gd1BIPfOC+zB9dp+mbJiDN5GvLa3RgKEmS8IrbZX4aMBdqdK7riRMIFVjfqq6rBVSnBh+JS2Z
T/QPT+NpTpJq1Ao8HhYl9aa/YX25GArBoJXVgVnV84mBYGf054CQFP7BIe8wBo7+mlXYc3JlMvFv
5nGNInT8P8nf3p+uFypbmWYzSHmYG9I0GcJW/vTDZpVVzHu4Q7FIlgyk6gsa+R4gyL/5zcshkUtr
5o9rSgWVYJsPOxD7xvHpamQEEl6VN+Dh2747WMMM/UgmXj6fr5dx+NBwTFnisUGAyunFHCsWX0sZ
EP3Z8+XZH1jrxcRl4GGBmqPVTiz69ewnG8ywIh5wv2+6imFVQtO+KifqE4SiEqis4ZrYCOSvo0Us
fgOhAeDi43nNmRXOey06Azm2Xqhgz7bMklpNHdBOt+JOOql2P0mOqTbGTlZPrSBvzFnOEWPKbyTE
X1yq7jik5EhvDsPWm3PdTzKkxHMpwF5iz4/q4ptuOZeFIst1PR+VzqgEjvhV9sVpVtWJo8JIDwjQ
h9G1yFrv7xtXToOUzTdSTj7DDUYw+vEGCptIICsDd2t88IBRCuEwbziVvXIiu94uOumQ/0ivZ9eJ
rhLsNbQVXVEeARVJfTZbAN/mQRxG1s7bJZfsQE2dHoBFIQK5g8gBAIwxHNOPdunzt6ARkwwKtibh
73mrugjqBlVCaV0kJX2daLjsSQaI/Gf6p4QYiL7pwtfYh1YlgleI0VmashdSRGPRcfS04zrFjDma
yvYseI1RhatBhKs4qFROLCXyOtmHiOQAuhmD+qktOXVw8Ti5B8s1hOx2C3sOngZRORUJtK6wpJhz
Fv8/qGZM7WgdPXrNVtOnizhMerFF9vbsHgP4ATY35Fs5LLgfuPctP3ImCZR0JryX8EqWaVcl/Mom
W4LTyiHv+HMbNtxJ9xq9Xiy+ZNGGiCGICTzQLSfDYd9XrHUSiKjBUXa04bCBjT3CR/TJCymtZH0S
bJrPCFJ+wU2c126DZeOFu3RAzgxJx5uc1UV2R4HkU/2lT7dECgAbNu6zR4ICNJX2FKYZIuU0H8Z6
KNHoIaQGkTaevAY7m7tClLsXFH4A42houkUPsLjjN6uVdn+eJWvpJbkRi5tq/hnVXWxnr/0hshG2
zWtNgcnShFO5Sp2udENhzBM+7ovPop00LfgVIQSwUgZ6I+90JMkIIYdHobV5m0+AESHxb/aLwuUM
5bQgV5CK74xppgQXP51M5mNtymudHYWQzsmea8mvRpj0Uwm2kmutEyyo3wXHEg+wC3tLJRA/sx/r
sKBVUxDSsz1jfS/DAoObt5Sou/cYm6xWDI7tmhRwSPnXCyDYhJfQvzwNga2phGL4Cn00ERncL/HD
+KMj9FdtN0QTOU7vttpsh5+9UxjqarI8lTwn1ZAksIsnysZxlRh2gD9uJEYsJ9G7Wdp0seWq6yA8
7P6hrDk8UrzC+TC0qqAdIaQWgCcTamIshwY28/OlR/P3hv3Mkc/kX7HecfCNWAgkITotLousWerg
lPUzG6wM/6MVg0swbv/pWTY1KFaCT+QrJiJAfoAC2jG4fap2N3I3tzJswVRlu5gnb1FQyd7ctHeq
V3WMzuHroGzYm1uO2GVegLyQnOaDT8BmpWinPw1FEH8zcQrYK7pgpyzGWDatWeUVd2saJNkkPFM2
w3F/pVcU0r0vGp2hD/tOCFgo7+DKYJnBYlMn2mpzMPlWgVkY+0rd9UFV5wRCGY+QIZS6V3NXziy6
Gf/QoF/So2QZOGE9ng0/wzgOOkryNSmAa01fl1N0YLwmbdHtlvcoMP0rZ5YaCbrpv8WU5ip7R/gg
qlEHfD5Gr+yHNuzdfugLByUav+HiS8Dkg9QcXJQX47UasOsVyuyRO51yZuTuR82zsSo42bltS6ip
2a+U1HN84Yg5gAI2ArXKEOM+7ADEIm2Y4vZULLK8T7vde18bBL6AANEMjRxOgIb/4WcmcQGIQIVz
gWO1bob1e5e68cqHQfrFauo5crBhdZ3jb1aLt0g4QtXLfIVYfmK+U8IvQ/Cd3zEpLhNFpMHvOkrX
3zF8wOxDk1c9NWa273evihNeQk2bAZMWDApuUMjh5bHiJjSQ4NUXUmCBT3N06UxJXtbx1nqSTWpS
gVaoYrQlta96mOftuAGoptoVpx3U6OMFCh0YQFSste7jSNtN1ab1IwvEhaFH8cqtBmd+vPe+CWBW
TMppzyKffwqAj+4H76uq+kXygovBwlmvMAV+9+ALKrV9S93NJ2dSgV5+9YsDcs6GbZYLyNs2F7Pr
N7SFK7llCVAUQsGVCgv1EVp160uqcgdpHtAK38+lHmLAW4YOzJk9nj5ADTPnFQnPw08lnWfBXvDc
laBhN/FKo1RW8+L8aSIgvMXGffSiDchm8/pUoov/VaVPCCEQ0rHxCSG71VtkquFYKdROn7QZcjE0
3X33SS6qcW49/l3/W3l+uMz8ZfxaNCEkG+QvfKst4NOFliWUq0AZU4LaopfuJL1vhwe7ayTKn7++
KKuYS9uyTLdhVtWV0KyxF9oaxfCowYHupBHtXVWMis4W91DvYwlwtHE7BubFTZKrPqyBgj3GXm1j
SHGF6Fh2lDf8Uisj44bJOwTQP3InoMh4u440iCMt7SzHnQL6jOEhKgOhoaMbN81gxjEZMnOm/bQs
YqY3dMpicNXqTFAGVwQd1vvapX53K4UaF0QlLjDHVUCYCPxU6Zl2O2mfO48OBjYtnRznWFIrFoWd
piGa8+5zmTnjvxrk+lGnD1swW818QQaBOW0v3iOTx4R+g6comHNj/rVX1uE1XbmnQuSs10XMD6Hs
Rsh9+DWvBNkMXg6699NNSZ/lldbx4HVtkllAfMuFu3bgnL5b6Bz2UcNJvNqLynM1gxNG/8kHGKkz
th5gM3WNsQWpfaPMVbXrH89IrNpADkI6kItCHLGWQyZRKY0sUBJyioyrdXVPbQ1abE1Q3AbsvhDQ
piI22qkQ60v1Mt5CIOecnQrMmiEXwiryLhV1TAWId4UoxrgSLXxp8yRJQ4GHCkVu1DOioonheOEZ
5tJF0BIFzj1GwXU0tJVeJ1InXTU+iHAie7tCI0FDNqa5yW9ss3mNuFU8/b2GEz3ybd2RvVdqtDIf
yniVWCrb2QyNih6XOo8WW9DqxD+ywcBvyRnxQVlA2z7w0SyecaI0l7F8Rp9z7yKctDxWTdyWEqcj
qpXFoPKo4we7zS3FEMmZP7DAU/BeqJQ8tZxfgBFZ7kMR5escMLVutE9o9rUmyUNAzdoA/ePV8YDh
IyynJCXpkLDNOoalNivgUFRS2z4hTjmLWBD7P4l+taD3B9M+dPR2X+HOkO91vYwM9f1TBht41Hcj
8xWx8MT25oR54fsLr4zZAz+t2x/9keYwxysJtHmP7GxBKTFg2PCf6FHq8vhOWehMJCZdg/uEfj81
vrtws4H0cCDazA5Tz9WqCK7ArqMowSkLGmyPUbqIP/uuEgMZ8xvz1OeQ56RX0o3Ir7nwUBk5/Z9N
keb7WUWiR5M9qI04+W5XsPYnVQJ6FJMEdgh+TG1cZD/KIdDhE+h5l8N+HRWl4lD18O3ktdMJO8b1
QUGD2NZGC1ZwOPJq0dxqvJIIwuSz6uLJbFiw0Rj4FQ6+ferKWK6/Uvvf7tH24sb/zYWoiVgseeY3
Z+QETGjHcc17DF1V//Qd72kBGelz4VSRGsu06zgUJdmS4eYi/LoFmMmbYehsJkZbPfeFHQu5mycm
znPKctT5B13jKm4KmTVYsYglcSEHCMGsI/n4cCWRk0ANkIrQ2i8XD8yneEYuDEVyJXqfUM9uBHss
o2PGBLc1h98q2KYTB5sd2caaF6J9nd5Dx5IlYR2wNWybfkBbKcArk3prLVuQjf2UyR+f918tcn4p
2vIaV0BrD+yH/6CPwJeLLgd1BJD6C3hdZ2eRhY2mg2fiEU4kCGMLs5c/qWVjOYZn7NOzU9L0qjGS
qDhG0uIMvLegIjGuA5kBPYzlCK50EmBMkCc8cPfw70dHG5zBgcNYvm50SNL9HsSMZ2S4dlAw81P+
FQEcZPg05vAJaeu+svUWEcPpn6xYlYWZCM79Clyp/XuuyVqFVe2Gg12/9MVAXoNc219CCjJrRTWI
Ct0YAji6XCoDsaWfQWAono+P8F20F2AM+HiZz1vHHgp5K1iQqDHq6p9PTua997gVUeQuMGP8+N1n
fAaeLCstilBL/G1wKL6Ay5/SOcO4E9F/tuP2mpjWPgr17pWOKSMY0iVcwc6hB99OJEuMWmP3Q+W4
Kh3oT1R5SKE+JwviDj5m8FGsivyYnEBih3s2yYmRKqv8SLPPIu63PbvxrhKYabEZ5zhl8YNTioQ2
jEG5uKqFqSua+Cim6qnJwhY83zeh9fcnie4I9ggKRUMGSqI60UCo/TTFhkRPW2otNmcFlQNARlNl
wtImTXp8ho9z9/1jp30q7MvDX02WcYQSpeNmOkFxctq1Jw26xmhmOS9NGEa3DiUxjkRyZuJ8m8XC
k8qZ/gu+pNzZt7hjJ/2V7+S8Kh7OuMdK6C7N7ClWYmN0k7GTL4W30MxGGhmqg96EU4Oiwc4Z8Mf4
CfK3h6Dyyl6cthuYZUf0nC8FM0YtJy7napqJOpV7IQnkIjwUv9gj6j0rIhqRXV5IHBY7OoVYL2qr
He7ua84rUuHpi0vI40q0w84FSUbGFHkk0jAuiSef0nkHpUf47wQWd/k2xd9BdeQDParAIV4j2I3D
HSIEmmV0zjQgDODGR/SSDr9SFFGV3IzvVGcvh/ybkJKfhnXLJa15b7zHTlQJZ/tNyv5NIE5BOyUl
QpyfNBl11Yecpt92ztvTSSuiio1Q+8xvFQz3MmYOa7s5tsHSy+lZFVbJoZedfpiaAQl4dnM/YbcQ
+FElWDbHGX0LbHVsiT37Ab5t6mryiMC+sS035KKudFsVlyS3SWFEl9jEvFgYyrPgTetYU4DPRijA
DTBVya3qbXvRgio1WHau+I0ClFc021atJGnrjBuQZk3wuNvixDJ5yQo7oA45DtXV/fhzVt2o0veb
805wn14y8wQC/QkcEUgp8gWAu6TpDB3I3+CeINUyHBc608TY/3F2omPF4BI7a9JXWfM/WfrB7z+8
TnNywdy+pCudG79YA+3iajL3kuY0TyjRiejq1I1JZQ4oIPkwZG9UWLJFApuHsbzL/KndOd+tm2/f
GBmycPEPOu5Po9OzoEppsH6TR/0bQD6aFW0nM6iqJRfuQmlG4vv4PFSeq+gmLXmWJo7zHSMa5nhq
EegaA3wr2JzLegGxUtBm0LafYP5wEGn54jdOAPrObBbIUlR2qYlotClir/hKHQwC0l8bib+5x7WI
ALA3+MOnXYE0IA+xlYWlhG648UEYi4b2QsASxolBm7zaLwBBYJhZYbOxgta7hlsfnpRPhbqKenR6
I/H1K9jUjbiLjPNcCOgoqduqwxCLk2DCNlMB5E8T8mt7wi/c0GAiEtTgI6XIOcPPvALfk1pFt2Ui
Rd+pFh+vKwFYIZBdHzu2s47ssAQqgg/hFyGuZ42ygJt5upw3pa7D7vzkuZZGp7kQTfzer2I5LdWt
UQ5xfblA977j0mvhd4oxy+EG6nGO2rykHu4ksBzCIsG2y7VuPc0d06Pm4QFibbK/3+gzdbjHhIiv
stPtWpeU/K4EZLjLmFN0QdqoS1GJJBeK2LyMImWPkyCUySQl344jLoYBO77kAZi8SWUCccngcXs5
yQbN0X8mk8EyQHcfxhbM3g12Dp4hmwefrSemc7r0UhxM1A72Dfrrlb0AYkcwZpZeIAx1bS3O6vFJ
hmPftTc3RoZSWGIDp2dTEpA4Uqg5HBZIJA8x5jJnuBwLZyX+G0/Bq+M+pBCw20Kifn4DACDvh666
yYXH7MGRcPkYh3OS1bqqmeHdKqHYVOStiq5AqhxnYAwJJ1RW6S+RdGGRSp/k1vqNIBL9tkj8IAsG
1WOOafLLS2IjGSoJwA8D8CFGYpE98D6sLaf2BHn1aE9QZbtRCdmLktxlK3cV0uj/ayoNdY410D8W
bqDVKUq2gTDQXVX2IETnlue6XGiGt0Wjq2TT0FPNDV9wffNKPajA9//Oyd1B8+okozXtmE22HPfC
ZaMNI/8UfHjKyEkpa+ydQP3oYmjNzoma8UpG+XyR1V4oYtmasuirZ2uIo9wYlgOe9Ez4jCZqcTsx
vXwJQWyzqyBsoRx0uAaK7PZop8oWiRjYxiUYZ7E2PnSSxu5sQWK/7RuZKmKTAAbRoCkX/gPNjolI
vExcgrPH2/orj6Nqx8q5CHCgO4X0OrQF+u1o8GTdL93nIp/YD7WZY/FnRm4+v6a+jBflHcCEOqUB
63pQgwarUqmWVl+c1LFtrZFt2OOwosU5liymW9RtrxO2jdj9mgN9HJG4tTghkqakCZFNDD9LjZPA
OZeNYoW3IX8aBdYHbfPDQziKXHf48Njuhf1FfXYPVnoaBXMwU4YVp3nhL6u9fqDzk9CfhzpFXs1A
bzHx0/Wq4AzzbHxcHhJHj1hWMulzRvTkErQO9pGP1CUX/262j8KWqvBTM2UgEdMhfXmFH1Dn9LLR
N7wXfjsjiYJgvXPMtqMMfGz0QIjZEqVMewBzI92XocAwoUBOEeOLXHy7wPONZyxm5ep1AXtUj2yi
k212w0OyAEPNZcgV/KVaXodGmTFDj1ErnYZl2hahIvihgIyyvL6orq3m3kKLSScYSLZ1S2CkmkDr
yhF1KOvPx8Z8dbQQpd3/WQxbGUvnt7a1aYphWQ7f6AVJSW9Ie0LAZdAxoo8UuiQE5qIorpIGUh87
frSoC+PO5a68zqDaPs9xMWSO97+2rjC7xUMAzAGHEE17KOZrwMlTuXvVOAfld8Gu01otW6s5KFqM
ycCxuWWRr24wfcWJdBdL7w==
`protect end_protected
