`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
PEWLNJITZPcfEa++ZxC2ipRisjsA9rhcFiMtL6FBLJv0R3mo/cipA2ZzvD7MLJdp5JHedwF1+j/L
3bi42sMuug==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LgRAWuxTDdhry9Ll1pWVqAfpA5bYCm1qOfGDj6Zx+L4GR48fvJglZKlK3GE5lGoCINSeeKqLqB3I
MpwCZwRkVWGxmuI+awGBq/Z2rv4R85zedQ4jJL4EgxMU90qO0Cq8BJOECLU2uNUBcx5ybITL54fC
3S+K+nHJsZi7iFMHKjY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Rk2B8RDUI1TU0nAVvt66Mr2HYOd0rlwk/Vx3reWZY46LUzdEMbXhGH4AVmp4/miG0LM9Uv8es2mg
ee8aDjlrvnCgi3UmyE7Lo7m0iK96IvXO0YWKnSbf+LLh1fuxBAgdMkLAtFJKPg9lpwPBA8qC3h5H
VUYxXbVTVEMLTylRbvTfs9tedHbiMd4VKHThWtzbVJQxzpv0IgIVCcyXJnisDvj3cbEtYFo6tcZe
axQf/ap6zgDxFL4Lq2E9ouATJp1chQ7MiUTBFO0VUgSz5AQ3Hg59cmlsFY6ch1+3RrBDQlmheTk9
VKP9fUO7Us5NMqveQbQisrVYlKyoszSRTTK3+w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LMacKgckOoNETGGDSERi6hT2Bd0/m4jDMMXSpaowfKKqN8ddSbB9tw2wOCZiLSCZut0gZ2QuMN01
/CqcSwj7yGe1JOfIwjfbpFYzjKF01MD9iEwJvDrPE5ZZyh/5ell2V7py6JsQPsnXlPtHh9e2GSkb
MQmbCvtoI4LaN3TNmaI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iGO5NEdM1XyFAEt0ahmqwhKfjgAe43ZMhkzztVUXAfqF3ncnVQUaUX97dNwp8nt4Roq4chfi3fy/
6ZEBwtJjp8VipBaFeof+5kVPNGzEik9DUoqKOWJiD2ucwCQ2Zkzk7qSlckBJ861IHx8CbtBQxYTH
A30Fzi6pO2IiBV7Z71ZzQ5kyz7qCMB2QCGrVXcFcAhI6E/l6v6rJ7hi2Oz8oUjG8ANg5BHNIJDdg
SH+Dd/GEqB0IVGMFmBrn/P7huVm36AWGc0blR9Uh3EXcM5JqBJR2HlODdlMvgI4c9ClW1e5lrxGX
6/Z8HMP/LETgq+hVCLmDhzlIzYMofTlmVFtcgA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13728)
`protect data_block
ALRc32r8UPoIZzp+ouww6mmZ7BTLkJ/hj/466PR/QIGl9qGWb2oK/YqHGhZ3ixGOFMkkKmP1KzQm
1MsMUcEulVLUPcwFqRG6mwdvtBJT0utHz/itINF1QVfUCGRAfpPqguXmAk5hJUe7xxRJsbjYciwR
Skvfh/RjCRbgrKRFo9Ngbd5lztou+QLMgpxftVHgv72okKATEof/Sn1Ax30reRU0OifU2OEdiD7W
ZFVp1UV+mZddFs/c6CM4las2l7SL6Jfffh3yNuApzG7sUSHdrTD7D3Wih1nvc/jEXNrlgDSd0jHz
lGa3WVBLX82gyE+rdhlvGilX6QLQvXAWgzO8YOKySSoATmBkTeyLKieZ2TndEhsRBAmTta5M700G
qqks9kiuW5cbZhetnOE2mGpWYdS/nRc7FNkxLwCsUzUpBeL9XcRhsj2MDENbTUp83857uK6Y++TU
/Cui7LFYdBoV88Va9kw7vr5xwr5ekzLWUC7H9vNS4sorbyx9CpnMOG0Iuxlu1vo/xp7UoXyrUDLm
z3AvbBoRHC2Up8lcAYR2A0Mr7lg2M+Y2wyaSBK81VzaRNJd9KFmzWzrZySh9VFMwSpnHY5cJ8Sfk
L5LXUPMVjP07nQ6u67jDM2ihll0cyCgqip5vJZQGh/X0+hKC2pCqT7qe3Dnic7t0wKyscu0763tr
CZKoZj4xnquQ7rMDM4urWzr36jOZgnw3UTdeQd/hYax14MVvN+t7lyL4Q4FewsQPT3z1zkoNDXG0
26zDHFzbW7xolftyrXQ8WCqkLsAP5ONQzQRhEVS/BkBKzxSExOWOyBCt3i10KMHDQVbuxghUFm/w
TjSNVgBtecJJhYKYtrG+EKE+rQDWplcWMzGjdEDkgHcQ2+0hNAJumLWUaajMBCMuxbt1AMfQoW/H
KcoPLAJmbxLwr2ZHb6ySoXZ9ak35vbHAErRmGq5y7NIIkZeYubiLARi+4OpV2NvUexjH0BJ6/xf5
AXKGHnrrsR+lB/5/ws+NNB/OoDde6/oWf2pmmt8DugzbJRiP9G4Gk/Qauo08dJl4bcpIr/Wce0Bm
Ipvc82uO42d0w3OT1FE04Y468MzQafYcE/U7VXu4xdKudD5a9u791a802qS7A0bP78rOKOu9FDHa
ptP6anlVKFnacF3byMh7jn4YUryQCAtAqQ2UaQtt5lMOOplNklyj9eCN4w13qsRyDaYwy1coIiQH
Rk+VIlmtdzNHz2hIykmdK5c2/WrKgJlAD9esSLABFqeEea/3Vh4k31aoET7xDQhu5AYNeEP9Qvo8
kld+jYGOujyuKIVtGrUEHcgm14GF+3c4Uz6hv3JrE+ZOi/K2SBBkhYLYYpfKl8oiioumOQ0lKs8F
nsncj62LurQzRHX7RwXk4sPkzJT9g4eGNWGe9relq8BlmRkdPTymco5EsrJJdN6SPY0sUasLCE7K
IF9hoxsWxuuS0iEIRsf9V1x4metTt1DZ6efn1UMKm28VWpSWaP1kHFgfBkAIXqL3C0/3OK+TCCO7
kfiQSMEolsNXaah364GkTFlSxjxEEncKe+uZXakqAnGORcQmHnmBH83O1TdwfZ2na6KyVhj34gH1
kiP9WriNe7audJ35FvlGzn56zkoW8U3is4UnBaZ5Fq1vNrvOihXOmnpLLpqZzmeHuhSg6P4XClox
xp2tDp/tRD+t7betQuwDbdkbMIqNaN0hhw63w/f+wwju10K6+cbrRSy9+yH4gLhMszuvQ1u76LVy
Vghels91yjKqLt9penNM9madP+8V0BfmYNS4/T3GDlYao+6FRUjIqKqNsAgDXochuHqizgPmWCmo
0D7FUHsDYN9sNCVAX+dPiEySjxslOXwCBpEAVvTi3EBdrnzaVgToZu+fjcc0JTSwNuvANvIXN0sW
+mT6xxJ5dVlAOQFaHnm34/yVz6LEx0gA+/rQhg3/GRjKYh0QWR/4ODlae2RI6W9UcunXVwh7IMRk
1UCc/m45SIthRDfZ8JP9uiBTRE6HL3l9J0mtSoJ4qV7Z4ynFYEov4tOSX+staA3dQuna8sHP3vYj
CkVhtM8KbadnjKHc0zp5wqvYAlAm6+VY3gb+74T6bROX4EQM6ejmfKIuNIlBHiqaTSH5L0WE+Yma
FVsL5gQfR86PZ4gXL7ybwcth8d9Y4NoCK5bXYRI2BxRjYTmuQWmEXdtmGdXNXGg+g76FXvsrkqxj
7/QYWWvSjaa/Mhxko71S4CuV1PjGH4W/JRgj6NSr0+vz3A1sYTRGBDpsVV/qg6/bwV2CYvFJ/ZOw
c/0LhQ92RAZkimKBYUOx7sPbtqbVzv97kN0AhZ6FgzmjddnRTBmbMU0zOcIdwF+JQj0k0ohFNBWr
X8B2D9ngclxwGFpJT6lJWo0VtPWAp36l9/YqCvYuQqvXzYIx0QXru0nHIjM5enS/7zEGKNNHyWV5
5ph5ZP7fBMaey9850n2kVORC6IDZlUW5edHGSJ71C6eApNIvjaTKBir2KkAgJhLJ8gvF+vZyJSGs
h5d4z0nkDljVcoIqjl4rrA5bOlr7zDiaPfE/gutMj+KsmTc/nDEPmY6ce3m/I5L6g+GwuEJldrl0
NYInvDqrGxXLa+CC8f/AViS2oxMbXEbObr9L6CAHtnB2gd1YMz5itFXX5nDxasVnoV+nhZeMcDic
ixm+XHXb+7JG3+aSJbFRx4oFV50ZBKfvWDI0yZDFx9Xw+GQ0S5U2ciFXtIUvHB+crew8XWmKorBf
qntOir9Xa8dWwe86H2sKpqzvsiYPeRoOwObiQWgcXnFV77UvWAMuXL7yKdAJ8t6GL9+Cnu/sUiuW
uO+WynFQaSrHoru08kpyunv+NTcqloe4LBRc4ntMgHpCKOr+3FzTyiWm0XwwH4hZubAlmtGKvd1+
0UZzPl3/cFVT0ZNY+faWxDptY1Iox6qHbixjuOGRx9VxP6SBFkd3hlHZp8gTtj7oKvJsO0jFc8Ce
umr4+9LvKKe3Ip1PUcPHu/6bLnWtI2uHRNnCI6d8FK/NDTrWl/KjhJJcx8DO2EPrkTgj3/u/Trsf
12H3Lf6NQYHTf1KhSkkgFlkUgYWETZMy9sOfXsgSg2ZdzOKNgHyBPrD+7BJK++SITtwqACE8yds1
95QOt2ZYo9hYyW8Iu1KEgsOEDBHGrvxs23qkVbMHoqEZGO2G8dmA34ZpIERtQfSj0sz7w5smqWMc
/ACnekmDIoHpGrsCMjpQxFbboTskvHZGs7kAaTrarDBssCdTwwE90PPCu38n45HVoZbB3N2vQvq5
Bkc5YoqUME/+1kX+881g4YrUZZHmgDWsXppU9D26IS2FSM3ZXFBfCqSUUSHgkkQvJUwgAp+i84Di
OtWL+2ASCau+MttlQeKgcC97Qr7/P6lhdTd5Op+mNeU4xU5ZeztBSPSznysNp8K1UUT2EPACLCMu
rp/7P/nwd0lZ6mntuvC4CoZruTyqCQRhTRsGqEL8HGE2JFArnlKK0VQ1fTSxJubX0oCFFmA/xKaU
Lh2TxiSzoXoL4GaBu8WwdmlZLwDh6rHK0izF69V/R7p39dqguFmW6HtkfTPg9XlLXa6jmYw+q/Za
bLQoE0JsLub3E7I37dbZWqEFQ3ZiIiVWykJGeTq1QIWeAiArJ1eiW1HYTWzMg0WqXUSIX/+Ewq5H
H+ER3phMZkGggil3LtVgkloXEAyCs71xfC4iRKCW1lMAnjyFk5rH5U03Rw0l7XhsjVXl5VaVlJiN
dwhFg21HetPMQQijYhu2rhYMF0P/f+Cwlncn4/rGvyqcnMMS+gXepEC0xR8L0tXoHooeSL2Z1hNv
7RITxSOr7EADpiLUEiukVooSS/Tys5jo1OJRVSnvv8RKM8Pq9Wr7eRvnUbPvAT3RtWbAGlDgL7Rq
ztapUVpfsAkxzGFWrzE2AhYEIk56nL2Bvi7535SndXHRwwILwprJJY/sKk/Qs53Z224bS5O1DOYj
lPtP8jrMJe0alsVYXhR3oCs2mGpl3YNe3ItWOEBwlzmHYY5U7e1ENlbuDOn7s5j6nVQXrAt2TIOL
GZvlZQ032fAn++3sLP6ZALmzq3ekLlxbRJCvSlwv1XePpClmcKjmoHsxuGCtgmmAUcgs7/MBwIUj
uTLZbNdsiWI7Lky4D1TlCroLJAiCM9heS5piL+csugfCi1lkkYyvr3xbxDq8anwsvKl0eHlXyiLT
0+55d4vUOAExUX6L9+QpAYFF4/EBIgyYMBao17Beviiw+Ay7uxVx9hpewgwTbXoSz5RZJSCyrUwK
iLRxuULME5D+Rn13q+5RuDUoewL/m3/LAunkRhNltfyBxBYSpJruY6ayUVxiXnq9Ey33UwExE8ED
pZpDWrsWT5Zh92FOLL0/e4qIT5Fz7varFEmeiO7Llpp6D90Hq+XAISvSQ6PbM3S4Klxigzrf1z29
RHrZJHNY5Ky3k+HjxKOv3POQxymgDJYuLQHfXSDGn4GiYFkBjjGMv56JT2MR2XWXnumCFYvOtllm
zsTcZjAK5JoOxV9gZpkdxWrmzOtwBUu2f46jDjBmHOxQ8mnap8TgmxtRHfUbHYWon70YOHn+AH3u
LVzTj9sTObG7TLwnz6kjOOoSR/WO0tIRRamu1NhuvSpjz1Vyo71YvekS0UQprXVz9SZdxO2YepZt
hhyznyKpyEEUEYGT0ZsQlVPOy4oVJEW5jxiycmffmIki0I+FfMjsoALU90SbG1gMIu54phaJi7nN
Y8wPuGity/p5ztXh/T2nmCay+diNkSzj7bWJg+PIX1b6uhQCMCdFoTGwdPbVm013Zqt17gTjuZuR
oLWq3uZkRGGOcFG9pyV7YLyEmacdr7Is2F4xKkFMz/fdxqgqALyhct3eMqgBi6w2wKaA/wbnILJG
L/yhHV7hFlala/4w2lKCmihpRW4XhEIIf57Q2Pzq3LH1bbvMkKRd47dowMLiKJzftqALlU+s6wL2
OLZnUCbtql3uWhgfbRbK0XPhtzR8qnzhZdz4kJNPYB5j/wRfk99JR2hUozhMqDLnQz4fv4jj4m//
27Wn+IXYYkmilNYPIoZRpkGP1pr6tDdvZrr39INydTvZ0AuyiYIe9vtymc+jice1h9IHLfUiABeg
gH83W1pAJgY3gLfn0UVaAACoqWbwlRc6a522KotAN41157Yqh3DrrxJZocRd40PnrQhJff2//NGX
s3aJ7zPSfOAL4h8Z4buosPkK76+fjEq9+lZgTf4864uIMe4stcoTou7/wYoQe/nCvDmxGTSWnhA6
62DDPm9PHbuxUbEJjlM4HIp2XqiGNsK4X3u2pEeKXau6o5iZU0z5Mi3yqL5liAvyPNogFw7MfYks
osHn5em2KfOTIkEaw6PLeLwWZqjjiDvEwjXEDL417NUhsmvuigCCNM2BgJ5fbtgttabY23ry/KDW
aW8QQjmr7SCXSTXHZp8ORo87XHT8gynVGtw47xKDGpTmMbrhQITNDdEloZwCU7QdOZVsE7FrdMAw
Sn9eGumebxfJl8KfY4Z3sq3SJ0rjI0s6vih+hPP4PEZmK8auK/rlVgOODieb4tnhuILkP/kQbIfh
Iut+1DRQV5lTLbmhLLW7+JP7JnJC79nak1M2k5tQ4B2UFWiA7wGHI3Pspc7iVSKzZtiA/7ZOoQzR
53RpXi9B7wkS/pNKIK4T6A4fs2ZUj+MjSDZ1l3RDHdZeQ81XaqMUPFqDgd8dyYaIJwMx6LFOaR5h
/RGyMNzEcn9QQqINZHmjom8ZqUX6/lOlY+4gBRb5ZPCk5cj8tRGen0sxAbVzToiG9VHUIl16QFdV
4QIvt3ebCLy1lYTOP1rr0DnRMgSituWfsqycZzJO96zHRyZ7zfBZv2rAUnLkhCaPjBERqXodLCzR
fI/VlgeDWfIgt45kbihQbyluU2vKLZ5hHkNra6NZ20Gd8ltiDEbE0kh3iG//b15cDjI2rDZXvGuh
G1PL6GW5wWu6MiZwnkS329Ug1CFHm4flh8wYzOv6T37b2/zroJHJVAjNuOtALPu+1I1hdDm0xQys
rxZZAeufcUpYAiYt3gB8VYz13NBWVbiMgDHSp5bCzQNeZ7d2FctUBNYzh+kiN1V8IUeHqcI/M5b9
hTH97gvCnn4el8IJMaeMyzaveDAenQduYQe7rmTbiENoHzCdsOegYYBturm1lUj72CPH+IZvYQ2l
i6xaW95gj4+oKpwlCJ4+L0ML7bCdM9ru7CLuJcFkNRVKSrIUJKWi75YwaMv55MAt0/iUDQje+89b
yjXNbo/5Pf3CENtKO3N+LLxSw9wAnikxc07cyRoLvg9URRBhr6SUJtrt0vHEDthFZzNSKhM/GZ4N
qCVocSf/6cIXzKFQiQSikHvzZPIK9aG9aJ1x/8LjPZ/L92/LjDzqlaZtpw0GmUrrr+7djZhmr/Dm
8dHrWmiFaFpWwZ9Vr5mz9cklhraY6wMvpI1RpezYNmdhpR3KLteRFlldosHe3d9WdksNAKimx/SA
zG+kqElrTKoF80UmhY6m+ZZ9ylG6BYPt/zJB/J5kgIv6Epp+qOQSCIFYil0aOYbLXekN2U3NUzLC
6oZSJ5DU1RIE/eQorgvuFHgHHQ6oFdrjyNn9HDRH5/IncwMnatQyLDmQj2P5YOyS6jQ4mawwByA8
k+9NupVsyLae24SzhRvuHkZ7RuqgOhvze5fy//+GbzdF5oAVclfNt8Koo6dW6k4Cn7QjyOtk2Sht
jFiK4rZ2FuriLmMO4GaMj2UbEah6Oo0O2B+OefA4TjsCFcgvExLKTivPBaWjrQ3ajN+2Qo3n9lUc
3ae7QaNuAwanKwWqU5aClUp+zu3CB1l/dJto0zPVlLhzVTYb4SaRccQ0VhIARv3tY5IVVI0XSkNq
w2iRH4Y3AhWwoVrAc/MUu5EeqgHwyLwa0UknhIR1ybWX6knGyiJOzq/wLa/n34KFTUs0ApTJ4LGA
zDKOKSRZ+d+aIbWDN04QzjxHubh9yyDmjcMB1/S2BodPWxApK4+nStLsPzjLoomlgUt2Bd9oXeYB
IIWsaCQxJ0EWdKUPOFp7cW/iHU0ZFqXbUWKXRhZbA3PLGbKD34lj9pnN3m0pKD47Xi5WQr1Qc2EJ
7TkEsUexVvLfoF7s7RZMI5Ip2ssquF00BYbdfn97rplrEcwkv/nMS1mBgoqbpWTOpvKxOYkI4IPW
vLEXYJrjytbtxlMivhc990I2bfjUorAeT3eT6I/04GVf9vQF6U7uwhSGBgRtThYlBjb7+Di4l1te
iyG1VKQDQdevKozcSORwH0lHBhDSZffU2ag5azqC2ptR65LubQBD5/Qzb89fmySJHFTlSTPXyL5m
NMNuM2+Wd5g6OMTwHtWud4xkuWzsFR7q7M3zc8FWLa9Yl2YgZpfrQo5nr+hm6sRWWS0QjTJbfWlu
v27+wT4UFgFAyT3lsshqgcfWnZloLskWkQvIeEfcvx4IBEd7qjkKbQJutEyLTp8gzpPhYW9mZw7D
yW0Zgwmfk1DdoMHNDxrHD8JsFsZwY5juEjcnh6URf/4r6ygiYMZtUozZnmwaQT1qRVmWixY4qgrF
4n3+1dOUPP6BELXdPl2Itz2G5yEtnQq5qG0wRAasRCIQe0Qr2sj8beBMjkJIInw8u1B7Z0qPRb/T
BJT1Av0AAIYrjdPxk8GJNadjsDK197zDuNsyD4/VtsyuVqiIYt4Nzhm4JYJHcvIfjW0+C9mWifoj
0uvsOmR9Y6C6WgcX347SYqai1yEl2T7KdFiemglP7r/7+9lUZ/i8BpldsX5y/BuZ9xO/EfFr2JPd
uTeI+dITJfh0beWLCABiL+ImHcbzHKOH2KNKNZjXcxlMpL8IBYwetg3eS0JMWHxxAOL+py+3cRUh
z5PLlD65ArnGlDIQEZ0Sb5+K8Dv2eY647ljfX2XQYuzcvHtTvwF4Et9VU794eHTgHX4NKrHTICbI
0KcN6DMabpI8vjDhOGXF47GAxZpC3Y7FHHDNCncLqENtyFVIrqIf/kDQosRJABJc8QorkY/orS8f
4CL6f/CaA1MLGWJXxXpUYDQ1FPvY+jl7YLMuGMFa/+cbI2uXoqx+8wU9nar5RTN5cYyUcz7wqcXq
icNSHcSsT9SnXScaHF0S2tbBO6hVwgKrXNfYBDuBW2U4JPoynSW5jGd22GktGj0W4xx/yNgQrVyv
qSUxm8sPcbgBW5l02yyIe3YgUbmjfEdpRGoaNnz+qOTPBUP/oZF0HAgxXdkPUEudQd+8F0IaiiZ7
Ova4EDSmHdUTh7vxkDSzBCfvJ4yjqBzQB/jipe4Z2Hd3sdZkomSiZMe0lOTHfMhIUUBCAj6YOzk0
GRtqaAftQ9LEMr/BJ47egQFhuzQzi7Ym7IozmrEyBtPqTyz44Ta45zBcK0SYc/tu56vnAJYGendg
iwJsnXd1Z0bfAkroYVKba2ngT0DipcB2b04kbfOTSzvnLtECK4/JEvo4BADRP5uMnJmFx7EJ/aMX
aiGaLwIcDh2kldrVTmswc/LO8aHK83VzJzcLjpmn8YdgGsv8sNbODYHXgcBJInB1BMWABeFZYAn+
Dk/QMj7MzD2/P9f2+Zvg3ImqCGAsRciWRtjnSOuhiJEmFgPP/pE8U44wdKiCNkH5ly0Dm1QNWy4a
CePldtBwABGnPh4X1uUvl1Kun6QvmWOwyhbqlB1znrgRYAWI0Z/h58QjpPWU1OLoAe7+KAxyWx3g
fmj38UIfmrjrAZqSaZJhINjAoHHzgHg22mSQSR4gb8OHeitO8V4cPY24Ah/YmGeeL2XOG8sB+p7j
rcOCc3KhvVUcObKaKcB9uSY483wQCvckvSrKM64tLO807Xwr6t50RscTRiBLf4iojN////PfAsur
TFPqBE1ViliEhKtemkDzggrdxCsPOcYGh0oLSfh0hyNelLU/LilmrCzBAU4AkVRbtSH3qoDLykeA
Yw21n4J80aoXap/gMF5jkvgHduLHHndLXOPCKNvUJ7RHYerkQ/KwUpJWgwPzR9CFLXJyYJG0R9um
SsmE/vQN7/PBGOx4jxf8pOBfHk+u68HmdYKCudhxQUGbVAZeHp88W7J/H0UvChskH8EjEbqS51cL
D35xSIrBYTDDNLty0Z1OPwW95se0oZNB/VsDaHkrWwCQT8WGFsUBQ+C5jDNu8lfL48kJ/J45D8F4
MCuc6b/h01D4NhD6Ih+/5Qg9jBXtsvfBPINXJgkMwQtzaCcpSM82FFTL+xuQg2/l4+trnTld/vQ/
z2Jh+Cd4P0GendRHtW5HWxW6bTKtAMzPThHFydPZ5SfV1VV3RdJjUlYmXYaRNRRoEnHFrlTZRht4
5Nuzxlq0RfGHlOF+qB+StvPJ57ZGlu5Q5mKjBuHYBFNOEEL5cXcTQgw4eYBxCjOI1XvzFwCKpi/7
fY2Hp9Yn33nlSQ5mU94wmsPVyUiv5pYK3HzC8LXUkArg/qpOPGaqT3N7E8YLtcF9r6FPw3y72VgT
ywKs7PeOdczx+6sNmhRtgv77Le3KO3/++L/69FM+s/AAMd50wXBtbPuRj7nclIbNDFrbOZxLQxxx
dFVDMrO5FBM1xKZ3StulXkqkxrEGnW5+dJr5FegjwZ05E2cwtK/x5mzxE/rw8SIk4iCI50Yo44ss
N9p2bqbT8e4S7UIyt5ptwwn68YXiFoPzW8hhiTHonOXjt3oabITyIkkWbrfbeCV/FjgiYw3rU3SW
sw7IAvvGtscmcPxtQ1pqlZ+2fffUaq09zyitgYj88D4VBbJrKwJNuDY9DQLAcU+8abTUATHmiK83
4Wov8Ne5qTrJVb3pOAgH0K+TT9zzddYeo15wSXbMWrgpVb8/sH7L+ArNytXaK0zJ1YE73TMVHCZc
58PrMhCsCVoLULDXI6xvJabv18QB5FX0kfr1CVufGzopw4yt2M8UEw5VWlZ/ArjVCwAtQa9BIDHC
FsUdS4orqPza4NLFczhCItbEq2hh+oUxUS1I8FoPSFZVhN8D/SasKrIPWnNdA6+6UCGlX3cquUAA
4mpyXpfDoS40Q+CSihsfm54LvGVxg8/TbSeOE3R0H7ZF9hjeSNXBifZZ3S+4s/+YZv14nJRDVd/j
wV3uuoLuO9gh1OsklCf2OfFH7/xKeXNOS7AX+94zbTQH0lI9QgaiN4144Z0MVObwngZ+dPHhPwB+
ZHvA06HN4Ip2wtiyuurUhzecjF2XMFkgN6U/IgCVvwWYQOS6bNDP4uJiChJNbjcnCRiAGa+N8asx
K6mLt+k0sz1OQyHQ+Hb+hd7sDI8pXZup7GisMjA4mHNg3vaDhqtsrKydeDRclo6YFnmwk+rAiYw4
pgLc2/asSO8L2ws1cAMXRRJ3S5+NAW0y9DH3C33KAeUGxBg7/curzrPnIoI0G/zhS+xr98feq6pa
fYb+wcd9rJRv3wZGnfYNhKspMS8MiZiomoQChLOp4Fll0aI6SSNjfB44XShZbmx9lTvRFDgIvLWa
S4m+hOfthOF29oA5bNymF7lBOlT+3b4VjgvyWlY0pJ/u8aK3pygQrOb6rtP7bptRmp5cJin/GU7O
d0dDJQBpWbZpQX0/ecJZ6JkCXip7l1fw/6EtL1XXPOQD0xZH2THPS3aGJZoOUz3PeK/6KE+wtcdR
4frtZT4MFdjRMLDqZsY0kgPKNcfI5HqNLEkhtJx4c7y24soBk9sP7i2OpMEffcCoXxnPqJfz0mfs
Sij0audR6Iz7kDkj3ZPtpOlvYmmY0VEFVIM/SFJUUbo1k2ZIyWRykir1w/DKgKcxQvvhUWUZ38TR
phXeYJoIc2fVdYeGDHQin6Uzlg8TaqmyxzG5eVqhciwF8Agp5FMjkoiL8bRrA96pj62i/jX2X737
ZsIVJIhJZcL5ngdsfe7hs1SNx4OdWyGagWHO1qqMlnxJFln+xlxXuiICdHDhbr92pRbR/D50axnE
Blloo+2M4UkAeTNGOSumF7e9xfw1IFmvLUrkZZqSp9toUP2fEzNdUZgoSrLho5B8Jv6IGvWa/XO8
e/zMlsrSAnN6TjIEeUTHM+Jo6JuPnelLvSJ+7Rn5EC5fc0BDG+WFkEqHaWYsbhAXC4wQlJ4Y6GRA
C9KP1t7TCRMkRMMg6zM6q4Tzgvq/Wve91KL+7ItpQ80LnXgrDHATGZMTP9D/AXToR7fxChSW7X3q
xINF1/bS8dOHaH6hh7hxMg8gT+jdGPqEKEdrGmGUc1il41ZdeSOkXSnW/HfiR+l4T0jE0g4hXOG5
GT7HuwLhwOqG87zL3cVDs/UKd48F5qqv5w+1aBiyX9sHbAQpSsdLPELP7hQMphFGa60dVcxyAV0e
8T4rMtpgvI/VIBwBk/zD209xCO/M8ycTsglMr4zDuPVMmgqFnqj0FlVK+0Ss4Z+kSPMGgE8mZPMl
KpkVGuZAcDys3LSZSDU47U7yhpcgJk/VPFIYPT+DiNZqFITkc7OtQXe1jMTxmn3Vhza2IhaSSZzx
CSY3wgx5rD/1hfdpz2yENBZAaxOCwzziIi+YhoXPTLEpwAvc/jRsbflQlVl451S2EiDkQ4EiZOop
fenLlWt05+cFhswF8h7QmxD5HkjvwwfoTJ/K+/NiQ6cm6l64Km/9MkE7RRh8/K1bpjljLaIvyoBN
jajo7MmJkwitB1F5kF/PYiilg/x8I2NlR+TFI7jbvss/XGjxYXizQvEuXdcGgfG7ZfzpMln7i9AX
qqJ1Tct4IqJuV6MOnqR6QOGSuk23wmM8JpLFw594AuFcr6DvudA+xdjbjaXUXzSHYrQFmxzcwtL0
Xh2O5514jUMHU23fRv9aN3ssnZ6ETwnKrhZXrt1qqLt7PYSsiiHti7ytKjwqfGQMaV1qk6Bvl9lm
8iWwpswC1V7iiuA3bf5OZwCk/mm++i6pGoQLbY9mZLBo31r/CByBM4FobptaruWuXbsCxm/ZPRzp
zxTEA6sePEXeZiXsiAn1i9bgQviVoFb5PQ4Gc1MOzIPr8ABbkHRHnUHFGUep/OPnfRChgnO7+Qzz
Gavp8spgJDwtGOI9+UuBd09FOUEI644u9ok/2z7txFx8LffLmW6ESjORcTMXk7V5cFpPPh15a/2C
jND8svjr7fX41MArse/t4chepzTA/R43MQmf+y3CWn3HSe4JAo6jR7+YfSDNAzG3lGmzXXkDjJSa
8ss6EMvG1btA+PiEUA4qcUaMASuioJeiLfbWF/mxNEmrXCyQSO2cntat33y8Zk9LyvKlMAfeZUuo
wFlDd1CbTAA5OxxZ2uGvE9fI7H18Iwgh+4EmK8yCvMyNXEAo+Zr74XFBkfMMjHzL5TSP4BFloWTR
uEcGqS+13cGeExBmtEG57Kh2al6lI4jRZeWp93fI1VLjT24clxsX53Ve63wyyRWLnBLv6x28mI8h
2oV0MVLta1COXaBjGyk48bF8tY6zWh9RwScmAwGiJFbaWoKvcyWPOPVliKFiuZzIScEFsK0S38+D
D46mMqjcKfbqm9c7US1LQ8pfQuiuxllOUIuZKXyKoqqdlQ2+cJhPq7PzQ6LkkcKlwXoB1EONsStO
RaP69d6vKOE7hZxWRraA2sciZ4DK9ZcVLZW+vCQbdt8115GciA460liSK6gXlq6vBdXG02gyWOIj
i49uVm/6uJAFp9S0bRxMxBU93mHQnPETHnA3GmEhpnuADmGTifN3douw5tXO+b5r6S07WVPi5J4Z
y8kH7qq13HDVFNpF8vLbAuVQ/MIsH5O4lDnuARkEnfQKLOm+pegY4JiP8yuN0CcNJZejlJPYLaYA
iW9JrTX03V5XkZJI6ExdSpLeBOkZT8AXp4ATT8ThihTwhm7MbfXwAwF1OLvrxb5iKZMkDvzosfXW
4orL9V1l11PJqi3HGE1snEBGfVmlnAN2B7HWTqta2dJNzTTMkXH/dhkKjn9MPmvAlUVSbSL5XY0D
ImxsJbmK+oxWsBQC9afjQIWPmnMhlquMT4CXnPioDPuKEtMXob6ey+VNorE47Woysc4qC79QXRvG
DDcxVrFzZbjSQicemlxf3rL0tVUq3QMrsMqdQ+2+SA5QS+7QbSLexQA4TfSzHQ3ga2jmlKtLUhK5
cyfrhGiB33n3TLcMZMvBeRl+H/D8juzozVGJTFazm95w3rfbI6RU9P9aSX+q+cJYJ3lMpVZadRV4
rf6Qm1RDXoOKRR+MEp1gIqeLucBwXaYLTv/RYGfP5FTzUgYQZX778+J9Kmdc+Mzncwl4ZG0ZNrmJ
7xHXfd9wNIo7EqCP3KiEEcFzbHnxWwKNP5k9M7KWObWNMihGh63eochSaittPXZcALCHr3u4qYoa
NUZ6/VT9c8tmKfJ17BsluHTMGLrd2wUTXyTRbFhwEhYg6ihu2JfY3fwBm8TOV26rDIhQoowAtwYe
wMpNBi7v0nKT8g36h0tc9F+hBwyXw3wKcVtgIpI8Q+iY0M/LMuR5qANyYgZJh5QPNDDQfhPUucOJ
E+GaW5HszSXTA3S/kYSCgLiwjozyx+heAjqN4ZH+pv8Kxxfm9Vl1RPD70WemGGk+ykOZQgyYj+mv
2sLFKdDqMdxv7X1K07lli8CL4v1R8CrsENKqHSLtsPleUHalHE2/uv993vB3p9rnyOOKG5sduS22
ebCNRPT/2niJRXu348nvhUMN3tR0lJJe59DLsEmifAzjSwbcria2986PPElmy8Pwe/LkH14tiXUq
EhqKaqyNl3O9CTIGEK4w2+SvLv41p02n0+lCDx0l2al9Ib1QTNpmBy/fjV8flUCsAZCuTtYVzWiu
rSeOF7gHJNtPjR0zFSezB6PCdrtDvwUKjmvLoumMeOD4fY7FhLSbcl7kXI8B8ewrUQql2GlYdW8A
aE7uWKuuiFV/0b1TT1J9CBH7gy08HJKjXeAMM0DDhlP7VasvIgjSjGKKUDdJLihleSsFigIXtFLa
oZSWudD1zyOvoqExzUXv7fMB8zcjDp7HIv6K+Lxrpk6BTRscHfEHFNWxDvG8Jrq3Nn0E2kijfrrf
jSbQRTjYn+GlG02xHQnWRJFOI3nh5msJdSz4Xb4KI5bIeeKuxU8v2pCVuAfgiaZ5NHy086JPLMUW
PtOvvIAJ/XMBfZrpJzKAEIzB6y03Xah6kVypVIkfMSM4RBX1SKCGqSWz9WPckQQpk9zRNDMsoIEi
qX1IANllRg0lvINVdOH8mCcyyVCRuohbRUaAA7jf8QC02AoDfFxuyKGjkjiD2I/vWsrbLs952m+C
GzqfJjOPBmxis4kGQC1T18wGvAyfbT6pTkRuRGE2ykYVwI0bb9yIJBWbtXTFPfsFsuAVDNlJQiJ6
fhPTl+piiMDl//MvnwKkznAo7RpevtcV8urdiN9OXpzrAFRZ6faMg22mqWwUyroh80jiLz9YTmLe
GXL964EEdc9XyuRBOsJgxDYlYx3JHZPc6B0xB5up3UywtAAD22kuoPhiKM+B7wx1JPgeKMxovg3Q
Zco7/elrLs1zdBYFcXZ7TpzRQprlYIB/OirwLZrNcd02Ps4SDM9aWeGhnQUaATyF+OoDf78ZnApQ
atDjWqukZcQ35CUuEze2miZQuxVRkDnuIdHSuNxbPTPHYLLZ+wi0UnlJN24Poti5MjYD/OqvBRyk
HXYPeHj6E1lr2cumFkPDD0vSLza0txZs8OXOCtnzigIyYmxXPtFKTkVM2PTuuEbPjjqln4qRt0s2
YObXo/dbg1wZDn7c5Fc8ZCntx6VMCJX3cza29R/sM3GcC3zhKvA6B/Uej1ofIHyFkxfEFeaLCg/s
woc4FZcwrF9tjK3tglc1c9GtQ7SQ35EXJvIFQl/pyXZYCDfOnQiQDQxofn+w9f7TJsufteGCWBds
+8N8efC5uogdCvsVfwnkRcMjsfLco4L06QtdUy6fuG3qWojN0jAuiHq3Ssbx24IBFxJWy0aEbPiP
hUakpVdOw+gH+fyZDCto+iHlcNdPYrlmtScOhEGRP72gFHSGNuL0ERtnt3M6Czox0tZG4p3CzaZ9
ISjFjSf4CR9e1PBNuNRf0F81lj+AlWhJMUPegT41ghyKeeuzAmC07QuohdWL+lhokdBCo4ZrAdCG
LVMkJqrlo5g/D076+nyys1oOTqFFwWZM7thb3WLFKoo8NAWFRfUySzIQ9GlHtN5miUK9dV7IPMU8
E2Mxxs0HC1zu6GwONXlPjr1M9VtdYdumqiHFbmHzF/xRCm1pfwm9Iv6n5MfLguan5d8476XfAcYF
KSkA4QyfcGTq4D2LkyojIoArFEcOrZy0WqYpEYtrJCHBkTlaRBJUGkQHG4DFm/OyuId3tAP4b0be
2FHXGI5pOLfi+iBMnCoB+Fd/TMn2/7XpsVAtZ/n47n5UhmO3KVzmAIy/aOpUIZTYdqi7SdcF195y
bHBXeSVS7Ud/Wl8W4SZj9dWFu8f67ByYfvriVert72kfnfyx4ai3+KkKw1UnmWjISmWb2yWXfwXt
jiT+Xl9WvVBbHfrGWyhmfq3rapNjjPqA3usVz5NZQFiVbvqlVg+PshSgnvkg4lkEMr2gLCcQ06yG
QlLt3w10IqzOkD5gzFsuv0/YsHTbjejmXjqxOVM5Mh4zEaPHO5qB8wY4d+G7H8KzT2dDPR19i+Qg
WopNrEGLR6o58EFtEu97Aj8l3H6jFEharDx/qdKlEO7gJA+Ul2AKqic2LDzsy26IvuGzrT2lyzgG
eY0TQlHkI+ZHJZ2B1drTFx7Mw0PTanWOBr7gbE1ne8tflwBaGCn/XxcvSpi1i5HsWlbEFUySIph3
tLP2O6IhPZ1zAbACLArfr6a87JMLSMkN50/CEe7XLzjimefaL6JuJRW1DcIyUhYC4GSUTim/V06E
DLZMZcI64Rz6BKFC2tmywnDGTOjYmboBDlqWo7bFjQ7YJ6uRJT42sUTqpJ+68KwWsne5YPFlEUxv
D3+8gDyCf6YrDQ5U5ONsWN/t3YsRoU2WD5uTPO58G2J92UYMYK+7169RP21eVY7qgtRqvyDctpLi
Iw6Jz2j6b68CPiKHeewxPpvVoNhCeLu2YaCMIu76aP6DT5Ry6qQcMNPNrGCaWNcWv+FtlWP5pC7U
HB3GLgnRfA/ThYtOkbs/nY2oQbl1t+6fuBJdb1WkwZjkIQdqIkfjhdjvNj7ZmjU+i6ZCCRPfBu2L
NjczzfjXanU/lop14qEn37e5+LAwE9LFZyj6ndL/7PgO0mLReFQ/fIruV6sjfa6dK/79r18GAONn
0HujIVE6L0VOTbY1sMyJC7EGL+Y8qdjuDeq5hgSwi6hFo1Aju+q9Dkby5Oz1SA/KPGSjSQBGCTSC
eMlDGdQ5lcb1OMO2wIsaT8TM9UemyFh97lzvbPj/SfEqVyBnZ9LBN2bO9MeLU1Z87Avq9cKcoTp7
Vi7Aw4bFbGCylyqD+zDQHlDDw0jEUtEmSQkFwLzVhdfbeyME/Ossgqi7Zf/fdSNOV5yQPOksQZun
EWnH4Y2S+9RTdu92gda/AZo0rpmUJKdEB6D//q1A4McuiWFyFYbm4K6wDWYElMXqUWzazsMq6cto
MXlvPt4jFocaDIavEQq7kg6dPYg/JHA0ALjIFy9jY94cxcCV9noP6/a9SvEETXZ2Saw2OJOyqqR6
SKtzfRlBNsOuAPNrlfwDRD1F2QXnMCk6vs4+oBshtvI/n36RHwrDYT3VDNVz6FO4ObEaanNhxjlx
/xjT3sYgG1jSX9lWFifAlzKULQP5x2ji7DuR5zXzWNMQo17ExqGRoUDitzlEbKgt6HWDyCnEdWZi
n19KtaGqafRwu/1VYeTT1H1fkI9pNdY9gZ7tr+NX9VR6Pi/bIwntee0PgAgpGqlTXuy0PXwA5L+J
fmHfA5G2fbhM9bCSb55dRrf3OwdsZUtTcyhgiAakh+NkAApIsbCgBH6ok9EexSLupheUF0BwrQS+
y7cE/Y6sgWu4M81Ijh+pOicT8llXZz5bOeopblG8jjGw6M1y5FaHImX8ngcS7pagLIs2uIh6V+78
Y7jMl2Xegczcy22yy/Y+SUn+SUvTmxTdTzjiUjYCeRzo139Jvzk4kpWlokOYxz//oPw/CefcnkIU
aJLtx3LUjfFwMtKPGszXBdCcAbOeYAPWrKPJy2fcdCTXaT/toXYZFDVePWaC0SjYbS8a7SLPwVfa
1icrA7MgzcdxUeNVB2LIz/DDGx3hH0AeFhj1XS0xSErSxbojG0l3kj0fZ7zmNUs+gC6rJ1RkiNxa
Uz4XBmocmhOdEukMBpgXC6obT6oUVSMIpitSvgzo4qyaIsIwhm+GD7YGmy/zDNijCBRCWEKgqmkP
8I+O8FZ1QQn++LBNaakhIpg4PozuERHnN5XTfIRe800O1R6dFk6UZp3mnvxd5F6R9dePpF+KobgM
ZGqTEHZ3hrEF8hGogRy1VLpLeRrEK2OZRS6j0DiktxTg7am1awb63Y4x0EMH9WIQFF1fdDctY6X8
YMwP8BdH4HA4vagxA0/2PdPsEHCQQGBX3Uf0hQMlBwfx4WZNl05v+hcfw6OpSXKLZfH08ahfV13F
Fz2a+OqLal5Jll41OVll+Jy6Gd/cBSOlSZWGvwYWS+sIp00q1WdZsMddrY7rtelMRk2JMXgGGzaz
lYGjr1gxtsa6lNNOLRaPrVthsth0xIr6JWBXyWnOUTjGOQfmjazatvl7foRBWRThn+wDDU4LReCH
Fuf8NIikcazAZ8WJsyyVSPBL9BPj+yOTWJhayi3whlTKa+sYeRPOjYlCAGmsmFZScITdctLxrX4U
Ji1JyvzD3yxqoyHdV+OQfQzLB0QTOv/nwG3pIzQYAP4yzXREjN8gYglYPkoW6pujJd19LksXFYMd
4jwxlUSsWmE2xw4dFCLblMQatwXAk07BugLzHm8xmBg42bHH4UpO2Sy+YMeUsk7opbjZoWl6AtFH
ljyvLJP7Jw/dxp5CY4GAAolJOGNSSTxLjo4EA0gZQXfuuA7aeFn8f/Rp1vc23EbONe9fx2UHboDR
6gGxm3CVrlI/bB3yVoeuOr68JcjKZ8fD3GRpvsh6eDNds/O8MM2IxzP+hjI9DKUZ3HqIRzWxueeg
6xBW0bA3fC/GONCTlCZElTq6QyrxcpKHrvTqM7U1LWzQf3e2hqqHN0ke9hL0aZYqq9G84TGxoyke
Sz5slphWdLlPKO27Da51nDizVl3yJsaj7XlXKYh56caWzqJQwlC0paTuHhCoEr0hQCtdKLhas7r6
AXiUC0a8QIebtK5ao0Vbst9G8mdfxksFleao3s8xOLWYCRjXXmkLDUZ827aJl0Cx7pjt4L2aw7VY
Yp3XcwCibDV5rwAcuPCY1rmG7MfQjA9wz0ggYdPFqCJOd2vcpwBPk8xSMq7wKL6YXn1hhOiGpvoY
jw0944+iZOiQWDpilhcgbQDims3etkxC4kFPDeMaJXM/S2KVRMtKN1JnCXY106jz
`protect end_protected
