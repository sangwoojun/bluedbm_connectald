`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gxSc/rVkw/Cf80Cm3arjjAoQlCTwhEWfl2jEPPVNt4KhuRmu9IphekQowQ+MrEBCHrmvLDNUk/R1
DF2l+/d77g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bJnH/vrXi/AXNHSsdKNf0oqe500n2rr+s3M4VDS+z1hNMYHjhzf4H/9EsQ10lT0u+lPlD6KhzkrJ
uc1f1gBG/1fZfa5YGqo/7uld8ihEWRqxJdk4ITEP8F7qCwLlyCQhRxAzfRD8ghUdkKUFTJGhMjcd
Dwlb6wToAnrP8SXi4I0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eZVAg7J9O80pnzqGaXtQU/BtH7bl56Fbce0FcraO+P9+MAIY43ouhGCqpgn8x8Gp2h7BAZGgHnb2
u04/ainwTfghFlVTT3c7MzLZtshTRXDP8gLcLJs90wbaGyvAV11C8XBs2rBtZbSX5aw1VwaxtE6+
2JApdinVq49GpgW2vHkVAh+LXKObHlm4t1z4I0qu2chHYVy9Ja4p1v9LC21QDCqIZK/qPBpctR4j
0cTFZzhOfhVrme7IoLA7EPFjzCwsDmRNN+pOKAfeOv3KNCnU87XaWCh7ZAwkSmlijJ6nh1gqhWpT
QQdpNX9YeS5kDN9CSqg/eeB51USufaHqreUJAg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lhanFB55e9zzb+9KISY7QPqyy59yC3AqHSLu1Dg7jJCsH1PfHUSdrYmJljHyyy1GyhFGoa8cPZZQ
xnDFlEZJVen9zfjRQW39LNliS10pq8G4T73qfP/M35uZ45uBCYR6MMIYwpyQjfcd/zeGRnjUhfMM
D9UhLlmtHJb4Yu0Zrjg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IWOy2ixeztzD95/O6D56sjdkzdy1dIWR6aCyZwL4zxkAYUm/CLbr43wnvnB+eopCTRQP7jCzyiH6
vQSt57g7O5x7q6w6DokiacYfpbH3vJljSuztgpEzTPeW5U6epvtUPWng0QrkTq4zdoiRLJLyn1w0
zK6/XtquimefPalWHriTvJHvAbYzFdovUFqTMPKd584j6+A8I5YI6xBYrVrcqolBpS4n1ggB5wMk
F8wuxk/QDg1TPPQ/5sT4ElRUZG0Lek+xjNCmhJCNuIV5AkAX/27C1ioHPxuCEd4OfxSPMYNdXnP4
GkDpMQZKgndiwSM8LF8PLWqiwSj/harG1cP1Mw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48992)
`protect data_block
xeVF3th21GUN9Bisd7UiAsKGzSiL7Syp/Mjbg30QdJNGvA/2KdzGD5MWsltYENcFCpXv9IasOvCi
Th49rPJoWkkamDjlOuMuEJ5N3QJeda78MOT2NRBmsf7VtxF8FlgqcRltM4MJRoEdVfQmvwiH10rq
BSD8CNC7zvM8cgYKvV6Jj30tnoMAQ/NsAI0ZgeHdD6rXx1r9PequhoFez1NxpjAp40AT3DsVV8Kn
nYqhikMzDzUwpP2FqIPlRmxz9GrfbbuMvt6xD+w8V6ZyIhiX0QRNeMSRrS3NrTcj3BmgzQSmDjIq
SFCOeO9ZYhFeu1lSFXAe1UuYL6+pK7XeOCjN/1FfHO+SurPDhBzAEt1eRnVrhTFoRU7EAzLQHqBW
fF3/9kZTuwzQ58VVKtJjODDm2pYriXPTHGTztk4br7Ay0IdClTM3oXgnz/yV3bNIwaW0Uj8086rm
mPpoXP6oaJUk0BwhX3/HTimF0BHBOJkb7L2M0QEMdO+M5yS4krg4KPxxlcnj6vygWJ5BuUnJwPwu
+/9C7KoFOuh5DZifBOOTsuHQrYqBDirwYdlkGSHzLW9lZKCI6QYyUkf4WcmiFYKwbFyjlxp5r+hz
Kv86ulbwaGg8dk4dwDk44ZIXjFxogNC6up+32xxdJg5eeZR1fUn1i73EHvvsQrKyd4aeHLAbQ3K6
bq1R3ViR+Lrg3iicnklERsMrrymv4m0Q7b/i+gdEkND2Vc6VIE+9z6U1+CZ8+YiuwfOuyHhD8W8X
wyJ3JlDIVM70jlO3zwY06rIBeTBBRJa19ROKWnCrsO920ltIg1gF07wumf6wCkaRrM7wEjPPlyuk
iN1xJk4rkjXerEVrrCn5rMz0z3ovqfUlmXhBIuFTX4Xwcn2hNVGCClU8+DZdoiHADYgfXUklTBW5
8nbk5FeR+S+RBmpEd4lacLOyYGXdV8G+Bl67/GbSbqbsMl+qB05Rl580owzCslriIzVfxzAVRrLt
4GgHM8bR7PdhtiU3FvPt/5wxkmKUJH0DHxWId8TCXu/QrG3fOPOH7WjIaUNHBgZThe4aHfx2fLIZ
waPJbBbzG2w6Se3S+UxsGIvFGMne5JSY9Nw5aL/Fc4bUoQTp/UVJNJKD/OCZ2A0i8sIuVzaycK7E
Ig+gElpaM/Kd2JBRoFdhd8OV2b0omzGZ2UqxN0x6V+Zhq9JJ1NL41mKHntE0h8bIsOpz6vcvrPnJ
XU6A9SI99PKg9UHOs7q/yhYvBXVrS8fAEmB3912pZSmc/5wISufm1WiuwfsYNojhfbk9xlfR1MZv
7eXHyAAmp9MwET3aMuSmJfCtJB8a6rWxHqavjSq+QDeR1c94JoU2Pm0AknG//4LBiN8UwPZ9QwSt
ReRHZdnSvhEK7lm1tuiZw0cH3Pcul4av1fD6y8pkZDnWN0LPoDZ6Gvd5zz6FLIHetjd0nVclWQe1
gfGk8WLJvmw4tNoTNe6rFYezIqL2RwThqnOTtdgwlhamxBYzuxHqaBTeNj2of/KjcIRA8Uzpwjcj
qF3FoBZqoDEt1bgVdRH6hZgtJzKQj8pKKF6rLxw8HHfSner5PjzsemwBueZTUAO+cd/j+kHc7hqs
jhF/uBCR9uSFEVchzqq5Fm+jUd+wlzyDOFrKrfUAiL5zTIT2W0inhznEMVntXolUiy7H33MUlAef
EEus9RuMYFjMCz8MS6pP4cLzxy/k88UPvDf43V12Pklk9Tcww32AmUts9RLTFEJiu9gSXQMId9PW
uDVRbi9ib2Eqn5Uhiw/l+J1GTcc80B8vEvkAGWO7/ysYoHvVFyDmlrJgmHjvAop87sKVGJIiYFN9
XFOfRMsErryVKosreznPeRIxVmU1U3RulDyssqz0BeeK1uMxJw0jrp/UJq75FVlb8auiih8ewJpR
2gP3OaoYXo9Y3K5X6hdksiMr/Bl2w+mF6cirRrZ2KKtVZbz/32Ucg0qaFfeV+UMKgwqPAV/D4vdf
z5iEcJ+B/kecQk21rLln5rch3Lg/v8lRIO/wZHDBV1u54MkWbd0OVz1yk8A/zueqypCtS0OXesX3
XE8t+lX+y9QW3RxLjKSHmTGp+3izBZILL//Rr/S3SoaQrJaMUwn09xyXbfnTDMn83I8RDkFh+qQf
6z+vrgdYUra3u5tfvm7biklimIToqGPIccuFB2f2qLef5fqTsW4/uJi9FrsWN6OmtktpMRFZLPLA
F+YJ9z/G06IO8Y+/4ch5x+Bfqg8SkLDex2uYK++dez3qDgTXd+I1k8jvjOQyxcyfzhXdj49J7Cmx
hydobVd/n4DSIp4HrOGnngTML3OUOBaetAfEPvHzj9PEazPTN/UKUwRoS6pFSnq3w0o3jIBorTlY
Qj5qFSLq4n4jUKczYdMwpsMjc4I8LL+LzzjNJCPo9E21cRDlTv0BFsXeTinpWlo+YESnDQHlt/Pm
JdfgKUc1C4yjUpQC1s7cGuHQBBt0LXcc5tQmYW9EfEAayhdAbAWlYARfmyMxLciXYcQajZpsVR3s
ZdfCI2qlGhev0prbSTFUonww63A3hb3kPvnFubhM4aKIkiAkU+lwm7xhunE19dNEGXu2MYSUiH9/
lxctpMAbRtciopoMUQx9zK/5EubvR5NL3035LrEwoLSyEPIUNno6xZug7P+bs6UFUw0klpWK7NHv
726L7i9IlA2ehyO47qaXoE/j1tQm+u4iTdu9/Qtqww8BFzRE91IYzs8fhr8oO/pdbUQkAc/cmmff
JaXO/YX0+qWJHcFoo8JDCDWbaSBUKzf3RmCHo1s1fYszdpVpk8jQLeZtP4rXYFsWfhkkXhIdX5oW
pZ54Vtz7A98QYYoZcZqpup7kDkzcoGMBSOVhw3D9ZCtEA5xHxanhNkEDhjkAxtjpssJlTiBsHpk3
4FPSb7r6WwTCCtTs86KQ/5LVZxpR9gajjbMrlWqUBnbw9JOanpw/cUw0KV63hdR59Klwdv0IBBEP
zza5iHTazvm1VYkkCXnaJOnT6UIvuDa90UUOUD7WPKXBxiL/en+snQOlVVWtzuUyBPEBYW/rVaC4
xqWOXxUrnUBivtGrJtcqvAis+Hw7Os+AC5eP3qqSiWWtMWSi0oXm83hTZlI4LV2EHp8Gk/ffI+LE
XRffrudMEid3RONVcx8T3eMXjnE7emjEsLWPmwROLVLejTc+uku4yJwfZU/5YO1h3i6rsghsFy/M
bnAlIohTG26sTOt9pOYWGrbdRtSQe/MQGtA3gEXd2dxkLNCu5c0PQJZwj7ys9u68PC3PqGP1Jwfw
38dYoz89fVcJsK3gvEibumPxCOf4AqT1NUJvVJS+5bK2hccLagjLkPsMgV1MKTf5oFKiUGBURvga
yiZAIhhpdoDAMHutdFqjR1FYTJjjIz8LWv8QbtNeebop5kNr3YSXRY/xdoqZmSyZPI2HiL8uEf/b
Fa6RMk/pVkYPAXKYWCr0dNAMEIGQdCnjh0fcs1iSNc28aph/mAM8HhJlAo8m7rTJ/KHFdFpTIQf6
Pd5XTPamPaboG9Qiz1lZscNfZ5yn6Q9jOf4fDA9D2Nu92FUJPpcWG3u+dEWAFI/GVR+hJn2Gv7iI
x9vbJf7rizWO7uagKMtn94UV3c2zuFEOfEaDKcyfT7/7hjRMxEyVKsjXJSeGlmmIkzbuMwBXm/Ue
6zlf6fcTF4OfTXYFFArLdNkbIOVW5doDzwHb6SsVuO+RLWmlPM+Ys+uvzM/YT4Pg7HvUznyY8AY+
GPbUcA8OH3ZHAjVgjGSCN72oqmRc6mIy38xdhIvGpsD0HWvwZ57RVRN01pKhVtWGbPdOfCiuY7PK
flDd5qjP38qxZUyBSXImtOvTAXRuxNZvB7zXPmCt2hEJCfKmR2HKOITBCM5Zvh6V+3nGBhtJFcOx
xZALHeYffNuA/kxpK3C2EmSwFW0FdDax4mTqFKXvkhhY2mSpq1//fqB80R/srZUvWqVRtOG4/vao
UOFIbB9d97ulGSkpcBKWfl/MvBAL0PN20lHrKgkoOgjhanDHlVCBjqWlCwZMVystoCYDmUbEdld1
d6rNN95G8q1dkxuCkU13PY1aqQzlHUrGFCG85ZKX/zAZQuwa6Lz1hLLYx6eQTUL3z/mZ6y6Jn8l4
NCJpIRS2zP1f6i77OgxQIAhbedyc4/H4DhKMWzCSDRNIqji4LM3+Q1gy8KnOgP1pWuXc2PdAag6q
s2m7Bp1BTgaypKE9Jkav2X37T1iUMk4sKqH04LaHesJkhp59O8UnTptb79FzZZM0t1RHAbzt94Jf
PNnEfpzk2Z+OnDYrUPq28panAGJNctsQ8Uwf97aGg02XL5RHC8pw9CIXjRnPjTfY0coIo2B7ydzN
Ic3Y86MWRFNQXGKyK1bN6xC0NxlAQU8Dik8+hVVUINHr18IrBC0Q5WCQ8pAhidoeJx/4R2nc1u1d
N6coNX9ysGl1yCAMCnjVFx1WQ9YGnZHLGAnxSXm7opLuJI4Q7LruP1zB2bNDQ4KuONOThxBUrpvG
BJc56YvvBpMioL6pbVtMBVV0JHar6O5G0ONB/ARVirrggOILaPsdFEeDGifyF3kKnJNfzB1pcYhU
vTA8nX/Bf8mM7FDeUo7JZKX9Q3SouJEu5bg5kQDmhVJwEgG6+PXGpRBcaDkKqf3SsTppr6QUtmQj
2DQDwJZcpdBFioaLkDFfsFMCsX06nDHQQzRgBHGYHKDDzI2akh9fd0H2g6lqS+Y0I3CH/eQ2VS80
0x/SuL6JLVyn1jjM2dvDgXG9QEL2aEFtLe6o5fjUDrrlK+jDqvdnFJQW/peXkMuxrUfz5nqyHAkb
CYFa36ZsafPGbhnof7W/7k6uR499MzrlPn+Agr5l+7rdj+ZMIi0wDqODmM7AWEV1QrwbFYeZfBtL
iDRQ0P7akZ6y+MbXaET4bx6MVr+NGHsd4NSQwPox5eRuBnCUHmqjinKtGVryW6MShshAOnh5OynR
doKAklDqQBkwXwmg/3cPgSz3gO3O66lgZ04srq3pjVwNZEyz8k08z4hx+Y+TlvkLTUv2GIVYA1hN
vb7jBLUSJGQXGxLgQY6+x8DNyOwACZ0dDxTlQ623ZRQH/K+z6yOMWhk7jmLJ3HnjOOfnPVwt9/jw
4ZIF2AWh1dwiFlDOYxLBk9pwLRnlMv+Azif07izyeHA/dbPNJ1xrFlrCcrSOfjOHiZY94pOM0PUR
RtgMdmT1ZgJIvU/j9BkCvTRpf9Hksq1tIz343ZMkOm1u7FKmtCleahFG5v841EHzIVEkkXceU85o
xbo9RPDw0jvGD2S5EFB7VfJt43kjUlbhFrs30/f2XLNQf5lO6S7ibKGHaNPhjEB6NQBE8E46xsHG
CIhTQD8PKWZ1yPyiSN8BcUCWd/zsOFcwtpqhumSUaqDwKq2X0x86JS2qaZS9QEMzqDFUuDXipf2w
5mAj3rMVxWI+29aPTth3X+YDpcSUUZVZ9SDilOrasOj3D6usbVtKVGAqYCGb60gIagQ7JwgGQVvd
oCBLFoYu7XoiY4+98sT2kplgbMg6S1AxF4jrnCZ8gdRXVWrbtthTjbnbnG6p5dPZaaRVjPUCh0mt
qIFRiSTTrV6y6YHSLtmPQ42+2uKOTtRTONahrlauxIklOdH6CKVqI8lWLzSEhDwTlH9mF0i6zd+f
1O64J4CgBBKNzh/w9npMPOZM35+R6qIp09g2BN3taJDxKMNAq+pL21Jcc0xPNgF5UJTvv2wVCM5q
dnEGHzfTjmEhjSKEC6mFPiXnTIRj8VDZ9OEuUnnqMs09++Z6VK75tf/9pC3oHVNq/Ih9Va56tEq8
tBOtQA9ulMMmZkts0SUtD/t1TYQ+UAHcsXpUcUvdKJ7PZD4MiXV8WZ91dKhMMNKlKlk865wfbEO6
8X/uvBzj+DEZQ33TgZUlk6HHW4kkW4qH9LmCbsD46BKDI0EkeFj+9+ZZSX0HdnkCaG7jOZcr8s8o
EGs364peZC1RPEOevxMGlgEg2ME3VcczxwxuaH0ceJVTJV37gU5G03iDUOqunzo/Ut/W3rM/SjTD
W7xj4JGoe/ocPSIoMHsKhkEqsf0mCISgS4ep2v6Dcq09QoX6uACMtRqKmo9GTlo6tXw56jZnsWbp
hOVH8BvSKoLz1rx1CSQVCcorJ345OhP5NhPGg56Wvexvr4hLpyS0/2Y5Ya13EeW1b8G0GEoRG8lQ
duCO0to/lemLy1SBbpNgJ0HvCX0b4rOVfjExfkNU0IEj22pNFl/zSt3pxgalJ9O+gEmsc2q39HJb
C0oAZ0sHgLilkj7ZvlaNZ49iAQRhN/hmdjrJv7CWL8+hxKUvysGX45nxEHRjB6CVlXFHIUM27pQ+
s366JqJaIj0DwWR7vgDnTx8gGl3jVDclY5JHtUp41hdhjlOSdOla+ZuN/UpfCAZVQKPUb24b4ERX
EPrIq3RxlEPZxEJ9bSOqO7rsRNGSH+eeAJ4BwxvNiP1pImXYiAzhVFn5yvCdapqg0vB+X4uKrI8o
z5TMBZnDnXmOGJHenQ7Ci7VzBWkfZ0D80tW/V1prGRGZXOTnPo/F5Bz0LCebOkY/JDweg0MeodZ2
n3xtTwIxAYLwW1pgs9Q1ko3Tz8+W+47MtxkuEiedGUQD6vFP+aFCzvJKJ37ugN6Y7lz6GanGcYT+
G5FSCDN3ffeHEpx/9k7goB67DQ6pIFlkkzZeTMiMQmYOu7EIU9M7da78xSky5C6YoeP1SXsaTSAI
NCdsm/MQMd9qwksVlgn+L1+PAYiwk4Sm3xSIaVTZxgRwTicmI4DncVS5KxRU0CAUmCbJXefhD7uT
giHorN8KiBCKptOS4Suqv4RPGLYA11TLVgTlBTLT2o1Z7EkxDFnn4jxzXFqzmngwqRg6tjT5CHyR
4LFPafp0GVQ/p9gDfAeeSxsbxu9cJZyJtVwL/zN3a9ACL8ATUR7+IPHeyNk+ULGgbNy3KbM5vKGB
D8r1W5kG2My+7UCoyanbodGX34PhzNppksoG9SFrYWtAfOJ+RvN2t1Alne3idoFC8fo59d4sGbVY
5UkeMXBJyRwn7y6XKlGiTyM6E7dKRVSg7fsujcYDtcsw5WKYY4EwO5a67sVK8U0Kykhkcrk8ZdM1
xEXoRNcaxnhGz7vuunZKpfuPJc+2PmJzNezZIRnUZxiYgOGSzLJ7NNQb5ZNsi6VZbl1q8NoZs1sJ
Sc4VyOrvLle8lhMbgBjo6/y2CQAu3D6t8gw961y64Tiu1J9BLhYWH2buj2o85OLqeIK7/Bylj16w
adp4LpP3GwwgN4BlofqtFTLm3YX+Vb7u4DpBdhFQe42CMZGh5rhbzsQ6XNTb5AqGkNXE3lqDpznm
rkfRt3kmggUajVXbS8e96ILjpFtTA9UDXMwrK8n2h1vSVQz3VCP1+gktgEonNossq73ddauXlCLV
AodMFJIXOVblbIi5MmcXXv/4QPP0GedwY60QvM3jKSANIOS4Pids4DaQbn82r0PFTbwZvU1RiU+x
4dkiLAzNmeltrJWskwaldZTh0Qi2nrKubDfwjndgi+TSNYA19DyHX6lyd3c25xdX/uCDAWZUK8lq
S0d+7q3vZ7/NUZ5DHrm4ZZoSVezxSbTm/dhNYq0SN0y7z+QU4queLPuHoWZuqyONJ+Y5yNs5uvpO
76Cx3g5YpYIHi4E0wDE8ZgUD1sXCj7cVe+U4RbOO8hii3J9Iu18tdhdv0bZ4xm8kT543Wfx/XkPF
3qnKhHtO3E6Ru9iS56G4az5E8uujq44YWpw+VdNRqYN6ut88rRjKLR6PZAL77suU3YaGe9hx0E4z
WYTcFpY0kKf+umrT0iuz05qahe+spEtOIwECVbjQa4a3VDMcm8kgSfvBMYMGvcr1xmKFOelECVHi
ErOks0cIzzCKeYhjDHZby1lZ6QZ5ru79WSCkRVKN74H1Lzl1ivtXKVifeW7H8pUBPiX5r1y7oBlY
XpmqE+9j+MWAdeOdoczrOT+59ByrcbWLaJKklLAnww0OIYJvjGfq4G/RZTmqBCUS6EJhLW13Tu9z
Z6/HYcFz2jmqIIoDILIBEcu0OWaLqvlfOEy9qiQL3gnTd2D09rETjJFLj0F86Woqbh1owovaQg4O
FB1HNagVoF3rjKhzYciPIWROB3Xo2ug3M/EOH1zda2JqiV/wy29/I7yorLJe7kdPKlWAeW05JYXn
kaWl8g4H1rTbJ7qViVh6yeywrsYn2YcxznCvcIv6rfe0Y9VK46/j+bWoMSgBKwfp+aRLhjlhBSY1
obIQ6DCAn6d0/KZmsFQuazpsyM9PwI8TxiBkg4zAF5Y4D6LDEa5PBzQiX0IroBdtWVEuCWVq5Vfg
vtZiykREFG3kLStQNY1iw5hpddh5tn4ReCFpJgTCpDurqQJo6zcCtBYfziCCwV4E8bFrtht18igA
AOLkdS8lBe7kT2k/sgQOeqGrxKITC+K3zJP5U4kuoYFjCM4USOST6AjFM0C3CXoaCiHg9d6sQNeo
HBOWIx8d9U6pIbW90tK89hHJ19x2ZWG57pN5XBTNvOzrpRrDhTlpJn/AYysHKqN8qoTC25wcKGZq
eSplPGrq0NDCchUAPP+5BJzQhdeW6CaKQpgnVTr2EmSA7S0apH9+mSMSnVAjv7NfsPbJB2lG5DAg
Hnwj4L0WWq472/QmmZlLTA+CQI9r5JoOEy/9xiYSJpj6u+bDJNsYIHDPjz6V9cBko3l8vt8tnFDh
ZXG5tRzlRPtqCGReKr6jpZQffqzQCxrfNqcS0jXskYoAvHGTXmddSXDYXhUNBhCBN9cQ6AtyIE9i
eA80rSKQSb7DmwfNOEx0WXTyin6YNaFhf+D0cTx+bA4yf37FF8oYk7dyphljrgO9H5QeXhlRnY1c
1slSRwtKKncp9bL+Y1LEd2G8I1Fad5+arT5EZFiCGGuA5R+4sB+ol5QPW7aWUjkQhZxYpaNzua0/
4DkF6UFSlXMwkdqAY+7es1JmPI5Y6syRvZQUM8XeXu7zS5K/cp2HwI3L6kd4AaltE0qCU9/tHfjd
/36PEpVg2g5A7EbxJwfx5uPwS7afXo05kF8+XjC62Dlt+fPpf+WIKhP5Tg6jZXjcwLmCNRVkz/RU
7/u2wKu/QoFYIEMhcj2WRu8kp2G9VtBlEm9VImbOoi/yaCOLXX6vCXnPHv73KtxIBOMPD43RTnIz
cxPRPCc3X0BkjuAwgRaXZeEawE6ENpU5OtrI15WfvKhaLdGLv4tWxjpOD4enBgmrjQ0K8WOfpD+c
4z9LxpE+rPzJ9dnso0lRiGWq7PxWsIsvaYhq6akG0r5fBB0rC/X/eAcIPoED0F2MKxzFPGdRh7Kx
uJtB3ugnoZE1E2v0lcZoTGjeSEit/d4/8+ZEn3HNE/DtDuxfmqGy5j+p308PMSBqgAmz9/oWpLFj
wYSUDQwgJ7E3yQd84LH+4STsrJeAwPU5QiHIdvGLz7yaP5x1qxqCSQQvL41rINUhoUN/Y9GAvV7x
ImZbAYJk5xmJsybkqGOZYBI25+BPGEDSdT+ge9QVn41gQ+e9s0i9FMdQEVGnBcaT/IH7d/5URvOM
LSQLEdzkmSWDagtNGfR3ydK3EuydmAKMaX3sFYqY9Ddd6/pBmRafl6oXXzsoEz3IlDn5AaY3pENh
j8aabnLYrb+ViRPAg66FLIDSXaJ7RWGvbfkaZWb2T3KMzdTbZCw5ZE0yCnGX19ihJJNnucgWfMVf
4vNds8I1qxgvJ8cS3dECwpYU+VRW+aX2o2nOAHCAIFb5+z7XnLmW0QlM57pgNwFavMZnntoZEq4M
J0lNhURPoDKVDnln+wyDqn+pyExuvoIiyXT72t+uld9ogZpnzR26vIoK9zKB2T889yx8ieL5KjMF
X+OoStJoWbJ57KsjjsbgSGIP53Z/RdZwVGdsx8nr7Blycdu/0fn4eibtt5aPwRtG9KinFbIDn0W2
8xHLWWAIat1KH3SJhLFsGue6ZwRGr3pYdlMd7kgnjxNJ4AyvgMVyfq7NhX1k+gKLZP9IcB2OBoHd
LpukRYaCqvxrzZxBFoBPc3mS0eS6Ld1BlLmr61nl4D5v8xBrK3NArirpPwJcNExPwpj5bhHK8vXG
x81zav5cAReuKOrzn+eeolvOsO+GZa2eqBQdz7VeLH+31O9Ibf+RfNGrqRcTJf9700B+mQDS5Hxa
PfJZirGszGl+yb55P0Vqk2ddH8auTEbS5q6ObNHGQAgM6eYbMmGw4s5udy1FCRdd36g1iC5Fm5Qk
HUzJPAk4IWIe+gJJetp8JjkhPVmNxbR29HyQwhe7zq5gL1WkY5x5/0+rnbe3RNSJV0UpK2KNU53e
6mDq4Qwglj7SCAGB6hApJ1mjg1VjQcgjDk0ReGnBLclR8nL9+w62y5fbr0F33YD2QoExoiLut4lB
Uq9njZ5LG8TbEvNpWesbB3E0pB0QfyF13i/L/3+BketKykHArtmbBEmbZwRLZD6yldES21wE/L/s
Mhrle5yBCqSD9xTVTZ5P1nUQ7tdZnf4YotiSMcehFPFDP7v9VYvMZVnJ6i7mrL8gDyR1HMpzdhBz
xtgzB0dIavzTA+QmN5hSCTdDB/ziWYGGcthx3zhUEWAYmrH1TUko+5+QukkK4DmIIZlnUUPwCbaC
hwydoKraW8ZZnB+SET57k0IN6B4/uQrKvQv6e9SsbxkjgWxyCt1BYKrp4MLtUboWtA/p1zGSnmcH
RjRHIizse+DZvL1eE7rOyIWPL2qKap9rojk2qNtr5Uf3hAiNG9LC5E0dD+rPwyxe+L2tQQ16Swv8
Nwe21x9lBZONWckUd5kmC7winG6wL+U53vL1jxn/y8vwA9YoKIpIZkqqy8h8BN+RrywlpCQCaE8n
C9OT5SuJp2E5IsjZW4NBBXQfsRXbVtAQsz0GtW64WF1g5leViOKHo47DUd/8XPKi/IsbE+qGDwhv
yU6fNVvaKbwq7+UvAqIfcXYIfcAayOBZmJPlO7cBM+Sn3txhtkaDHl7r596uIrvk4QyF8GG385tO
LwB/RUQwW0zgqx2nHHxLnQFqQwR3IFewf3RGLp4raN/A/0v5oECMJk1+aybz9nyjmEKdE1qb/DGy
b9Ed3XTm9VgPLsfuPMr4GuVaURPNFeHj30YarSnyYk0crTG7kMpJwDjydMg+Uj5Dv0TqHyPBPzFe
SVn+IoDFvS0PNzVJtGrmw9MeVTm69Vfyl5iIUPDlwIMxs0wpo1pGrP15WwUPh0/bbVPJT30OPf2Q
2ai2JspWUKpjGSqXuNJIQSaFqCchDKpKlTiNEjRhONlOt+USTsjgP0jqP57OyytM1uVqSRnZVgPF
t+oNysNmWk466CgqDx9s3LaZE5sbYf+wLYFysgyC1mNPwT5693mugT7SqChogy6VAV2UsavonPnJ
y/XwCj5dOflzOziIojZGpR/t65sFCOaD+rFql64djKC2RHT8fJqku5fW12jAFNz4PGlHzSfXwzUO
nlnBKuWXLeps9CyN6SrZqO+TXyljw/nHr4TXUe2g3b1VIh3VjjvxJiTWsnGW3o3lAF/Aa6wajtSK
s6VyKiJ4M6bAqnjMTQ6oufJe+KvGej1vt0IRFkJUpO+E7JRzKKIIIwzRatz/0sy6M+i9BXrOSyuq
e2GaxFcGikkBbSAgk27iptmM6yC+Sud6k9p9z7tJB3EvptoZEQNGA3tilRzbLzQckv6IVGNPosPJ
1d1WgKCvaQAdMMOZhdAtXFgfamnrob2bKNAg7b3MQ4jNKpVgtE5jsuX8HAoeNU76fzm5IVyjgvou
Qzh1NVn2tbPrXq1bX6bwcGHLjd2fmABE2i5401DtxWJ412h0YM41pZMjueU/yWfvMYw+GkGU0OzC
1+O5GCwUQAQcpXujqPh79HJdj4VX5Es9Nv0v97z/9ov+GQR9hD1gzQtMaDu67D7mUsn1FxcDlTyN
sJth8sFrrMYEyz7/Z8U1Qn6f8tKJA7bq3BFCIRIPgxfjTxXrqocdEyz/vJljcWmPOHI8DRtOECof
WCFFkTHxwVqDJdzyhWfRnF/4QKw6eqnQ+PogNm36EJLZFsAKBLdG9K5J9f8nXiNTpWd5xvzyTyW0
k1bBDiGbm7YbIQEHu7L/K/b3b3Fh47+KLC0g7d3nrrVWxOAGDM1nGrjiRHYJErHq3f8hE5wNeYOk
Yijo6F3wX8KPgEnP3uQEHkqvuPxsviI8wXdkk5SOsnSXSVav45zZ92SJo/ukV9lFKPdCsQJgGEuN
LVtrAJobyR0LaYDaNIh2CoPOcqpFOZ4juHnAejvtqdjf04pDzfQkyBQJrr0LVlweLxw8VXNcuiN8
sUvzBBVKQu3LRcKFPjAv8dG/u0uF3WJVvSC8/CkWVthttlZodUxFC1SCzIY9VAVddjdInmG5MYn9
pi3Xw6LPy53C0w6+gDgm5Mxaw0Q4cUkjTWKWCjoGs/XqjwRmaU/W8HwdIi0bJr4/KNOLfPDGgLL4
norz+D3XPv9U00gsfhH92Q7UEythFL0WcytYMfAtPwlXLXL6+oWDlbvTqe5ObNMQICOcS0SliFW0
YYTApQ7CP/ikfSgT/LdNqHaPzxqwQG23zaBVEdYeuWRla0N3M0ZA21+182K8tmmuBYlNiQvcimM5
Jh0CWw+vkvbu69dUNqUVaucCi4aU9ZUqlLAjQoMJjbCuO9g9s0aGPN6ycbRvEmGjlSyIO9iib7kV
zQ3sdMpYf08JNCbyGhDg62IY0AIF0+Pa4S8LqZ022ChjvIukVw/pmeXMpDMzM73nIkVi84Clqqdm
GMMQZ6togy97y06f6MQDs/QczAz4tr3dWygjT5cmLs2FXTJUjbUEmjcqDde+KnG6b110PBFhiNNL
cJlq9Ivuk4ozVv+ZF9i8LwtRqSHQdOmfktCK91j4/5Ki7YMnLgjOoDoFBhOY3nSgGvyzfvWFIije
But68r9QZgIlfIl2ITkYMLXFHHZbLThBH3BZ8b5rnqCh/GWjo9or20XTolEf7C9RBvlupa8yatUD
BDI/qKTo8BCaVybcBNK81ES88d4ietelE7bduDGlgUJPHPx0l7HXlGb8fh5sREVmlfWvlDF8h9v9
7ZqEQA5HdZn1oGXmBcvB75e27bCR+m3zdNkkfQitmUy2bIQUHylhTMNU+f8xrzLiq/lF0gEzTHxW
TeTewtRFMdRanI31fwcGH8XpEVUGpWlAZ+q7n6fW6u0z8P2rODQ6Wv4xZn8CLNwRXtn/ghHs3rw0
ckJ72ZLDGr9ck2mfRCqy3bTVdOCFHbyMGj5pHwV91QWghzDKMJCx0HPP8i0yqRlpTO2DWk8xfVk3
b8CKNh50UKhCGGReStd2YBBnk0qRZ8N5ItLM0Bulg87OWjzzcm8GKL8Fd3Pswdk7Yhd0lI5R8QBN
DTATLCvic2hblRXzOGLqUtQ9Gk0Y05mS2wW1tqn10u+ThaQ7hf9wzdjtqfwnoYhu326wyJ1+azy/
g3NxWh7NYdKKefeIw42XEIGnIeTJNKfCWhEct1v6BtXuwBiEiiNbVqyO3J3yWxhAwOe2T5TbXV+e
5Jhc54EwgHu6Jp2PPXaViX75gqTUfYzUg4NJIlLw7klJ38I9/MVg2mw+zyRfUdwrK5QuaJl/ro3T
+eGCLXcgVebx5OY/TuTzMFUwvtYlw3MNTNOHKq25NqlrOfZpk6susgEUT1vz7/SXCmzModeTcBsR
SwGiVuzf2j9bIyfWLdU6fuPRKuF76ggtILgK4gtsTSDnPx4gMZDnPvwul2NNVU3fCwzRYIPkbzaz
aw+kgDzB5NMGDsS+vSIXsZk8f1OtlYwNYAh4JdgVr8vJEba7ESN8LQDA/9NtG506luorKvqMe7jx
alcXZxQST9l4mXRSQG/emGFx71ZeI23mzKxXuyxQRLTCEowk4BW5vPlRb2uPE3qReuU2tCTz4hNS
17/lWYB0VN+UxF440qoj9P9UPgYj0i5EQid3atE2OKixqJPZkjXpeeMfkYbF/ojViPTG6A8496M1
N3FtoYojU19wWixDQ7fIJTbgJjnrtZ9iBaKPxSskdh9Fh+UyHMvG2ea74EtKsI/qKRC1nU9Tfyt9
cNkWTuGURFFrhaJZhjQdnrpNTqDcQbeYOwnwcIGl32a3e7V12lvakAV2tOP07gWghav2oJmNogXk
nLEsSl0NuzV5+n83rIMVAX5kM6ppedhVXEe/VEl/XgQrdfHgTNKYpM253SNkNBWgBKyJDCinEBQV
YpiZOVIclUIXsG/WLrqqkE50RFQZOml9zYWnWosE/S4Q4uzXN/+9Qf9F7J2zlvlFtFh2jtmO1WXz
94WX8qq8BKZlbVbPWkQPQd/y0hqfWNWb2T8HsGTcLM4S+T0GEoyTqff0KaD14Sx2rnzF7vsoWaPc
kSyvE9ovD0qTUzVkZJsj2nQFH5Z9RA0BF1XrISeClwKM42Q+8m889cDGWkUvUG8r45bVRzgmvvVJ
dDO750LAYDb3P297yNhiDyc9xjgRGXLrdNLX3mcDvULR7LwXZgugVvjzxRav7KzHS3nN2xy5f/UP
uleRI5Tgj85IGzOq0FM9HMcqmF+ihFPPDZw/yasD9UnDFJQmWPcmJC7oxSPJq1Rw4YL32mzbeza3
JiD1mfZMUOml3Afb5lYJ3z9Ge3Lx48AsUo1Mu3riAhgPdJ/ofjP7fSAVeN0fbgvWSYJi3pUI8Yxh
YNSE5tyHmIUMn8hpah0/GVzey7RWwNMsImsrANrxTLxx6BHmS6kLYgn/vOI86HbNaypRePIo5FcJ
en6FdoTFxrgSzwddlEERSsZxlX39NcPN1OnDouQQFZo7wEM0Xm+TwMDofyDUj960IifWKqL0+Y7F
vZDXrMPC994AeJrE0VVTus6Chhl+ztxRUJuJrj++laFo258+RIP9pU6u0NlP7sSZH4ZWsnLxaOSn
mdAz2qnAIoZ7q28+oKV196OvcXrYIWiUtlVpDJpmQQxF8YsbCKv57AiB8WRwcbdQSuFbJCT7Qwnc
3nQQ6qF2l57BH9KdJiui5hNd1abMxTiKPv//Bd3MSA7FJJeLxrw115OYbRePQF0XtcwFLTY+SJ3Y
0py5BLq8VNOomeTOmVtBqa4nswPFRLGtDVjBNSJrKsL2UFxqcsssRMar3edtTKIhzGqrax0X9g5w
lGtgMX1mtLzCUMWAuIEzcB/XFzKkxwGNvpTlew03Ofz1ZRcXD89JizneWOsRI5Lf9PkvJNblRHxw
v58icZMhOjnFHNwCxqz5FEe6yVY/OL+eFiIoQyobW93mIjF3GuCG63BrRMxKXCbU1zOASlJAPR1y
iaWoiwd0y7yOLjLhh4Rl3lPvOnzHGSxAVsbqq4K43NLO1xDceo8hwCOVDSvicow91uDvk0ble98R
PG3TzDHUQUnuTqKSV7KvcHpxZiAGTqsmmz0P/1r3Lmz8Cp+tXIEg7zuciaE+8fgPcTeywSVNxgMi
OIqPg7ckAxPNLltMAPY6i1UicIiHbfg/VusbD81Hw685UIbuL6iOkCGC8WN0LAMOrnkeG5bnTvHf
flIf/XUGAUTQAnt6QNr3ih+QGXobhNzBLlKxUj+Eh2jtPw7ZXBAFiaBpxmJ2h4E8J4D9u+nbZnvQ
kbM+Sbwd09eT9pncRCV9ivkcGgs1bioyj+NNkcaZOA8tWxKfbLNSfHcWjUW4CrAkjgldPJgklan0
4A+IezW/VmVOHpgr3i8HSJnmUzYiJtsH9/WrdADOT0lx5J0jhX2MNHZLiykq0mDkps02G2rWGI6H
ws/qwlarz/5b2wfpSVwvpPJPz/+e+Qzby0GoOLeoGZmg+WJdUlvDrzeKn8V0v7q+5XzulwAaY01t
jsIGMHt+vBQ1e2ybD+PJhv+wZBS9xYuNRX6sNzhW4a4LLbOHArRuW6VBVOGVQsP/tbUbfkjedzG9
BI/LEiZUOdFMZeuQLJ44bYytjEfLGfOgcNpGz6IX/HI8wsLBKoUp5F5yeqEl57CMso0d53oLYno9
ZKKk/xQCmp/bVii+ZbjXqDj8aas6aubjgarLeNo3E/1Vh3ouXy849SdgGVYi4vvuK7xboOp3+zGa
fUZaXK4rg8XZMAG1zw9o4em10GjJLMK/XUuZzRxjhkYu6wqT2/thijfL3Q0hFZFKYmqPcXkcGhBK
vslikS3rfd+Iv7j78872JViCn+k13sZtzwEpAlcmp+k1njUqAi3Ge6XPEyDjoWs+JSIjyqqvxhO0
BrzBXtHgCZ5GH0ZA/dAaunyrGWmENb1obHapf73ThdaUy62zx55EsijHoViAhxncdRLRtiWJvmyT
Cp30WyfbrOILFGImXpH20FXM+SvCI9YkPrWGZY/lGq7xzoqne2Y0FR2dQRWnL1pdDKLatEWBZpPu
+towcMEJC/fkpLdR4Xv7KCbBlqsUcyHMFDOdzJWHz3repEW+5UDISMzlPY7flIpLuhgkMN6nxqiZ
wq5HDY7sVOiCebAAC3n1hn9lsi3gF+A47x/C7hPUq+4UmaeOZ8UlcIHoOVJWYisgOnt0bA9xub3H
NoUUNeAyDDJqm4jKWlw6/EtuVOiramOXlefDgHZ62AUeRg7sgwRrIkDqDWePFlypwRQ3k41dD1m7
K8CfthPCYwWcrH7m3uwefyZO5AmtIlpD4XXH0eVn/3A26ggeFHVkvY6fC9V6C9rJ930kADu7QKBv
FlEy+5ZZ/a+sPLP65YiyquNr5NUHxg8D58hW5wL6ZOw0LPw7VCR+WO/ekFKKtizQd5MSZZ8gRBj/
HncfiSevrtHu5k2olHepknoOOEcCkjjki4oek5zNVSX1pmZgCWfpB8p0sKmXUNm9PItITD6Cu037
M3TeXE43uIRvRVgShP+3inSZEUQudZE5Mcd8qLo8gPviT0cMUMwgHPN8iaaF3QKw7nx99Dxs4K41
hCvGXWy2RZ06uoYej/FuYSSaScbDdGahD6ni5vOKRO7q+XGD7vWOOhnXvVwnmN5+RC20EyBKgm7o
YIx/d9GXBXHEE3+rwO44txrFjttoi4qwHaiFdXZ3VIF3WibOC6WzmLPSEZwmcua3+F7asa7Nwh7t
OOQQABCp/EyoOoQqP9rz3lGJsGUMevALthpD3HKW1248VN/z/ANiFJ18dKaqUvTkJahDqhBGw1Iz
AczXdtzzIkmU2Npuk3pucbRSx14r6a7lQ3MrxZJ+QKrdH/Ow87GQcpO8i6Pr7W4DdlyxOsikAY4V
1aM+fOOENLN+8PXYIhotLT18Tt4INCyOTBltsPLg4r8aQR415PJpegbPPDDd0RS4sVfWMlygbABS
xBVBwAu4zQIVWOLXMK54/v0c9XKI9Y8Xd/RdAkgmWM4tffZnc2qD7xnKCe3BYYagwAvEHi4g1Vyw
ZJQ03HiH4VkuMuQWIj36zNVD1OlO56j4MlwU+ahogTHkWqn6P/xNTB/d8zge4f8lBXn3nOF3/z1q
0q81bBvCxQnPKJYTE59wHn3aksIWUv6kuoZwHV2MNIFYolBVYsZD4Xggkq3v5sVQaRRS/P6JVTyd
oO5jzsdxubBsKfouYE20ylic2dS5rzba1LgLCue40+WeiGps/NvcmrLYdfg/fHz56Sds82t8RtPs
oqJGfzFHzK6AthiwJG6+fc7Q0KbVEujGK2A7F25iODNJy+JJ7UCn9AjZ2mrISD7t8g+EvNkRp8nR
nA8MbPCl3kV6uBK1IlSQmbO3aJKolTKU1pGAwK4vh2jgY7czwoRQoTs6dr1G922Mx/W0dW3RtTzQ
xBxic0lJu0SfZYzgtO5oDphKeO5OnrEsSj3YafSXcH95+BP4ixxPsAIFk0KSWl3NbEVt311b0ewC
Lizwg3ADWWmTnPXaDekY77J13dg21XYNwNxneGnwyJ9MuzrLw0dOemcty1KDHzAoNAy0xgUAqiHC
WTq74uvUautENuBc75IRBCwazUL1QVdZ2XtMUjKCLjSYCL2A9Z9sRA6cteLan/gvl66P1m8omzJa
jvYq4szfvy87MYBS8Mv0fyy55oGgEkhVdnFovvhdyju65wVH3L8OTd5jesqW86JAZmcVyTbwDEVp
u1zA6SCFgdhyniq2u29uqQvj4zoSV28uCoFCHypEldwVTznM0d+KPLtXXHsZDYcRqGdyJcqe/Odu
AdMhmcKl8CI8GunGGiuic8xCxtH8iRovX5CZXZTz9uqye2IH7XzlQ5KEb61UrXaEQ8Vfngc9mB9C
eDgkUhB2dTd4B00jUUUJ1rYjnrHjKcD0d2dGLaTp2v5/QGEYvx5/o1YvYsCuBF7QDSES4qgZC2qI
3mviGza1FgnsDeTEsqHtwLxSkdgLBWCR8LkI/dSwdRGMGUC9VzEU2GuzBPx3owXlTBbJHwcBwWSI
1moOz/mVoI9kd4dQ92iKwe9S4Q1eV7KI9dZubhJbdJaPSvxh61xF56jcp2GHZuMNeBBHelOzhNBO
i22ZnKfo49u25XFl0kBXcwBBPw6w5hbdW/gfuAbmaTsR+WpBKAmYd1mSrDmiJB9NIDtsq6XC6fz9
Ewv7jNjjdXuCsoYzhQBnd8bZaiur5/xcLUiwNL631PyFtyyrP96CWqJVgMAWg8wp/yaz3lNfLXXs
1AQkqMGe6NVF72A5/83M0CZ9WCr7N85Fe3HeifqoAL/KgSxH45dPfzKNjfaJmaEOoAG8Jei9RtSn
OUMALmI/NB6+w/tfdWWcYAUSPvdn5GncjVQmT3ROvKUb9vHgRCvI686NntxeyZYUB0GeKS2iOu8w
WmYb2ntsI37FIZaIx9QBeCPes41L+xyQBX23N54IzTcJq+24NLp6ZoFoXh27U2vlQqy6u37PT+XE
EEAyxqnpm3IkRexcHF5oOmalowIY9twBzPg4tXgQU+VHz0hMZNc0TDzjpLKbupBH8x1QswxVqP33
peGa9gK5XhY3N3xQ0ZTts1TLYPniqpi6WSMQm/vRBNftn9mIT0klGhOXgXzLAWjY+YDMlNXLmpAK
NPV/9MZi6+qImgFT0PTqKGtOhpyHFYcw3YoRjwHpDjYUeRsNPklT0F0r9Qw/ScBJlm4KXw/Mz8e2
sAGpH7CgjR6w5A1xwhCYB7tf38vsZXqP7JAR+bPqE/PSTeBLTLl2WasduNUx7v0milQHooPZJ5JW
6ut8xjz6FtohweNRa4gLMTAs/0XWrdmsGzgHK4eTX/pFH1eO5DZj9baj4FqHSpPayOBCKtm/g2Wj
CXpG4u8CZvMef18HuQm+/WpVeLS97tyEYrBecj/oCIQxdFnQw2JPyacFVqv/dhRhIIxonb4b4l0u
/0SyeZ7CK0OVrnvXUkcCeglEQEZqVEVbrtDQ5g24zYyuL9+vz8y2kYRy9QI3yx7zN8bOl+yg+esg
ouISPST/Zp0Vqp6keCCtNGsySHymAeh+x4AOja9uwlxpzQ2NOVVjglTGoUtkkqJSDaCVChT9kdaI
XKOIUnTGyH7V8Qqr7qHyH534P7B6dQexmpq19KNS5e12Dt0yoU0JDtID62tZeU1uXNo17mNNB9ov
EZ+HqU9Tz+dc/gXpeT/tO+Rp668KS70Z8yUVGwcWBR0RXzhh93pJtajPN2WKaKQPKBetJkyg+CNE
PPSgwH2wBS77kkZA8ipJABuMBX3TBv1RjzsRUAY2EmwEuaLpP13avo3WLiH7NLh2xGkNais992qQ
48SbfiE8SuOvRg+g0/k3ucrKFqTpwyxfhtpivFfEnd1mguWxDe/ByL+RuO8CgBAo80IN/SQKYTmR
AYF/Zv3ftIXS2ur/CF9svvzmetXSvhqyyEI6slMBkh4dyRCpjB0g82UaXbcZd+sWsJOsskvqXA2W
fqvCuC5hQsbpHifye9xxifH5hQzQzdFm+L46yaIUj75FZkXqE3+DpP0R6Agk6iVqVTf/r7SyZCHH
CNLHS7ZTT5VcpjsViZUN9nKYnzJ/4TJSNUKPEe5rt0jBFj8/7Kg6ADeUZYBq567Ma4ALOs7yz3dN
BlEwPfNCy/NDINNf3DnZJE8tzdh147VC3Mtmk7URwSijUsWTtzfVM83on0B9md9+U5lbePUthFjw
bS1aNx1pH9dKz+uf0GM76UpNAXsYagL3lc/zFscNwPd2nzKm5y/JQWDhkFJpbmHPfjOto8zh1HCs
aeT1NH/iEOVk3tsqYwms1hPaOT2v1mG3bcHSBapL9u0QbV6a2Iy4JNie4Mu/AlsKdEKG1qNuWYjj
rfDMnQu/7xkUbl4ysi3YvvCpeEqSy9p9lCT+hNSQ2gVO1FSwx1g+0YdtuyoNQs5/rffkZ3+GSM5h
WgdhDH3YY0h5irDa6OMzTZUkE+pn22NNt+8vkqS/BFKk3cMjFsCo8X4xYrPLMw3h3pWAsZrjSP7H
1tEbqnCwJJd45FP47CeKeWmwkGg8yP6o4gA0qtrAD3SRVpVQsGNnQgkQ6onKm+uke9rWg4cwj2G/
taUdHItaN2hcEnXjmZtwqg3uY9pewpiFvCgZZVJxGacrZevhi6tIKnu5ILwe2yVGBwt3V+syGrFC
JR5FeKRKO7Lmecu8AVBmgwrTNOS6jFg6OnvOv6jvu3bbKV3tlA8ClNKw89y6R97nSV8qCrWQhhwG
uJDDxezlHbHtIykVBpoZa/F5RffNEx/BwWazZdyb/aq31gbNFljKO9hJKxFT0lT0GCwgXxtOc0B2
z9iTg9iG6GsswIwMx+whC7hYocrxPqST2mSHMlrc6KfDCjv53Bv7xrbDf1GYQLmV8vzbDtGFwi5I
bNRiFTDLUcjqqT3dsPomgwoAM+Jinj3a6u6isNcsA3lcy3WBf8PltXI54fEg10xiGnvSeM5gBkq/
E5GowNZgGy8KbyCnwE4QmGynmFefGlylmjjpdUjrT6GBxb5Ztn+Q0LxTIU2CrGgSNsO73IdCcuSI
dCbHVW/AvpzklbUtXFHBXOH+LfNO4OELx2y8iBf7yuF3wZBj4o80g5+ZlP62mMMfhYlb9BEFEkYQ
o9fxMqcp6eykQScGZJ9svHraBr+yBFyxXcJ3iBp4N0JWBxrIGXdy7a63jgcMuxYZklFsVapkhbyO
/p4DgW0Da78pRv0ynoPq0k3A9BsQcRSioKPziEZ+yStKeJtCoC1+EZYzkqzJzZh/PLfqNy/srYZS
SXBlpJY225D7cCSq0DN6frElgTp8VuG+qfKrc8dZA8OT70wrq9Lajx+NICjkCGqKQ0Xy8TKqn2Ad
LIm4mwEVb7R8JBB37CadRuAVf0RsHtws7jCgMYuIFo+LcFVcuiHQ7khlxNWh0gjMy3RLPIDYiovT
+Qir4iCIjF4heQamrGO/vCTKCduPqZkyJ5PrHSU5fUR+Gw5D4iTheArzhclYzWfOb/u5fKb1/Isq
+yndL+ryUhZ9D4Wtf/l2KhDcXbGumE4KxOcK114xRCq6y9nAT7aJVI3GIZxFd62M1Sj0dUayxQC7
xGfLoVyyXW7udUkkwl7IeOhkfwhG1gozQN9iYT1KRCGYgBPmjuVlQyXU94hsZi+Gdu11bLGjPE3D
JRqQqWWstm80SS9x70I/hMJzQklf9Gv58PiEtzp6HGh4Jmbkq0sSoULDEXlP68ejGUoFBtETG9ZR
wyVLTv3C4pHNw0B/sYCoLhpPof7/3cVliY8q38sOexCXOkNLT25VdAgU5aJ58atGsEvqDOce/YdU
CUV6ckQeMcXpuVLzSogjQos8s9PxVmBcucqUm1gv9XcbpTPEyL5lcV3F7ucMwO0El+PjqH6NHTW5
dofzE+ELzkRrD/KyLaKoU8Ap1Jv0TSgY0v8aTWiSIZTzXrOZb/FPe0SMpcR26NPaF8u7oqyEJHB/
PsBkVa+M0KiZFN4zTJ91ENb/SYHHOMrFQWyEBZhvx7mm1v3lvLIwIgEaqMdAGMl/2TXfCh+ccF6Z
hgFjOrwTrbA0E0GO68LP2tFFGFKiDfsX1m0YoPrnPIDuO4UmGEloUm9Q9SfJp1np7bb6ucL4Ur/Z
PaST8jP8c5HOCSKtN0voGEmOurGahckcXrhzNosGEQIrP3JADp+GAUX6PJk+7RxuLuZwnv2y5+F8
G3ffDnuBPn9vZiwyrkt+pK743Cc6Jdbr64eiV9ShMquzpC9Am0gHUOGpWPwiY/KDDjbRxbiQnj4L
qmPvxnkUPOJY4pOpaDAmLossvt8v0c7d9SeJxwLmINQVxwRJ8gDAAeKdRW/URvbP5JU4qaZe/YN4
qbw9ZGSTOAUCwNj9jl28kZZVzY9595Up1GXOuEZ+MtGaMAHIC2E2ywhRS8nq+Td9EGgpcUPBPenC
Jzd9GQ7lg7yy65eQByB9BpkdWqj5tdUS9ecpvDgA4HkAppIt2o+76PxBzcH4Y+U8pbraPajL/3PL
JS/eYoIwx8TXqdTUix4pyJ39AcZIqXBfLrY2/0qvv46SNXGrMYTOvFhyxDWoKzM4wlKptATOVMpf
AbytxC8Hx9CeKYtzELBSKSj4NVU+Q3lW9fzKVAy34n2hc2Bb1pdaEA/sLS1TEjri4zm5Kdxntv7i
Uik9pr/0XLuT+8FKGo5MilihivKnABpm/VLS3LAVP+D8QjacFwJdpD+Xv9dkcAiBrAPaCQdN5Y4g
tFB/cwsdsBPYKxDUaX6yiytATm+W0rMiztY5yJ1H2Rda2cyloLnGIC6YaCQXgwDHFVceZXVO1qLU
9HtClwjb5NhoseuVIaph5F8u0Wijw8WBo+HMyO//2DmJIX8wC0Ge552G+lEKALID+LNMF7X8kBu3
rbmUlQ43fWwSbAkUQBZDkvGKy+pjGiNCJngBUfnC5c3X9iVoHDyUoEpQTjTlWRg61dBffkIhAJwy
K06g68ZT4/C1LE/sny/0n/6m8zSOXaNdJlky8pq5Mbj9k7ggHfDnn0AJE7kNC1oxeBYin7HFXvHr
8jtMUTeGZgeMOhPNHmPfXzvRMmoitLnHVi2Mc6MVu+ZuNl0XmMXJOfhIc6Z9bQrqajuNIsXXnrXr
8i9HJW0hFEn+2OHFUaRbBKG5uY+jyTyPYnf/laYxKC3ZisKAThRrw03X44xMPp3ywvFtkgqL29WZ
nnTb9rF4su1oGFtTuY3e1cupaL4I9LSnmtyYQLVOtPDt6D0RKun3p+QKQkDp0N3MwIhhM2uH8ghr
Si7mrcAc5YBQEMxd9hLMpo0nQmWW+ZHBQprnVfTSZrs1N/5jmAvjACWIWVjzW04PVM0nFU84dzP+
ZMru7RjVwU/zkbxQLCQSbdxcEw8XOP6YojhQeghzCIQBvu+MhWtnEpiDrCZqv2fXWN7g29MDp97b
Ca2vixojtG61nvIwnf3f9kzMivoHu6K3FX/JaY4YDOuM97DYb+uC2PZwXtLo2HSX5YF2LeVc+WlP
N0ox3g4A1kS7zfN0RbhlBDqbY5FMK1C1RK+YNhnsou7NOSYB81ByYRy5+S76uT5uQo5lVIfoJXYc
lPL0CPOMWYm2+IaTgPSa5k3IQK1gBqBUneqBPLNKdtv4X08t/qkBbFw9RUnqwpGtufDWU0PXFAju
9TZdeycUrOG/h/o54yw9kkrS/HQdbE/F8QbSAfKf9gTzSZ/SiED981UA7nElqC3xktkF0G9ESv1y
0pG7vC6VPFC5DbNMmZhF4vbvR+xYVsWBxdKeCNbwtbSpdxKpbFJvnD7hRpnzvv0Im6TBJxvkRX2h
dqozGKr/jp1G6+GxIJxAhr3D/WdPSlQFObXnyTM1dOo4k9qTnSTx+NOovdL4W6PGTBI2m4b06VU+
HrUyaBRmu/KdY3tXjGxtzL4hEYVukdt2TuIdkhR98vk9xORypZbGeE6owRHF6lc1nfoP0y5D81fm
+e+GpnBZwXE0Vn9Gr6VcOyLnOTa+hcJbnZCZkqvg5rwvu37JMuKCQtlpwTS1/suSCkox+rzsRikO
v9zMFwUqtiwaCbI0UeeoZjS9Flmc9HrAITEMrBEqUtFWRgshTWv06/opJEpOFqxGpVOJEQCymu39
jMyA0RWCqt2VGdvOBMer0Pb4HV1psC1hKjGgCPbwGOBVEmRuhcEfPnmQHFf8FF3+iFuayB3sNAFs
dsik4hhA7dEwhY+x5Ed8WuqKa6H9PhDQ/43iYL7S1Y7+nxiqgrKBnAdjyb1f7c/K2vu7EAoKkSuR
51L9ZEwaTQwv6AeaMh6Mnu5zxaErcZGyDXnrvLgNwdCFGAY7kD5nTAjOwWmMRKuTCw7qfMD19cjk
2nV72iLiUEemHethiysKCzx7333Ub4SuHerpJbxlXdKmG2YvTS0FhIU1UMJuiiKKDXSeunF38uio
o/QKyBAPPAE6mxoElEYAoXeTZlwm3ifhrhkoP1RCRgpyKbZ5rgzbOuOml9QyRVJd3jv5mVkyTu3L
FbU8XM7cOrakqrGsYpzjcvuBi6EZxkfhWk4LGrxaozeCDI85M2wddJQkJq9fUfgk1+DYfFDvVmKg
UU2mWZL+PlQMJi4aa9Ekr2FiLOLmeMFjJenZ9rXJwr3Tu1KI0LFJvkRD5k178eqJjF//XlidC4G6
5yREvNmSWOEoLvYqKuZWFpdu3emzegASmUG+TG/PTDeAjtfR3PxIZHJ+Z8YNTM3ZkdDQ+D0Y9qnW
/Rf8AyV2h7Q34hTO5SZzVE14ZkXDNzX91IeilfVWOWN8HcVqZfqLY4iWgYMBGkQCd7rbI54Ovk6p
tUC0EwuYetVtYB1Q18U8OCf4UOKcSzDY3e5pLnAaaP2aP1fp0IHhOqX0shm/an4XFB5quLliHXC6
BJgqEjJccbOFfCg6M9hvDrXb5MqlhZFq86MdQek20p/HQOqLPd7GY+Cokkv03+lfGvb1RcwCFI2e
bsnCYFrbJBCEdpchBUBujOjXCnvYJ/DsVoXnHa77kN6WOA4L6YN/r3o3Uh69aEWX4USsJXleVdbp
ksU4qVVqpDFWenJrYX/01+evEIpzEo7GAC2yw1KN9vDRO9Fykpey/UfmOfrlnRKxL8my1tYg8OIM
foer9/TQ6FMd+qDRlhHKNX5qES9zjIZ8P6hf47XX4UYCHlMpdzvtWkMUN1peJmY0+qRc9tMzmuaR
wKQqJYzSaGioFjOvAGde3NEh2w9y0XFs7c43IWboppabyQ9ZN/V36r7jQ8yEuU8gXE9+/X89A6z2
ZPeRB0peSB/Gs1YAWkctdTu5oL9LcQ/lD9+Uxs87HBOQw8mlSKaKlc5n30zFGfCHPxr9bs3HNngo
fvtRsjLoD3yDu3guh4HjMhIxu+qtMevT+2EkwzKM5A/kO32ktt4+CcqyKTrCE+jTZ+CkGmFGmq1R
BssUmQD6nSorTs/dMF/NNz0yObLYztphxCXMYM9FlyxvQ8b0KmkTN5LVLLsDgg1UUcgA8311od6i
m1sSDkG5Jtv9gj4rgc/vd/OM4D4wTWapTbmlZzl9TTvj1qUZk6atH6ZwrJXomqyplP8D3Eqmu+kZ
HF4r43Z8cIJvRzBUMI6fGWPZrt0IXXeFPX/cCggodQbH/PYbTaO0W6/8ofik3r4fe4hzttMRxIUv
tppGO4Tv0lGStLJAiKZEmTWemtIE+LUzrSoL6bD0cbeGeyQzPtR28uIBgFd75OnIpjZjfuVpWL8J
wGpaPtbtbW7Hu/0DzkFYNQnX0ZP3RWP1nlhMFeyeag7YIgB2DmQo/SbderTtmU/udoVOOYpcoEp0
g9RFJJjOvicT9I+3wh1MUQzLY35CLFC0ekUcnrvZVTcdTjRjPKY0cqZw8b01fw1W+75wB12YTFNF
Vbu5jAP1GgNrzMUZSWIn3Soq7ATrt8dsKPNRp8aSFRxPGAuYP0Lq5q+Z0usq4weXkZupr8Oo1Z/0
A6YJ5jy3eW5GfeckXShPfwaYAiaM/LR/2w7h4f4hJtNo7tQA5G4WeTSO6Z2ta4hDxsppkR5/HHS4
BLRGAxj8OEAhsTLWxlDDNE+8OcjHgC8whTVU6fPGGSXBsYsyElWzL5OJ+7uT8MRr3vg2itNNTIdA
G2XD6/QlrTwnLKBjRTdLRIRmsnwDQuUOiLtjzp1aKAhUuKaibyUu+Pv8yEHYuNkdQWeSFIcRaAxg
6LgboinmTpJBE5brA+gdpQBTHDIcU7l9CRSzpYAvgMwcWxEaXW4WN83ErZ0JuWhEJVyEmGISBh3e
o0KZIWNvD3IBbjuGXJbm9ftkynBufWyxNDVpJB/AMod5154/qcTff5DNc0pmWCK0WGwq/+BvS/x0
l/kjSLu7AXTLc2pk8koAd2AMRJJoi9TvsNQm0ajTvckhqUeSvlY9XHZL8W7jhzkMr/jkDIQktdSt
P552ENrpPLexNUEl0FWRDFbe6PP+Fi6VrI0nsTUfXIMadDFpQGhzIgLH1L7Lj90/la+BUKyB386d
9DeFmBuYEsTKoG6oYZN5x4F9Jigisv8MGlawenrO79TwEB5bJMw5S+HH/CAfAJt4FAcGyxNsTFlD
ZUJWoH96/trckHMeN5NymZtEEkAKiRz24ENQO3LgvbFnKKHAuYpbJSMiGLsMEE/PfYE32d4d3QQz
fa2GaVh8lvTbHoX98vEsyEVRsNluh2RvA/EjTL00hXfM2e2KT2IiY17qOi90YA88Rq51JhjqOb8/
Bjd4ckL+5eob9sN1jgHwMhKfc07PD7Aai0etv+vrSr4S70IMcoXgBSZYtoSilZHaZu1GGv4SGM4W
D+rdjYcqJ/7VNWNLfuwb5a5y8QtwyVP2XY3hBkRxnCkPO/UCaW3myV6pH4h4gaWS8bD4uH49RhTG
1rzObBOWVh7c3N6pbxEkXo5tbAeXXecyXCxjZCR49OSk7pTz5bk1cLDSfwKCdneojhWy0NGkfXsw
A3Xsi6/NyGfNFAiHKj3vYGzy9RC5/S2nQP9MkFSqt2ZN9+tTUcB0CXEB8Db4ts+ilpnBySlVsJ/+
MFVqL+kPUiLQfhnLllTdsCdaSo1yU/EhJ6l8HMM+5lh473t5q3foCyJv/Aw8zfCXmwpZvPqvAvTH
IrKwC7bWcKKfSjyzmm/GxzN9aYlLkHThYgrZ1iqgmO5VbXF5Iyx0lYqgFf8JjWB+7QMCEqrdTM/t
GREA1RD2Zbh+f0YBoqmEj7cz4fZG25KCJXKazPkufz1JkPov2BlENcbMg3UvB3WnIgrSHUKg4ahc
6kGuwtQJOClCvTbo4mhxDnnVIQqH2VMGG3VsgCm8NNkS2O+CxkDEdM5XNKrii4CV7lQmY/pbIdXQ
Dg6CqK8kkqxA+RnfAIVzOG0EI3P8QVz+ft2AlHolOZ7TBxOCOM7jLzX5wM7ZQR70UfsMwhAypVxL
jFQ7odIHcrRyrH4KT4vHgJCIrcxLZpdyTDvV5Qkk9rjvye/qk8/nCRgAZnknWFdCxVr65u2a9dR6
JQvyJEgK1PrMBHvI5Ha/kGTv235KiKo7fsEv+9NCMJVAFSETK4J9RPUabaW9Y1Ooz5HgCh4HOB+y
C3zHkYeg+y/5Af/rSdOP1+OouLZokw8AA6pxL524dwgmF/E1/UQQck9/oQet+frJrJbmpsRzELCU
p96CkreLMp700FFRI53QpWDYARO148MVg2zR30Cg2AEDIUb19FybZUkZve/85r5dCTiH2N98b26I
xI3n6BXGI6pDJVn4q+eFC0FimJhyW92jXLwFb07umFEjzDKTyHTCHAqWI28rEuxSG4gUSi3AdUGv
9l3+2IGReUdKYzqtYRF9iP259S2KtsvmjZ9XQaUrKT+Jz5Bl7GsVVjDGAAQe0/Uf6pvLfBufOXZ3
7OAxQQaCMj4U5f1HSjg4m+WCbT1GEIOwPmR23KwxxzS+Uv07ChENqbbGFQ1O3rOFfFqGM8Ul64VP
8etEZV5QCq7mF905XP5pLDgWgkQh7a4gbPJ9NEAMExg0j1OaVoeQn1XI4WA4+MIEyV04ElwhYU1R
d/oSr+9VueSEx8Jiz1k6Zx8kkZY83wmoCZw+UMrO7mg8kTzxi1KpufOOFChUqgUuW76mPbbLpmOF
ts7WLN8iVKLAw7LJn2yNR9u1EeFPxr0Rry22/j8+dl8XhmYYkRCNW4DVoTtk+ThbaP0QbGv33e7F
DAUJmcBzBXvswcDO4Mygma+3rJpI2Ypp28Q0c2DxgUYSDPp+7Dmdr/jxdyC0gX0u1Vw2k+r5B80T
Pyh8fxjtr2j7tU1BWDpnYfAtqZyePyM8HACK7cOoTESRnLUvCYHNk0YgCbJv9Ox6o0HbxagBbh2W
fQX3Sgfax8DeiKR9s5qnHR7agkAx/oKY+vhH4mVjO6VX15TaeNgkpWq/3dQY+dXJuFUV58KRi/j2
Qxbm8JNI24oGwB7KnRQr5YY4smbMeEvgCHtCKT6FhGMaK0apdwt3whLofeiL7N4XVDo4N/PeseYl
MCY/Gqnt+3QO2OE4h2q3IYgWDAyxdBbMKgQdkkI6oPRB49E6QjcW7GOhlNfpJQGBV4OxLosKAKc5
hNE6HqdJTjlilTyienqUKdw+GXRmUBk/n9J/EwUW+h6O8Ptfraw2K4EUKRyHZbKcv4EaFYL2SwiA
jM5q1+ddNFrLurVjvP762q2yAXqBYPEReGTqZIwyjjEvENLfOLVEVFHGattVo1HCdYN4phjN7L1f
jrM2NvrkzdEI/qY1qRNlrUxZSyRPxP3R+1v2QpeITOU9/Vojt4GwBPanTFMA+upYBqkooXHPAFxF
i7umcDpF0exk6ov639IGABSzreLLXMCayKZTiF7g2hyemwP8xa6iosnGZDV6A80MGpBXaDN4MzoJ
hBA/BQUGkPSi/Moc84cBe8o/Nb0CZbwZHXHL9wj9qJsZj9oTTYGZRFGOPiTlRGLdNsoeXriq4Ifi
Yp7YtV5Mrj6iwNDcmKyhYyyLefcU5achHrpKVWVgofy9ccETGyKJ3yrU4Cxbz+ZJwu+Vhu7nIBJQ
xHWxNqU+j3ZaliI7JVbl7HPA0u1wVGy/MdJeP0gdGDABHar69scJ9IfT4Kj/PBsGOA3XUq18aeLm
aKBB7Xk86ZNswUxBRgBDBCnnaZIzCaWJu5JpetIF8ybpjTgtoXMyyn2/Y+9l9hDf8Yzb9bUAl20R
lrP73oAOIFHgKka0tPn5bp7tjFzsgCBnpgtogpaVe72cSeI+BvDglmQI182V7sFJ7gVmFiaQSP+J
Jf7FFiSw1yDOIdJCJYpazOpKokwOokU7RxxzU3yopm0126HxoApjXiuMJj6maogsTKEYyBRkZ7G/
DkhXMdCzrg6c2G5/OAwnSwmJJo+TU/5Hoh/owHIrRKfi+feMUdonmK1kiwHexqmaEUylfaJfTm9I
BFGJIGd20Hp4XtjvfnJdXX7oyr8CgtdoZwR6PTQlrQxvoMManmFx80PHiUJpVNyUOJecQeUIOpQo
mHdfn/FHJVrGPtfgPi8Sdd/kso6Nbzc0YHCggkpccSRfp9lFJKuv/4EYwtFQsiuS8uAKB6dPDoQx
qHj764sB9AdMB0uHfEe9xztTpTbrmyvomjslPezqAfOf9gDzkPgORQo4iFCZgwPDDEhsuJgTokeg
4FZUno4+GyPkV/suijE4dM2X3hngBJSKBe+6Rtt+68UtjPcA9ekDWYu2OZ1lAUE0a9aBHsAR+xmi
v+DcdDgmNB1I3hJijXMNVPrO8Rf406xogKvuZx5GZ5tqzZvEGmtUB9EIFQqXuy5E6rIhfvot4T0n
ZqqkJh17v3vwYH9ZenpofxJ1bFit0josB0PG8soSnOofBQS4gYhGtOjthHKNU3Fi3qBJxadjh3Rz
OhU0KlJsbzrLRB9QI7G4cdqwtsWmXj5TqnaF/3D/JnZ/AYDfLEp3onZM2vOcCN7FCI4CQznKAVL4
znv3wA8IC4W7K+1uv92Cxb234KQnAXk5PMqQ4LwkL/nRZsDxjiowPXjSuCmh/rH6MbgVl/vWL6Zg
AR/C/8nxFbKHRtdMLUPPR8y1knTHHW743oAJArW9+bqsGcx6UrU7TIWSvlQABbfDntJP+qmlD6HD
2Z5/OoiOIvqReshI24a5vx839CtuVRb8e4luVbFOCXiRJ2hMsmKizO3ckP5AgKZrSS2Zz7eFsq7W
WrngArZqPmq58vhNjm/pp+9EUUtQdbPVHxbT2vq4r/meR/fWzFpXFJe+zJ51Hu1rZSZmD68orXSR
LtQjH57cql3ROoZaSRRizh/PhmM/3sFyHGrrAX9nMSNdugUU0p7zLKKDZTjfkyS0Z3qOnIqGVV+i
NkI5Zg2fXmL1DsI3BDLuYYxQJ7K1jb9EgzbZVLzvwXg3XKjFedNOwUInlhAUNIc2Zlk+JzOlUo3Y
XIQfMWTdb7Qtusd9CSaJPAf8mpStvKZ4j7Fdwq42uqMPkqRop1PxIZQMeDBiAr5PvRZr0Sa4cZ7s
DXEJZD6UN3HUypKfMmZefBWCxnRFoIY+eef15BaAv1ze5Y7NwlL/N3JAmgDjkZc45vaJRsCTMk2j
eUWMCFCatjLexTAuaE82JMB7ENpT13A6wrwojjhGusetiGPw4YbwyzU7Ih9kMfol+YpmRVLZGBuW
oD8Ah2nppOC2YFktmiB/KLTeRYP5Bz3+XKSyRHBQEF6v/F5lYXgw8l0kfRtuLFmIM0yCnQeYCEWK
XwhAhsG3bNxTO3K4l4Fahq3Wqa1QO7ZVw4ZFv6zdTe0n6IvsApZKlU/PPMpwQ16tXp/xLg1tu5AC
zFH9MnfhZgFXtAh2b8bYiWstuQbcC0M9Z9WXlbMM71gxUmM6wtBgvquVIQ1Tviq9TmP1x0k9Urkl
um8d3Bmjij45wE2u3O3dqYTDNLJxO8U43c560qyVrGtUYEqJSEXqmawtfi0Y+0EUVAC+lrrSGca9
LMmWvl4uQlJIEc1+/fEMbVLBxNZhA5/tHkmzhHK85VnNiLhim2SOul19u6yC6ODXtGXKVMHVv7/J
VaLztyHO9o1em1XyHsc6npRW9Ty46KMIlN1bYFvur0dDB1BkvJp0dAY95v5gjKS6UIMO32rU13Cz
R6sGqj5JC9z4UfFBG5hLIC8NEKeG7WYHlZJ+IGV1+jbyxIGTABalK0Qe8BsygGniY/x6EHLvbljd
bVq/15xXlFJtudvc+KxUYSrz619yyDA0Xd4aBUTHHCJd0dDolbaZoH+cKYwY2O3aHmxTGzOoYpLR
pWy7ntmf6zmup4aD6vPIuu6EdX5d3METamz+rTyjOPDsh+D4bzibLs1XvjO0ykcJSB2uI7ioBuOb
1C/v8IXkJYQybDKI/gtnZeGwrisOYgwPSJHA2nWBh6VbZcac6w63P3ghuntoXlT1HkP08lfgNPu/
BVyzl6M2q3pF4fXvnXIPG4o6hhD0t/ofNv1nKjd2cqL3iEIjtDD+56fpMXu8FXnRnE8OPAwGrlXF
foOyztQdzQP2EXPezsJ+Js/4ZFyPl/CpqkI6ze1HrV6qIlLvWABLDDHXEM/BqAS5e428YtYRr1Do
aqZJlcTFroSFu2JNU4U2HIAgBnI5Y2CQ+XNN7bnDasqZNm+OK+fg/SFh1Q314lY/44epVmUoUz6X
PSi6tvopQGwrr7xJakPWjsOwaHtEuovM1KX5JBHrN6k5rrWW8Pn2ZMtbtQw5PtJuF+A6tGJyFW28
zNQnF+/+m+R+rKGElYkcs94XpCCxTnJkvPmIGQ1m1H430W+ZXhqcwaXV7KNehPvSmvvzNFEdiNd7
CNS1cP71MTZpENSLQxJvjj0kLZzgwYx1QuqMHS3SOgZ3uQ0+uKrRaej2/zsJSS/H1V/jNpDAIL4O
Fy7ZUpBZHs6bimCUv41i7CegBTwNkRLx620+ez1ZYX1znzYtCNSYMGa5uXja4r5knImze9QNCbnR
WHbfEtE+rxIbXAdlQ1JcpwJl11Ua8yOqGczvohNwbK0Xo8i6kDWO8Go3fCwyFgEjKxdcs5VjKO7X
zEX2sic4CCrNDY5/6PeGqcFmhzoSWwFTk4iAzt1lK5HcwfFkaMhtj41EJ8hTWn5xnkJiPmyN+RXI
cINTh2Q9AoB3AVB//kUG9Et+FiZe7ntLFsCptHiaebIe8nDUW9dXjSxg50osdnq7F2XmyR11eTT3
O1UoYLW1NzO/SMtqrfSOpHjMKU2fN2PnPFyQ4YjRxjqGra2r4RZ9slWCeUPafU+UM1GhmGiOo/te
GJgO/8u6tdz7bRrmG3px8cy4ds4cfz7U+XwiamXLdBE5dVm3V/utCzpMcXx+2mLUYDdUWq4/NPU/
HCq03o684dZIOpvoXrA0qVKlhtda1V1zLSmMJBKEaYGwmaW7AlB/ZvER+3+aVY2wO4fQ3zCNcW0c
5xVCjwU4DHd0KqkbZeM5mBYMH2/mUQ7HJM1RxcZq7qxtN59i94b6H/kN9TZYZNxoSpaARo9MXTHO
6NqVpXwMZYhDxGMn60VzulElcjgbRL2i1RF8lt1AGQbqDynOxWSaKhC+kybpClqIfg2Pj3e1Z62q
1NBNRarEtBgU91QQEcdNqvywekRLHt1FzsCd07Bc5PhoyH81akIbn7YIVNwrroIQhSu4sGnsetJ4
JOGptP2D6vImiMwoEPq73pK72fHc+Plo+nLfHcoBnsYALU8nWovAEiXY5duKUlmH6BrzE9KnM6yd
LdU0WYoQXX6goVGHJU1hcTPh24VC8Yt8x2Lc7BMkn+krsdZWxZbmX9Di2pUxeEKkQxBl0WCJ7alc
l3dp95HiLTZd6c05zqFGJfHkVAtpDY6FT9eIi20nBuiznhjTMp/x79VYFa/prgaxYLeDpyQ72kUq
oSsJInHBKJYxquE+vKRe6cSTS79q0PWTok3zaedN37ZoyfgQaQBJHO+QEH3eYqRQUcq8kPO9JOIs
w72lzL5z4cY/jMvVkJg1Tl7ZOZkq7hV/8lekyRK2FAb7dcipLJKBF8Vt07yaQTzuspRBguxp86dt
+eC2YwfNO+Rc8R98ik1iiaWWBJaemeVTfPk1deOTbqN5qTJDxOd6tZKpofKRFUclhyzvGlQ5GnNX
fGnrVENVqFOvkkLMrtH66HOsM0HYCGh3Ki8FS6JnyRWAqv30nN5+zj3BCKMpOBx4vSkDkFbk6zmF
e5War3knQoK9CiXbJZTLv49fvfMYCPR7C5QdXwuTu0fBULot/DTWkMXdnO6mdlGEvdPmsQUYBRYH
mvTpjFeiOCyvLSqlPrSgpcKQacYVa0hcKSKg+V7E5WZyWs96zE/GkPzlZrqgmWwqFR1/zrD79UoV
WELv3pb91xdtnX6D30t1YHBZvjelG2jhET2zLILhtko/NTO5XKqm//8XS+m44KoI+KuyYUEb497l
E02kE8JlqlT6P5qr744FlQ4ystFz8LAjn1NOu2/1IdmWxBjVNIrQY0UQ4dLw1qfA5W1EFcjHU0wV
OSa8wtbooco7BOC/FG9KzVo2Lz7zdYgpHpnMJM2wi6O7sqqa+o8+1e/2+KukvEs2N5WJNlTenA+r
0N//QxrqhcIiSteCcWgYOAyEl7w7jnvXItRrkUGmgvey7fnIPSz6T2aNa5vktirH6dCSWhK09fEf
0fZusSY2m9tUDKYc02tf42Yp5J7MUrwXYiExvxf8CAgH6B1s75qyAAY/NLCUwSVi9gmoNQwiNIYz
pPuOKTUznbT2YDchmAFXojQbppIf1Q4C84m0u8OpAJV5rK1N8BaXcsLOwUwF3S86trAR3JjVIBL1
9K9ZwGDtyDK9Kb+/1AMqbhHWjU9uRO+i10mpMRIcp0Dqt98ifg8r0ijMS0m0QYpxGUBJxVjUwvOq
SqM0SdHDD71YTJQDUwMGtyVQGQJ0FXI9g/KUu1QqTpfPodk2KwvXYOIFrNRt9dDYIHGYHjQXLCFQ
vCafIMMT6z4WgX9kWeLxfhURohD6OU4XpA3dnKDsc0TQ9Cf/FLGlvY/FCSZT49wM4ax0OPAUgoDn
ZuCAxV4fcCGgENEeB8rinFtbq2lM0U2fq9EUA6xACWl2YpNLhfcplcrDh8ic3qjCQS0anyqst9Nx
cspIuQQ+74p412tAKgfXsdh6BHc9/UVajg7TbE6Cc1RpJV/CALYDoEe+30kUiF+MQuOjoHLU1CwI
2aD7Fgie4sScxNaG3bDedhsIOUGlnWUwThW+DZvSmqalxCeAnlWJu5pumn7gpJqQGcO6KVjvjNIs
OKGoZqoCHAsJguw8nkRoJIvxRfot8IIXO+rC2OpL7lK/212UKt0BEpDmksBxtnInxCTjdtzKcBMr
yyMKWAURVF/kOwbJ/EcHaF4HthVSP10K4D8DkH6dTT8qY/4IQ/C8ylT5diQ4693Bh8mVkIL4UUL3
1/ErbgCPUIpnP2ZAZRjvzF552b0XFEiuj1Jz30nqLUmZnMV657EKICs3PDfZ95lk7o2ZRU3ZFQql
iGVQeLpOMEIKyD1fVr2J75uG0nw/HD0EBOiSScF2LCFXt6iaR6hpqlMh6r7EdYBaHWMBZIUH/iEG
zyV1J/vj3ZtxX7QVaJXIK5RN5f2FdNlOEWBEiZ6keJm85tJQH+U2e+aUKikJyjFeeI3lYuR5bn5+
ZUhzGPSvXy1FhZBCRPAQwZSLu7yf/TF8XUon6GayTwxVcf8g8P8mczv8ZoE4MSbCOZ2bq0AWbrYS
2TkgWnVTwE70JeCvQrQGH6hzKj/RA/PUauXirZk4vUTlDJGTLGha/uN56ofE5Qacsg+5mAi8Hh+o
2XRrnUD534mhXMo7AFrLm4QiMR8w9lfZz2vJnMIKh2lZyhAxFwcm4iCenGZQUvoO2qexeFnlbBB8
hq3gKk/JdGDmOgSFOEBXbRjVfDFb2sHi8xmvIlEcjN9ENHebsAbptKIgvCWDu3AorvDYN43R4FSC
N63RPCOZQX/l+m0BGYvhS/ntez229vT+buAg2TAWsUAANhFp5r/BRc6X/dptAANzUelw9G/OalJL
iTraQh/xxuVi3VmRYLShuScsioSmQ9D9j+ZQQep7vbNk9Ci8WTzff2/Sd+4FUDXQIu0z8F97zVK+
QYgsuP7NO/80yyzrfPsiCX8j58+MB5veBNZJJQryW0hx1ezhI2wtDZQkgmg5UkLKJlaL7RUp73RF
SE76lzaCLZkb7eZBHs7mSGQ3UKQFrFZPkYGSEjR+mJRXb62s9v+VwRZN3kBZfpEVG/aEY6LgsPfm
XxI6/rl3QVnXHNTCAjesju1plVsg0NCcB2foWDHzZ1JKZIsJpyC395abhFDtAmND/cPo8LgExUwb
ZvIVmnWD8ivhaRr7qwsVFh9EL57mlSiUInTJzoBrCbJ4K4Smv2k+tQU7wwy2QtABRyoVz4/AjgDp
FRB34AJz7RmvaDsPV06WiGH+Cb5f9G+0Rjg57p1uZVEozngUyBQEzpR3MsePOhtbcIuEJzvnd7N9
YwKPTaUyv4zH7ei/vSEsnuG4NIxHYXjTuGib7jU6LcoikMxPj36ink8qsSPNFoZLndUmBh3rOgjJ
NZJ9Ix9oVnqZDjRmRk9VT1FgvMEFsMrhVmJG1iYZAVY0tD45uCyff3KFog//4ZTfPzd5Qynbz2Bm
kfgk0YwXmR9+ZzmemqaTtRvf/iOfWlv43Xyawj0/AnztdGirStVgc3KGhPZ8VpCXmNCeIx2wokkp
9NUaISgOQe9ys+jRuwyGjo3FCLdKfoZ32u3VeH6UKCWbAj+6bbrqvZmfGoLliCGv/5A4uhfosN3M
nhMtNxz2UJmMLtJE3PGAX9CKCajzn4XrKpUTHbRXVqwbPIxqHF/Q+vO3IABm8nhuC34mZp4T+3jo
b6ezHC1TFgs17wOLdzDJZG+Z7zecxszzIk6/PNF0bS+CuqRSmP2Kipf1TUCpIxCFL40mufyv1YNg
nMwfv9ZbSDuG2Ft4dcKiEGjAzmI/eNJd/+Sxnuz7d/srgbqOFr1tDQfZuHdpsTdPQep0402S39fk
s6SGB1A4JfdR0sx29C6nlbjJ+PArZCvyJXigqDTgL/kr5+jhkhjGHJxEz1mPlee0Hrh8qqofrdmg
2zF4YCUm6cB4LSdjYjSPpIMF7fHxRRI6tDVxCCoFLfYbfH5yF7oepa6/bWAlA3LXDGYhZzh2/iIr
2Ai8MPHAtrhJUFPGX50gyTs35Gg8HABleR9vwA9afntzSxVGS2A/wXQy8nLQSyfR3PkwUIRLJM2j
AljDCBZB5owt6hn/JCmqIfapb3eKoTWZvPSovum2gaBqhO8WfyCaCoDD41ob3K99/YYEcli6dFiB
Bce9Jz/m5P2puqLFQClknCELmi88ATF36idClitidDfTh6IB6tmtK4BqdW9WBeRC4pJOQDJt0uYD
gtzSJnd5291hLjFy2u+CbI1CJFrsvkmxConjxSXk3+1n9HCGWjSdQ/fHyAnW3kEhBRo11dr6k1zC
OZLcdcZfATuwrOSy2G8q3jZLog3LztvuBHU/XQbgfJ4Gj3isZ16TdZ16R0bMiigFpvDJIOCiVPIG
kwL08R6489fPCOUFlNRIzkwsIPLtUSFsMR1mWT/woflYinylLHnYTxk50grv9v83ogVnKhRvOEYi
ZKZYNVlPtyQPI0uiJ/vaMl/qSKMUYggPlRM4FjXxlVjWHyx7kzwA3Ay2JA1YVIn+iLxP+7Zw0z5h
xS/A256RhkvEK8gGIa8Ht2ZQBQVcbbe1EogjnXrAK0stRgj9Sbu7NmGXuOF2y2b1JSVz/os3hUrU
Rg9RblAFMj0BDEgktdVYpOq7NQLJOiMT9LOlZtvctbPhJUVbaytyMCB6ipfM3tEYzBCK2HCgkdXK
RhXhN1l4u6hyRWYb5KFjFQVtNrZ3aSdGiI7qPfJx2UqQIYEiXlgtMzVLjhlg0UikHeS37/fdERwZ
nATIkkkRlCwOQNHz8tn479A62xzw89L2ZwtA6O5y+ubLzpbsEb43+D61YBab+pJGW1R/gJbUnVrf
JfOk9mzbaQtYbIlsdGynqZme0wnMChDpySoPdZcHhQ35pFOHJhP1mIHPxas64Obl1NC4Swjq5mzh
cip0jRpmLVrJ+ZarFrkwcaXEQGEHObiT+VMgauf9/AUu28D6qRrc4uNvwC7fIasU6ZkUouWejkUI
7UPexqhVo9Ue0SLleLYTMM7My2zzvyAjBSSOgyrJgTRVFB2URPoNwsdo4fMI7Bns3psTeLIlG3Fg
MkU2Xhb3n/WCXZeVdlUPAZHBig6V0d6n7emOrTnb/3FnZN+zqiHWoj1sM/frhvcSjGmrDLv73V93
FDk8d714Gcyusn4lWG4WIGK0G5V2d3TUL5+zJUghxptivFanWRRxivC203DYlI3W4tnF/zS5754S
HOeCADajoUGUpd2cFi3gCsR7V31X1k1Sp3bhc2sMYhIfVqFVUye8fc1PN7VQsjnNgCr+9oXfW5cH
jP+qUd0/u5JpONp2GS79FpL5fznhdRzjv+y6ZNoxNRW887NGiMei23UfdnOp8S/+t9Nu7yclzra2
jP7+fJwfjKDEigQa6lZvi5yDpYNA4bY0imCe8uBvdyW1pQp+sgJvdD7OlN8dZGiwdlxq2I8J/X3A
uPFaeFSWpR1bV35C9vFjOlBxDCEUdQPpeil8hc23uAP3Hqf4/nU4PmfWiDeT1AgZJ6A0qQiW85iS
xquwqshOlA2TXNh1lj+ED7zI9+YTBlLaji/ey/Wwpehv4tzfG3ycMQlSTMqB8lDhyn0bkVJdE32p
zpumfE9cIANl8ipWlnsDfCH9u9RuyYtxYfPKzay91qlZ/cyMf1gBOmdJNavEyp44b1/8ahx7tqpA
NqpG4eVK4FbEgVa0hmVS8hX1unfZ7cmLVAdg9WhZHsf029eEUO+iwRqS2IzK/ri0WM/H7JUzvMGM
czRscsrkmYqVOcDU7/GQ7t457yGFRdS+qHJ+XOgAWt901msnb6CGAb8Y43TgSshjcI/g2xH9LttD
1fv8q4O6He4EKWC/DFeWq1YYAyOZ6P1qvssvd4HkhcFvQgBKYfswXKIluvmO0I/QmyeItVYX7ll5
UfnWlyzshlHBrDkcV1FfcBjMI/6TbWG+KBoqFu5eIHaUWKh3AB4NwCa79Jikdyu7z/4I/e4NFFnw
qZO6CLZpD2g42WCHdmxY8rgJvfx9BkVk61goh9n/8zcSnNiAgvhoxxh9Fimum2m572kDNvQrVYiF
Fs7RJR5Dpeffbfgoypqs7NT/jUSChISVanbOEoipJN7lOjrFMH5SlaTKaKWVMYdjYYXp33fwqQ/I
6E3t2c44pO0ujhuEoU8SJOoAYBb+Fbq2MR6TF5eowDsQn4VLS24NaEF5weg6DsVuM4jyiWpVCZXD
AYGev8c9DMzYJZccM80US1vRMRk1X+JhSOCG2zTp429WT5KNGC1n0lunykFDLjj/kw4PhLfgGYm/
RBDrqVyhGdezNgJje7wNFpwnLxtTcCmuQfINrddazVOSMwkyyrYb3FoXWbdW3z1LOpeB83CzDOT7
b2fsdVGEuWLbn9P3hQU2kx4N8oogj8Fym941hJhfoak17fqTv0NzNRmv1lzuVd5goKNxTFnO+Fc+
flt+pPTuViJ728PCyojjUqTiZJBLxocTo6+K+i8z4sjX0bnLb842VZjp8wYn+xC16uXsy5LBnvJ/
q300aU/T7tgKjkeyi7ql/Wmd+HSCpwKcWthfXpd8LwiJSEr8SUaSazv5unC5am2r8gH5pNif+tCb
AAKoLSskPepM7lbBp5MoE/SAYHzciCcxVTdOj+n5qNahqm8Vp1m9rHjHkUTgU/nP5oZAmAroHzQo
j1LqTqiUWQ10mtJhVSQzdwIcC5BnSmhG8hEpG0qgjLi+pU381MngxthVg+2pc/yF3EJqw9aCp6nb
/c2BhoQK11CzyPpeoAmGtqzahUuu0mTBJxZ9/W6jfbdLKWxZ2BKc4gPc7gRtd9xv95ToFG7OI1fb
eoJXRfCro0NyfN38+YrNPToUARGqkMxUI44DOYUKfs+0BEGFKwLnBbW45hKDPWrKOp8k9guodie+
Xy/EYd2dIJo84NcOaREs+GVFWfFEgzGlJX4K45nSCNxqA3CC1eB/4WwYCsaV4/8Adf77HtygNwdO
xVKs3BmAhm6hQkoLTxo0nBhlg4oft3E8ZNDYIKkMEN2D4XeFBBHkLHwZLSwJ8kVsO1vEpHTQLw7h
y80pKI7Y8XvAcT1gtDPdu8o/VrZztLGXpsonr+XUIscHnw/vL8nQzMXgGuuXtKtM49Ac3oB4oIQu
4SJ7Mt2knGx14ultBRimDh8qL5XePgLp78NaNOqDW1tQHN25ZxvfPT7DCgJb9RyH01T924m8FliU
Bglm5xx0ROqYCdEe4x+u22EUmCRuXn31/mJn8kOC4AibSIsQBgMe1W342fRcx/fbLc/kxcr4BmBS
WjOEEOIfvWSQWVuG1h9m1XIWDMmLWHwsdG1EkVokrpAu3mwW7Q+6drTxLAzkt7M7oSRsfoL/iImI
X/0mB8oapK3lHyeRXGKxdfz2M2fhq6ZjFxmscVbY8gdAkEBXS0ZdHEoY1t6P/0D3VVHUacJmTOiz
zkKJIjUO7G2ujx5g/kNQMoXIrIg3zAvs9Xj9I+hsW7UZ+HvYzlgBLRzGHoZi76Qli9wd59JMS4Po
927hVE2twdIdDC9RaGAhLEvxh93VggLyWzpAN/ahfAu0kt1TKICsl2jmB56Zugore/V8EWFEocqE
5o4iG0YsXGopYiXQKzGQfYopwY3wm8JVI/TmkE7AHTZt47PEzTNzhblc/13aTmW77YgYRuDftDqM
sqaaWFWm3D1Hu5jQA1+h53MWM/Zl0FRI+yd/QCJ06k6iCvSG1H6HAe+CYoz003czEBSCGp+ZvvF6
UP17lNqGq40bot91zi9re18dltCDV1sFcwkBv/Pa1kTEFEHtqg9zN28oUwLNTcSa6kU5Db+OFPOS
XMYMtUbAuykUTWa6w0xyTuVgIzodKovNUoUtySNmPkDoIYkL1gGqm/0TEFPBq87aZvJKQm3mkQOY
y7g2u8qMBfyjqbP2gvaXtdGHbFBYdXJRPFYAQdSq96Zztr80kFNvptUbj4r/Z/kjji5QbMxvtBGu
o0KrRGUWmKXEeV/Do/1/o30aUT0G0b9J/TjiP3P5sdeGN3syYCI6WniksuD1usFTDyNM5WRtau2W
QSiuTKdVP/kOVSe4A3nZJjEbhg1CaIBOQqfjX8bXpCPNEJWyNPmzCrENuLMPdFlHlSrb5hSfUs0h
c4zKr65eWj1EksJNRHJEMEAthnMT9BDVYxXX32b80/4UGzs+2haL0KK2do4fdkqA4kLLNrrO/f0o
mEMOLG0FfZi7IARHWhe0H+ym9nUUG4oS9kZba8Teg0bFH6+5ZCRQKr90iuWJ2P9XdpaCkx3zgIGA
lk7Upb/v2cxXo4DpRlRgrf9IE0esc+ugl8lbp6t2Y4RGuKys29AbAY+xrAPzYeZbTC1vFj5/Qrm0
EkAEqNtDBM3O5k8VOgRSOXv/Bh1ael7dKhM0vB7LgpsSsOy4KcczENesAgJqNDQN3KTC80bfmu/H
eQ5X3O/fyT3NvBxRqog3GZ8EhOdkJBB4uIZ8veT9jJzIKhXRrtKzlld7GRCYdcV/3ML3Gvjl6kLJ
YBMd7RdJV6LaFWq+M+DWITu6C8szmQxh/EO5ZeX3Ew+2yErvbzhDNPcU7rvHT6Xh+Z0K/zl8stEp
e2Fz24CKUsf3NCwdxWBEJjz+egEkmOribvrTThwEvoCcpco5lBpeKZhnyR1W4y1f1otmwbt1BzfH
y1JYrkSeGSFGtMRWu8rhFNAth8wm82FUyb+H15OhkHXjqrhomOVvUe6exg7Qf78iZx/8Sm6VSyjU
iSm57Ma3vNFbOi5IWn72pEIafI6cV4ZE4pKUjZYc1jQQqhM4MFRKfkBW+v9wXck094E0NNrNALGs
S5AaEL1/t4QHHxpKrX7WLhKFgDkeZZw1PP7oE9Q/6XiNHev+Iut03UNDHLXHxEBmjvHhHjDsiXI0
C36lHBQLOqZ3NWTNdziQqrZ+jOK4oQvV1yseRr2U3xpzVxEhrbEVFFb8Y1k8gpiNcCA2Xf+7/khp
9QCOcoX4mW2WVC4lqouldiTiCfRZx/8l1GtdhihWCpOqcvmTl3BjHAAxEkgRmd8iKgBeaNCY1JSI
WOOp7ykcCD/h22MhXkQHL2bIR9d1IFnRqIWa1H6r5D2s2RYuCCLRKXTCyZ5wRTEYeAz3ZpM1iMlU
kSKpj7ScDuBWgdZi1CR4aUwXX4HD4ojqUQ4JPmIor3plHb5kSevrHDbkJMcjGKFWdCTO7IRbeRTR
32LycvCQvYnNr2D1iBL0duLgTlUQISXhTQF8pXuaglxOnmAw1+V/XDwy9xigwsVSpTQqZwv1UvJM
bDFCoobBtPq3AQWBkevgypW+Sfd0aWYSZeYlbfLuixg/MKAKZcVBdtMBsXz1RMMVl03Xq3Mc5VWp
VtlaIt6SzGzb/ND5aCQkDM/NEnSHV9426OjNxd+VuHjeN/44l3aR4QqijGxDP1z1B5Bt6p8L+07A
aRNFljqwNFfT7gbJ009PVikqvMG2FyMDbLk+v2+6YMiyuDe6ISvoKP3CntkY1yAysQPkhlqMHvpF
XP9hFbngVmblirWLon8uLqGDwNHA9ZhDNO3HVHcbhAnGOA3YACs0s0Ty/ibK4xbR0NX+THG0BwCE
t6u+XzfnNcBJwz7TMj+g31yqhHZx9VVabvOgV4S9k3U6zIbIwouNXKxLYfRZt/CEcKnSHOG0fIWx
5IU4BDJ751Sn7byhCBX15+G3AmZlCml/XPWoMiYb1+w+qUnnMLUGUMAlZ0DoS5Dy4c1P08kaR+yy
V7UTl60jJ41Wab/Ga+M7PorLegy03hfpiagWqxzB7mX0HUfss+YoW9AuzHB+0w3AFuEVFybZnB9k
Q87mtk52pHksyWHqHAG/8LOnhkFSY54oOE7s3DpSALHSwGqBle1WBIqIu48finb2gNyEyIM/BC3n
D40lvo7UO9j5twxafxWBSOiSQR6aMTdLdVrsSQA6qscN9bBhTRq9PLtWbRLClzuumqmPMK4m3nAj
v/ngw0XnHJ2H6CNZ4JJV//QNF8J6CmdA4QNk4/69nrHUMsmTz3KnzEBX13SKZgqucTcouB7tYTP3
HY9vUO/EJ3eF+8G+KUM0H+P9TikiRnuFCiXLLcmiTkhPnrh5gKdmG2RKRNHPcAurvQfWQPqt+Nni
Dj9Wiq455imFYf5Cr8CVS0AyIDTiAJNpfb5kc9rYd3GxpDXB4pI1A4++WQ/TS9ZGotMPbqqBMj9u
w61mjRCDd5Asrx9PNH6MD4nSU+0r0C3g0V4HsTLM6vPTzWRM4J01sHNAfgydWMWKlxsm8i2XHvTx
oqe+svxZMHNsHJixVdJrxjssaDWF7xIhNeaBsdXPAjwf6v4+0/rAgajoPxZDij1SY7GiGAd2Z5Y2
7IuhCKfIN3WsMfhx13A9ro14kesVUe2iMUHf0ZsTOjykAbGnpUgfZ808+sQk7Zv3NztTc8ZRjI91
O0VxdKaq6b6uMqh0DOFi1kRCKL9+b7zJjxo8pGiE11/Vx+x1JIj5b8lD1FszQvrHIc3YkQ/a1jor
oMpE/ZPaSR14CfM0c7abWPop/dzVystBbk+97gZeI8nNMSTsU1wAraN7zoFxEjpBTySCFQ8eGdDG
SeZ9D33y+oMyQUyeq5slwLGVYCe+4GvkfydEMAubhMF8j/8WwYnWygxHI/QoDzJ0yyZmiDH3vti5
7PiFaqagyn+hw86uDnH8mi0OlDFmRQxM8eWadNfGcQFq8+1L8NhDVgn7AzWpLIIUlTeEoMDUM9uq
1cgwIe2e1zQHKJmDfAtBwaPgOrjC6G4fBJ1TAP5zZl/acbvyr5+AMJ4V270HIlSgOgbT4JRWtjCa
fulnGc+Rbnj2AOOI/rFI4e/XFlQ7v6aDoiT2mv8VZY3eYdy05G/vu3CGdS/Q9pTDsABvyWoMFs1N
SGsk7oBlpHjsVhA8XgRFSing4In6s2GQbiKUGy9TJ5b9Tqinjw1VUMxvXqS9zgIsLRPZcJfiwn0/
ZgWNFAzEbc3p7n5PFECSXvpA5ZawGLbKJFlE9GKjU8GnJabMiGgk8JoHvlJwBeWqx4azApkIWQFv
dajWS5Pzzk+9hiCqODgplZ34K4LYEihWn8QVQCBOscY/U29Y4OU+Y+Ccc598anY3IY3qqA14O9pF
r8dkHPxyAVrcEymcAt76AI4rEkspAGrwFF0WspcP0k7mqY6Rs7o4M4TuqECDtkQpg5w8OBzkUj73
Hx0waUqJ4EUE3Ghn0jhSLpnqRIpMyKcnNmiqh9vGT0IyS9LNCTNblHo0NY1IObdQbhQFnowpDJOt
NI28eciJ4jKcmhHwDaeMyKcM/S6ZnyP9IfJD6IiR4DWmsWvFTP4i9DpJZX7gHXCBMpLy2at1XvzN
+r/JUQvYWcSchALyyXA5oFb6S5zCiyFxHjzONved1csXE4lmPkLUzloBFyMuNUJgvGxRG/NmtPqG
gmmYJp6OlH7uhkfk/Z76+SAlHmQnPrSOIG5BGuoEzNM5nuHxF59DFXuqlyUPJEZkxFz++MT60e7o
rLWBP2b3NBDTriQ+2DVqN3Jjx2azQwhaTlEop1qINQlfcQPuVgYJydJ0ZWe6lFIRpIreqpONerw2
aGxQxiiML0CHiyqm93RDL+2zVK6g+AkKODrqZkUnGgMQN9a9fySKdDAlw/8KQJ7fHUv5Jx6RObdg
q68ZsO6q1T0cX/Z1vj2BPSXzuU/EaNv3nq0ye9/R8Yxb7bg23yWctbVj7NVW6m8ks8eh2b7zss5e
nTJ5oLTg9MN10L6pT0vKLdcQE9G8XpAps92JAazPzhjFDR0kQaojR9cd0CvcPayLntdaw3WMht8T
/IH9qJvyKvZWEctmqixmXREC0biFMGc41g9eJ7nRoEPalTJPL9kTRdkd+yYJ66MU2fI25qjwCfrR
Zx2+TyVxoD1vUGOeRoUoEcro29qAq8unWJS169spKQAT953GftUAXkFRwMdAC5fzY+WbDl786BBz
cn/Zwc7GkFp5aWgpxDgt2cZsH/WH+ZZVXSgSxRVVq7JCk8bnh8W6Vf47D4AxHxbMzfQhYVpQgMiJ
KLST/Lvjnw2DSmcmE0tbWTwNlMoD/x+jE8O6z7nbBJOsph97YzbVW53s80xKf/MbMjOqq7/Rka55
bCcawjR3rCjG0Gnm6NTnknxLw/ooJKeT+NUcfZcMlD/IHgQkV6ihQCfHwL569KKJg+CO1jKqTBpg
Aod4uaUYstLrfyBB0y4BBRHTvmJsmvQ+m7W8AiDiQt7S2NkBZ15KV+xdgS2P/3q4/SrNzhrmn3dC
gmwf1MOUKJ+m7PPNxyJ3q3PQCvawFBb5/oAxag8nT0VUUo7YNpER9Mw/XIgBdxAfTGkqMhB5OZf+
OT5ULiK+pFtCfPAbFum3iSa2D64GchQB2ZfEWoX9tRU7yYn4fkKKcS/goMMZlLoqNPs5+zv20EH4
1CwPqJ4+cu2VoW6PhtkKMzYDPQZ7LAwsSkt/n1eYyElCIHRAYFQgJP5E2lReFeqcmX/5+IStsfQM
FozV5GmARJTowTNwGSDP9mmYsVtGuf87nDUZXnpLi3ob577uAb8Eo3SmbfNr9EcPxgis+xj+JADl
STY6VrnwhH5XgSUnqnqqzQJETijoOs0qEb103VGZnk37ei55cjVpM1+t+IRYIFRDm8yHLD4RE8O3
NqoAJmhCTxie3Fsi+rlXCOx+lIk3p8R8PLcAMtlJwGqfIMa61iFKRB018QJ2gXmuHxxYDE58OyRg
BNheos3NAxcvGBqe/AU0uG7/sOB1h6HU9/tnyqpqn0Wcj27yt32M6oAgA8MoqjWzjAMC/vuPb59i
oZQ1YAfOGus9esOghpq+Uu+2xzBasZImld6ljn+HqH9bnVfFpaTB32lO8TvceEVHwQ687Hs4Iepp
ruxibeHrBjEPYNwP35k2n9i2EVNEp1yTIXgeIi3RyIS0xHXxp5wABqoF5v+uUZL41HxjtfQCoYA7
aMTUyX+wKcGQ6vnFPjPpVxardTQ30dXkjaQvduOkXRuVu0nar02dtAmrl0aLib0NlGKBH+bXdxqR
MTLcSVSm1gb0QSOsE/Id+y9JhAEK1MGqBsNBx3rw+QOIfVTdIBl/YIL8UM12z/vcpg0TY/lInqx9
ZaRQ7RbTJMkaWDAxvY9MjyGq+ZYh9zVHYU2vT4i4kAx7k0f/cHQ/JTSW47MqohC10TogZEVg15RS
lP06lxQ+DFf5lOztkyiF9BUkvTXoTL2o8jpzQmA/mkj3Z6PYq1+aU4+MyBLVAmkX8dOnCXfFRtTu
D39Uo2doiMV9ztbjWDop4zjwTSMV6dr45Iaq0HXywdzpyb5otEdFu0OsSwr6wuOIAvjGBNnQwEwV
dHYo4fCrg2JDxvINdsIRCyZSRr9Sz/kNDzACktQNQMslCiYloOSZ5kqSCSbJ1OWkc7BrO/LI3wcC
k14v6lLybjLeZ8zcdloGXg8p680aPZLJOurhLualtkBX+8p0ABas5xKv61Y9gXAloxUY8eATF+Yb
EF3u3MlLDE6jIz56BmlAKDygof1ErS6vstPf0JemyViOF7AZBEGn1q25GMjg9991l1Gd37Ofiixn
p9eo3do/hNP+HZmtkn5X1ga/TkpK1H/Xzdk+dT7wVIwpysYI0grPYf20iip0V9v1R8RQa0AH9ivy
r8vTEgRrBniWhNakULs/ScIWpl2B1EZqQ1K4/zuCFBMuoW7ap33pfVLR2bExdltMfh8bFxXVRB4z
4IuoUwtKXJK82jj1dFrO++ZM+Eii8sq8HumplSZSkn3HOtqKYM/0QrJNQdWkj0w0swlTBEhhmRLR
Eot52eDek3j6s5kHxnMcdcqUzGNBVProaczIflF97D7BDYhLmMricX41UYXkOtxKfcz4dffKAyqP
9yeLj54MgJa4+E7IxF0AiQkOMCRVwZN6WC2owK56Pf1x+JxmizvCYQ5IuXsHwUNgkrxlEfpeB3JA
KNh0NnlQaZYw08fhbk/5xHTZ9jqlO+3GfQTQAXF7vQiEqmk+l19pdLhBP9b0l0Z9GR7/diVNaMOn
phd1HKvY9x9rka/BKwP1QCcBfwOKGTtf+Nm7sxMXz3e1ubOIZ7SRefOgEWsuhezHwnWXEE03CTM1
UnpChzbE5vbr9nrIxlmRqAGDWA8w7X+wcP4v/XCAvN+6utEgbFlXJVaaW+iqqCEJXEcVQdSQ8FBL
l11DrNb/xoKYgdIHJqBJASIC2czSgBv/fQhLa17QbU7NMbs6pGlxHxuHyVZVrcmu+yQA28WV7a6F
abzYgWZOkqg8KGh5vj8OT2eQIoGPSf+PxCKEFb7Mr1S9fkLSfXFaUiRsTu91jyRKeVYjvwbVsRW7
axK7CRPP6CW0Byr3ZOl4TNC9whpSUyQuKS0XuuBl8c/LwRLJnKL6rQ3cUaup2DxILALoEDnB208c
yIgP7QDMjXYv5frq/aeuLN2Pq+uAzyK4Ymcwzaw7KXl6htdVqWvzp+XUvvdri4WkN5TDsOGgzAFw
XmF5D1YZiY5HY2fobziA/jqt3A10IrYyynybn36D4ZXwzxY8kmHsqZq+MylaDZnjmm/h7s1ruTOE
llQPUYGqXd/jNMos+//NNKCj6AEAlsY8IDRgPMdOtcIbtXxiHi2j/PSSEPnb6+YXZPIsG0sGjBKu
Hmskq+pRIm8OVBa/gNqr9W/45sBNgSJYpCpz9i3ddWNRiQKS8sFsovC7OuXt/Wz2/HMnAbcSNaL2
clJNkEwrKFxBzRWrfk+mXkw4T6mBiuctRrUo+O2C9I1XBGPrYArOAgHFv/C7anXE3gxnxpaERIOX
Wt1kG+ARGVPziniW/OYz921YN88QBaruZPaEVY0dz1qWCrnB3vjO0NwnOMHcfdgEjR1XXw9US/b5
rOUHi+cHWA9WZKl6coUHt6WXNrNJmcF07bzlM2MjTv8jg1vj4v86U+xcDmsz18t5cMzH7mTHjNve
q9wq2dAbEWCDYuEgFTavThyyoivrVvXgJad+4fZ4mRgeLF+J8WdqGmTvQrQ7O+jYb5TtZOJWsk1B
9ndoq3Pe7yiikvV7Ad1pZcqXENcv585KOgjiI7Riabq3o1QY+c0kYlfMIeDVkm2M+EQ/YEZ4M6HJ
qAmQkpyDHeQ/JRluf6MB64D3OpOwHN3XlrIApdPeKGKxhMXnL7rj8twN4DLskvjEKRMnqAhEpPTC
fksoAoAhdhFZsOfmxIYDoAGQCvfH7Bd0NnI1/Nb2tC7MYFhiVuW0X/RgQDSXmDnsvaLVzgMLXzEj
hThWUAci6AEHfBpI7gWnSsJIBMGB16UdB+Tn+oQ1okDEwPpgIQ2sBWE9l//r/AHEkVYpmQ2+KQpa
cf9cqzO+PyXF1JNluST9g8/wGkOD3Qr0Iri2gwTO/5mUlj5/gmBQ6DgPN7gsMAoUBUKqHavVrck+
jEkVHiVoQ65WZAqDRtMlMxII5hWWSRbPp98R8HdMV+Ay+8Df6+N9imW/2WcsmP54fg2WP7M5Kb/t
lMZBEEFDhADeDapwh2tRV0/xVPuvHYpJRv/xF93C7i8ZfGWkLm3gDhmpF35Bte4Qtc6b2/dY23GL
Y9RFqfOrY2OtzqL2zH+byFo58EkMcG9aL0JY/OsxJkmUh5m8RhzYyfGt/vqxomcQ4YWmLZAz9spe
iKNAc9kSDGhqjxWQ6HjXbr179sddojoI0SmsK25wNyOhBHptG81Uya2VjdFmsZoKpf221JnCV/yN
9kzAIpz86rGHFZ3yZuUTWatNjwLhEClfySkSSNC+4VxcZ8geOwJfOGqXkwx9H0LgK9K122i5J0+O
RjEZDNxNV4fS+ncPSzlxIkvgIAuJF12k9IrZlGy6H7S3pr+YgydmjDz1HOsCHWo8ExEnG6xMKg+a
eB/GL+CGRPhLRyDXerYu7mCbqQalrNM2YK23Vo8WbZqrm0WoUy5LIiCfS+YCFQleIFVUpN9hrSga
9tLGWENyWBlj/CvlUVvfLSApKGdMzufdvxAg8cBebOQXz1B4+XyD+s30jDN4I5O79/DdHV8hzuFL
/TvKmJDbbxYFPTVM285nGBcAZcbbGXQWt4VH8Wb7NaY0a/VMT5szLeZDzoxFDVi47X94Bm48EyRu
G9FaqQZ882xFecz4x3SsTBnS92ba6LwTVGphZA7/ueOsnYN1MI98uwppSBOSGuljRrUinpBm6laG
F3T8KfLv/sCtZxnuAs7qJNMeRvJM8lmrF1HcLGIs8h/CPUigS3LUYaFkfQs0+t5SueUcqBI9SdUm
biwUIpBt3eq8Ljihdq7CJ7Ufsf5pZ6gMuBE0r8dcS4h3koQlz6UT1q5E/io3FlN7Iatu6/AjF2n4
mvBA9Pe5k9rU6BxtpoSjZhn2AilxVHcI9bukNwrasb0AjJNzKCBuv2fyHm0LqKW1KoBcyx4gMc1L
QTK1syhMp4E9wnfmq3iJh9KA5MOYTYn7rQdAHfJFPHdA9AmjOWYhDVnJeiVHm/JgHp5VX3eLn3LL
mcvryLwRBgCP96HA1SiyEkHJITn1TpvJh5I9D/EGPBMGeibx/ai669wbKjJQBF3/henMsTxBb8ZU
AdT5Xg+vTCEcabYkHGsdxyOXLzwiacZgkK2m+P0il4zISxHTETbn3kip4xC9M9xqx7jgN0raczXa
K+hlPvsrIWbKW4nvhHd80JC/DdI4s8Gww0VJnpqdVz+QjCmS238r0I/AxhzI2zA3plJLsoY6AIYv
98Do82h7ER/LP2+GR5ftXc3M4rRvYapmBWWc31rHdDUD2EEjU3DlT1/Io8t/8B9o6kVNN8vzVlv8
Q/75c6LMKJtDfSh6FSOnW2GK5mGDLetFNvU3+4mDfeBu38w0arU7Cik+aaP1Q1+Mt1tDnl6hmCN0
EE/8JPMxzsqNtFkulxcUKICYG78ojv3zgJcINXXmhWFePfT2MAkZYd+yt+HLJqFYSl63wq6jCA6t
cinBe9ktX6z0mf3yvLfBb96m/zb1N3zSDh3jRPc4GS5FTWeCwmGhhfh4hHvltV+i3rBgElCsjopd
a7W9vNSFApzSNHvECANjo600uxdigZtxg3rAR9QWGD8QkNtpdLVtwWTt1qNI4EVyAxdqUwhe4n6s
kX7bWqCHaEQCv4Rhp6oHafB6UAOCP/+LQs5h0tOT8zDNXKumuAfBNhaL7TmzwUf2j5sYJ88fg3Xy
9l1HpNPLbk5KYQUcPZyHBYc/Dr7my9wdzm16RiBUDFn0F2Q6lxPOjcS9BL29OoJcqlKXhR1L765u
6l84Sez0U138E2yx83hWtMAMNVEhW0yDJcd7++mUj0hXpSeAegWB1chPUuyT/OjUMWKlPGukSgf6
jqif8zJlZ5QoO7FRc2pZDGHl2IdasmGFcIzFd19pk3hpADy0JHGRLTgUQTiCI8oEdqbHCMStfOA9
voeNJtdks0TBmg9wfURXCNf9P7ZFezgrrj6cOTxO7OzeQJDtruAGd22wAB5I9djWUWtlhk6TV88e
6YhPF577NrVvOobZW+EJ67qhtI9XzHnfQrAztkP4/2yVYDbVaNZk1z143SlA60D304ZW3+j3BEYr
ug70CK/xp3mAnzHroyeyeZDE0CJD42+2NcZEnfWP9eWZca9PKbEkfR0OvLsYAvrxl1+cD8Q2q+AZ
sC+YDAYCav2yxDZHftDuXm1frg8E20WPM+lKLimCrTV/Z4mtpIZuAaChcrG+I1701y1aB1sIEKbJ
wTlidxxyOBvqVsbkh1rgXc4uuGV97AtOHFBYfhWZSDCUSPF3gny5KFqbgR4UtxlhqJNPnKbulT0F
0oCklk7dn7VfmrfUnI+mArOabKn1yq2CHNwLZSd4d73aIX9xrt9FyygdvZ79sg7ZurffO62l+lkg
LDFqDdSjbk9P+FGYOM/ZQu3trlyEs1G7NFTn6f1lVzKh220nbqgIWl9W8qxjrLPpFkwr7yXLTLV/
OoPuGpVd3FdnP5VIy6YEXouNYOHZtPEvhuH6CNHz8nnIBHtf7N/nZSvERUGqfUweC0v7ii71fZ+h
HfK9xs20g6ZyiyYV0Sne4ZkjwdjMGh4MADz2TOpirNF69v0R+/Sov4WEzbMEeFqjyzSQOWPjNdCS
mjWJ2y59Y7SZxEN5koiuxWv1mWbk5s/1RXMJRWaAYj1gJGoFvqKNPu1JVbNgTRfoznBrRyshcSko
jp+qH+6RhNxgUiR55C6Xm4chMIbLnRA1DqnmOsukOz8bBDBcQ1fPkecNOuM8ZTLB513m21ITS9Jb
x0NO6m3Al/fso7WdeE66lompQlYOIWPlFk1+nojVisl2a5mdvLkuxD6wl5xFJVDeYq1sGJoR3EX3
DSBmKVI6NKnkUoWRtpiQti1AcXuD1CH7i4jT7CFO9GIt7bBGyaAYj8o94883NjvCfCp7krX/+r1p
wvq9ZLS1Y9G0lqol/gknjNpgPOEd9tr9AXNElhwxzzXuA0KJcqrL6rikZEgrpidkfUxRB+VpNo2y
v2qkAh8/FYcKUPbEoIaHGQK1DaiWHVvmqKTvoLBfMN5ZZKWhpoTYom7Ohc4YW0J5HSlqTNqv8xH1
LK/UUe8vif+Mai6mIh7E+ahlrix/allFGqmu38XLbARbhWa0+IEK4ddGQDlWb6bB8reE03oi8msJ
mlL9tnemJY+9rpn4BDaHx1p1qwFB7R0teEfHMUwVmDOaonbWE6OL2tOwetHzM8CGJgUl6TzXt3Kv
i5RdRGZrzadRvxn/eaHoRkrHF7vD55bXvMLwmYBXPpGMUI4zytUl3mlYyrxs6B2VVpYGCu3NmnWT
YmyN2iZJqw4kkCPeO7AwlXjqyOtDbjD0qdhLuwPfyXgxtKGxkK6zn4sDSXuKtL1y1U0nj4UbKmwm
mKcxsLD59eANZUmj9XRPptRE63qUdCpYH4AuBVB1Tx86dQOP2GcpgQajekM8hyus4kgCSqS8jioR
WT8sNMEsSDwd95jiVYt1i7vq3fDYI43oIlVNxOR9RmWSWP2wWrVinExh0RdSgbfvulazmhQGOMTt
scW8LGf6tsMpe3+kTHu7jfNZCZXB/v+/AskupujLHf5wDil48Gt31PfraB3fnDynXp0ZlffnWD4Z
YKdMvFOpHAA/9fh23LfEqgxtObgy9ecWR3YzFP/GOKsuRWf9TVnxqyDPfobHrD+3rabN2gonQgTj
571CPO6pq3Uq8vxZAMMRD8xwxvH8bQXM2Hvu1yKTVlNdUuxfo/HevF6I2T6une1Vl9is+B6n6KIh
fo7L1yNqddzl4FoGaA3qwK7Fkx0K/cZUYiT2ca6v4cdCgKxqDqyn9XXuXizmg0Gf1/kpDc5cmPwr
yUFAadQZy3x/s+pwY51iVtazu3kBOPSI19FnQbEHoCCD4T99vD9p7auJZeoF/tATqJfc/a9Ib9Pu
WH5smZFF3XA/L/tZJFKqRnb5cKD+VQtt7mV/f6IxfN//PBdlhpXTci6n2j39T/1/63vleTZyzQr4
dAcOmPCfS1jM6u+g4Z00HqesbUBN0HpTannyNFidIVOrfqSNfBAgh5eF836zuP0Oq0yUZnC2N4pS
0tL1k+K0Zkt08JGXm3f7+Nh3lftS2FJhLa0Nt57FQFzebytI/Gm4U/+ZC0461UMqUTNkld08X4El
lamr2jcD0qY5sR3tRufnTS2etJrbwzJm/2T0YYFqrVgdnI5dFD8ulhp1G4atEGCJEnPnqbhMsyas
4HeJjwFfI30/G7hv3uoxPwg9Uncibrvxfv4B4P6ESdQ4j/jk2Zy6KwrGFj7SAAUCB6hffk8pl8qq
7gNFw4a6icWgLAr7tsNnW06cgYQC8JHpFdWUyY9VviJzpmsG8z6Pp8axmVWx+PK/j71RvaGij7rg
RN2HJ+iP1oXsjZAyQa2iUtkr2ctvenGTPVrqDzaoavLTqQLRBiJcfQzP6Mq8M3834z5vD1V9tgAq
tUJUnHqkiOD4v5+i63+n3Kg5RFWoChkB6gP4AzQofRxjmGx1jUIuNJ17pgGQE3ItwN+YG/o5uqP6
YGrCTKAnovKMWqe/efxxt4+HZfMDmAOBxkBxwa4zhpu4R1NMYCdmFFKkGm/z6slpqCg51cawylFB
p3I8pwQdxqQfh90b2DmYaUCZSBf3cQEc9YQyx3jRuuo6bdT+kiM4hbGbj2FHEU+8pBAPwVYh/eiy
IpQ914HmAg2NJ8ieXGiCCAk1WRaYg/zFtIH7jbKmwIz9pQyFzyIYpWtn/mHm8FMIVGBJehpIZLfe
PeYCzDJfMrVdpHXBVz1rDH3nRmWh2u41rc1I4oyzfecZ1/2ads3vCFg8OvDGJBbK2Mu4Lp6dSsA7
wBUjizDqh/X36QNlNae1MEmjLLgZ78YhoLp5LKf1cu9p2Y/KSUkj7AfPe5ghuLEO+RPSg8LlCnxC
Ml8zoilaoPtrKoX+5kSOA//c2GBofajQ87Irw28BgLVBtxL90+vviTkQIT02qQUfr/zC9s9yXGCW
ymcE976e3rCEVG4g3KqTV52mHsH5iM9674LyEkf9NZUGngRlKVCPgBBBWX8gV8U9ffpirdBf6Hrb
jm/CBeb9n2sU1PKkOBPSPZn/kpJuJ2Or6xxSlPchYqkOwMQgXPUiUd3NpEfXhrkLsL7lA74+UOdE
XA5tP1xLCWKixSd9+zcxqmt8siM7M8l828kF/fifAhjCUBr6CJcMmsLEzlksgJE/ysbknSvutQd2
/U65mRKEk4hIIbpX7j3qPhhGSVVC58I9n4ywTiJLF8pM2SOZ9v7B0PhCIguz0/v9a34atAxTTiRK
vGCRHsVNjv2umvK8QMDA5UebJnzM83ds8mrKkt6n3snKzAn0cOUTCBn2qXPrRxCGf/geFV7pbWlr
eKkRPpkDdwIZgeLJfJmWaYFzCIF/FNHw7R0LdnsUVszd+zps+BUkZFdduArv7Dyh5pdYFhvhKDo4
5e/tpw76j6W3GGRKFWVr8rYsPbcHO2A9zLjqfFwA5PvhGwWd+QG/yo+Ns3XzkfeR7Pf35Kk2x6tL
BQzlS1Sqo8WMlwUhUUqpWETJt4L0+Du41nvnoBVMPQ1U6X3ucnszD4ob3B9EPkXswae09Sd8sHAq
iW0YBReZ8Jld+ynR5I4lkQDQ/4Fav+jGK5k2ISvTzNj/w8j5tb8hejyFKHmaV/quhunVDP9toUcH
WPg4FAYWP3SVZIkp6YsCJZdn2WqbwuwkyI0gZyzJ6skNSc4ZimBLYM5AKHkHtWM0xW9dhYQt4Elw
NYZFigXonGQZkol6XBQTldKn6ptDiruFav89nPYwa7uxnc70sqkyh29BRppkQSthNyFu0sQAtal8
YA6jNGEFNsiKCUeVo/ZzUbAvvhESude9FnQiDu7z8fNlSnc5acHvYBh6ddzIb19xYSj4F1SR5tes
HeFQhJVT6QjNyoq1TsGTmDM8qwjqHPYd3dpQxJWiykSltTFXT3Np7LkYx7UkWomB9PjzZWzxS4vo
WJ2h6X5Qwhbkp4glZBEFx7UAqwhfj0/WzptITUXv+sSgnzIC3PerIRqYrMqtsPHIWfErV0e9Foh+
I+m4WN/wS2FYgOybsw4sqG41yEtIFPSBRZHOHgXhZ2ZMSx2BMF+sNMJcVfMHgygPEf2defQ84rEw
JxB+RHwgkmLw0bCVMb3HHLb6HFnynl0XB3BcrhuyVVxfhlmHxq4gOf6WS1yiJvyVYgUr20VQuBAV
mPSKVydA6T4mPbou3lICGXaro14+a6h29EHWhTPd88WNn2p0bXIpp8fJKfAtxCweNHtaxFQuQp0w
LFTzPC/mZ9mp9n+rnW62vQqbGB3B84eVwghuqxGTrxuGiJ8tLpEK/pacpdKBlAlONXLwkKQQLaA5
fR057zb13vimvYAcLx7mfhWDTasg0fdDrSGwKO1i/671HJrOg6SOjC9x6K9+S2673a3C+UxAw8bm
yU2jJtNkSgnXqYK+cYCNTwEFfkJIPjeqJx+Dfwqr3z9WxTMoy8EyIKwF1XNgrJVjRVeJgfONZHt1
qkSVsDFL+dKfw2zaXQ5aWLxuYS/RZTjIF+4IT+P5Woix4AX4NTd4iuzGVetkxYGNV3JgRxOZqUhI
f5shxwOT1ckvUQF56yB6Mczs1z/GD6HVDFnHHEfHM1EeufdWvLMsGlEbsZt15lI8JofABuMQnmCJ
d2FWm+0edZdWrEi7FhBLWsRy9DR3s99uHB50Bgob4ku6AXc0bQygyJVU0+uSfCiygkwAf+4yMXP2
3s29NOzMF48D5fNFiHsfRxBYieZcaioY3AMTV+A95jz0+sfJPHmKFAWz7swjvXtvnL27Dcl6JxQR
XiV0vOWikpV60Z5j3w4vu4tq2gaNtn/b1ObWx3hiK67+hS4cYh9U53v6kBaC0TH+FKoDE6broxKs
sNflCrSYUtfQ5Yb53tx4SyjpC7yTakfeXTmu4s5GHSMOPgknHYckcaXjG1FKO0m1wADgTZ6aDTrV
eST/0URlwaxI2mlG2g/K+u1j4gMWlzkPFPYbcfLfmZQDaKMsDG0LlZqGHwBmI6w2LMosMaU8JL8v
Fc+Mz5wpYRY1PJ9Bc+tRK3QCJ+SoXKojDV09xifQzL51Io+HqJ/5ISICzTZTJc4JxaMSG0I+jRF7
EpYdrcx2Sdy/uRD8HnGOKc7+7FigDw3hs9Nn01p0rII/8BLFl2Beg6GEyNbAXRSg1+mWkBexTmRa
pi3rAHBu4aSpSt69DEiA2Z9a+ORspBQy6uYS9yXNiCU8d1ByT5d6yzBc/BrE7RcgSeT+Z1kBBA/R
2p6XrRpnDAORGCQwrhVkR8JPQr/Xnp8iMKEZkPZZTXt/IUybQPQYP1Yn0k/sTqJhzZX1CWWGEAFj
PEDxl89WxtVVvaxdqMhknLI7zRLPnFMmHtmJsfFHBZcRItLdml+oGWEr3cOHovykTZW9rGLbFaDj
q836yaGmqDAXQm2erOGLCsDbjyUHQ6rE2YLKEep8fxno+tBUQ7ZYKtkh/DbHUyW98DezsgnVKXeh
Pm881YDiQuaP3ewrpwB3lr8O2RGpDEGIzBn6boumBvfQBKKTJMjvVPdECNI1YZQybHkoXQgV30fB
5u77kntcjW0JGvIoMVOnsHztevZYqpsJUMOCAdiVaXoGlxhngbFFksaaH47a1qVQiPaJ9QkHNQZZ
0KjxeqOTgjEbryc+PvF+9pOPef9VCh4bcMoS1fsR2umUBzL6tXWwl1XxwdtEEburYpGWQOOD2hK0
odD7/1IULWXAkoLN5SU1fOW5xudt41qBkTSZZAOT/kO8QHnQLA+Kxt8M9dsnIu5oflO62zY8pSBG
sgkW7EstNPPPvEOfNzqdw+SV0txNXyffpBzwYpZMNAWUKXjjAoLePCaplpAVFL2FVzkNKcGlnW/+
RbgsCNuhYzZyDOz2kXSVogwHV2UNYXYYPCIqjXJMgEMeprIopqN5ZkpUbknIB066mpQwzvSPqWth
sGPgdp1oE72VRXJ1cP1wMoLRfYCiMFZ9TS+gevIH7rYO4H2Ekl24TCFoHpTVJks5BtQaPI6cMCbG
pVpSffIxSRBUFlebWnhSpoG7AABld7v8WI9rKOI5H9S8MMNXvlJafUXpKEMaBYikry2Kc/QxMGc1
t5gSVnN4ocwt3vklf3BKYgqeaDhgf2IoMaNajt43OxXQYhFHMmV9TcMv1UTPCEW1H9MHW+IBPPmr
pr70gIDLKhkmTWEwcZedJuFKW5gJb6vFQsU4BGRbpHg8aYoSNHWjUkIfPRlWebXcK9QTlmSDyePB
xNvCcKkpBuIZoTKnPw1hWyZo0k63fkWcKEYxqu38jpWDKJd6XrHftKCD4Y1jJslzVFmACfZF4scU
cJ5yOm/VcoNlei+YsmGhnqpL+193gMQOM2mWgi9ZjkcYmgV66/zesf270b5FgA+djVFSyqFsHyU5
yE18mA7763LcS6HWFpZFtgNy5+qZDCkdI6moeonRBAJI36bg+0KpPTq+x/W6W1XDqDKfydOR9/93
aSWkCNRtJc8rTlKYP9jHBS/ySUiImlUkJL9g+y/Z3GGAXhi0vYvUMKnOwoMRs7DUuuz0muJVzG84
9LSOxOLuTKWA+VgbL8EFSk8rAfMZRfLujhoDjtPfG4O5gaadQ7o68hAJqoTiFmD0+86L7GsQhR0c
zfKpH/qqk4e1P2IyEvDNEo0KNrHMRt8PXSiMjUlcPbaHRFfMCsT0+V1+ruxJ8P4PsPv9ZPHF5zyX
uUNLi7tT1q6gEbfyjBoZmPRBJAf0rUc3D2tLg7ebKXZOYTSwO1dwRVfywxLyPnE+2rEfhX4ghaI/
ZqW9bRn9XqN1s9AY0V0bAYdmQZ2B4yY2kKMNplwbDIDQQhMi7c1ZYNp9OxzrBcSJgLhCl6g1qlFr
jRPVtYXjULmO3TIYy4LrLgcFUZcWgU1aTGpS5LW5Xd0PcA/UwB7fsnNVaAU7Yxu01S7l7ddmJqq2
PAak6VqXualQgbL6/YU4jLe8QOXwKIT9okq98kIlqx7b0mML2sX7T8IB0ExbahPoSk/A+Om7RY81
uwTodUXSS6ES+OGa0CjebTm7swPVyMoZIE4PsiHGjyqsWmKNmw2l3j+L10E18vM/bwfTtPSawfg/
+8x21XoDmi21PPdlx5LZiV5yZALkDh96iRuou5N7SvUbvYcFe2dJ6AUAzgzPzna8ghAPUHUmo+x7
inFzyfpFWtXfl1l9jlEKeydIdgpl1PaQRPu+xGY8OqYGIADOjoa0J1GGUAV9lQyPbPwadI96kOiG
hcLBzvYVnT9UH9N3C9hKvLRQvFOYwRKufGLKt/Ee6fxzUBth+yKfHxM6gqGhKPFldiLKgZU8J/L2
7opt0cnEbQMyrhgDQ8l0LD4IL1jL6NyXCCPBOUhiLMPtXhSS6RFilOYBkjz9nyWJHM6htp7pHeSD
sN6cZb7ayPiOZHrRY0l0QGXfx/CNNJf6sKiJ+rzcy4FcvzT3HbeKb3Ca9bQMfFgQHZlOEt+tRY/I
EHy8DHaaRWBwAiWqC96TqDE9M5t5BfMCAHhDSViUWWOKF2tEKW440Sc3tnKKtbbdKIk1P20ZVsSm
Vdv6TvU6AUXZiCgkPBSHyoLC/G9Y7R97UbowKfEAw5wiGjK/IAYMPMKOjBFOXZoWTrsLuHp+uuKN
OnbNjBjl2D02MdCybutnebEXePc+PxyvepF1So6kLez7eWbnuqQR62NL9JM1eAAFZ8AFX1WRv98M
Uk4VuTr04xFLtvRJ8evgc5kLSuMstyfr3k9QSrKvP+6TSWCbVPgLdxptkr/O8u4E0658mz1uv2kf
oH+MiuJgPz1RGMKiWNLmr2WLVMqk4z2AKGv7/QG0qvkyzVwUsVOobphoAWJDh8eRzhxoYvqf40d4
zRTNX6+fsz1vOWqrcahRwkWeVP6X9NoLIvKRU8fQoqIXOAm9VLy9CnCa8Q2lcywkwCszLQkroW7/
giOieGIIjC4cbTNNHxr3nntUeHGOuccmqZ5bD2KdJYAKIOJFd+K0fMLCZG5sTMmGVolHras6tNSO
3zc1g+cRK8fGyEegGq+4vtp6iWPppINL8AZ4DRP1cRk61eIasbsu9yXNUeW62wTYFJ+gwWGlbnd6
8SpbzrWnBWdyydOeAL10yB1yJn6q4NnTc3JXR8xsr7XINKyEw5nM8/uH2bSCqDn0xdOiX2uBKz0c
Oxd0zC50bwbnaxukBH0AbVc43pa+Zyiv2XFcNjwVrBiT6h1Ad9z2i3a7DE98wWflRoS+9wBofsXx
/KNZREBTnRCrMloSMyb0nZXojuHo7oTK/ye8C2FCP2beIBhllcUiMcStJBu9i0P8CiaX1TRVZbi6
6kC8+Esk+W7VwazwcrEqa8GpNCgkbAob3hPK4T0t+XKJCwLIHZPMJuEVcX5e9k4+REG7EPqia6gG
4AFEFiS0nXhSzWSSy4LJzDoq/NQKlXEwxPajyckzGj9Bzv7yyMxmyPYVFvep1FWDrtnleZklfpup
cvuN8bSrBwcsPha0mOO43tdZbR66bJXu5mnjY9TXCmGDrPF1nYkFDGNnV0A0SOfK/u5OhIQSHzmj
AIsS5FjDd+SV8xVrRfXeAa6el6KF2bojUWXiQ70BFQvL2HRUXDu3svct0QDZjgRXm5Fha0uW7JPd
6fT5LPjTrqpl2+bn7fpbv0MWMxxNa+cDlH3gRIeW4DKp74fcCFjMjbVMPN7jHAZ/QH89W6x+i/JQ
AcevQMsD8LQVys+/+kqNmRio3qaUYzx1drLugYORqYekVQPrxYXS/PnP4gyCuc+hUKmaOwzvRhel
Iuf4Xk6xAtSrXTx/6769wubFft6mk7bO+t1lEqWmsKUDTqrdJ61xqEUOh7Tb+HCrLlxssCvr0LWC
ByQ4WPmEr7m3Unjl2bbywPEraOrex2oSs8Pxp3GyXTYCRIfzWgD3WiJnL+rQ/mLgyFmSLTQ6hxu1
uxRifkT6mRW96ASnPq/9YkX3iCHVBViV0L0tzNoyWtV8Qvoy//JOVcfLBNWAd+YyJ0VjSU88iPOc
pjwMoTl9EAAnZ6/nqlquCvphv3j9eMoPdKf98/dxMGKp7KTYi/GZSX8/xWhNmJzv1Gp1LqRxgFiW
Ow5wvzurzRpzFIeZH4XM3Lz/jKc+D7/HaUPl7XmiHVu2/y6mrVPlzYl6nm8CFPEGS8dej1/UQUqT
qCtjG9l/4ZBkOR7yyE13wGlmJrqKfFLKhEeqXZM51/1XUnwkSumVvNs6ehM6hE2LgMKz6dFuWFWE
j+kI89QUFDH0HoPjSb0h5JIp6OGmxWVYKARNZm6zMOe+kqtSrTcXUJFKAyFKYyQLhnWcA+pRn5qX
Ykr9m2FRd8Lr5LGtgUFknzTcMnJ/xUgsfpdsJ9RUDsQRoOJs9AMCOep0sEcEFf/F7GRxc4UmEmH/
bY1jQ0qmIUnifOrLddXBHMmHLY1RTT0Nj3vPwnVk6z3F9ztQmaR0M09GIeAYwutyVxy+jMsaNe3f
jNC0wYhdRSMteGR5ArIfbyWj6c5WvjqMZL6jSa6WD+uo6uNND6Uau23A30vQV0YRM/LLwpfY6Mjb
hP8+ci0JVWoCqDH2mFWncK/9AV5/rIcfhs3dr0wR+RgZQp9WIE5egCODENsqlwncVuFIV+nGp8wl
EQAN7boTyj/yyMeZdxAOtESFLQ7K/76CSQ9lU2JArDQJwSj3beB3tObC+Q5EG1MqBgRx67LmrnOl
fEGyCjzc9JZ7tKRcgwqiyfnZznYFUCkcOLIEGasDuczckbs96UPl2XRfUKcuMAywxIW1BX9CW+6E
TwJlzJYwL57HnExY5iLYOg/qEqLq3Af5oUQaqzkt2kLF5ot1YJowXwG7oUlvm/fPVxt8ZLu0vSfx
7AXAi2eiHrd8q4/Kgf6sEmCh7IcWrIvd8vgtALWws5G9nepG/irdMV17GLm7oaD12GUOD5AwN9ha
5SCjLmhPVn0Uv/eF49fwNuem1YibHo/G8/85w8+7AL4oa/3pfQTfJBgpYToMMDigL0H67sF7eMOf
fSBzeJYd40bliEy/pk2TzZN8aibDZAH74hvjUygin3bW0kl/kn73pvQKyZeLmy972eGT7S9s79Z1
qnproKc5aMcL3Kk50HSNZKfjrH3wpZbgoGCcrtXKGwpuYDHmE8DOr1lBMcYQogjZRFzrVs6x0+9e
T+MFLtMr/1nGEIe9Vs9zon7Yr40oU+DzWByAsGpiydodrMHbnnpEkZzltj3jgYOw5Re/Id4tmhNR
MaBZUp1vn5OM7a+rcT8odLdm22Y6l9Ewr2c6KuM1fFj4cyp9Jtb9WCOkfEED4oK86S1kWwIDc3pd
7uxpXuv13e3ck65sDhOW5+is/XD13viawgv6ZqcZmSaONcDx/X+zH4nkSm3+jzJg0UL7oyVH2MOC
p1rNyDtxkiuPLPZoC8zHigrWYSAlZgAARLyp7naSdyaIJkWyT6ycjWBoD4VWYxc8/Bau1B0ZPAMU
Z1Ato1zrYZhpMdHnYunu9PeXBbNvr/GRK2p001U29wdE9GhFxpaXhOkcMz6hHxu2DDcg5Keg4u6B
3Z/xuLDkklGgkd4jYRHoW8JdJM+oMQphrE//nCRilAZ2jIkbhpoF9qeCPEBbOlG5U0rywM6jhtJc
fpAPaBrtP8sBfASLrTH34vSlcQZWDcKsSar6OKQeqOkpGunYcp6fI79KZnO1DvoMbkH/Go/2cBy5
7lwYDfrjoOxrnyq4y4xSLLNGm/2AHCrj5MTmMj/2Yuh72sGenX1vHp6d2WIrNqAvTol7NCsaIZJy
IDMgcCJVvos7KdxiYe7eTR34LMrlsV/WF7YqXOAy5yKaksl9/xwyM4CSroOIYEP7SMddLMA6Ir9d
9IacLY5KoAYS8U1AfXOiCVPZsPuOuYBaRlX0EvuuL3gEbEuUdl1re0d6T/4IQZ5gn+irzZY8dr+m
qcFxcezVadNDk72qfNFHVySeq+/AfY4yx65HiW0k8MPCgqnvkOURAnTLjoNvCWnkge81BnlujWn2
l62XTykYEdciZ98CaZ76JetisX5zp8kDSRfMoo/ERkjIVUG7SqMQh6OyeEiNbPSMiEhw8jLH/h21
R30pn1MrXwbS2yypZDJi4yZ1q4VH67Z2M6GocL2UVTg1d9bmCJtMO4BE83a69/LpRe6KHag5I6ei
yauJqELZauHugTOe/xuaVoYze9IOFYxCUKlRRt18ddErpuxXMBh++s7T5x65THk79Y0Ur3IHClq3
gQpPYkcfXAMVs5pDDGxOwnbGG+fMhn24ZoHq61cra2cZVzMLXXNkFT9l1a32xKEREXQhBtTAnPg2
2Yl/eRHcPog9rcH+BBbvG+qVlme67mA4mm87y3h9xM3vkGdu2u3ZsywhY9WscjbYGMZ4k0r7pnO4
4VXO5DzvFi6zRcH3GgO20lpAe0NhjhIvWxA+DhOqaWTu+xDLSpPjvh/Z90sRF87qmBEh8lV3pzJX
Xv9DPEdtk9tc21S14wABkjG0DjGQJ6Z80y2/aVhK+tnYZb40I2cwcaZdMh/6+YeZ/9tLIyLBOar8
0EZPW6a080UkKKImBnoCzJa1/8YhCOzWKWJ2NBSYWZMzSRDncL1mbv3XgeX6bj61FjvxdWUYqkEj
Z2pAtWSIChKE2XhBbQ7SvDmAQ0+yFeALGM0j7uC8/bHUBDhgEkA5xJieMO9SBE1qBAL8bLIAUXZC
qeYVdWGXe4LZO0d0kvkMPuBF587OkMXLNt4vxK3+V8qpZ+AvtNWfPgMYHJ5aCHaOnpH+Lz5Uuvb9
6eaGkTA/9et/WfTujJH96WFle/9CaX+aki+ErLJDFscz70Q7nNaupzb/4cU+wdl3O+Y9MTvpZxsn
j8iJuVzoKg+5qb+m76+fqQ3+IqBUahulcpuEwtvrt4TWrF40WA4nHHHa1NMdBkmYX0+SUmjURakH
Vazei21cCgBeIpGFMR8ziQNMhZq67RDlWQqOwb3PJI61IFpnArMg8F6fMvEhbtvlqcHiHPatvYnY
MM4YxQ/u5wHnpJ/8BqNbc5P28S6FbpS/hIRkNRofObD352K2GHj25FYM8dCNAs7RzvWtuaMMMxpn
OHnx89UbEcz6nGRwluOUeFs9n9VVL8NO151hSZXO7j3Wm1fjI3YMCxP5UIU2FbzZs2UKgEs0Cb5X
f8GCiYD7Ztz2/i0Nkj9RltwpUXpLxYTqVQVkd6LE+kShyV2KBTbYFfEsSzRUzSrC4LELcmBbai/V
JFie65C0jrfS5ZmUrg2R9mPbhturBGVeheq9cLRSebTg4wjsvzpaovztBziOrkkMFiTJvVN5k1CT
gFu6dua9KtmVzXKNUEzsf2z+ghXecH67BFG3r9g/wEsbXiflRf/BTFidEiKjDpYixFO25Sgo1vcq
9/FKRcM9lNTEVGrdnktm4MW5LjsaXdAAHA033Eo3vb6VJOv8sjFaDZGYDp7zmo6QSVHSeDKZ3Q73
CkI/3/BEFXbLFWEi0lXR+3HY8/9eESdLklCKyMqP+qq+fCOBcT5HNjjc7axBEJgQIQIuBgMYUBak
zbsQ4bBMzaR+UHwwx8ZLlkxTDX2dSfwLlN1ePLORrtRw+XBZFVcsjq7nptlBukLyQ3KA68LezZgY
98kUx3mDS1F4nmqdCNLwvEfHs3e8Tyk63VzpaoRY55jnzFr7IBhQfwkHVcZw9uqZq0dQt2AZZyRo
WoGuTTMMEjKMQ93Del+2kE+0c4Kx7pZL6EL8MxaNIzhqchZD273BZ6ox+u3zsAiJRm+DJAQJQfIP
el6MHRV9B2o3ei1CDPe0f2jK74r/JhRwjzaJGfYWPOOJXAsWh67IxhVO0hGbqLSiJM8HHwU5BRsc
OF509VQmGxMUSw2BTGPZhb0a9Drr2Eqk3+wH0pWaqO/p7dC2NdpsOalLyawmaaLBe/IauI4wSTl9
TXajYt+fsZyOXMTY5J7UjYM1kSfwhAJqgYDhqrrskwtdi+da/HNX9h84pUmv+i0bavwgGBpl8xTR
pqpjoAOMs09EkiYwTaTG5oadKWD+BSURZJ2ULCZcURD3I/y2HWlCWmW/frcKBfMNuLxZdpeHMTKG
dIiopyAfiXwdqch5c4jvgLMEX2W1jfm3F6eZ1B60RhNeO/Nh1ctKeBPwqZTg5pZChGBlI01RZwof
FWbhEPkN4/Bf2x0gqGe9YKTnjQEZJtIt1eSZu0IanCyVDT+Zs1sASvaQB+v5F2nVf5L5KGwT/g3J
iG7lzSAZPqyuzzqhh5hxgZy7BzDr9vmPO0CthyS2ojdC9r/9RH3/CvhhgomO7jHN9gZT0/fUCovR
LF+7GFgAEbB0h4AIgZM+hq6XFiri3jtNisqbrFK4O4k929CLQUiB6edVJ+25sn2XJXYf8TOpSUGN
e1oCN/jTJHfZvHUYZxJvw6fu9v/whGfC9QTOfQUj+yJOYfPGcWp/ouWndrgVFMoubYYyZmkNQZmr
kTDPO8Ym/WiOXfW5fsMQ1n9e127FE77W7iBToHtxAk559XWkta5YJcaKAJiobNCjmLlaG5ibI+OX
gB9MUUUWb+f70+xKUG2vfKPXNFryBlPO/I/eQi9TmoAlAZacYX16/e0bR7bursUPJNveKEHA7QlO
dt+7sIQ17qe476q+thNfjLeaQAR890MwZU5qHNtdZbJ0NvJ4IN1Yo+g4+UZtgfvuD12JLWRSfFTw
2aH6BACWfmY3J/6mzuHvKclqlE2LRxy2XwVC58gxiLikFciAKkGgPqo3chMT2VN44iUmzutyTzpO
RVS0Q+xjBhtIS9ol2Q33ny3OQU5VuOm5hCEVel9qMZ4c6dG6pX1fgdpc7oX6zcSPuK2o86K3AwA1
wokPGA2HSDjBbplRBqRw2jTcx2K/QYXcmWUfb57u1SuwJzIIAR1SB9+5NK9yWtG19VXwM665v2KU
kPDTf/sdixRqXtKaEylOayVoaOpyW1ITGdap5oMElN1bqmu0gclXwsRprOgFnPwK+gyDwlOh7yAr
9pMF7ypfXQEtEPH5N830Z44tJPV/YwZ8SuSuHtxm1oW/7b1QK5b/Nd3ItC7mg7KAxlGqb6r4v4as
kPxQTMaktp2dBOF9DA19CWNg3aDDEORdmV4HJ3kh1cHRx65pbjH37n0DVu5eSUijYbBfZBmX2CS3
E4L5pAjTRDgOEUa/Y/5nFvwTsx1l7kSfUvpvgRCHWbzTRaLO5ZwtgLLJ5a0oQCLY8Tz91kcxjvDD
T022aG3QpcIPQxACg54B+HLCPYYSOpKKS/BltJw5VwKJWsmouoZf7NIflwtyWqp9QRnpx5Rf6l4r
/vM5H9Plm7ZActnNUIDCRIP1vFzjm+fcU8douCgE8r//2MY0R3tpwiqK2ljpA3gGbFhi3FG2yTOo
qSkGgTczxoBTeuJJ/NSVY3iHZBALkNu7E6XX7wfEl1Bt4dR8drF0wIzjmK4OXrSSsLxWWeY86iNZ
3BjtR2mq43I3Ot3PtD0dYt7T1mxPIKLnR1//G5DteP7Jz9CU2s4EtcraeNcChk786hW0PpDutau3
WnyrPPFPDN4ddkQAGPt+hHlIjZQoSL0a1lY6D77F1js6Kad6P+ZlX1guTJAVHRbpPohCEVwZ+lgC
s5c6qppQvyib9bn3tr6dhFGVTZjsXYSPx0Y8UHwTF4sgu3lZUROZ+dZ/MStkLELHGZE57Lr8Kcem
p/TPA5whI8AK6OHID30uNDLiKZENg+Bni0Dd2RYb2cLyjztRDeHBFVeIDXGdQVIiK2tbmiWb+4D8
kMFKCv1ml8a6GvqcM9ZPpgRWUWjMWXzsUD9nrOFYXuzSUaML6xjpqxDNnfOS/sADRlRn+3PwDZiZ
HRy/DN53uT6EyIsH936WtP4bb+lx55mrvtEQ0nrhQpRVJbLMEUxL33tiXRsGGPzIvbHiHKDf34n5
juyvrA/eSSqCpy1dZZ02Yx6dCqSJcyYILld8DRiYZJbnWPmpwGbiLjeJyDFUxnrRLViS91qAUcpc
J0XqaKFvQRRwRcatK8lfK1b+0k2GbDgOc+esblVw6kKg7KneBlmdzCSSGJe0YVY45jORjXTmXXQM
zeQUMsxf5FYg2nJg6kfKqRi/TZwwWP4T4Cg+7kBfIu4pIJqB+V+Pv5K+CdK2Fd8kpUEFY+6pULkx
orMWOorM5W2uQj/RzSVTOaZdcqe2BSLzslRUfNKtTWctOJ5LpUoRBJrsKMYZMTeIVZ3trriwzUM4
eCWmOTy7b942vULEK63A8K32Bu0GAI0VPCRvNElglRG4z3NzISlmL44Jb9+rFE4E9udqXYdaSWgx
EyO/ldgR4lF8G2XzNxSokWsyHDxAEk3jlyDGLntpfKFi/KUHfHlyWn+CwKII8ZT2AId2UXOzFoJ1
X4OlABEji3dmwSl0O1husvJEKi8sSbqncBKL5a1VTmfrSCTNJkD+OCY2o1v2hLeJZbHP6n91Uc41
ANBpvRxHKZe6SISCrtgS9a5T5LksgllkdLuG9xsYDi/lVJWhBn4qhKna+PuhdH2dLSuxYFXauTCD
fIAHdDKSTigPYx14C3w81fxYATJdur9h0zicOpyYBSUT8s95rCsJFs1V2ATOzkhZ2DI/MlM8XRii
H1ihQMOINGgCL36RcsBDg4DZ5ktjfsXW5U9GZIC3Da7Zd06K2vUupU4hCG+Wny1Y0H9EFZRgo8ss
1B5bC8hxtaPz4OXIWWnvaeceAvo72qa408RslcT5nSdo9oAmAwEklj0rqFR32Op8IHPDDvv8XHAX
wwUK3egpsuGr56Sx+4FR/x0ckOYnNk2JAjmahaIQlxLWkDkyYPNRDZ9e1QW46LSrpoVs80M448B2
cfr8PFa3+cnay7G7awlzYrAn4jV7ZU3xvshaCiGiDsWziJprusOONde5Xoe3jVaaHOgdhs/aLfZy
uwUSnI2ifjjI0p7wyWhBhImgoPewj5lQYdwwHk9l5k8q/R7vuN3XZQDV9OmbDWuGoFAjlCcRm8ru
OdkGKy9mXV+7+oXlm9/Osu+tHiX0aE4nez2n0jHC8U14yH0+RAwGW+z0pjaFw1szej7JH12bfpiN
UftC9eyQDbFoqMCdXZW6LISYuSldqaWNFCgyMNyQICYMOiQef7Gyl61NOsnjQ9LFcJRSJfcu/2lT
ujlkAWyIHpuBpZhrUo4TQCqMDsueXOihD67jjdyhPqlIE1bg7TMhQ9rQDSYE20cgaWPyH3V2hk5B
Fzev232uLTkUeg0XMTWYei9Mp+Ootn/Z1GbIS5X+7M7iH6sFvGpwhtm/gAjWfSIFW4EmO5FDiq0b
2LnpfE/vI7LmiPqKOqfzPI5rYgoe0DA0m9UTX9U=
`protect end_protected
