`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mbiBBUsfqc1SGLY7a/gq1nRfo9EBTydekPlUBQTEGHJOp90YH73udfzIg5YQEUB6HoDeub/m3eLY
3cfJtnAUYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cD/BFw//iBGOWm5BAe5qjMggWUhbsheOL/t0eYjiZF3YS8HkeRHT77riAaMjwD3UyV+wWMnrHKzu
7HNfWBW4kkRUPB4J2DPyUbUCRXrkGQClwK9OttT9J3KugHV9QiwozfP1ByZ2pI0w05o1tnr6F8Wz
UXZOnvAbwD5e7DU5TP8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M0QEm9soXR8UVwsZd3+1TmFyW0B+X2X3J1d3bxUkPejZndE7g5RKYGCXUNTVVYVGWdJtSPKXy1WB
xFFOi1bcMTqPr6Bgu+vmF6pFDv05fw0EeEyszEG4gFHuZLn+icGObdE0e9cEuyU6KU4QCwbWpH6h
DcNZ7xriZwuOolkUNaRJPf7C3X69RUYYLrfsPPBANRsj4V4/nfO3b8pXe6Eeib08tyHxmXDEdnE1
VFqOyPIA7bDxXyVaAviEME71ngSGJcFjJfdZdL86yELm7khwt3RA8iNS+j1g4sfIMZZInYJeApJ+
n3sTJPtEBjBXwXc9+Yx5hwX9YFapwLEwPZGJ6A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
svPBaqpf6OSldfu4j4p8Asg+UwedAfikAN+OulpYtIJTWdmRWdgzuqobRHOvGuqa9vjmC/Ci+1Vk
YmUbxzGAwnEokmmsp3z7sDtJlavSCzKG3RqSYrdoGscFBuwhZGLUB8gqLQIvCZmhtGeAj25rJbb5
auJBKmQRQOJZzjhSKes=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
l4aZSnVBb+9gHXXwaUcdvWmraAog0DlBwuis1jmnIBTbvyFP8/m501XDc+3iVOyD6OM38n1W9Wbe
ciUZnxGe1xxwJym56P0tb/BhYPNAYu0ephNZkvRMm3pc7w0UIJZMtSuKKYBDc2LpZ3zjC71Rtpxg
L9n33wwM1GRbYducLIqfPxj/YU1LYavMX6sELaBdbJDz0N5NVwffWSuZpSXpQrtOrnBlgev2MnHM
vMahBfNKBJZtQGrynuwkigeUUMOfWklhHFE8j1lVJpJDs3Q8eaS3gDJwRedmF46J5tuNk17SMywX
crijhDlRZIbvfbVd1G4qrg1ohMNUSWZBbMiZLA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1517888)
`protect data_block
XTtq3y6m/YiVBuV63+BcSvKEAcRTPTIB+cbq13fgKGrK8r3QJ2t8Z0a3GTRdNV8R6KXmg1rZ/qoU
R7cRjynPZSfHmGID+AvAKP5H3L85s0sBtNLF64HoUdM3rFedJtnkRdTMqKG5tuHejGzLroWTr8J4
Gpz8D0bLC75lpcITfvfPvzuaOydV/36nhmrKe2Mmb+BFxXrTAaTyAhaGcsbqJhWiy9MUblmotW7C
KIo76mIcEWnLul0D/O/lfE/heG9PlFhpG3lJ+bi1vVIKf/yXUhxx/+xWh1nw+4my7cd1qGDO9pKL
1ZdL5/vTsC3HS0EWLO4pb5Yn7iQY05e5uWGP2KicuI9AZ81QxTxOz+KUFkb7rUpaochl13fAnyPd
thKW7oEYgdQOwvQbUksHUls7mCBfXuR6T3qkgdNLE3Mx9aA3j7dVaeYrVzU7QCYjyaVTLCI07eZp
NpRKD/llJHl76TS0MB32iVwQs78JHXjRUpv7P2aLYtGc44mDIBJOTAo1T49dOBUxl9Bj48P+CllM
4rYsRLjIwKdlQloszayP0T8jmhCxVKtkLGZ3mGRbvaWpg9w3npGELd05JdrPZWy8E9urKoO6bSKc
nQTefaNtX+KKktdtfKZCg/bH2FUjhF9z3QSEhMlVXUOmmkvPmifNqFFP3eQR3GUmTss+ZwyNKzNo
J/qdcKIGbHB4VY1+ufh43heBlhmHb3IoWvgx8QaD4mvJPSUNJfCkRdrjqPd7Vx4XFzmE83CWqLt1
kTY9/mmaqkMTAUmu9nbMcnvUBhfhOP5thLSQttJ1HOLrx6xPqYxHMB37ktjqWDflbCT8IWAT2Ai1
tzgwl21B87MSr2DNIkoS8pcZGyZkexa8MtB9Lo6EHWccWG5sqyZx4RQXQyegouKxn6rlx3GWqkUx
WFMGW2zWW6cPuEFs4/9AdHPelI5MyQR/vkEd+U9ZGfLupwo0gNnklWUNC0nV6aLCqWGj1UQhZ6XB
Joxigt0BFHVSAXimPq9niQYl8vIbKkuA3DPoPpMtcFi7DZWc/YxrnuvdoKX0swwGUb9bGZvYKZdp
1q17Ar/Yhd6pT/giHhmwUZoajorLdEYTDG3CdIhoOJCCW1zrkt2r8KGBS0npvcZuRtfl3X+VTXOW
3fCyHNozJaUApF+sLVcszBayQ92y+BAYZ4HXwSuBJZOfStZwWB5O1npG/a12oZ6l6+vYnGkZXKQN
sUb7UkX8Dvl+hxZmU+sFPnSeBm37+3oE5rJ/Q81kuypCL1Eqs3hxSBntDRf+SQR2ilGfYxI9OaCS
HuGC3yg+nboJyRqOFjnl9gzSnzKeMg8oAyi+8R3ZNzC9gqaTE1FiEKcijgbxN+3VnWixdypTl23K
/0//dCkla/oj1ECaWU8EF/GmgBtTlWvRB1wDyXJqrxH1sfm6au837lCTia/tAl3liUUhVuV6XdMR
lWtAbdzit7g0bW8dapMftkbZA1t2xPixDUy2PP1TlB+20y/jqEYVo0lHR69wH+5S5cINbZUh4lCG
/I1Qt4X3PDrXmTo+vHZQb3cVkOTf8pqSzzhSKCX5Sil0bclkxdnO/Oq4zxDraVOBuh4kJneKlbuI
gFC0JdIctPJuv//n+kN/ZL2UY98kQYJZ1ogy2KAHYjd9yCph2jfErNuwg10wJ20TrwDNVvgtAona
VmrEnlszUZAGEUkTF3zt++dO6qJ0Di959qutuyL8/wzZSfQEVWevFdTYBrRxG7IkKn7lVIAcuDY3
5ADOebYF4Pjj7kouDUqvBk9p2hykp824P9SPGPn864gI04WaG+5u3/hRX+aNYdhWY+46AIGNXoL8
kc3os3R63YYIhAmGz7vE2ogAhTnhBJrwSU6Sy1/ZaKzGeAn3wLGp/6Jl6PCyqOqsRo/VHpA3YI+4
pImMMz4SZh/LJnvFRDoPnGG7nhNy4VkJnNeU0qQVLiyOgR1mt3I+/lkoTaGjy0BzAwS74w1K1jQ9
kCxYnTRtWdgjMeiQhPdcjdOcpNjl/iuPUP2xK4mGN5pn7r5VCiMxd6qCRCHsh1z5hRVU++3MMhOX
xd8W8TXSmiabPo1g0v+E3odoq1U1QHq6cTSj5DqxwCe/lA2veg/B5lFoxe4oVKDvsM3ET2Sz58Dn
X85qRhwdYCSF3JK6llb4P+lv6IVCduz1HO5H3tTVBhTc9WmRxE9cFQohK79y/w6TLzWLzCc1VwLF
puQlhcjEsCBMjfBKWE01tyiOYhZv/gYK7VfejJL+f8iGT9bQ3eQNERRg3OmsikDGSaGrM9ETPJmb
fYegYIjOby5bd6KIEzoog3q+JJbaT0H+Ol2nV+GQ+Ic1anmYnflYox7Lr2JSVNa0vOz2FGG+EN7k
ds73YvXC/GoRyqkBFmVGP1FsPQ5tXYTsstcVRfL1SAAuu69lP8dKgcCBMIdKrWyJ8fzJoDh3sUVV
Yr/+gDWy4/9D4cBuEp0ti68HRCIe22Sm3d5TGytnqMN7MSV0Yb3v2KDNudIkkEwwYboXfaTfIvn/
7VdrwO43PRnbAm2d3EvLfkc5dWah6Jl5DJSQxhelQR3G2lh9ka7RFeNAb1dC7vxVYFaU+wgE4DkB
YVYaShqOCYmzl0jhQRc+xI3mRM4NFHmXcEY9iRvGwkvBmvB8XHZgSijZLm4AGaymYnaAr5eO7jtY
uj8lrLoKI/zpdVrYlERtln1hAJ1azgv5otY16bGV3aqZ+H9Kb0coB7n5gtm5jHP2uuQscCKVuTDh
25aI7kLaVEjM/jcQ9cJR2OzZn9Z1xDzDE5Ewvt/CI00txsnb/K7Sry82dyNwrj8h0oZ8NS8SEvo7
9Yn13vE4V0PxYjduEhovaH5Us6CDP3TnfGWJNhKVWmjeE2d1PIcSuhS4xzSBDhqToxLbJTurMEIO
WbbrqTFm9lwQaq3597YJ2HHoEp6clj2kDDG0QyjPA06E9qnv+G+3gvTVTGprB5wbv12FVe3eSQqY
2zRJzBSylrsam1ErTsS93dyl9hauEbmWflgler7Riwme3zZT9M8iJlquZaDn/ujajaxxkdINJgx4
QLEEJdZc7J4/Qlb4QjbBGTaFkD2dQ+xnQVouiz8KfvoEzMGKuLI3RIhGrZOMD+Fk0vL1Bk8F5RoA
9fSkqzMoPX2te2lgMABjbxN/KHtO/FNMX+K89gOWgjFWlRduASugFH5tQNsB5XXpufEtSoXh2tdW
DEkePIUodFlQ8PU9CXPiUhNuYW/Lhluht1/CcG3yxfWHsdmV/TnmLBqJT+HkXjFaTvLVAZ2SfUUj
RLIViPR5YZ5prAe8nKN/LZVbkdlsoUfPpoW8Ru41riw8VH2cZZiPJ7y7B00UFpx361HpzYa4Z9ef
1pEGEdKp9cmgKCpWctkRWMk38LruITCMH2DHBgwlq6yCHjsZZ7hqDMdC0v3/Bf4obUaufq6RyFrC
Ns6FYOcHcO28nXEqgEr6nYeIIJnq4xkX9L2tnKAt2EYZPIB3AE/E8n2eHYk2eE5FOXcBX4s2pYmH
yYmbqSnmLRz5yo1x5/kovA3L1L14MWrR2ECsODdeNxr1y5bvimrXecWsdel8LtZQcGLaDWggsrXC
AZsEwdjqI+xesF9oS0Fpj8Xor9xvDFWbG9xKEy7tfYiyUNLd1neEUI+iixE3IF2egYCO1LNQ4AXo
POdvFfb3v+zt//FFWrpzDE7S5kREq3GCoLOdzrfsL5IySIuh0BWQTAuzNwLAN2aHqLF6DSblQ5JJ
DW2zsrLcjtkxlTqlWn5EhrtVqw5Y9iI59LzCBGf/UTqm83PgulhW+hEQ3A6Jh5HDThDv3kuGjwQw
svOG4bnG9IBeVSLEhYYibZk+FsCoSAgvASSjjfp3fk455oHcPss53GgGOX51wFQ1zD0G/KSdUFAv
vzHimv+M9HfueFGs1jRviy2ylt72Ccx+0Pf/DVaGUA4PeTJTUPQTjbwfff3YHIXonbqP3BZ0uOW4
hIFGKcs+0zCpfw5pKlwLUPUq0nxxBM/p3I6z4/XLj+hoSkkGgTfNeqzsFjxUgaGQEESoC5IgXk2m
vzosLacrVn68hiV/HIkV30ErvwedpEhYsmcu2HVTaAGw5hFhiECI2RHHInFQfEpBuj8oEOEVHBSS
Y8S6T2Z5JIMKa3uYuD4VU4KUeXHTj3XCF5PNzaqlOddSnYlE4h18uUxFbfJWbO1yr20qop+lyf23
YvAcSv5N6mjJPfEUxkTxmNLzrVW2ZB6oawznmIV72mSAXp9bOtu8QOAQrfR/UbrChCCMXGcyCOHo
HhaIsgqhiaZsHnkJSatMmlZcegULABnrmUmgaoD1dF+SwcdFoZRa0QD7c8quPU5+a3aN8f1B+qTE
uuoXZ3Rj8sGLDDgvGeTCuyDIW1qfxQgErQ6JkKM0VbpLkdt+j3by2fqhuQk9b1FZ70VuTsD6+lfR
k26WlMweXGkScZBCYFRXhgslxAeJ2ZV3RZOOoNphc5AvMw+ZDtDLp4t7XBU9XO9SXsAKjdi61mvo
gdwxlORwtWwCgmyTcfgeMW6f18aEyvBbYj/LhCOWQSmUV8/QyG60vgTJQX/6Wd0853hN2yzBwzBt
OrijlDTZbazUP2nwqrnuXn8vkPy3kTUAjN9/W0yIYBsm+Ki/FLXd7sN4PC9ldz30KZtEo1/sRdtr
K1D6+mLMi5q2qXNImjZBJWl6h1vdl+OQslrlpTlrVboFrsijTfQEqkoA5tHkefkNxvGmjAC0icjY
SR6QUPEvM24wmYy+Rg9h7X5Rgx0LremwwNJrfvduTZAmCBwEFQFseNtU0FZgA8wKEOMDJX+L8Jls
78ieSqrDyOgVVxexTcS5uYT4554FsNim8oC2o6Qz7mjRWExRNse/QRjrJ87x9YHo7EHV0cORpMZ+
tbRmnGYffDTWdEOVfTePp21/2G9X9LS9ZQPKqQnJvkRuYlULW8Jh6aNa77vgVLe3DAA2GFi4mJzF
+QFHClwe7tcZ4MusGIVjbmLHNCrSjMbVr5SY8LVLD4OmoxFThjq8YDnleBHzAzq2nzu/Gc3U5rlp
QUqZT7xJxc6IQndCFOjdFbVxPvvrXxnh63f9MxhEG/AmpcBL2praBYaFiokw408XYW8HpSd2wXgr
1KqMtetXuIlP1cg9VgcBTHVNWV8Z3GfavIYX/76+NeY2mylOT4KjIXmbENFsy00XiUc1YBVccg0k
zg9YaQLg3LfJ7T0mCUWnNZRhOdGOYYnNWn/8F7HtLPmV48Wzjb+ifM27uUh+bc2wGcr/8LLeuUJg
GKR/dLqex2K8FIrRGTIf5i5PsFbsqidtF9jz8uv35qNTB0hOO8OQE1Jtn7npeV/+Q732ingggyt9
UyU+5EjNkQwHUyIxMfYqsKyFW+pe/p7p73Lv5YwRHYynkU3vMF/f/cCJtzAeFnozGt3TarUoZcNv
O309JPVq4qk1jwAcAJeZcSs+aTGeVWn4co6sa20dMs1ioH7CF0ItOVXbdGNF40/agNSILgTx1q0D
KIm1wRKgd6efCKWCxffxXOZXkD6J0aBL09vamCEjepgIwJJXdB70UxQ/+XywSMRt29KfDkWO5Wey
OlOBDRcnUK+1WvldpAFxkQ0YNYNWQBI8J442Z6PymbWR923pwTjKuGDuKpb+9F0si8UI9gd3ngzz
ZDbn4uBhOhZJQWudQqSh55eQQlrAANV8wdbVtqKZoYutmcUBaoPwzSn5/giDRvYbkCYnBrAF/bey
+wv6IfZYqaUMeSFGYPhr1pJWsCYX9ItTYjuFqAfjbKmuiF8HB+Ol+pwd+bwyBhqIynP6kdb7Ya/6
dYlZyF5Y+yo31mCfBvmrIJrORvtDuoNKDUb6pNwNnHr+VnyI9Qdt7qSE2HdLuCVdATTS6nzgd+5c
KHlsHBbxPTfbHs1z9IyoZkdbw6OF6xNDDsGkcfhp3cHe1dnmE3MIkiYToHkHARX0V1juX4WV6rYt
s2U5CLB2r++Q6URFHtJU4sYeHe+XT7ac+thDPUFtlcaAoYXRcZeSC6woEk9DPDcyRElz3EqiXj5A
WdiFW68d+H15kTQim68dzjA1EX4GL4A7XXMCy5Ii1Q8a+fm9NZ0O1TUzJja51ZEYCgBjRZyLiU6v
28lHjM2Znx0Iql0G8c7T3p6sXv24UmNrQyQQtsyeM6WpSEYfYxbpu5chgy6HYCpbukllAbYkUxLg
WB4IAEXjcVmNRQ4mS2mDkvHbRKvjv98wpTyMiwBa6dnV5cjsS0pqnVFuh6eo6Xq50yvJAUtijTdt
10I57KfXC1zyDJDtGqJUhj8dVWZS+P/WPKAR8OEOSfS9k0o6fRn0u4KBPPvPHkYIOjf6dAGwsfjB
vaF9H6u/30R7bvuhjtbCOz8IVdp5nZIi0EY9Ht+i1FFgjlYiENhTw0yiwO8pCpblplc2cWnBxsij
l7cZNFZwX/EueRePg+I4Z5oRnv5cCKG2WLYp8X9eWdu22cd4CGDDXme/lUDBbVCHw1truSQGPGzn
mGyFTY3dzXrEFyRfZrnt6YcuBa7HvQAq3gfM6gRlP8UZUpDt3OSlkEQ0Aek6YY71zy35N8Id1if9
720G5toVMk8r9FHixA5CmmjsC7vLChnSrzrjrzSGnctk7ubRgeuewTYo26NC4F2M8hLV+5TqpXp/
0qu1NA46ULujO5tzNWxLjALjt7H03u8LvV3mQyIAkmMdz78tG6JjnCJ7FW8DSO8n4TZRU4eaPqRx
WIyOquO012TMhD3i9EfxkpyzR9BeLAKPFTlcbioP4ECNba2PvV3PA3lts6kGnbWqsr4OETfuqmHO
YDifFq1BUUXpVOtJFIUYd/P4ooqLoOPfzsIoFi065WO7W6TiT2TUFYWI7yeXaaWsjcGQt3Ns8U1t
8OBic+EbREbkTyLUZFN5ojxszC3QrxqmdHKAjo14ifUvrgAOuRhEswcQzFjLiFyJaM78mkwCs4ea
cM6j9h517cDjwtQ437TBJdBkBmmqBluc3hk4J0EWX3hM2SRb88y1J7CdWMqHYEqP75UPy8dghQJb
vR7Y5NJ4ChPTMLBHlORJ/2sMeTNWo59upJ+83NoalmybbtFs+Ts8X3hVs6MKFP5DbYRW1FCdGk3Z
2MQXrBYrmyCWxRQ18xGFFcISM5M2oMuZMaPSEolvvBHCJm1CLb6w8I3wnVMBYNPIyaZ322qMD7Dw
JDRlzUT+2YHwsjJoGGkWD+LriPWqe8+F7xGAHEfT85yX6sDghn9HTa/pXzRFqOCr4TmV1DGJ7ndq
kCRWaOKFJd5j1EvBC06h+aYRK9vonbKE1noaWqK8gF2MA1Fr5a4boH6QkmbtGQ0lEYFJSrPZU5Cg
HM7WxiA5ILznL7JiVNWOVjg9u7kcWRuYMnADBRqzJeInFDZHKV4m2ee5rN+33eQCOxH32TPYaAJw
cuCyE/ouB+i2oh5DFiWH0g+4WvSlbnUErI2KJXCBq8+O3o8zrqkC/OlofDFgdmrDLN8teeghY0Y6
bRGdG0SMyOgZVnMMc+sCbvxFtv8JMLtM29W9SpBUx1MidJz7ajRrkoF5OWB41dR0hrwc0fLrIuIw
bChm8vH1eHuIITQxpnOoZbD92Ez0mX+yD7M+TVQeYoHw4qy4/ZpAXxN/3uAlewGUJg1mNaF3MUqc
Yb5OGQEsdVCe9LdA2OKdcXo+056oRT15dcWWxZcasZuxHXNkB+fFJe0Mcs38QvJrDm3fnIzFPrXc
uGIoXGmxJqd9htYof5XwcViybo81DPttMsOZ8MiF5m2ecqd0NLwDGf6g8x9jyCwFsvD/3ruC0elg
Ia2de19lJ1xnGGsLE7YjixkzoDQmTOj7CJqvx8ojAoxP0yPF6Ru9itczFGtfjjzSJbb4ddO42CB1
BSLvCXQepuvEDs5Vj/H1Cr2rwBFqrajfIbU47GWdYUdoMVIAuRjUV0SyNKiBWl/roEKeowGRZ+/o
lA3so5PCfGJQntHhKwb09RiYXXCmAWGco254srMGOXZPBTgFOg6QMoEYsDtwB9Wu3CtvvKCfqHs3
oXYDmNvPfKQkLoGtDcBh5Y2YlZA+uJTE1HbJ5EHSYzBZaG6cB5+Fyc7lo3g+N7fUlKuMs6a2afek
YyHfK3pnr2B7NcuTFYdIgPa8hCHRPQd8P/+yq3RoYM1+bhPMCSPXunp7i/KyQfGyrb4kMsu2PMoM
iUAN7Ax0vM5yG/dB6by5fm0IzlzZ1eWCdT24gK59LdxIohp8UVSWvwLFoFQRJAc6aNYacgAvulWo
ql36HXNvxG9YIK5tFoxq1mlM3S885GYF2h7vvfFSqdXkYNP2iKZ74koLHdkBj+X2vLaxCHdHCGP6
Hw2wJQWzQkMmpeiOlcfsXZMDwu9oNNLiyBMeNkXFQEhsX83MB6pF0xCcEEmBvQsEV2lJQ/+bNqEF
AVI2UM+9B8BYFygKVIqZApDk1QgMrrm1QDQ74bUzPSZdg3WFK2PuDZPOrmH0UiFNQ0MU/0N9UXNe
XEqW4QxqOGemWmVB7ARFgNdQHt8NCFaykvbCHIBj8UZfOt2rMocuHva2eCuhr8HFjv4EiZNhNO21
wjcbl8zHBA0+NUOSH29UaG+dfpijqgFdcQ7SKgarBV73EqKJa/pVRzS3Z44BWfaG9YrCBMGG5nzC
lNXFqVHfG8WjxBUlyaxm3j3T4pu+Ph8NItb+Pfdvsy8cQBnUbnczDTlauBPVuV9Qs5tr6UHb/pm2
Zbnfctg2jutZqA63M5n6PJtfPas6wqCQn391jqmin0HUPGRQJgezm4zbVoNkhFX69/amncrU2nWB
L3T7/ag5EaNTPBkdj9wapaOzi4+OZLoL2XCxIfq3Ig20MrhT/O6NJEoUT3uUE7tdIeW5bYi3jgUg
ZGgUsneOE2FeHJEq3DUkGXJVNdqpqpmIIIFTjUQEKGDGLN4BfSlsbYuhmteacVEYuIIOpQZ+OzEJ
fW2eRhhrGiN8MP48OtJnLjTYn8USHubV254lDWWBpOqwGfZEYyagFkKwEB8qPixHG3LdALfVyNHN
Raknn/COHTVs4nhnPSrCyf75LhBTExgeqhVUAzludZtGNSaBDMN/zrBnkuuWgkQ4+FjCQY1kKfk4
HnDJslPT95QnFBBMGn4gePB8MvH2xNTeTeJT61C+vWhff6gQitCcIu+qwpd1qMD8h8eQXZT5f4Ww
uHdxyaMbVSL9Dpg40kOTiFSkE2BvjAdeBgI6lM6fAF0ZSpv1rOA+vlzAsAZw2K+ZxnTfgssM2lq8
bVb7MGSqBsoIwoIqqv3E0OvwvwcQ1DpRrq2EKOCyvnMY9qLl+T8xWvr3snIM6Y2Qyw4uloyfCAkk
i1PIeuEQr6Gi7VPGtH9eNjSs0cUbRnFIKcYHkuxxwVACWDQSRT6NbnPXSgqZBFCm39Q0+eN9CFrp
pP59hyuw2M54/N3QgKzlHdo4YH/Q0x/+056SRduG3SKk33077WilDwPdUkom1aXUSOmEfGz1nMkF
abfR/6qRiUJfXKCrXzbeZBTOf5XBWrb+kDlZIFlc9RzfsTMvNAaSQhmGUbEniW3IPI57hYyN60Za
DpTDZSXsravA0ciCZsu0uHywNH1CYxUwZlVXZ0rCPng+7IAhYTaH01+Q4AjfIBB0zAHb2AI37f4K
rmrSjuxBfm61byp6DdeQ7orMwbCy+ERkmSJnZbSdkQDr3OOjnPeeW7n0K3uHhcfnc20QRQ6uyp/o
Njz0MQHi1grixA9D3fzGR1QB150vhNSDMEHWOf03JGI7Hwp77MTv8/er7mXv3Dhku2jE1r7/6Kp6
J3GOaPV1dujTkTG8GdPEiUf0QdcFWAYtxlrNNm1rwBFY+CZ5cD0+ZuLcEB2rsEl9DDQNxK3KbjYN
LxkquXZrNxcUadQnz8hf1Ei9JfRNU4XPPb1EpiM8WHOghkFM6vdsyMIw6N9+0p916R56FGOCEyYE
Njzxfj9HaqyYfpyyls5yQyxX4MsKMULDE3+LbH4J4neSzzFveHjavIUqZU9oy3TCAUddWqcthpyd
1PK3OOoW+Dr0U3Ki1hOQHgNZeRNLtM9kCoTpWT7jdRzDN4j2M6r1DfP9pbMCt6BmZ+v13VIBE5NC
/qJOLYfqLdiJY74KsdYU2ASPNn0Hb8XqsyuVs8vdMQCMplz/I6inVIZ3xDNk5vAWp3GV+gR3hA4A
r6uHygvuCKEtSn7rum4ll2wB62PNyc0tFrNvkOuiBgp6um5MLEkUGi5OqpiplWioMjCglbCi6RoG
sccI9FV88Ft962ZQgGfPxscYuWGD1WrUQAjYHRKv3vDZLFJ8fEfiXGLV0c7u4KZ5akgRnGIe5JJT
WJ1URet1mL5f9hkescVVAP8QVRqWZVcB5bO1l1/uUjey0QJgiDS/ITZeBHILrgLj1Dj+uQb/xVtG
uaV2pINmqLN/lJALRhXEJsW6L2RMUEsKB6GXVu20mNUQGSEfWuOvImR3ABiZrMWbZsUhUJIxmwqA
p+/qVCp7Xu0aBrsHlg3uqomlAr9Bw291ar4TAwF1Iu90ZfEv+zuWqH/a+4Sy3pRVIIWcpiBaBlkg
IIDOJ2E6NyyhJZjXeByRiXWZKxJ8g31ihCwPOWWRWK1FIo/oPbrh+8vWhrE+OhnaPhaepAz7fhz+
7jVpO16drn9Sy1bAxjb0fLQ6MB/CyKwq/rRxA5UPt9X8Ex5QzHnQakva9eg4VH0V/Ji6eQTsbpAu
4KYsYIRhL7GdwoYt61tee25aJGz3UrS0t0X5lBCdB2UIOPPwHW5o0GLEXmV7UaQKEsHMOoH4uElH
KzICLC7IIGm9hYMYPMaM3CQTNq/79cxx3UlivPv9gz7Id3mfKeXkX8T0A4h8W5HFOpDQkK+a+NKo
CfBl3yQUwEPO1InewmMtQFmtWC2WiWaypUwc3VVGTiXoU0cZCzyf+J57MibwcOkH4wi8cAGvZYMG
P+xz3cprf3o3M4JJVAIICXo4rU7ikkkcneAupZ5N/BfrFiFWh6epIN/i8FgOvFQ+RkBOXLRntI6m
9zztQ/xdi1YHAP0sCBC94kZPTb+0I6g4VIgjD1q0DN5GQBK8hXahJPKzyHl4pRVfDGVIVJLyhYqV
KePhHfmq//KIYA3SS/zsHECZRJAvu9jvi7rmGrtEOANUXSnQ0LVHrm5oys6h7ttWJcKai9a3sJAP
B4aIvRkzpQsRDTMKJ00TDJaemV/OyzNxg5rs2sS3X4bWZFNW5FFgiyEMYGOJE3komsFxVDV7YO0r
98LxyUr7Ht/NPpaItx+Txl9H8GpHEwYh9VxKpuifSGYeJGr7EkAVeMbHRQBd1gkfH0QOp6Y9YNfW
qt8iqtc1dUlv9wcm/vhJJKxaLabDZerj8lIiYtdy2NgiF4waaEd/apBMHE2ItQU/85L4aJtgX3S3
m9nsNQgi2LSONbPU1EvPLz6DJgtf27+0C7f4EfW7pcGDJp2zNsVSkP+UpYrY7Na49qJ+pSt5FW8c
hLX9jNQTbdLfyMTzFpkqq28non9XVcFjqP3onBQ+qqDwOdGRf0PIgiYszmw8wd1UFhw2hCirXB2z
+TSVSTzbLbl0/aqas5SRAnwrmNmvWelyK+mbuRcKKcTFsQZVgka+9AhSNLVx/fKRBTSoDC46KdSQ
CGGDxLEhl7H92MkcNBnkjt344sTpN2PrZflBbXFTX/pfpkgOJzXDsRrG7f8ViRbHNvTy/xgpUs5n
FB73P1rLYd2K0gi0vu1IlOEqBjnqCkPvPLA6pFRtmqkIucEGWm1DBiDuhSDA8zsYuYIbM0DZ39IU
Waqfs8mQI5WP0H8hyzH3YuiPmprYYBrOK2Hwxpipt1ClvJcyIZeLUwoU7udjwIgrRLst91SNHywV
VjnHQsPIVS2PUprZyWFoNOx80PyTcNvHvU9GysnMgnpA9hb67HIat6dNmeNnb0w5jtr0rnxutoBN
h6UbaAg6qnuho9kmvJ3kKXUqdOI24a4VAyUipgvCvQDusEQLifdODqoXInOcFVnF8sLOlKpxl4Ss
QSEsmo4xzIFShXgbKkfxk0eWG/mv4aUFW/ivEqklGu/dthd0m/wZjbSS+vFnq5sQ+jsmXRvKl0SC
LzPUPuNxGwFDKu2nHXKflr1x5ohxQBLP0uUPvItEfxQaaz4DLjxdYxN250CoozhrNm8YJs2K6Nt/
3r6L/qFEABgsNQu4xUBgFUEWrm+NG6MrAKlVCaBweXqTTwCY/eA4Lg2pkb9XX7tGu3t4YEZWbnfl
HXD9oG5vLj551GZRdsixesHkcRrcRqrL7d1sVaSeKfqxCAFR3xErvZtEkAkYxekelfY1j6bh5O07
WaJiDkz68SKjwl7RrT37is3jh3kyCaHj3T0fWmLvIXAN6DnnqHGtL92w+KxdhlizP4LF28vR/45q
IjsRoeTCzmn9tdfgsg5+LiFKpYKBZ2N2asAWMuNiKvza42MgnW9kxYxYoJA/R866olEc2Vdgss04
QZdIOVXxx6wXYH2oZNpvHx+/Rv/9mQbdTaJLbP+6/wyVRzIIsKs/KAEs9/VJmvt3e9ILEtdjaHt1
8MOkSRhp5kSMX4UuGWd6Dusrop3GpeyzWT0bolyw80viUEuGyi2INNetvxBudbux2qGjgjz/ZmdP
kkm6BOQMN/tvPtqSs7cMeftNoWaecFaO6Y0+R4iedZLHdtAdkUkGuWJiHSajiAsbajQj08o8H6lU
IjrtGoAiO2IYKGv568zoVy7fzhG4ONU0dGb5q+Vfs7aTA52yxkp3GaWe3naciLjB5WEOv4AZLTsj
nfcvk17Tv+3ffVisLOda2rzeapBksR3gwTUFDx+2xxMh8t9tkmyP68+VEQ76eQSmH3biOrsqjuas
iX6FjUd41jYYajFLU3o0LlfiVHR+LJpYTWpxZpYGdPqaWOWJJF0kzhAKRwpaxd1KH4z019UjIT4T
wM+F1NVwLitNlmlVAw+vuwQ9O+ZiUtJXMQyACex0FQsZq58RrdjZwdsH78iA17JAVvP1gmULgL6g
2DEkbGZQrzWMm8NhtMzIfKGsWyt5O+Z2viPXQxpjlPZZcBUq6qjJ38sBc1IBsEYPtiIRFhnUbe5y
RZeKvkQ7gCFJV0/1h7zBBUW9brHFNd5eXI1Fo4flalYYXzhoE0nMZFEHzHDAGjbActm3eU2DlJkG
tzBGPmrdTZ+xe748y/Ea/jfriYCFAYM/xkzAoTPqBmL2uKJU+Ip8/hGbLHbYwZlezRlTOBvTUJD2
A9/ciSrFbWuSfELgNFfWVSxfoww+DEyEF82YohWf6Y0M0W9i8HvICWjpjWCr7hgshyJhlYDCVQ/W
I5kBS0fooWyD1M7/T9kbpPUy79iyGATDYWDpf41kgdzuEKj5jp8XVQAfydkGtpS5MjRAG1ovk7tf
0JhcoD1ghvmpl92tIIfiyyp1aje82/bSnwAW2CTwdAmkADwQLAEkeoH91VDjzPoeZFwWJy35ib52
ExtbC+AqeUUG3IdAKn0L9C3lGH94rOg4Mebe6ooPU1ThfHLXZXSPBEc38VVA+wUk946nHZiD1meW
lN4auy3aTneOIXRd3GnlnqFxCul/6IYro9QbRLDTVXQu6dWmE3BYRUDSNsBf8KWFSCUfnZlE6YyB
I4uY9EHSa2n8JRzvs+ONzG8jZM0JEeSm+P6xZVp9Mou37rdETXoIh7jiAmb7hxBQIGCEuSQJZ4eE
3WlzUlst7cqBd5+N8/Q8mza8CSWd8R5hrCfAF9hkrv1RAE9bwmmCGcDRDq/PI7X9PiTQts3taPMY
N66aNRFv5ZCtDj7zywvxctHKahOda+KitIvzi7guHN0U7H9ZhbBLBQX0yTxMBBnoWiPa38hfWkZe
teNoUbdsDfdzaI0KnQN+A8qFc6r5wd/96YL9bPkAto3WHjCmOc/ahYx4ZpL/loSW6PvK1KaZnQtr
39OXFsIloleSzsKEcOfqwh+s2UEgoeZerY5JsYpuI+ybBLHs0VAhYFmWH/aGXhs5JQFPwFZKGkSx
il+F5yNHNhMO4jLHEs1VP9EvUZIXsdZrlgwti+4ntdSB7SEjq7s7lUg3bG4l3WVrpbAy/qLMr6fh
fpDJ0AT6kLTIhel7AKc/QHJsTSJrPLUsv3khqV8qg0/X7fxMSGBTcScJwsQ+D73FW7mhPpxQYR7a
IOc7UJxZYs8ZyNTCKm4Xq2otWYbVTV6nx7IcR8/2HWKHXOv4o/0CGaXTp+IFdmY9HR7V/7As2AjH
4JKuMR4BxUU220CcBZ++IDob9WCqXX6e3o8qyaz2tEu3fzTbfzFOOmfVWXmGRw++U8qWN77VcMXC
gFuuJDJ8PIfpdvh0RG/bUkwNow5jzivfU1k+9opiitBSpGfiqgUWR14gzIGTF96bKLctKZ6zz9WT
E5wFDLEXDmdAUG+AxrlehfOD7151+BGnfX/jw4RTjsm6/Dpx3sb6aq8jAmYQVBNiBtGTCzOpdLTa
DpawqMswRWTZV8rqcQf2ZreQW8GfDZp3rX5P3LD6ix/VucYRGGho19evmmI8PbHNiSuPFunD1c6Y
2P5pdfUuajHSWZwM3oKnW1KnYSojM1TJgKinYYzeWC9LroCiCcOJ+Yi78rjYQkKmN+xn/zPuklD5
q+HTKlw58XF/Mn88DknO7q7jPIKyKCxL+O7sGahJbxof1PwRjyp763ZUuGPNwzOLRO5MN608h9Di
xRJ/m6nwuFLZo3GZVvkRCo7PhwDDqOuhRLLo/GIoBDaV6gPLkKY7dfUPKZOg64IUZu4xzSr28Z0f
GMZJ9JefjSERbCGcd6E7LQr8CQpaeYNhE+jtmfBm80cZ7c06mGnRlOQXDJZ/88xlBW+c7ziTJ6yM
6s6LYcExX+56hEVkg7mFgtfvImEAwvWxNV0sOK39WNeKEz1flI9yD6VaR5YIAKpAyL8BC/15EW0K
ohBMZ13wocAUevL3Up2CpoI0ZE5tcUu/GuAjohbHF6ofb265MtTFlV1TU8wfaaG5S433FNJ5BrxH
tj4IsrHzhwwPSLJIDRf+vjjioXJeC6dZnUP0ihRtFJeq9HzIP870jN3/Xl5Qa5G1ucZaW9IwTlmn
OrILYflKP8zwKJjFiJl4BhdPsJl4B1jP62v4M21Qd7ot1qbeFuOQheExR2MpHW60dX5hlhdHvv5l
ZVbxkjgF5cPrFetePEpK6R9nvUXd8msVgbNtUU73t0uRkkGKZVVvnPX5FjkUJocnc+82TwLbVchL
FqZXG4dKoBG4pQ6jXYo1M2nEdYKzaQ51q8vktWspui3Eyu2mzeZcnT1xyjCAqBHf19b9wZWNqS2e
tViCkDn3pRUQgkONnXbiQz9Cu1ZIw1HCO4wdBk3R+0kt6UHfHKItr1C1F19kW8r7pZncWiNr/v/4
yuPD+wh1z6d20IYxuitXA3wkptxePHZkf8zdjZMZ/LBMb8vrRBe05Ad5ZubuMYakRADbruhjsLdY
SBdJRBfEgjJAt8yruzjQB6mczWvLxthUy6ARDCaPz7gtRmWRPN01MS2zYN5zWj4qoQTwxeaZe5Bi
mqfcYt2QHfgTj3ijcOe1MBn7wRE3460dZKSm5+ZGQJZT+B+LSL9HWUlVxNl2Quzy75B8JJ7W+1kE
b4vuBK5yx0BnLjlni/6hs2Brj6siyWwfUVnTfp71YIHtMmN39VdQyIeiF/rKc/8u5VyCKR01ArhJ
Q1EhYNDMoiAvyaloWxnEn/QJN1vuRtHh+2jOPzGU5NwEVAXrjaYlsTibNJwEKjRTXUwNi1LY/j0U
JaurF4ICOiHF8caTyvz1KD1zRk+VVE7x0Mnl9ek99RlNfASO5AUebUa/nzjHj3EBIh+zanlm+nXf
ckAdWuw1nV/WMpUqu5iNTA080YC9gu7DbpK1OUG4PNm2Bg2tegN3bh7K8q46juhAs9G+JN8yuvEw
v0Gj5pO+MVUz0NZXDATBP0OyclJeDt/PXhzYvFseE8vdVwWhHsnFYZ+b6kqUc2T85LKqm89+thLs
tBjLK2sPmmvAzg1ukar4Qk8AxInMNqyyTTkYeyYmnkHQIg/10eTeIkq4t0EuPrQjT/6V2yN3PrXO
QbLy8nORFCA79WPTNV+llwP4rlLGu5GqEW1z3IeQhKxMRQZsgpzuWDZwcAncSk1aI7zXcp94SNlU
x0bW3+tLTUQAPH6boHCRsHFbY4vozOlZcQsXztbKmy4T4uR8iySjQHeZTPpnMFUZWVZ4qZkXesFu
AlJMV9GETnWYM++frHsHYVFW8MilNT67dffvn6lBZG6Ao7D733EYNfq7X4gS8k9SlTaGZK1LM7g/
z5AuykeA5hHVfTQYGN9WVhi2SdPcG/AioPgZ96pEnNd4zJOUF0Z8HtQ7QL15FEwKU5ecmiOtaFTl
Y/IJ0xp336+Aol3DSw4NI1GpKda9LbWvBhpnPgrO498f6FcAS5Al9WOBCQviDsL20wh5mae2Fdhm
UCIoFqWEIvDP4A07B0x6McKftm1kadzWH0ShsQrf299Sel07obrqhawAAQfjowp6YgB2JuYH5bAX
tYHx+ez/7w77DgqJSLftPc+UkTPehIFMot68eMmWDZqHC+YuvMTM0ANTsfKh6vSEcUvyJmh1spt/
rZvIe8rDBN+nyjd912xAQyUgP53quZDOI9VH3F4yBQwSQA1SP4WIhieX58aRDTZ9QqLh2lZXx9BT
O/w2tXth159Ic3R1LXccowRUEqDzUcO4WpsE9SMMXrq5+zg4Y/ZdbebgOMmesv85hvwn2dMzBnGv
KG+n8z0PdvgoD6J4/7RSvKoWuMLMBFSlkeX6REttSgSUXGGcbjUfQRlxUsEYpH9dZutp6s6qJBYr
ld3+1pILRM1VEpcdFNAlSVlDbbEURb77g0QNRQyblodTnepZzKLW2RSQHrfUqO4mK76/Tqn7CKIV
1yBfpLCJAme8SbmHeiOUGbUB5drMM8E1o6e+r83ekxtGPGsEo4VomP13XNzQUw2qKEfd/egF263H
dQ5fa8/tuxUqcKJOy82BssLZGJNmdW1Q/WMhdcvivcnWhtYCenb7Q/BmLDlLiMR+nbFvrkSsdsW6
PXZySVImeo1FvxBDc5b+joqK/rXcpZ4xClzlLBce4laGPiLwAYDxAeOy/YSaSsD7q505/DYiDb6n
5R+iSuYga0hs5ClGuKeZBnlF0CvLkHFv1lKrMWwbpv3q6wxCvbSqNQ/kVdm+2CR9t2khdBK0mXUQ
pJzge3PhiVmEqTSp60ZySyCRQVBTpCI/3hIrqrgYB8WzLVmBLUFRpiDyUc1sjQta50fVxsaVlxPg
YwwuNcf4NQdyznoqOuLR2FqZzWsSr5ca0fjqECyyTSE2mSRcyA0ClVou5c8JByGniLnbwkGssk2O
2miOSZpIv18FI5HakrozWdOdBJYG8Q3VUPry7aoIKBxReC93l059QQrlDGTI/4PSK4hz2smKm7j0
EZIkUH7ABANlFdbSY/pALF/SywmGtWP6jjyMX1AWjANH+3OZ0R7u4tBwE6C8D/dyMKEK0h7sZ/+b
vqVA2gjzkbOkz0N0U3T/uG8y4kHEIoQV2y9duP6F7dJwNy1opI8fANcSrW/iepl/PZZyZ5DuVdKC
uJ4d+p7Gwm8GxiZNaANWfFEHnt04G2TzrPkoN4zsDtT46+GVzoupZxElrwmTo0M7/j1xJ8DhFMyB
znp3RtalHDDriPyi4ctLKOxrgRt9b4DZUgCEDXJiBuKP1Henag6H7UoCpppf0jhoXW+im5Qu5d7b
Cw5EPG3VNFsiJDzXlJe39jNEUHl5+9LJOWsa7RTkvJj+6LRmS6JeEl0rJ8ohKozyuB4lCQVKPpBA
lTv+bsdV7yqgiQ2IXWT0bockhay7dwBdCS8IbSuICwH9nNrfKUXCsC6LTPEM7VRaUUwzqwCcBe8b
qP45I01dCBZwVoQmr3QfEuprq45ph7c1y62By8hcYCeu0daXairaQ9iE+l3A0OYlSbAha6utZCZC
mPZjCFzk3/Pn1aXk0ABUzfGy1z/4iFRRqv+4JChvr9V1iIfmxYCO9UvmfagbtRBx+q4eqUIU2FGc
p2J1tA188f6S24sIjQhsB1/SKrZ0a9vlBhFbuH4jVi83O7/EHH1qZbfAYNmaiOvjmieLL+sLPs0J
OCKD/hcHMD7s3O9vD89EnQqEqCL7O35VL7E4yKZb5zZtSb5oQSXqlaFCjUVL5PMncInBADYAO1tU
9/irFBE8lQBNv32N8WIV/lh4D599BFa70pH9YFp19U4PHPZfa1Iva3OA2DlAgARbRAQdfZ/5AwWK
kgAnKY8iA6ECoKLhT0HFUwM5aG6vI9RsL9oJK9Yams3h4GtU7AONodrfdJ3/QPR0ygxEr3M+/UfJ
8QDUbudIeEiL6ucG4B4jFv9owPhDvc47++TZ2LrR7sQsd3eEI9PzaVIx8+2Bl+ozWqMrqy4lHPt7
9XXeIJGqrFgiXMKLW3kA/Vz5LFjBaUI5GVVnIVAfxrPSzVGbGeR8y2tYym6Fbx+F6PqgOJ1ZWPxP
JpHcbKZwW6dKu0WIwXeJH8Y0JbWdYNDmNBKk6tIYzCFKzde6YW8hDtY4+Wz0tJ0EKAmUZOe1vZrN
MkE5YTFB8OC5kSK5hoD4SohgIgW6qYYN++Y0q7uVHSQDwblXWDzuqDxKxvYGcf3rRCU2eY3Rmh3U
SNEhGW0gCfwoo3GI5fnLnSNUNU0AHAk19iP3bm/+u3lOYmPBX/vSLrWWqCyeC/NI5g4u8YP4of/A
aHlzo7eCJo8M4CJcSB4OnA0JcyLsWpjdXmHcwLJ0rS+Btpd22lBx2K4CD34OwnhDXNK9SMOzjbTk
H2vD3qpfsEqqqvQMkk5A8BpJxhti1OSi0ufk6uoIgGotwSqWJ9gpQ3PvZJIpcnrVNMPnvI422BES
VSglertm2PHG8XqDTIlcMo6TnJf4KGH/uSwSl+nUom8equOq6GuqOnxDuC3BJNJj0VtQTvz5LdME
HTRRAAkvmLJobz+rXKfRepuVtCMwbYkhr+CdP7UzR+Jy3TUcszK5isN1agigWxcNiw4E6O38/aRL
9VlDjWJnaQaCzDEQns0dgDy1xeLUuN61jobI4fhH+hS+whChiev/qItDPnDfChQVCxGp80BMcBpQ
5OvvAsYK6gawKl6Pv3aF1W90jZ1IIOX9x/U1wMII7p7lpQweoTJHgFZkrS+03doyG5KmCZFC1ZMv
DP5fPsqAjNYvFaqDDLK/c4kkNB2oGet07YBhgG02cKHxkN79MiRRNKKOiCXwIZrMzk7oLYywDECh
/tXiVZdxTjnpwSu27qojBdGPuXK+gnBbOsKCXqgCKHPQfjEjeMbRRpt/7EdTNOOrFuN0kaBCJ3ED
afnk3a8jxKkxZ2wsvv+5OVzlMxgWG//PkSdFnPrA8gXTqddXNHHEAl6/CcjbFxTraNotClbBP4Vu
IItv+CcK7OlvpKEnQsTLZmWunKDXifp2/8EwTgM03nTYukiJNp/JnBqvRdyXbgnyCvmYIIZiDmA8
oQ/vOb48wKDgFELkNakb2Tm2UfOeXgrTrNGzLx71u5Vqon2BiVT4e70HqJvDtX5pqbBcIxRbUkqo
haqCJKyQpvgOKcxKAhOb/0FHMu32JZWEIecgRWWW7PmKCvayB78rQJQhm/NZ6afFNnlry6B6tNry
bMpetjOJ1+s4+OWhOFJpgTRcaa/ef3qDNiRjcVXuR5jp3pjGsR0/C066o/PAO3bsqRaBlVOi1PWZ
EdU3kYdTzNQpHy1HiW95bjj+fUINL3w2nJiMv7v4jCh891YdzxtE1mSkcexDlpKmrpbF9rGb9nVG
dtPQRdEh1w2MZaoP/x6KhXRpvXzrUZVKv2rYkOiksiuic2WLJ51KC4A1crKF479ZAqZdIgjVaBh3
ZzgRKTs6VhkKmoQoNFyqWekWssOgV7VYbNHfS/x1q6qalzmH1gxjKfazkZWE9CMqMyA7XpYLfRtP
waeIefUP7qRe3+O/I/Pf3PC2KHRlDxDt0Gc6hkTuO7216o1LLKqZlfaOIYOBfkbaUNMABS3d8cxD
tAePkEpjSGQFdiOIdqseT3mQ94+5pKk5RQ+XdPnXq7VVsbw0ikeadw9i5+9JBwrls3Ev6xn66ixB
bcSqRJLm0R0zsP7DAnyhj6rS5e8ewvnV4FwF4ddSWHxRGlGcVoYYIpFj8n4Ycanub5bP+RROaI0S
i1/Q09p4pTjkhkJVrtVclF0rBoZEgkkeFKJoHDI9OgoohGoidzOuTaBNsD4Uw28W95RjJNtH5OY8
EwgMtOyJT7+ddiQfz/3lr/ziVLGthwf4SHRJdWMpz6ev6ZHAdIjJAXcXCcaysnKGPVqMHdyZq3ul
j2tRonyEfnfxZ9cIr4R7+B5HpIcW2oQ1FGSgPFqwPzITtvLQ2LoaXms8/XRrH2JHEE3r5HWgrRmW
5N0N2XLXhgu6P5Nmyxx/6lk/UVNqk3o2czzJPWN559ochBcyQuODHSFwIFSjDw56SvYDyP5KWYAT
0TkAxUL1+9ONpYh9Z+/hGB+UsR+pIY0w4T3eami+K3T0sbXxWhRfbpPSKNVX+dC9DHKrM8LIxvvP
+Du2yT2YUHFL6LLy7DdjEZXuZNAmEmf9CmIAC/ByDBHhWheIlcJXSwynkjGIqIxUo5fXVQ4e2MpL
T5saIRW7ovdDYu5lpTRcV7t1HaKr/Rn9S7pov9LKJAxvOxi/O/ffCv2zB+/3hk92biBkLDJzStqq
KkvsIJcDteBZQFGMnXuN3+Ba93hnCtqN6Hpijuo3K91NN8/qtLOXQLYm8PwMAQWKjOvhdcY1bwHe
kA5lDSRTuw8HyZ31URk/2P+VUFNyF8hM4p3IeLKManQvkzbHQgXWxom2dYOecNktwTkzJoe3Y4WO
E/FOGNwbkfHDrNKZTmdHqw1h0SfgDdJMI29Hr2eosgzAZ8uE9yI5StRFATxxKIWeLhRPJpR24kRR
g4ayJSRd7RkT6AUnCyPzSg0R9f4QYyy9C8Lh2TXTIw+X9wvuoJw6io0J+B+5LjvXrbUZ417/1utK
QrC7Zu1pkObcRh2kyiPUuQwzwaB7OYoY9N/wuIZutM15J5XYy9KQUw2bM1ywDKmbPmbn5rgoMqru
89JSk/v56J3Y1sHegkXDT/ThOhghZ8Q1uIDjQA1xBfEzbeTQxR6fcm9Lo/gKsHTtoKrwdH0Ku0xp
4ZIyR1SrMJ+sOA4zZeA0CgreeD2CnYi0vQsIWuGGNSH2lWEu/zd/q9ZpF/gjLym1vtZswywC4hZ/
GguqmFfZJzAt/IwoL1ewxWHcogshjVqDVgtnXgWxZYSCL2gkBjDcCYZBOWRFXaWtLwOTxV0crLHc
X/XiX7XT2d4Ab2Z2IRaXquEQi7ZxHtgD14mKDL+qSRY4wNBB7OB3bqqCVe+OK2dSJs3+0ChWT1c7
WRKgNqlBSUhFj8kire6CTwQ/6NGY3KlI10VtKhKrGuKlUgppProQTsu8uMvuprENym+gcPEOtRkU
ApLaouMH/GsCNq+ctqzEYMIqJLGwzjsJSJjS2S4AWDDSwBxf81kq7u2dly0gAgDycY8zfOIlra+k
woR5x27JxjoQjnRTIMDbg/2OmOrU9O2kZJlz01tpExTV3kATflEBbD0lUyDjOM2kdpTmgUwCUviH
XlTa7w7z8N1KZhMXtSXhQGEoe2glGt/yXJY1OlNR7HRGBDGSBmWsWPJERyHoSfzkTPmtaB0ULe43
004FKnqyFOQXb/c65V9I1we5uqJen8MY+ABX8eUlTORI131OfOkbkV4gK/003LlEKL5gb24/DcWb
n6YLZHHwjP+fnqr3I6zyhMkLI9196U6sdcKnvdPeyq1OA4/VhCF3IG/m+Z3Jq/tEsINQH+BD1aPd
WzbTg+75bbmL3uGwq/t7+hwLnmIOFxCs+O7iBEeGnUsiTUauqP4FZTEbUZ8tS7OxdjxkR/b7BtQ9
Xiu8MXrhqACv1YG7mVr8qqXZ1rJXF1nzme/X2dSsCWJbE+yKEIR80gqWiRBR3QacjfKIYZpGQy+1
yQYGm2gEsgc7vWrkd5DN07POOeJjc1zn52WHVBgi8wO/41VGwMC9VWDC7gdTzOWDj1TvU168aVPD
qgk5O8k+XZkXsJSrJyZJpF1cqnEnWxRqLS+kUjtc37nvhCvCR9rOycZKnxLeJFgG5CGslRqerGKm
UGvrJCP0vGmDxGoaT/OVlwggTlHQU7mhTosOx3ZzvL60zexuksgYgvYZlda4vDTCJVljaQVeDOQp
fPjin/gtbCDfQa9l8rsuvCyFOHXX9IUYoLlzsPy9/gHgFbDApUo/3DmyCdFiDB3Y3CR8sJGhlYFW
IdyGvea8THcFlNMftKm40fP1GmoW1vh3mtdkPXgmn6B3ufwxHcxoAOgAYEQlSXSN+S7BtpCThs/i
rH1t6cbiKU3OFGEbyTQV7RDm3U8UHCFPJ2Xs0Zfp2wXdG42+EW6qFU4kGHu1Lb9K7EUfLVLyXEZ4
EHmGHhDZ7MZOxJDWNg9w+aZzkQ43QgZxO8g6IFh5YQky8iHubFaOG5gN6El4lC54wKe+KjJ8d6eM
zHqhzZhkCo2o5G9ujO7MtIiI2swsB9h924iK11LH+ylc7Q7lv1K/fSaR2RTlg3nlgMJf0bmse6RP
7CG5eF66PB4k70mlyB80EDXw0bP9yt+za5ebVs61cfw1SPt3L0p4iMHcklH8mZL2VqjykAkO+sVL
PCrr0NjC1Wn56fIANoQFQCvtCv5pQakMdC0sAawiGY2Gsk+Kah5SoHLRFu4Z1v00LXvKrDxgwY32
iqoLuQgl/uY2eIhc3KBeGht5xrAwfTOfa+NMzCBILkuucL2Ze3R2u9uimua+VIyyWLAd4DaeT7ez
qE+M84vM+QazooQpxVorYxu40oj/YQEN3GSNCLfgbs2Ji3OVX9SGhf+Ln4DTfzNa278XY6mz0zgE
rJRAlX9dMGJUrDPr2wZPKPRPjqcfnSDtyQRslAey+LeRZ/10ax6D8nk01wTb7nWdELfQVaEh3Dvl
Qf0/JFxq0ZxPl+wEyD1zvABEfJwuD5EpotG997Hufr1yYwGn0yQDGBj+WHdrg7clXfgocpzr5Jmi
PbEonROgvobMRsrcbGOeGXi9nRvjyLnppnRLJmb/OcPj3VmuvxFt88pvXEHcbir5PePRnNgumcxL
pZsgP43vhwpQvZLu+40DwK6bQs3iZcs1IK6Jl99yby41vl200pbjdp7n9EZDrlM4tCH4kgTnf140
/UISwODZB5iHs2gK19RzPUV7T9mb0FxkzdzvSXZmfSoCIwS1eZxLT0EDIM8+gJP5mreWaZ3KKPxg
t+oFE6R13cKu7O57hZKtW/f75rG9rSQp+8UgZrciNPYUZqQXuE+RIBYaLCewxfF667SvBTkBHe1p
l4E3+SBKZHREJXy+TRPY4ZXf5F4wA85PQEJ3mkwKIcv474Zout3axMSCNDtbVyzC0OrwFOcWAaaW
vCGj0EX7shTRj1Z2CKuoPXrmx/0w6oQX9Znn585HKJIOB5UZeYR0tKQ6q3ftVY7N28Nq1jbzQnKU
niTu0UJ81LQ1MV58nhexkRJyPJMxujBBd4nwwrYar4ehGCbNbTTEpAplTLIiAKbq4hQ8qU33d3Iu
UUwGIS9+lpqlA6r++R2V4v0EfDDsBZlV4eNICGePWO2wm/Yqg+hURfvB4bIE9mbA1b24J4aYVD1g
ZMaq4kmwh9SEv8Td1L+eZWvymHQDNvbdn51FrhsJKBqha4Y0CBj1a2kpScZNsFKbOyYnir20pEqq
pzv0WakfRQN2oITOaC2QzR1ENVWINl/Yhftij49u1Fe+ba1eEOifysQsP6F6C/NmQNOepaQ2GKSP
YCLlG5JgKj7L7XHnOEFWqdiUOkKdjqcKGz8wTwD2IWoUoAv2xPv+xuzLzMNcvpehYE+RSS+1PCts
eDm/afJy7JqkWsfQo1b1UvIXDTrV2HF9KMANH3XZ4JTauYPZvN083HhDZI9SyUMSbUAq59tWMcxR
Q02KzYipYY6tM59aqIWVoX1Q35nts9R4inz5kHv3BpoNTIT3O7YQ+eUTvVzZCbnkNCI96y1o2eyo
BviuYu5635nf0uYBgz/ax9Vvq0bisD+LhVrebmd6qycJ428kkanoq5wjVDUcfFkSEm+IsfbgqAjl
ymWMgyrP1+6Svxdl1PIZlJYfpjO5bHgTinbVZs/dTN7hJHVE+subrLBhSxp7bDtfWdZ0k41IrxXP
NeaMdSp8Rstlwd+UOJp3rO0CMFHnPMWYA/2oNzxeLk53AKa9kvS3695ZQqS5ysg5E9qAAdBK7NUL
lHsp2QNGzvRP6S2r04kVt7EicqMdeLNYw76+EXJ/0dJ+WNfCXWO2fv1PE0aq6E/a6Cclt+5G5u+S
tk3akqhGtNS01TGQ2xinwUVNi+onUgIp9V9cI0nGTn66CCFf2WIcbzh08TMI3gFZBhKlE7hwC9kd
qAM+RCEqAfxsdRSp6rEF7QjRVGhCayn8097MQhxlsF9qTw09lyaS13XbVjEpGaPjx+ZSVy3afiTT
tmt66scKI7/GpEliZ2d9piaUJ26LPXT59v1Nv9LM1uXJ0ftPVg0v54Iiir4vx3wWGlryVglt3Ij7
MFIpL/td7wJVN9UpTM+KdDzoGlDyRlFbkxAugUW/m1ZQ5tZmR6YQtNWZssrGEhemGpEPfKdFk7MJ
i807EzbXEAfc5Ymb7Rs5IpgHM6wjLt0cJC4d03jQ6yBxpa236VUMky916bnG+zRbVlNU4leuCS62
Kimnv2K1FJrKhVltxgiiG/C7qOJd8LUtXzLMEYF8iJAKAVhSLRk6Ydkf6Z4+gG06QiJpPfYrtkyR
9gGyQR0QUElWwyDKpBMGsNjHxQ25S/im3aycoHRgliI6JFFkG4P2dYHpNiA+qFO4NAI35TDp713B
cfU5gZNhXdS4BrJBIDmCkELdhhKve3ItrSKqbrvTQTmmNKppykqppxfxiooekA3kW/g/q7yZF5R8
Komp1tpPYqSVO7w/7Iymcf7bg+b9hre3d7xW9e4Pa+bP4cL7DBxuRpeIRLUVrTmtSFK47w26dO9F
EJnDH7Ve0Bw4yiIvTx/IB4S2c3DR2ZxeiBQa2e9rS4ODZNlR9IT5fdSBeJbf5LhExoK8kuKbLtS4
J9TxysHpZlrS5j8Z8nFWtZhu0mi0xy0+mO5NshAWuSzg9kTnG5QKX6+BImbnlJTPesvHYR0wIv3T
3l1THP0TvJq+nUycZT+I6KFzDBh/hozGzvLVzT/BfW46+t/Gv4CYJc4K9S065Y50GEXaOcq4sniN
rLfUBCoIooFwLAPT8IhsmfTjpyBs6uuUZZNZBnG+NTEPGhrFe7dB3/HoPQlcThc8Qu5nLvyJh3Lg
yjM80gvfNliHWK7pbHQohY5fU1lE8yhpHwGKCjEind7Tejf+GHpkDBJbv0XLUmYGWHeQPwyZm+CO
aIR4WtgUtoDRZYKpGX9tzHfI0OsFySPpIUJPKv9le+TBc4xWwTmTu0pTgfwdDQGl9rHx3Ltt1UNj
a4Rx5dnX75ajRCxm3gvUqK7jeeWY1732LWsSP96xCW6b0ApumpoRf5kMuP4UQJ76WqwObp0fPr1h
KV8/cGqF2mfIm45p6tEnDLvqsN1TrqqanLitGf9wC1+PRcY6ynicW/TmnsPh44LZpKto59ma4Anu
9JWoEoIOAVsHG5xNk26Ja5UBizZ1qWGaYBQBgwOtxkC7xk//qmTXCStmxiMwZzrRX+zN1tDVp8Ad
1prVzyxPLM1bHOc6xMvJZW8nQEB2Na8pl9Rz7uW7r2qNN1/BhDWE+8MsdxhR6CTmpULZq0wF/KzX
dIxUMnTClfEY3K6pD7u1+a/vkbnMWfC8+M4ihvYKIi1lOvKPCwHuj0zXESfeJ6cfUH3UyOFOXj0J
yekg/K10JJ+3+gORF2fQjBBVJ9uwzmKGuJEahtMyUYEpi2rH35U42XP2Imzw7V16abDiqiBLWy8C
sK4ePADRb/px9Lv7lUqrmiY82J1OJe/S1JAsLBJJKgDrc8TXQDSn+9NubEqyZ2LYnS1rQkvbn8yu
68MIOzJPmQkZ4WC6FHYTJQkaA1VP3iMXR/6+8pAYs3e40BVT7Zop1krY4VBm8WEPdpqoNq1ucK+q
mTsCnU/K22+WMrtVAd5jxZhTmvHRNEZqEO8psl1qTfSDC27ToCT+OoJVvJdryFZJoRDIg4TwV5Kd
JS+Bw6oQt2fEjkrzydq85nlqziFZ/7vrXC8JPYHZL8QaVExY6bVrilmfvhAXpClLlTL2cPkf1fdc
GJXVHAkVR9O8kDya2/AoG5IGxSYJhczvcXznrXVl9LTSmOT/lTBtJUj3s3NqZXzI1fTyvA0wE7g7
l9Jr+GXnP4OYOCGlzq/iK1rzcAMw21MxLxk6MznV9+ddEroXB/SV+Dv9OCIXlTeR67B8645vIiW+
Ng5VmL0ApSdg4dD3dU0/jgfftGnRnXspZjBdghTx55ls0hNkznuB6ik97bMeI7mjjhBQBF+VIHvh
vFYGh8vaV8jyLHdEiDcnAlSOSjt7R6DtlrVcxl7DCk6xGmUFU88Qt7dRTUVZWHkXeTVouXn5vk06
Hifo3X2s3mDm41LiuaR8yFzaAdK/id7y943Lcdjag4S52ILiJz8ptDndHeSddF8pITwmOwG8qEvk
gWU/4i0eJhCjR26eeyNyWcNy0KynMra6RrgwlI4LsJvfvgMgXEz1tXUwna+TS6h7SYygrmGLaocr
YyRl/whL1uoTDFnA96jAJPWgIYwqXwnTbr/BMXnXOt/l2OdSPOKTyJ3KS0/nGpD2S+yZFTCKGbTG
95zUteHgCtfcov45EJ8wo3UGAOLdOoHSNmVogxE7dQb67xulKo1VwEy6TW756hAfY8MP6VHr0iC1
Vo7burCjqj9SniPOBPhinaS71+tdgw5ThCYu01tafmi/omd095l5QqWVea32Nnv7eNIsCYPDEw5k
xO5Rm+IawEkQuhbQ75tRM0Xsbcf8PTEP17NiJ3rphs21VSfNt7fj6wO4Omg39vbZpnkzPT4V14GM
aC1o1Xqvl8CqgiFwHd9tYTrXAOW+ZWgwaizmnb3TT6vwK0tUFnNedrJhWSKohifoDzmirX8EuS0W
z6v3cHBMQnw4wemlrejUJtBvwSj2qvAhZi/Kr5/6UxbvLaKcWlmQoS/JLYijkSethiYNZ/qZcKdF
3reydqA7KSML4ZuSe5c7uRnykalWgI91W1U/y+uPUeLfr+CHN92/PCimPKrVD+Xfa/Aec6T9126U
qgMlA2ycNNxjaW6bfJMYp47n9M7NPL5b5A0oeDY0vDUyeq/MruHnoMhpgk0Fi22tjtodK+8+92P1
Q/gGRKLeTDEcKpdq81t+1P83lHt0Et/iXNL/VKf4LpH/ugOAGoKChcLfkS2MQH47Fh0ddG7L1o3/
pjzFh7fKJP9TElpwnjzmSo9T6cCdnoc20mruYGbDFtEdZgLrNnbPD4VA0RjU/olRiZHzrmtCRsEl
zaC7XrIuA1Mk8lQcbojXfN3P2xleaYH3ew/GWtolBH0kUP8th3okb74Ap8WZkItTG/MYxk+q8jay
O45fFZcIpy4Qk2Qu89OKDC+ZTSoaEd4iRuFGxs0NjFSExye6xn5Wq/Sqp+Cm+lVJHXlCZb9PiF/k
xDs8dblfOYq1SNCdiD9lELfmeBUYW49M+i0LwciQHosyjvXbcjlr7rZEpU4omw65jysDKK1XqSQF
eQ1G2MjJc88nVbq+FXuqRVDbTN58/xIkwVV0SabCZvY6ekZtWhyqQ5dAQ62BW+1r8XVjpzGhyiNb
mdYNnkRby7niDN4N8t1UaUE1BGAJaY48eoAF4lj2qM0tSS+xhBtrv7wYBp0fNPWnX2Fo21q4RR9T
9A/akhQC0Dl0jPLsWL958OXHfcRRCklYDT6XhYRZzuJ8Q6uiniabSYdUzgOTmNB3qQ8WhYKTtG0/
sW7zzZivDzjuI6gN2EmAezw7zmU+ARZqVNGHHSOJg0STIP23zfHgxQPQ/Uw84wSY2szfauqiuhia
fQIoH4n11MMGCHIZRD2ME7Em7QCz+d6tvGYj5zP/SFMOD5BwqD/BDqagD7YPvev8kyM4/ldkYasB
9IILQUDdjsuIfAowk7Zq+4e/DCh1LTm/qG6RBMGiwvXkOk1c8BOawSEs+fAG/8GDFgtcnM9tGMdg
4KnulWUZsQDl8xZL+BVw+aSYSfeJ2yjwjcdrOan/1jTv7xMY5yCDdgtRAnCmmbw+HaZZeDQB776A
p2kY2zQCidT/vfzQE2nNtBUB85+9isf+yarnmo/o7ZOLzIt/lhjX81hvmeUd3M0f0OUXnSCqtDaW
GmnhdY8jwmFDs+ij38inqFyC8vZR9dCDDb8hd4bWxwOGsXFmSV3wL90yz51Ya2ihjaVXC9tn/ksv
yiUQWY3oZH+z61LKKaj924CBtwccVonXkGx7OYdw4749MpWNhFBR+wwN2xMxpFxSDtwfJzhY48XK
+QetuTE9iByTrEK5ybxmFJhIvwXEgbmxgwwhBSHrJ71wG4p08a4Zls/ZkQJ/YYPePjKHMyYRblZs
XehvE73JFN+REvNIrUyrCmG86XERY32zsS/DBFCU+dmI6ynvUJoNirbq8C9WHx9L4VGIvmn7PF3P
sjY2A/1iYccPvlQ0A1OXzLiYJLTseFM6AH4Q+edcm8J99sp0AXLGAbHyJ59tPdkhacmP3Bci+Djz
DyetiQwjwdVfSWliMJeY8WtrtxkghgjO8e2pteejqOO1H2XTfiuM/zQC5iPNMm6UDY0gZS+RgLGG
sI65IQRWi9Prx/8rZHL/UiEICWeE7ZPoh+duOdDvJBWsIbQHxZ5g6nV0yaLo5/9wQJ7Ycg0u3Ml8
FJOF30uISFkkDr4xL+Gk1gHKY/PhHM8FKUnMn0rkWejl2yeUmNMjHZ7/XJZM316+CPjYapD+8cIC
RRb6LeILmj/1b7FN+GH6lDZoMLc6LgsDWZNjw2o/y2r0Fz137nE20PJXupAZNY7kYMLitPDCjycR
X07Edn3aLi+zj1vSlTo3jBLfJUe33ueiEAEsnyIONxVsG1dzJCsHkZIxLIPyhFnM4meGGj3xk0zW
gKQuR70jQugbIqPL8AtkjL0sEfl5qev//8vNQ0dxYgCXy9MiukqnPs6zag1xFLtuyn9+ZP51a4L9
Z3g+WfJWtu3cmmMb496sOl0IPym9hiSFKno7cIGLQNtFvCx1acreoQXGXjbVAxCLcJWLyqsZDzxY
lyv3a8Pa3sA2ZF2kiBsh6V5o8Z6aammgTDbP82GaVYjJ77ODaekAu/bYn28ldbyr9efvJqbMg14U
QGnvscHWgyY/BR5xXT6Q1HkCwgylgBz32fCfJH7ENMyZDdukkWkwODrLmfyLS/OD3LmdDphpV728
onWNJgxWLPGm66IVn8TxhRAKi4sLNwx4aUNpisUIAtQ+1uJLjAjgruTcZ8waB1iL1nKX0EVpbW/p
Z24iVKOJEh5dOy3jjkLCFuyegOLdn2JB/eRc/zDH35L8NscIfxXUopYejg3qBxW/jEvJPcC5o+sC
Tn1SRMP8o2Q0VCrUkAWWZkbmYyei/wQDP6i/BP301dSukFMGFd9DEUhejeatbw1MOmqjP6w3hpBo
hr+cKjjFwUBZAoD1RtnaBfUBLuhLe11sjUNK0hJccNcygVPSQCpsoMpPIdqx1s/DmLULVB61orgX
cY9+sargwXzPWJkU//2qSFfELIa+oQdZsPNp7u9+6PjcuirKOgZ+5hp0IOTjtoVMCJ+6a1rrp9wz
0wX3HOjnABbVKlrnZYcwxLDs5V9UCj4l3czLZFneOvns/rv0cv5nqRYPaR9xBRu9A1odOwfh4bUu
XjOxqgD7pGoNydTSbyjY1fhaokqjl5DmSpt70QLgNTyjDi0umYXNypyc1uceNDyljx2TjLlKWFxI
o5OSxaSpNe+fP2Hpgsqn9HnMzdIS/W6POUS+e6qQU7aFKxHGS5va1Sl/M4WLm6sA5hFY03gtc9RY
17Q6tyxSnCPyIX3ngVcLHyTc9nmosTntL7KuEei98rXTxZD93uHHjX67FZzzRz33zd8/N5DnpSt9
uomcC+YZtpFrFdxpX4dP2Dor4OjmPvID9fWDBJ+JI9rat4daZ3aJ5D+R1AIGSD0r33qHHPDX8yVu
YncoGJsUw9QUWYP+QZsMOu76SJyvOjJOKsiBmHQJGiUBZ0qt93C0kQBqn4XpDtL40Yipu2sA4xzs
Kn2kjCKQA/afDhUy1vrvE6lrk90lHM52Csv4iTWrJ0mJO1NedQaOvRlQtdkHtzq7iYz3SDuS8u0L
fFiPb2wUZ+4Q6QjMdvATfjMduTD9zMvoeAxrQ/NqPDnFJxYPh9toeqvbqRN9xaKG6DOvyhV9vvlt
0qDIc3d3yQEj24r6GJ4JZs8agZDx71Q+iILODae1jZ54VgGxMcLQcTaNRCnOWz9GgG3Uj02nG0ng
M4M4O+D1XnbWQUs0KBc51AmjVQBXYz/vv8dbO1uPSIc/qmTmMyFjGljy+/VbSBAoKAx5nIA7PpDk
lF2ehaxM+GipUvKIByrWtSWPdlQOgAuaLdyON1fZJuWp5Pe9A87Pb3wABGocXWDpxw85j357T2oV
2P0iE0opKkaW1q09bc91TzLHWoINhHBkdlRJRK32wtbvS06415eNS2Z6wtPBsXqz8P//XrZDclhL
u/eZdLUL69XMF6+072Ga7EOP5ky2cOQ6Rnuw4lok77qoLdRQ5M6oNHd6ivV9hMWnU6Y4CobMQJHu
DL6/Id0jzbNVyse2387F3orc1/Do0kpxhs4cUjm9yynV6yqC/xj8Ht2memqJ1FLbMOhEkMQO6Ae/
tAfhxEPfnNMcOnnGVSaP16ijrU/a+V0iz6iU7VRcDofx9CWoH+zJz754ipHY6IL1onKV9A8jTqt1
MLoew8lMznzpf6BVQ4p8Ovox610vMyIactF1xBp152DXGrv0/tHSeiBiFsgrAjHxeNREeLIGstZl
71BDlSNzAkgvijL07bW7qsGk6QMMxMZci+d90OReXLhWwce5yqpOKlnlUGNbYv8Vye0HpMdvRZXe
snX/yHaPDqbU8pLrPHzoO3o8N+prIYoybBJa1pnisWePPfA835hfn9IJDmkLnQApcIMOcBeC743a
WJpsMi2fO5h5Ckaj3ih8T177uaZOwFVx09dJmO8mlLqEK+jdUtR2mPTl9m/YCv2GAnVkPH5fhUpC
AMU7WcaYQZR9rdFHnthplvTCc8R2UHa76ISrkQ7OCrhRwpJ7dStWf0BC9ymUsPEyGMvKX9e46AhY
aN7TR/zDeWxXlSFIejoMbSFCv57FIzR7cOyhVRdPj2bPcCCGo9nOo3V7CLwgAUn3B+X2yHywb3Vz
K8flKJeFKUdifQw4FppFI3zdd8k/Dpjf75QsgZQ4kpTmSUnqDfC+EhiTjqzTzlCVkhICNyKNCDJ/
EEAJqCZ5L1+MV9Rgp2eWcNQ9PLpF348ba9MkdAguApxf3mKvZQm66QY5ZHrOsJe2qVXtsxLoU6JC
BnVewj+Ha47j0jIe86Ba27DXY2UgW2RccCu7pY3DjJ3mt6xRC77cykoZnEvUuflU5uE+XBp9ATWz
K8h2yFOyU4uPdmjayRkhj1nIeJnkGgoHzUsxhgV2+/B4UdicWmVIMjsbj5ndW1DsGhuq+mvHlOED
Rg0JnkGUtF9iM485xADzBlYg4c5w1XzpLLkms6y4m/0KxCNKx3yZGytsnzbRgdBUWy6PuYbseEuA
IN37wylv36gmzfD5+92GYeDjptRQxMky8aZyrH6rsLjm6Ewsk3SuN+endFTyyq9icD31WjwNJuyS
KkNVInAUop/aEETEhWpXsHlOC2bvfCQ52Io1rRgzQULvfE2iw7iNpnzCpLLoYMgnkJqdRF4K61L8
qLzYKH2NHH1IU1hS9S4C62ZqhcJrXY5LEyVaFB6MON7a45DM5HJzHIhjk3U5QEmEcBHT3VoJPirM
cJJUZjK6Ez2R8oKFE/t0AsxNAESduWsCCAeD5BekdIw99PatKnXie8H3lVvJeMFG66mt8MULy21t
n4VKKEcMYc53w/BFfFLCnxPQFO5sVVWUv2+g+FnrWKY0iWGCqt0Zedcx6LQWxlqhZGGFZkUVjN0T
0WJ7jEnolIcG6rWF79cSV+xG27T16Z6J+eW9kFgyjM/4Fp4c66ccuQIDqoScn41UKEz3xk/UIC5O
1uFqlIGJYoKFjGu4af4D9urQFvGM/2LCt+TbyEY4wDugFEPFk4UWLwFJxoANM3ZEHyb8u8aBAKmC
VzVnhOAEhyU5DgWDf+0h7hi7JATqCddJKL0HXBA/o3L+kgVjGIRUxTNicaA+xeMlVXFpscSBDSSP
BXx4aZjhcdoFwIm8gYPWoMo8qXoAFPmJLU1Wzw5C2KH8Rjsn9qGQ/6FeX8YX9pH4LXCfGMwjMD9j
CZEptWup5PyWr7TW6k1F+vUhPjs8NsF40ZVdeY+HeLd5irrvSCKYZiGeHkuGimJrvWSWBKN9Ks7L
MaV5hEcORUu8KZMCutx14CYztgmmOSr/E7HFwqB+WQA6baWwfv1iGXjwiZLpacsD4McIxq0OGGRE
6cfWycHZbbj/iP21FKgvdSgy6OEJEDNu6yfTfhm7u6ntJ5coFSd/su/LanqYPU74vaQDPZ2J1Iis
bdm36eNsq8Zx7kr9KmWm7amoit4kmI2i5JslVDOWqf00EResNfZy3pnccUnVRwplrqKm11Flfg9X
kNgnmsR3xXpoLuThQjaDgWIoXBN9ddkkHXzxgBie3WubeDjY9Ztmv6ZmHzGTicQ0m925OzccVomQ
CSptfU+bzBS8t2l43hEReJxSciHuzT7q0CTRd5qWUoAAJdMfPWVPf4wG64U17t/ruJn/NWi/q/+Q
iMOfcOOtBH/yEOnAoeOKlJeY4ugEnT4YrvJ97yOEBSjtaOfF6kT5t8/oIf+xA3zzI9nGGDrwgw9y
29in8zDOjKuZDYQi/YulRDnTZGRHDA3fvPNwexdSi1Z4fk30xbJ3qx+2qmrwrZ9WPmwTw1IwVR7G
LkHDdUH9gaiZv8Ft0DLjq/6ZLxLr0QLqR90wcbZgwJAxdmtvPfAnSlLmTqAsfD8HB9kLGOoShuTF
PI7zbb8kdyu/WULvam709LHSRgSuO2ibuB4BmzsXYOMVifLIryarSrLoPsPbE4+TMK/iDsYiYWFp
bDVtYWvPsi+os7VLLus5KxyeyrffxpD41gThwlwAMFOuXm3YToKO3AtxqOJYKKOqwWCwr/2Z+JXT
QEkLwtVIIOcbX3rTnmg/TiFkQ015R7i+WUoapySmZVS+b1L05GRPKtgPTbaaF+FT0m7njVrbEKRw
YjJtsjoxwfVn3WXPZDtNfP7KPM57S9pViBiLjrvOCcwlPJr3Jrupv3o7DwWj74w1agK3cHYOl0nQ
TVtKGhWVr0tpwYd9ZjlZZg8/1q95dsYvQe+YWTKFek5Xa6WGkkiMnlYXpG8dxLHY+v4AN700G0ss
EYl/yGWUYA/Hr5DuyRGROxBVd7a3jqONZvDcBdzbPvGbOsVut0IuXnPHM8JsesW0TAn+g+up5chi
zyPq7tGkLbj7WiB10XLY9KK/oVA70cLXivI4U7dqJpHRA+jhhcIII0SLEUxPJZkFNeVckkAhff0f
BfhNOijKwZNaqih9vMXAXUcOOtnsJ0fr6rpvwXt0c7fkGaBm4krsJWZL6djaQ6JKCgqnWyfx+LHQ
kpgRkI30pGTyNIR/MwALCANv1LX/zxF7tWOIonA8xsi5GV6etiT7ZNkHsnnGIP3K8gqVgFjzMsIi
tL9evSQ0eZHiEhYlozo3AmpJZR6ZEBkKfbLPWKd4ybI95b5caG4BNLpHC9MI3/aMEpzPmh6AxOW2
JTebgO3DUZ466S0iqvEYTDWJWsEDmU2QMP1SmSph722SKKOjuDvS9H7CM1M6OOs57U1LEup1Lf8S
q3tn9u/PppBOLRJvqH0NWpuoKBd2NVng87f+euzxgyD8s3KINvIKzYlqNZGlI2VPb/k1A6lBqbeX
hnMWCDbJiKprHrIExO73wjTqWk435vIRHX2p14wdVfzW7TTvIjd2eUB2uIaeB3H78WtC6QKqLWJJ
4Ko+9q22aTPDpjzCUHACAM+aDwE7/S2Mo/0d6Gelx59OMldXSb2awcD25JOd3PuQTlZJjhIKXUpw
aj3y4o7g6YDMADcpcBHIKNP8L9q5jm9p7/fzpjE4y/sAfXpv7ADvRyursw0Amj5RDw1epWWC1Fx1
TeGfULSydPV8eTVbGqiubC7l3oGqanFN+WJ1yf0+nXd4Fbk4XeMMQzZ87qgN1oDMa1jbjWm3o0MH
HuvDsJ6oiQtn5UJ0bPhAknzV344mRt3hLmtCm9Gr+A2pdtBFAJ9w0n1M5IfWurzdFmVu+jkumEE3
OHhczZML6t7/nTpOC10s83akXHd5vLHBfkEzvhmWvsa7JwHavTfr2RcGlBGOML8BSByEgAKVcb9w
Lmn+0/DnK+YsVfXwZNergC3Q8TBNHt5fGFQOtfCe1xL0g0eplxFv2XT9GJP2mKOEIDBkFa5q7cL/
CqlQlDGqgPtrvAcinMWUExEMbECMryjMmlIlGJH4qTse9Kx0AaqNtRitxij9kUzhGhY5HaaTNVTT
P7/8z5k0OjrAiwphOzOKbQakxw/h2xca2Fm4yqSrqsXJXfeqYjgKPgU133htzlxsSkBwWdskJX3S
VKHWt/pEqy/dmuBGJIJnt+f1hG0uPDNbbyRf8/7vVnl7QxF1xGikuMFrLg4GMAeYR40J47aD5Wyq
4PE2kqA/5IXfs68bytmXWntQA995XPo5ds8qWZbhMVmUQLsBOYz2rnWJa4/wh8fmqTPsjmDEB8pu
R8lbMThAFmWtTg0kJTdSgIL1Qw/15GlJ3x+aBE4SiAnlD+IDjNCw8KHh4nVoUXKnnA0y02GGF3Ca
v9Z+vx0fjmkcJvLGkEYgl2TgcqkCnhgq9MCPs+dANOF4TAJ/JEJycxEuUfBWujIN5QZE9HGcHGrj
0unbZHlPrBuz0PPJfzVrJjAMP/scmvs2w0yRMi1XIQJMHVPyT4fw0C0D5HA1+E4xioyXGM3FB13T
D86wDU0fNV1OOhsyZIdXG322xzuwbImLLVcxQeNGIbTzaXdR4gK6kaDX0P5BO4WQQkmHWvDmeZDS
d9FYrLOzIGHaTztNYDoKeNTcfjW3MSBZfu++YJg3eI2XGynM7tvKQGzTrttGlpWF3rBuGNQ8x4sd
dtGsQHTs7l3QWo/xzakYwkE+d56WoT8J4SMU4pa8htYJvlb3nyJESJti+wW72fsXWQXoAIziIQd1
BR5VXQmvAEDYTOcRhsp6hzh6A7R++sUA3J9s3EiGh1pjspHvAodYseP+KtCSxLrzWTV43s/Y3p3P
9EsbxcZceDP94G38bBDNLIuOec2j9ChHAWO37jdtQx30G3Z/w3W9CoN7QZbWMr/fMoV9rVnpMtqC
q+yihwD9C0kEUl2N6L5x+4YaqYY+qZ+OXeVQd28mXqWrJv6b9d/medu21WkE+fEeCrXYFqEYQr1j
dDzVa2vgjYaLbFaVixW5rKW12739heMcfW6LIwgMVsMPIEWwHJYaI/kCLDkGeWUFEkWBbNn5g/3K
1gD/LY6y7ksFirSQgq7yEOmEXDYgIG0I/UePsok4ebX23h+c5oL14EH5+9GWAUXtibajhMR9kfRA
HNdQzP6OkNsXnOsJ3niGLrMmoo4BsARai2WVJ/zDCz8p+etDnI5W9OVsy4IB+Z96aTWL2BPVvtEM
jjIbwXTBdKdlwr1+RMIJeg1HQjWsZzzJDbcYJXLeXrFXcgzrmdaeTg5lpGknFlmPLsys70i3KqSR
ojjcOXXmPr+ik0D3mf8DF8cuG7Lpf/3MGHMxa4uAj1gfxOeUZi4YvukvTi5Ae1Dvwy8XpwTdTJEu
qxm10QtksOWroq7I1Qid2yeMhcDDRMz3fyE/nDbY8GD0LUMTrtDtkTAHIVzy9xIzpIozKspy6Nq8
i7+tgvsrL14Aqz0P6I2PV0UdEY5GnpmCmuja7XEFbZroGGY7X511TlDDx4QIO03QU75WqHuzSPJE
BJ+DMsePkfZ9SucKmBT5NxVIA9+JzCDUOBdGHknKbIMdZtnfXDpF5I/rEXcCYVN19qVYRDhKE6iY
iESRvZfGwfEXUbODEOiXarT+VZuTvMo/0MOLCukapOJVkfqJtQvwfMNFyNV6DHLZgLh+MmGCdbXD
5ZnwAyYNMQXQZxwKC4dlPmsOxrWAPtYLr9aUYIETnQ49e+AjbSxYz58Efb0TiTBqZ+bMfyCntMKC
21CExa1go4VfGYyokq75zLgnh9anjTLVyHhDd9c3RfOFp0bahhv5XPUL/JCWtnDmSFnB1LhZlt05
fYvq4Yn7UkXnT2gPJNzY89boer9Qqq/0OijCzUiWdmRHz8DqF9W1i904mLiAF/QtaEwYmQ19h2WN
4h5OU9uPM3vioHV3fEKFSm7TfHbdaTdvoWBXX/j8mF4a3IP+CJz/5WqA1bKQYfxpG6/EaV4PCPQY
WZja9SBD6mKIbPikWmEGW9COEfZyKKRvKbMentPxiULTshCqojIN4tiOaELxB2bU/Jd9y3LJhoIr
DC0uZs3Ahi23tB5SXlAo9SBXSDheUDiakMRt5pbid4tV01vrPiAOaP6kOXoh/UuTsR1z5CGqrJHZ
064ZOQiR7tHAOw8Hz/Ua5ikSNtpliAx1Cak0/qeLPAVHCo4vqzWVsMSbSJ+a0G4DaYuluCi4X2AI
1Y7gdclHx4YfE5hw++D9aus6cxgxmCQnZ2xXxw0LMCLajGkfSv+NOhhA/Mzz85V5UPFZl0LHN/UI
+gP2t/9IgtwjQ7MxH8Z2FzpeMmutsECdwu3zwck2Qk+Lbj3kkqpIH3KlLE2iISyZDzSP5ENECRWU
kgmFlhT/AJcKgioHSWq/U8bJdxyW1/Xo+V8di1CA/P4y1PGfLx6Xq/Gc/JyAwbcJmAVjOA+PuArW
YQ4QFoQVH99/74GEqqvMHItxbQ73s6u15LLY6eX72L+wWT1JKIqnRZqCn4Gr4FHFgk0JGRi11IDN
TV4k/DzRM2fpg1/CxZLLBMnajwfsyS34QT+l9aDr8fFhPNk1X5IYAe+fY9PcJYulr9yV+i6Pilq/
0dh1aXQBWefEGTFM1gEcwxpklnHuVC4Ej3nQe2fgmvQQ6KY6JI8oW/M3teJ4Kc2YTSbud7bddmxB
jq7YlEJC2XzfkU0L4xMDKvNTX0lqwhuShVWUFrWHDpdxiP6J/bAdpvvt9wdXSjbDKUpLGpGKzT6C
7JmLPfoMUsqTlLYwcH2+JhtLeNv9eQ5iWmRZ8u2lWojXXj7v0CbJituyuR4TcA1Kxg8E3DHi/Wmu
kcl1/GiffTnAUW/0i/jY80SpvvEPqnWPARReDvi4BNV60GSObtdkHCtzApQun/nShKsAjt/Gtmc4
ns0sbWtL7X1Cn04COT/UAtDU10N2NulGbd7Y7peonNkU9gHAm3+sahOr+CFDkkUXKfsqLCuRYEUp
7YsGGwlV0EyX3KNZMfnKI1V7lJocmxhKtkl3DXNhDjKvu+fvt3y5g2YycRtC+gsJQEJ52iJV9S8l
h29NtckhT12qEYRKLd4JvXJd6KQZTZGK81JS+JfAZ5q+mfjz6i1WeqpgB6s5RDckvjnodqxFKpSk
2I6lCgfyH7M5zvK6nluNjwKyT5EW7+iYwB6ojVvfwWNGZslx1mwbw4t1BNKOt9L9P9rz7Je1dj7V
lnt7aDjDhT2SDpLVbpkOEdIqyOL6Ei12GD4p0jPjHRZh0KpRzCyh8Tivkv/niGhAIEUZhU5YHFGd
udP/l942TY+edoBNuV1I1CZfYRyi5LkdOZpm2QJTPHoJOk6tUg3QsGB/qKq3XmU76MwQoq1dbYR1
qdFZQCXHEaLSdZ0CiyI34OdBKo/l48PsD57F4PxzvL3T8BKEpH5YIqxOdji1/jjPB908rCyHQTW2
Ic78eNtrHWy+PrnrEKnyhSvvl6oV57qENAf3QxP7YfkZukrJlhPc3aAXHRb1ojP2R69cQNciRnjW
a7ar+f5KHaFbWsGd6wItq3hK1Mu6tezXEWNSni/ths3OnDROnYPgcIi1wBLuTG7rMtGHtP05DoZT
BQz4WiyiDQRiV7jo6GKSJbGI6LuF2/Y5uKssHdIe1gM0nHfHDVMBfkmeyaLOTj2AM+5Cl0gG2LRa
SH6EWvixu//n7QRE22GSGTzDz6XFDoYeFifqQlWeidtVyKlgHzpGX/XinlpYCKJqAJe3/zta1aj8
PfFSjbMcZFTuADsswUB/YmAhsKTqplDnIGMmrjzeLuo93v+PJHcsLj2tGtPVX2rtNy8AuNzouend
hOBGmwtL9Z1gsGqMCmlNp4YZKlWioK5ZOuJbsxlzvcr39Qn6tnyizY/4JS6umilu5++xxzuczfKF
Y//pSLybEyCTnj50HRCjTXjEgU81I3gpmavTSYxeHq/+2mgrJW/dS0wbcUBj+uMSNjxBe6mWxmLZ
44tLviZ6eBTXkHBjMIAbt1m7Uteb17NpwO+7t2BeXgCbVBADE9sByRJF4AYZ6159BD6NG3eo7I7D
OLQM1WasnB0NMm6xfd/TxHS3bSpaK7iG77NWk5afoPHMrDE5TbkkhnS2soaE93nTK9Gwd/NzGoJI
7eimYGG5yVDYq0eJ5ytZKMj3Y5ub1IxyvgjTVFk53+idb/G7qoMOMa+AS8qSpJX0fmRltZzVREzf
oZY2jFdBta7OZwJd43jnLxdxGV8dolTe9x6ztphmrNoGojRjEXrMqhcjCg911Ls4CY4tCz9onFoP
2atzekgChDs/PrHVaY8DGE1N4PqJURQBFiYT/vg+zb3bY4weOE38eo3pALDSJJEwO6PbSEGyF3My
wSP1OL0Gi2LMy5z0EwsWB7ySvq3Vtgqu3KQLilV+ELLxYacLNOf94Y55ZtTFY3KObT9yfExw1zEs
rYOtXMsQ5zKiMrCLFWLkBsPOU9h2sd7NjY85YzCHxv35iz0X5tUoOP10ixiwpl7ouRJzzgyYqqeS
xNr9YJdeqLy7lymYcMUdL5Z8JHa5hGjnSDR5B12+uYslhDhN70iow2ucsTWhRPzktwT5VbrppvaY
55G2i3KCvFV3IX671RCTTJ5pvgGJXOT0PY48USLnWAucaZgnAZoelGcrftPm8wpsMfnJlf6PVLH3
uTKoPYY8Z35zch2kbP7DuxYOEY0PM0pwBLdciXs3TGCqDNGZAMglIYn90qleAcyitWIHxSY9z8La
RVGOchiMjo+u9pWUoP7h2QpOyKWbsTHaDWFwOraYa0afQ4sUoMZDH1iZUX4qz9phI+dalJdxbFoP
LnrX0DxOQtQ+gCWE+xPT2GboqvpwlTvVN2eRReDg7rgTJ5/Kk5eHYhnxlTL+u883WY3NcXZtuzex
zpb504a50pCbP89jsILQRegCYwiLZd3+kw2tG7xFelTIbsAsr0CNchLR3HgYuQN9fNoHQlLXqi6C
2CdbA8vRXOkL8iChFpPWuQpDOVFVY8t9K/13uBFlw3Zef5X3v6QJDiEUnrm8TLcKziM73oAlJUoN
gmwHWgudfdmuku09vgYdgvanuce1/PYtdbNO7F9gXWN6JF+tMC5UQcZTVRdg/N7g7oV57+fobekh
u3eghIYwWLxgVIcRGEodGGFM53thYL1HAdjNdzdT39vmudxN00eOj99u0VqYGKpfl1m7y3tnR6UP
s6z2c1Vo4Qb7z3s+jLNzXhdUBfAr6rbR/8xlYHc5mVrG8/5rSo72l2GPx+JqtVcUPw5+ZjRqR3+4
3We4kNj1EHJz3PyX1v/hcGgGeCjusHef/DyKL4atF9FF5kxTCl4snYX8vfDdRKOCDCHaBoCkGj15
r6uWF881ADXE6CmAj04ke+tGI2X26tM6AualhSSNgOUh/KQlnWjD9YgVgVpMlU0I6lE8xJZ4oVTQ
0u9nh9OlTkRjHvEKtVjb4iYiIwwIL+XrZsBr9XnJjWFa9CMGo0YSKAhoTmqzVb7LARLINSZotokP
0Jj6DJ7M734YXRe28fPGdd2JCDjmYIJrqptSNMAlK9LBXoYini1Z2LBCQPp/CdUjeAmo78WlWPKd
xEo05moCbdHpF9BCUzub1Z+jP2jY0B6iG4psKsqrbGEfYsw9NrYSyPwVJh8DBGTiLQBURt0kSyBY
ozMTuEyMOU06vba73UpMg0NawjI8O4G+lgeeQ90v2+q1IdwIycHJXLYK3K8l5CihuxSAYGS7xndC
DmcJqJqKHYDjvybOciVqhy1pdTQBK8LpVl80TvbYcuMTxN3MzfGF1XgmwbXyCIkA/z9Jxjam1Shz
QpwnKf1OpDplCo6WsqogEXjQdlFXZpu5gEXhk4xETPvbkOhspAdDNCy7a5sfi9G6bXQzSxIrVvTh
r9dECJHfzz6xV7BkHIWSHn2gz9AzAzczW04iidPwhXnBBIvGTJIS+H4c2DWqtxDopn1vkRNCv/Ro
D+G9wMgtgYceNyaNfvDM0qJcJrCPucV2WXd7GUFF5LBeJ3Ws1ngOy49+nD4qnHwIeCX4pFMuALXX
vYTPqAccy0IN/J4TBCZrgIzsg9FiurM1YMM6E7AbExGrt+Zv9lFy+8+e/ceejozb6vf050X8dfT+
S6eu+B9ov67dXmz4k2Kgl28ozY+q9B4lXK0KhO1Krmtlw3SKk/VDWwFsk2S6yij84OYxJiy+Ws6t
M81HL7bd7TgO5KvI4KDP8uCg97SI5hj0bUn9xtaD1dfTOra9SYbT8ItYdfIzJB3+VePnaHDgfQH7
eZlTgLCBndZ5vcYb/LhpJ3HPOy7W0CTH1fDxQLMC3/HVbOI6ApZLgrChn8rUzOYRIqhnV+bwgceM
R2vKi0aBS6iVuRxs/zuNORCXZLxhFv0ODrD5BxgTEpwZkRpFh/HOlN4ymXa80qUOGZZ/Q7jyCOGp
qZYHwlIVghgESxKHWlaq4q5DLVbE6JPWAaGb/Z1084GY6mVWBt/wvTxPGw6J/W26fpNaFqbE8Jla
FVEVyUZ3+CfeSOyYeby3LGdiZh/o8digeChdZ/eCb9VREBfm0S5T5V3ZuQ9O7HRW4uKc+JrbEnXp
5MhTXlgrdBNwRKIyDf4wF0NXidyxkga7D+wk0Vgxb/efh89YRjlTUTKxU7XJ4atxgKup1W5MnRtT
jgqV6GbSVwM3pYsNq0pyTj/5F9Wm3OnJAN54zfe4/mj3fVniL9zBy9Fgmsil1NzPpijUYjG8Y/GM
av/VKWENvGpIJJE+kMtYqKRO9NGlXJtnqeBQk5HDyfZTbN1N/+hbqF0FJxtMx919El8JJtHtMXjk
T+PDBKmpQCyLh+fmb8aq2XJ41hqPFqrJup2icqYkWu6OULcjjd1FmtbsLg72wqn47TsfgOthl4Sz
pUV8XdMHNqikfSu+YVWGBmmr6vaABHZDIjdi4mK9q70P/pG+NGErEOOfhXCV3MlpeSxxnCvXUjFO
1HlZcDZCadfCtRz1v8h+ttK55IMyzlgqBhsywETdF1AAobn3lnVecxcQwmJ+8SWFaFRCmmTL4u8L
xb/bQ+YWtz7xM1UJlcrKWePDuIV9/G7z+jLxr/YGh/TA0bYMKhVZFENnPvIPyG8OsJyAri8PEdax
pRivj1mmzT3+GmNru/p4LrrlnWe0iigecoMKuRK+v9Ky3NTxLbJiPN7bI6sCvKzJyjj573uV+HXi
mkj0ecbuaaOtGqprXBmvGS4X9ziirbNVjl/tKCU5NSakgkuWzhq/fhhKAAeGOf4/3SHpKCYitQP8
0+2wA+usNTiGs/rKJZxn4co60Vunyr4DGFbt6U+EOO8dVoVKL0jHyBMl70Po6vQxmHAZj2jHsjbL
4FaIUiCCGwbrckLM8dEHTqsG+HQQNnEx5uRGZVdg/T+NY69MfLnGqb9vxhgKgqPuVyxqjRnTv82g
ApUWQvbQzJK7PnWRkfweiGyRDkAUNjrxsxVPJdzDiM7c1NNQRaHrMgcmQKFFYMZKlWLo3Eh1TweQ
7+pM2d+RFAuynfMGDHfOipXtOUFNjnqh2uaP8ZO/B+GWQufu9NA/Z3wyTTWLLCPu9A+X1u8Uy9Tu
TMcEg3Hb3YXQfWXha1ToZijH6SgYhf0WaoWopWn3I4lhmobbUdmU1Q0s4yzJB4cRaeub2cVr6bIx
4KOx6XxAnnrIwjNfaRnK7LZg8JMvrPZd6J5E20ragij7lieMpQfPTcp14iqyBkpxIJe9da+trUnd
dziYHEAUCNBebroHSOHDZMaARnaHaCAaoTzNpiBOnNDL/QOnvq1iVzuNqmY3UbzOS9ao5dLecyh0
uUw3sygXDjSdx8Fe3/E/PqPNrPE1Q3GJ7iMoyN8Y467TNpLMSjKbyAJvDOrbDcHnCvJ8dyeUH/iK
mNDBUU6WXcgTRB5GHV7NzjyN0NmSZWdd3cg59r03TAf1QE/WrAcSX8yjqrxGkzapvCByGt0rtNTN
9HM5aZQvtBCIhHO2mtxJYd9VU6xZo65XezjDnx6xJkI5yWD6NyfZpKy3WzfzN34CP8guG19NcKkm
aOliwQQX9IasrSMcn8u2ZLvxj+kRElmB0KeQ/MVMOfelcxCW+9mXVlYZ8YPqo1LpHvLVPkS7qa9E
0gdPaju1TOvvDdhzqkTLtzTK4OQ3XHPL7PMYaxW81odjJ9T3q1qyKtKfEJ5zf7yF9UtAo0OxAP5u
RPWAMZbKJZyFqKFZ9m4++3FCA/g42v7ByzYWcCfCnvaugVgwXztemuKQ4clX7zV+UPOg797xD9Ib
F0hSRZVJ340Sd4DF7uEZTeutkgqK91wWLWyhfvEbrehXcsoCr/q5zJApL8BPEfSAEx9w9x+j/rvt
WDUbCRrWYreu3lPRZeTqUz/YgVqJ0Sgf+66xTHRhkD5jx+pGzMotrkq7ouKXBT+YRl19PmlkppwD
l0gZObx4pV1EKYEHDqeVwSxBntbpEVeor5EhSIF0px5GLrZz2dAX2FFXpaTD29IyTNbZpeD4dnsO
eZ6HJ4fkKtsIUgRbkL/y0ZibQESg2oUPhkhC0DZhZCEVQ9/V4etWa/75ItaZtAurl1necL07ov1w
U8Sv+g2LRhpIGG/qt3QQuwtvqCvTAERtlhkHpzSwSqzdMGXgkSUR32bf/9cddxYfoaSFsRJca1rr
RaDX5K6oty/gT17NGTdEr+FdXWUubICUfUwgLyv/9pntsrQ3ZnFZUj16zgbq064vUkVseH64xKyb
fJffJSePpTJPCWYOk7LHodLPlzzhhAJaCM2U5jssGsFnVYjcdnlRwUaON30vQz2Uu7y5N8vtg/hU
8KPy939/1FTi9mLsI1jckvWmpfkCnbLkKSnuPv1exoetWemzdBGuwf4rW4jLFhr0Hm+xkcSj9tik
wiZDAxTdH1E01M1nLwyN+TwvILEFq/zoiDCfNMTUjqJHeZTP8khs7nxvjJ1Juseh7tcLLlIVfMa+
9jPRBSDKehinN5n9FlJjCm1dDW9ZlSsSOneB3SV4+RkUAwuRm6NS5WqDA7sI3CbTS2fsb1Lp3n8J
u+spRyvEsB3px1tv913kjMrVsiQixYkNybZBF336NCnPg/Sp6XeRjiIzezdgLz2jZU7llB5cd/io
fwCNDhDBz3PqapScn8UNavKWzLHsq3BnLT77B8SBtFvNVSbI0lHvz2I4p4KMUHYewrx18+yJSv5d
NgIskdu1bhk5ObXhhK3r4j6E5maf1FpUWu8xnyozZpaE1sKMFvQ+1FPdMeQTu+J5Y1Ei/NA2kkzD
MG9Q30Z5+TFEFgAixupT/HKFt+rPn3CLflq1DGB9r1cTwaQzmVp3LmxWqDDsmt4xy7GCMBcj3oGW
vvU1G3oo8dabSskIB0z/FZ78wlM/u8jiw7hgypgxnJpCgdWXyRTGJmzYAF7YBXJ4scPV1knW6XeS
hzaQLg3MrWuGFG2SClMmYI3p+rqcCiwLp26EPzZDDtxWFpA3deF+/mbkPfG2262pyndojSFWXZo9
TIrAY7a4bpTAiPX4JN8xF3kbS8LRldqVMiNJuEiBewFHUFVJesgebWs7U/QO+dafiEiPa7BAJgLE
2C1+/EOXH7INoFFXavRLiSFxhhS+6N6EkitmSA6H+XnePGTb7+TAt5dTeRtPIui93e1BJTpdN9Vq
4DioXvbon2HfkSthdZpc6UsHusat8RUyb7Z2BKvMMYR4RbFzwyYUHNLJnI8JV2TbA9fuqeWufYbx
dDsuK9ruMkwSVXrYWrg6XkawIOUcxjoILqlHiez+6XbVBMhgBTpMUAuJKCyb1lEY0M9JppzXTvCh
iDECnDhnLteziY7Lf3O5l1loS/YFz7FxTdQorjU0BhtrrM2TUjoJvWu2U3G64XdfJCsj7EyUrRns
XsbzZktNpkWvEhJQsluAn/+pVn2dH2hCiCaUQ2teiS/JFl6f6Eq4rtJtdzkBCWivgrYzTVm5GoEA
ElPVCNyG6wyOdgbXzs9g9u1UJBCw/jj4MRS1Ty0+THr+Ed7qzG7+lgEwsaODa5nxjiM1xMqvFPqo
Iod+Lmyv0FL9RViLgZqcEppvAnGSUvQAYxU9iLdgzF9WpjH3TMDou10Yf7hft6L6sPFfuKcrMEpe
Ljj8oyPj6x0kvm3TngbDifr2BYTbHxayoaCdMlpOOUz0ee2lkCjiy7xlW/d7nj73CV9HPx6SgLC8
Kc7fufm6T3p3/7O/fqvCer2rIh8QtiH1FgvYl1a0+U7dWi0L7toB3dTcIgkcxubK7cc8EqKaofsi
mcMmmnByfxK8eJSqTwmfk7yDWBf6mWcKUdTyehgC49Z0CyG6wAlJ3gtY+fba38khUhQ1fWMZ8fgI
WIVkHzxUk3rLi7dvpGOfnscfs/6eHZ2UHAgZS3VKcglZp0w1uT89t5+Wu2USq8DgJtDon0chvtW/
sxlsLcC0WPdn+K4Hw0L33oP99NJC2hy5eCqROTxqa56pGFcfVbPcX+yKZjfiwVXPTulv2NSZ82C3
Uld+AXvl6mFg6m5MgufVzWH9XWFRm1rNMSKc6Jd1r6saI2ojLKG0X3dIaJUPLgC0pRVPO03P5Xfc
DfYK9DNsyhuw7kHSG9NjJi3BpDWRrUamV5ABlBG1K9pN2n8ovhn76yhXJkGwOdr8BHqc4/8Z/qZi
YENlGfdFxXHcqsIsWadFq1ZyCnxuuq1HhfDrXKy4XTOAFo8QqaoekfRSGhbYlroGH6vL0hwzhzdF
1VRhsSp9J0qY9qFqHcOvGo8vPKXIOJAcHQZ+3zfKJRLeKkoQTJNRLilhMf9aXgcN0FC1xfhqqMGS
e3NxwS40gMvBIVb4V0PPI6+pnD1fT8fisR/hDHRpz7VSBVW8RC2mGly9Z3pSYsmxEM3+NJAQQrLn
2VxmyzX9xGyF+HmHOlXDRqPGQ39Asw105rqQgEnE71m4BtpdiXCMsgpMtlLx5Iqq+Qm6HEsNKA7y
gjB+9qyWDdZ53Fo2QB+MzBV0LwXvUUb4LIaXamEO9y9Yu4hmvpvolJRV0qMm9tRd8EuK/8AdULyK
98RzsZY2pnrTTaPnqP/+eqpZ/ymGWtUDll9tJ8QLhI+QEnCwyE/93e5lX6aJVf31nDsGFj75ni27
CS3pc1GG9q2TREfy3Z1eWEB7UsDzQDVZHKz+We12TbNMb2EnrJuRGrr9joOwgijZjIsVGvzq4tOk
D1yGLmNPxWVa53Ns8mkmyURrT+zI8NVQTMYnfF+bBkdfE64Wf8WxfQA5kpnyBM1GIT8k8izrLkW7
IEyQt5SCiqwl5yL4YZks003FCnU4EgcqYEw+9yntwFnFy/dNGaT2nRd+6Hj+pXdgOq5h3Qq0mF5J
kgQET3o82LKDSc1FeVfCor4HcEkvrgTU8waUwZ5w1nTqbensIh2dhXqGMpeRYpMn0oYd8jyhdYK+
tSCKbGH7xOBC97zVhWa5BmVMTpmDtdeQmJBSKi9Yuprq9EbtXINCANQ2PBSWuKvpYlYwOwC/xOf0
xitH3paYFg4ngv1nk1Jd2FImTtHEx12M++NXJ+9w94k66WwxfTyPrHMhyP0xGcI+HU0Xlz+P3BoR
7umtqMTmiUDiiG46Z5oZKjpvjXw1pvjPt6nsmoesOBfkewdxkXxvhCtNkfn2Y9MHvxnM5TdLfCcf
uezH+Lo5lYY4OD/gNacwsgzb12qwx3Syw66hMC53ViGTKLLay0eUkcYu8LAfeooiMo0mWn84HDuT
kGuKKwX4Qo41CnZgoKQesY3k2NqSsIz/nG+I71qfW1oFZ7kOfv+KOhQjS1uxH9TQfZdt2uqz4Xq9
9aYdHZyaKDdi3Wi4PO/q3yuk62hX5EzI5/K5lUOKJ0y9BtDN4C9hgOI7ELCpV0iMs6wrfjaW9Eba
+M3KIEptVu9dxxClcn01zhGXKGXv2ZB0UjXeUnkFfR46R/fSHBetdpkRTzfo+byX8Z9SWJKvXVI4
6Bf5S/avANO7ihdG8HAHhxkFEpjO60ob6UI/9GXQfnybYgVhhCrzf7T1CunWiUBzlUx9jFD9IYj/
kDLFvRmHQ3XzX2yZIDWv525TRSqRd+FknOkhK2DwQTVJzm42XJ0QhI4xK6lnQ4xeWVQ2lI6lww9m
XOgjWNkixUT+HgZYrzJnDH7m294Q4eb9X5AI016Vlct++I4cwetLprX+j1u4mkaAwPPcw5X/b447
Acww8bf/BGPIgKbw0FMhkXHR9jloQxtg6/Mykwpkv/rNciNBM+Y/+SZfRdxHj3JiiL6qcLX5ZF9R
IDwQvBWTGq9V9VBKV09qdXAqsgjLNavFO8ggcz6s43toG1MSpeSRE1KgUVfzurz27gwPDhe31gvb
DA7UDJqtowzyg1zGci1lUFq21leAdv3u7xgib9xi8c9iIOwOhjMnparPRYr1KzUfGMNstjyDtsRY
FGm5ErmoL0v1sWbuqXRLe+dqs3vk3HhQknAB3BBQiYi5aXqwTWctFgZLew1jpxBbOXB8NFqIENFo
bSmlaZ8em3+l9gh1duVaYN0z36HJeHdgiZOz8t8Ga0fJKJ5sfMo+O3ryNPwycxlxA/KIPdpQdxpJ
/k4X3FKWxXNyJTAIIqGvSHjLH1EUC4VIuOar3bkhiUPngEPPlAFKyOgoOXqV4goy4wxB9WUorVdQ
xj4mEvK88qy4DefRBssoejbWJlTl3B7NJr6hvNgtnvyMtnZxIvIzaXuzkqpTMOjsy0rNFVdlbMU1
yNjg6RTFhHgv02T+J9pCrzTu/Xjs9rZQ234LhrWPC893uxKmUf0erzgA44ZQY2grgBOKXTyORz05
X/UpmcC5ION2hf6F4rgwjICAtRzjp651FLbO0l0MLfBYgmLKXDWTmvkJuF4YqymEwBrmIyk9WTLc
LiBriA42h2CXuaeQvvLzxJgLOSwe8XBPFhLxXoRR47u28vOMQtYGFuQ9PxxZHq58y2EoEqPc23LG
Ii4pAsGAgZMqKwLJJdApBW65Ljly7XFUeDJcztso1zj8y8G96F9r81mA+UInT2coMncxwgO0rGGY
YjHunQ5jHMBKUFFCzMGll2XBOsKVye/t6Aws3Gg+E9Eh7e3G6okl61P+dQtpVvkGOM3PuVvTWXck
Ixwm15Ys1/0vm01+5MJRt1a6IFA6jfAHy7VG7w9fGt1X0RZk27XezmN2OIT0N9fLk7xrBBMZbP5j
bfQs14wF9Tlt5zaB6GPhmN23UK3n5+qAjYH6NVlSfmqfEKdBHAK9yowqwoou0ADEKEXQzLEtYx5V
hrXmjbobfsRwIqTFfroq0jRY/fgHOCUlE1TlHcvNKZfvKaKXeqv4c0LBy5ZqLZvLA/ZNEr2iPQEP
uKh0mdKLecBZMoNSdut/1E9kIDPKHAK++P6r0Q+PFjWAx34PKOLGmKcWG09p3Q9VNw4RrQUK9stv
zu1UsDB0LL0eSmF0qbSiQnonOF/QxnPnPy7XWiUcveWvht0pwei0xoZDllR4O6j7xgKlB+yAyV8t
ObkLRc6xrtW7KuFZxnrY6yEerwBIHOy365hHqJEX9xn25FQFjsg9yoCPBE52R3aFYaoUBiIqdk5/
5WW0tnPsrPPKgm6/9o5CgCajCbSKBNYdgPIk0+kTkdeqXytNKR60F0Obr7J4FKjE6AxUH1tUqPJ8
u1UgHvegfb+UpF/vQLL0qf+kqh+f1YPkKX6GUruZyGnt1Dr6crsIu9iOEUwCxBFfLBDA8QU2UMjx
XEbuOmmi+m771IBG6Htu23Eigzl7Soa8oJrjFRB/n0O/cn9IxasyXaaUBCH8ooEZof5p5Qx7vSZ4
CENcIrV+NHS4pN6DbxcwcrT7V2RgcSxUk4AKoeA2zmaOuPfBHFcJVV4HnKjAIbNWMrpGJHQba93A
q38Q5rwpeF5hEqqfR1R29VICb4iaKBiI57r58+N5RB/NJEyXJSNGwf75iS4hV3+ejBgj8S9M2rwn
0pfiAnWEGtXpAiIbH29IGhz0a1Gyj5/amZZVIxWAR4HJBWrMeY9rNbIw9EiOCmIkuyuL+yMIGjen
7wWkYRVwoTzZtq+p4yU+sCFKE2rK/iNoGSngVnoW7/4raOnNjKZa1Zeqd5GyjQtO0Gi2h3LfKyXz
WbqcU2BYI7ihI7tP86HS1y/nX/7nB0Ekddv72XQCOSM0oHp8CzTKZ9JU26HR7ayik+aeoHjeMk46
uBhaEJS61LvpMhbZGY/walAAWE7CZX7F9o3rfV9RVNo7Tx6LtyPKvXy4sHpY7wuzW50qz6fuWHJt
SqFvDqOqJCPWIx7oBdpKQA3ud++618EMaPuV353iB0j6+C//WAHRAQYcOMa+Q2sPPDMpuQ4noejf
JfuuMR6ICi7KZp4OjQjTbxoNWtWGOQBvsqWBzYiFNl2J6RklIp8UI2lm/6LWU/teoXgEnCuW/6sp
Pcn1loEoT9eA8AlGn/VxcloRZU08M6Hj/ty+2VkLNRXcO2VTzfV9G+JGArCwWZ/QPDmo6+6UBwZb
XhO4Jap0C1euxG2v46FMoxbL5p6uXTcx+NY5hUEJRYd3dRBGRtYvDACZB6eYUEncG0hGXmgTXMtm
FSqBelSwxm4typOkoy/VwLAatZEBFwfROLsAsAGXklpz/TySP3B0miLeyIChv0erg3hmwta0p6fK
hgl655QEu5mfJn7hKX+nPzhoE+r+yF1B0lnhqG9xNPq8N0YiaRMLIzRrKHEHYPGxGbv35W/9JNAW
1a5nBOVU1nPz5AoD/+5vlSTk/JAIj4pvvCF3KDh70rwxkimsAgsqNavBHg/ivbknDUoU/mAtdXkp
cWXVQ3sBwMP9DTaqe5UGQbUmMUiYiLpoXZfNccRkagKHxugeSRjxK3jjUx83CzManARq7hrPKq41
rLak9TMC5FQRmrU2dPo9DRqtDRJZOIIPDc7KSAkW5U+y9WMLc2VI9CfJgObA8H3OjQibL5moNKoD
WREoHKNoV1hxEEyOMeX1Ig4dYMXbvfWedz38Ak3F4KjGFD1uPCKkkjMJ5PT3PtuBwBLrYFA/mMPj
bK+XLb5ykpJt20vPugRDlJCvM++eP0aZWFzkFQh61J1zWWqAEYyLeTih6icbvRem/lJ/y8vctxOD
PCWpaMR8AEXElNkmXuBmjYEMRw1L04V7hTx+BaU0DaTF8f6TozvKqotD3v9QJ7sUPF6zPcOYbJYP
NFAN+rJ1bc3a9RsR8SJOesxUFMevwcXqAYPa2cg3/+keAY2zP6rV0C4abrXJNUgXteMCBTCBNuL6
IL0Jt/1rnWRJFHFW4YiRqcWC0VgLK3CYQ5dEHI7LVF5uIOawXwq+HhFWUodriGy2YeE6V5MSwcOd
FDOTe+RBaSlCxWGUbeOCrtpccW5IiY5XAtlUadmvdVGWdsQQgR2jZGDVYOho5nO4LASfsr/sycLp
P2gQ6pLI0ux3GsicKMeh9VyQhobhyyocYhr051IUZ3qO3DtyZvr98HXSxkziNRGr9fKOQoqJeN7e
iz2JhrcufH0IhwqfwKPu/dIui4nXvG9DwS42shy12bSapMNh2sfyxWbpoznNNFloHmYF7LpPPV2I
t7bLdzX9ZK9qlEdANkMYEVSv1bZQmOhDNbeq+me1+epSsPaK8PDf7Fczk2EpxZUgSUBM2sdbQUhg
WV6VE79hmDpH+NQP57NKpFmN9lFhi/uvH0tJ6oPoSMmK3viXPLEb+ca2GWdnOmc7zk8LpZL9Gkyo
pKlbO59mdYkQkKOs2o1d5PTpCYTtazoTCvhYlXPMSTLbcnwm8jSUIWPsixDCejLoh5E3IKBMWbZG
aRA/tPlsNCsVNdNedAjBKbHJHVbq6IE+/2x8g2D+O+Cr0m3VBhkuchCZAXYgUxiIfY8cUvKPHnOX
u8SIogowMr0X8xgTisdgAguejNxKqh5LBW7eEM6+lt1SiJ00qI0V9j42i9PQiCawmKkzHBSvciyO
d4Mx504OSJUkS9PYchy8+jJ471y6GoxXa2bL7XW3oNLnZAjJKyl6eJA3rGGvYwuRaE5lBK8rhjcm
4rzZoz1l0SoZejkw37qLPrtiDxJCWBheTEoNDatVwz3W/XzXX6nzxEgy8I1YgAq9UBiP1DagcTPh
plhvZZrN1bKjhYM1l72w8g9NFffcIU0/tcp6hQSIhu87KrTdarWFPNQLbEW7P3aDc+7aIXfAzGE5
AmWvnEf3pewcLp73zAAfVgiCOyuBGYosumhg0zMJvTwzX4c1B8jJSldm74OnpL2TANUNZPjPAUHb
SjcrMuIf1HV60Lk6+NVdC5xR594Cf3JikGc1IsvCmVUqgm4rcomBbD0UoB3FQMMSrM8zT6WrLrft
z+46b1vv8pYIXGzVn7a6/tvyUUczSSHXSWTVeJ3s+pYcnHmJj1ONFTCCNN+eLB0lzOY8H9ceM9oz
/PsiCBMGx6pG5Hw/rCXG31xjxkDK7ULSRVVvDl5VWXmFBefncp1xO/H80HfZBfnPQqfXysShyXaq
TIow1eabRcXSCDCU0cV1PPhRoSFSS0Lqwkk48ry5JXE7rPuLCAeyPBfQALjuizAosN3Pqx8iEtQz
j6qQSb3fVbr5eboX/cv7xKwz+HBV0riAKMizbTXMxKKoZnYxmUfWLAEvyl5kIfzds5fueXbh5kF+
gwz37jkoYNytMklm/tf1u/AsSbiSb5p9uc/BZqWVtOwETnMzBtRKvyTy+/8kEY++68mKsgjrxKeK
+a3mOl8RFb2dwXjgoRNYF8/DgBGVJC9p/vZQMH9YGCft7uDtNdWV0s/ynn1QWgynJ6yJ0RZqYcgI
eLv+m9fHuLK8mO4DMhVxpi7Bdg51OggujGFqclGd/gZmO0vko+rmv0WMqTWGFgl9UTjRwW+Yvbtq
LEpqpyh45U8ylFb216T5eGk07ulOP/aPyMfZ/roLR+pySFwcPVK/gzJscpAL5eKXu9eg6g7A/TCy
/2iphdRBqANjPfXJrZunT78MbCKFPP8eRuga29U+mlYW820WpC+VdxB6jaVdpDG7lKDjdsPRc2mY
OiyCSPoOD4YCvBiYMlz73wgy812bKTwGe000c1AHQWQG4EX0sf+ynyst0n9Cf9mLVN8CTgCEVIgb
7v1w54G/j5Sa16DUEG0b7zgfOsdveKc0b9qHQsXjzFA/1yA4d1eCkans3YHhwFUYaBKwCdZHrWsv
9xvSSX0Ed4Bs/UxW6/HaRduG9AXp74jJmpk2s9IRkZscw44wCkzVUG6pcBwrxfhG09taQogZvPAf
XsK0wcj8fT7lxFghY/reeU7iGE4kzMKOS9Mkxs99nxqKeFCAFWc9iaci+ZqGAeZ7p3++JOySXqkG
cNXDxGVUQqRBUFkfdAGMtnAgSuj39xVet3RuFPbo3N1nPVwJtWCEWeY/3kumDD61cn5+AfUMOGii
jdIPiOHOxX2OjVnA0Pb9Z8eDmPnt2etvUx5PuQuBONvvM2pnqYH6HW7plRbIGMO6N7oGBYWPJTDH
URkeBqLs2lJpt2Njm4Hv+OvGMlWa4/e+aEHBUS0C8hJJSlmP4ZSFSi2TZpMMnVwsud//fVAf4dq4
/PA4T2lNqMJKui0tgTCembb+c+QnQBkFUnam+frGATRPEbWeG+9NAmDzs/c7s3TgFyPDj7Oaj9+n
xXxEdMJ/+9WebQQdKoQ6ZM9WGj8MFcQelFzar9glpGzHzrKvbT42YTQgMqQu/arAwiUzxzqBpk2s
tDZIeb6pOYckAHNvjxPZjRiaQhuP8G01UTxmprbZ/GNlQC+f+f5pXqR0dTLpGig3TdKQsSfla8Q3
FjYP+dxQhIilyUKoKAJTdpKCI+eqTgHI5koDghW5I4HErBQ83H4a8CRPSZpw99bXnrbFYz6LvcSR
PlLESyEZb6eJ0vB0UXI4I5p1iwchdSX/m9rzBYOOIQqgGboF/Y8Q1hRgtvVBV+lvdEzKTO2A9FmA
ponQ5tQ1JkPRTWJb891nWf2NpLnO995b/8rMBQF4Unu1GrbIawGaJGkxcecdee/h4Ir1lKA8197+
bPbwGiNSl0r9T5Svm+UO60ALaC25+vyLxrbMVNd4FtpNfO7tu+iTqxMcK/DAS4B2cMZ3I45p1MwV
fe6PUzdnrcLNyQ1zfEsSdpXS5J6Arr4wWK921io4TfDTAOaXDmtMCq/a/bwUrsnbagiHYSG8GMAr
gqdn+HQUEfpBM5+bnMvpY8ApgUNqQ943jFCuoUAvNki/rRG3KOnUtENKwZuTm7QtJ+0xQY2V8WvQ
GaUHU0Rzueoac8Pyy3VwtG63gKY3JnSoaXWa86E2uHZrCDAIf8WXKhrwbfT7uyhDwLIFjVFbVz8d
mpB0Hyuknc97B6KCII76JmZ2xJdiSW3sQZf6CFOOewg4qIGAuCFE7/PyWH5pdOPGCAymO87SaYre
Z+y1lEQ8N82YXIFg1ySjjsK4qlQQl6RJ63YD4WkBYl0pCegZpS4oHzukN5oGGcVFam+r2wO5XWfi
WPhWXydmtq9VK+DFo7thibYLb6ne0llRu9VxmfpCO3sb/4+jbguDbo6W3aTT01Lc3PUaUGg+rYoB
6NbzZgp3nHXWEpas+Ihu8e3PfCyzGKHWpksPGPzWyaptRYFyYn2kKULdZ06N271QfdfTxWckaNBn
v3ebx7CXArYwk0SsXNDZYHhxZAKkjCHusebOkC/DI0quAGmMYBvt1QEf7Mo2O7f8AqAShefMP7o/
BweqLq4w1NGj+AEDxK1wbiaxmX5wQ/BPV/Yc68LW/6v5MbbSHUq/uP/P2LouCyPhcUGo0BXUgfUO
9HLjuItizy74hqP+rr3xns/9KxX23w49XKOEA2oVuVBkNipp1Ubo/dH3RIHMas4LKwN3bflGpMbX
7+tllb2ZqfTkjg1dpyDS62eS2S7Z+r7Eg2vTP342cy+4TpNT91TmPddySGYKtsRmWDiE+NiZhyhF
A/GRKQfN2GEODB9AmU7zBXb9TxeGHwVNZU8jIHXUHrjOd650BBt61n9iTf/C+STAzyUEQgXDPIfy
QdOUKwH7pQggo51eOi75tbnLlYvvMEO+uO3RicbhTkJvpW0OQgiRumuQRd2jh6LnhFNA9mi/BbxY
yGCmzAUZt64bblnvUVGbych2LOSHjr7uFAzyLM4DbhgdxoeK5ertx/R/b01Se8yFZxDyOD8yW1/j
er2wuXrITXT8iSqk19iulVTe5DMdcnxEca/Eh6M/KGxIoF8hAdxIimlGb7DCwqdVEhyaJ7vB+ImZ
eGmAGV7hbxvM2AFCfWPUvwfuDQorba34lYOme8eZeCAkh83i/Btu3o0go/G6hhlbcGpJnRnf6VPt
IeYzvJpEz1vnIQ/vGkpcUFGmS8uPetwmNdLmfgKgNE6wIGNOlwh3ZKKgXNNcuZN5yRsZYrvwhoJO
1amHvObB2Qpmq3OChO2teYe4f6/A5KuKZoTg3wne8zt3lEH9ArPuPciNk5GGADA0gofEZnfNnhqW
O8FsVUNXwLgVNIfMoxlqJfsz6oBvo4YcpxiRJlQAbP+Q8R2RspKYkzGCZijFPGIJruz5sSnxED6U
NX+3PFtFk4oqAovPFPpyu5Mo3wC4Z98cxrTKPyBKKtk3TgBQm4jtp2CC2mq6K0buLPMpKbWCsB1L
6SRNXVtHOaM5CBecBJc7jwenMesQUfsE8c4PGTSEhY89AqGuRjy2d+6DZVO6124f/WBAjEATFPOn
fowENppSB4gM6HPcR5VdhznOXNdRvDF/YlbyRDiAT/gqTQEWqnPp3WUEvp1BhPeITwZB8xanIp1K
WlQOCycKc6IoeyWIM8QFHpWJqqvR4uHneIJaZ2TYHqNaqtGPkNGKqtLzzZ2uvuGfVmlzXijOToaV
n6D46jbLlWNGYYb65A3oE9RBjOwJy7GwPGfgfjiLtokh+3s7MNEYow8NbKr87CWPSHoZ8mQ5G74w
DgTYyeS4gC0EID/Bnpm5MYMKkJtDEzgZCyOt1VEKbZTCr/nhcSgwIiVU/jDh1qXx9u8ZhAs6rOoJ
n27uT82QEjQW8YXLq1/HoB21GYwqioB8PktwJDtD7HZFvpdFHkPZbCiGfAsqib2gJb57vWgbfYs8
D3Y4yQd4DqQAwX6GHYrEkipN9f3c5xXkLgg3PNdQslseY7+nSls950f3pIPLqvNcZWJZad05eD0V
DiZ/WyccWh9+8+TmayB6j8eEOZ/Qp1FpV2Pi+zFl9lQYhFYHXCH2NdFWlBhvPHQ1UpnQi7MA2uR8
rpUr1CmYTT1xldqEh101oKYpsiug+fMAeSSG3aH//EVYbdlJsZwzQCn0kYEfMbOWipUW1fXY2oo4
h+1x/gI3uKfb7qq6prrfW9gGQPfpeyon5urpF9wvrIw5YYuytlHu0+p/4qPp8aQiyxuq5ay7XOdw
7mqfpBPl8z9WmDFoPs/pxHUFr+CQfBw8PU86XmXGsPGIqASl62S0a2V9pBmDGafhuXiVMdmT8xdx
1FPOpzpHEiKGfcHoKNtuDHI60hDd0CikQ8jZXs0NJZ19RctNeAwB/eLnV/Qc/r05kMR/9EuJBfcw
MPse3eHu9DT0+6wHMgHRy7S+Sb9IhpkeluCEocppe1ouZHCCqQk/l4LIh+8xN4HMjhhSi3RwORWP
B9Fj6r8BDe5h//pVGU7eWO0nDifI9IIWqEXROAk241+/mpMOITr14SfnReSNnsqpu0ycyxim+GWy
2rVjLXmwaB/O0P8NXgZPhpVG7bFT+8ExskA8gHBu0k9HZRtDw6IpUkC5vy7lkRklgGy+GLmQa07H
DLU90KH5d9boSU6v/v+6VlVLJDdJdjEdKQ2utYTZ+TxW9h8UmbZfp4GtdyDqfy4Qdn0JAf5EWTUu
TU7EGGa8z+Ju1Exk2snztU5z+3ErRANbfABYD19Yen2o1pHUB1j0Q/+0ouxRhWvfrsLr2vFkJeQn
jYzyKGlI88LUOkxkf0RChy3sz6nr5mvW3/OYJ5DzRFXDwZbaw0W3wPybg2f/sbCdSE6Lg4R3Kd8M
9Wzakt0AwEBK7indjNFT9CYWPk036TLMrLyNscbB5ATyaaOaZAM3IRld4xL/MFGlCyV4+WAVj+E2
r6kGgDE313gYZPENOm2lj7rj1PXJmZf6dnk0uhy18pRO2AY6YX/0LKa1+UyJtwuhr2AjdJ19FkbP
tjxhFB1c9/cTFZRob53W1DyZbx/2tzl9YSZgM579ZjtADIX03w/G7HsDZJSu66hou8f8UDEwNdeI
Csa0hv7LvUQC6clkwGi8ar0C5BGfeH7qHnpKGme/a8VKTjlrYH/0TkpWgHBZOQPnCapQ0dmph1ve
4Lc/mkpeykXYgBKA4Fhw8/w4mwJM1WVbx3EUUWkHeZQPIngcCUPTW3IwA4j5jSfaVzpacGeD951Q
Zafk2USzzitS7a1YiG1Bg6MtJCTzWxo+teHATDtd8WZ96+IF/H6IKe3HU8KXOJwOPTunLbPFdcGc
lyrfo24DbbtxYZC9Ltuc5hBOLbOSwcQqaxxcssIgu7F61i4wJ8J1Hl4Lk8nNk1dBM4JzJyHAgAgO
DwmoUbsTK6vJeWtbVAY3GYRY7E73qKfoOYjZx75ibUAY/9MZxlr5bB9h4d0kohiTFPBEDVQxqiTq
V04Tcx9fg+SeNfLQegR/k9xdtoEhS5W7pNTjdSa8surF2kxG9yfwFgf6CvxfFp6ptu8qOseJ0E8M
KD9JcbTJvzewhKv4p1etRhh1DeaQSVr7TGYdZs5d89lu+7eOyJFbpKSfXpgVN1l9btaDM3Mqndzl
2El+mx5Sv5s01AQMOAuC3GBvg7ByMghdtXBhtTUDikJT3ZD+ZwLmORbpzrq4sZ1W+d2gEIbDvmXN
UUWHyvy4VqWngSWpWZ01y+fB+Bbe2p+1ar53Q2tD0NKNv7TOoSgBSDkLVY2CHSoK5LbJq7u3R9zO
1US6Jrtwdm/XYAxWpay2rOj0fC+ISTWYtzgcQEeEcaN4OrqQzTP5+5gXR0MmtzFThOy2cErOKJzm
DItbxWlGs3kbuxCxztXUoKAb9BuypidSN9R654XzlpX97j/3N9qw2WfIn8SqrZIm5bIsbIBnz1zb
QJA9YonuQAgS0oOjNkDfiYqAJPtdsccw/X27BgPMwRVSYy4Z7RX645R9Gywc0EJQz1Gg4eVScwev
LSdg8xyQ+xGjI34iqxS0yKlZVDc3sUvgT/CIf+Fbr+tJt7ZDHWPWI9YQRlny5IxS09KGeJf2N42x
JU092R9hjbKQV9xj3YsCk+zZQGMjNEnXVbA7Gm7axW5Pvmy5YT7xn0BTS/Fy0OtKFSrdk9lS8ijE
0LDLQN1iN6xftO/tUJb0SuASaZZN9qr7eyyV03/K8y6h8nr0xZQINEVV5xPHdH/sOKOvDBZd37FD
Mj66XfbNMwlHERgPQfIN9dHxtFh12HvDsY/McC+hpbceHe4aBKpcvNB/VdiLG5dzMHhdrJKGWznm
BH04TtmJblZ27cWsrz6tbq/pf7J5wfLrQzmarxw3Ek+zkikJ81tft70vb4PpQak0d51pd9nrBdyM
4p1Cn5Qj3JrvVIuVAU1sVLYS1j8mqDBptD0lFVw2fqovp5QmSDXTtQvD64mJ2zIeIzWuE1WE+i9E
Hqh3ey2gpcKkW23GiK2oSG/8ubeacETFYustrq68lh70yGEjpHsZOp+Kbcrp3t2ur2cuvvx92tVw
kd6zVT8orzWu02oA739xJmPshbpTjXC0xqgl+IqaAo8AoZ5evLCXvpyJK07sr/xAKPlAScx74gG2
Ib2So3BGps/p12tTIQt7UrqSRl5Tyh1V5ZwTOsnR+RBST2p9AAzADcdn4oKCgwGrL125JG4g0Tud
0CL6ofNSJT5nxwRwrJusMtg/0wE9asfnj+TFyieRmavMJ6TNohUvaVqlLM0Z/cbQSKrxwupkaV01
iHleA66JslDDu+zhaAFkx/Op1TiZy97mk0cJ1/ikjtna5KD+qLI5gagtOSPkKou05MEwKBIuaTcs
oNS8BqF2xodtHonEO9Iger6SljWWl5/763454EkIa+l4jO1yx4Bvmap9Frisic3dNIor5mekYXWI
F6q2FVMBIj6sZDtmPEsz1h8Zu5jHu52XRuCpWlsPHN4574pZP7DfyiOYYAcUAZb7xoy3QmjX2jSu
3QB5toPSUiSjW+eG1gdESfoRDyb2Q+c/RSirEQrxQKLNHtryZaYAkacsQA/nLdOT/8BL5wYxQ7jw
/nql4zaevonWdHQYkijvhUtDExnT+wGseY8JgXDZZ+HMROWeD5fpVEi1ExghfG9zavoHGhIRjHP+
GojY+BxuVgE9y4YUlfsfyPCCGznLXYtIQ/5VdtvFYYe8x6Q9r/2s6arAOgYnI7W3TbK5OMJRQpik
JC5AvHDdt6r7zArB46qCLuFQeYUQLoxV3NCriz69Hz3Phemcmx7RhdodBytNY0AgaCEJoG1T5o3G
mAwL3mls6yNbf4XAwB0A5QJQw0UcoEIUw2O7tlTeRgCnk0bdfwO7B13k7vQipXL3DnCUIvY5j9DH
8wY/LpBd9eilYDkfsJ9fMeGtlJJyEeUkp6NxExr8m5yMr3th10WEmc3PAglC0hioBLDOVd5az5vh
zWXcAwn5OYIbHjSij5eL2eNQePasAF8v/EqQiFBFXTZ/AXfJ85scxFe7/v5S+9fdkmVKaQSvAubD
1N+MXc4ItzELTf7ICa5wRTPKd0VaQi+6ZZqTOhkKsHLTMKwAtdR9cwu8nfL1AO84e22YOu8oW1UI
jPiX99nouMWZA/SZrNp9adFwtGEPleJZStpM14h9U96PQP35HUnpDl0ejSS0iexpOCclEv5JBtqQ
YLu3Lb63UG+2B4/QpmIfvFY7c+lKM2yeX+oW33LG39bzM782Ivhzp0Lj3xsyZCrygnaY4mtk11f8
A1XEFAvouKw5ZWNLcFc/I8mMqu76ItDu1fP1iPKqOIl0Ew8aXr6bNwc9MELMa0rYY+xRdvIcYZwD
9FZDB4cuJifsIh1TpEPNb073YA3RoHyT/xJ9MiQ6Q+Qfke+9LwkIAy6NcSbKaaeuk+IEK/tbWg1C
p1WlhF+JCf5fEitCscVjjlLKJTjyt1FnW6AT8tNHH4VcofJl/jtcQKHPw3CMLCLMCcIbZzb37swf
fhYRPIeLmm9CctJQZLrwUh372PTBuhQS2Klwl11B1s6k97MQWdwxRS7MUoqrJt3Jisc0fYCp9GO3
5hNFvA4+ZkTsxIr8HrD4swdPFu9TZnb5OEd1LERdSsdJFxl4Isr99I/0PZePu2kXvVeRROyKNn4P
l4KX360HHBlOpUJJh0J05f8CDxos0LKk3vYeue/gWtAfyCXGDf7AwbrsltbCCNASYdEBS3/Cwow9
wvzPlEuAWN28RPFSYvAZYWoaSLT0rJjM/KpAmjeMZbUn3yrRAFbfW3neiARiF7sLoUcawtMbxi7b
0XDeSOnwk0gEAtg6Vt6Mn7lb6BhY8fyrsb+JkLTYlTwAs9SkCV4S10uV19otMvD3jNj+wBts2Fom
Frh4Y8wO142MEC0u8aK2Tqr60A/ClZkmHBxu9bo9+VfKdVn6+8ybshj6UCdqtCfA1Niz43u0vN3q
1RGUHzb97QCCeW3dqyZ92c9hVBZ0wJXussDuC1IeI+PYD9WrLLKf6eoNBgUm2DG4NQlng3vr4qKO
xVC51AP9/zX47oEFNGX3Fn9h8hYI7BTQsPZug4E7muMifA08ij/Lc+XmCN+phdk70h+ZlI59ITR6
DSyyR6k7pYRJB9ctU5PxEBwARZi3SabOl4B6tIByGlCeahH9NQac5bqL7UIC7FpX5Mt2tPaGhx3L
WKNmk6dZ1bvna0XpuArsbCnu8rGy9BH3neRtNTAAtH5WtNRbd3UrMpUB9L9fDoZiPXOxbf4Li2ha
QQPvHD4VS7lpzKAoOnQEit21TiWv5LxBHAX3smFS+zu4p4K/eGMHVRCI46QotW70BCx5ziE6v7QL
LyV5jHNbzpaXC1wt5aQiJVoJ4DSE+zsu58XWwZh54UEqVpNFEtnOXsOvncs+d0hJvI+Q7azQhvG7
Pmgal5wEIsyzmmkfYn2q5nJw8IEuEXvlqNEEg+ZgktdmaXVRbIteA5wseHtl13+HkU7PVoX5QwiD
DCm6SYj05OaCe2xdX5t6JIk16KdOhuLm3rhcMKy6APxl411/09FsjaNsfj3+dOrLbZv2tt7aa4m4
jSzuYnhKatpDiaabn77gflueO9dqgp+Y3kvV/LYhU1LxlnRdl5y1DKKrraDAgRcz3dEGW6VJ9VgY
WDzKVo+MMlzAvKj0fAoWpRrhhvHEc/pwsFcfZ2uTqixIzkax+XbW94nrTEVOvQ5mYeftbcnwv65x
YH3imO43FOn19Mpev3iKrFWiQc5/ohdGoine9RWWvy20qHUFW8IzlkVvHXxthlENyJXQcOwxm59D
wOI9e1eAmeyBnBn1Vhymoaou36ZJ6YYe87947/UctCtxo7dudxjAGZyObdHxP+KyHfHz1sKWMNwa
xKumnOA+Drnfi/nzrrRBChKlqAf3blFaLXD2Fs0/ZwHbFsvfhm2orwpRmE5q0jr6FCqNpzi32E5G
mJaRAFCpkClVFWWzjDM1JjBSgZK6zUf8WxnQy0S5I+XV+VMPAJ5l4a6Ga8NtpkP5+mv1u5NqrYLB
h8Ku7w6aPL9yBExg640rCGRRLnv1ARp8LpJEOR4ao/pVzwxco8gfzNvrOIpri6VdL1MBd9TjPzY2
EPMOWita9f4jQrJVKWNQ4cjvshaxseezabEwyP8pZvLkEBDuUcg3kUeDZx19YzGHx4tyBkm6Jppz
klzd6UiaLMSGjYumd/VcIw88O0iLe1incDotCTFiLsm4NgCREPlucZm/L6msAo+eN2uhsTX94ZY9
nhebWWaQHXktAPqwmT0LGaFY8ofFmsIFr/dGR1Vf5NWxpKG5gAFcfG359jEzwX3HZrJ5AnZiMTCQ
xsdbQnD0SdLs6vQU/1cha8Calol+wbzZMUUBEEUjuKBScvQn9k5XhhOf2ic2qSaaDACnMAZGd8pt
Ot4QCpX8TfkxssEflSfbcygMlBHoAmzOFQdi82btVM7pld+0ii5IM6vwwawJP41Jc3xAZptRW4nq
8uwTfQ2oOHG/SAETQVL9alXorY8In8C4GD8VifmIuIs+XplDiHiunez74WK3885sNX0Pvyw26I8R
u3/2CeYUcwEVTS34PJFLBO3sKNBCx7QfuattJbrVvPOK46fcvltSBPwYu2dLe99KASUhVoverjUS
yjRBWPcPk4Hxf6j+mTZz+xZ5RVh7p1Xc7C0K/tdsYhoKgFdBFMU4UX6W9gnteHOTUMhpxN8XKsrK
NUp0uK3Wmil1ngo6P2+RHwdqw9hcyM6KclvnOlEfjlkZQstX9BJ58xpPAXfPvicdBFdHg4mBN8zJ
pjE4hIqZ4M2ZhzEd316zl6ZL4RvIAViI7/UIrYlrGhyngAkIzBvym1TM99ojxVRDYkRkvZf81NoS
eF7Gea5hIxwu5qXLbhD6FApuQt4PUB/zps+qVSgrUfRK8o9LsdDZmV2IqGLyWWlPW6LgBGPwUhRm
4kvEEzVL0UihuA1PPrWH8DgoQZlngFX1iO127PzHvDJsb6vQDtRuKhlGCkWZ00UPUnhb5+ZWMcj2
L6YPuM57qseuzDHi+oJ8XkEUJND7o9mBJ51jR3+PRneiTU+fRVXWLSDHm1dAKnN1WUbh/iWy6eQp
82r+y/sWTazMsdp+r31zsCVG45K5nbjb0uZ2MyL7T3jK2A9FSu/mxSfE4GtkFsTbg1ybfQQY+ZRj
Dg3i3fvup+kJS/+LTyfjyGf+JHvOQcY487Y9Q9h6wt3pCiOIMjhuu52Skumo61bsTFf18dkk1yyC
hKYCl7uk98v5RT2Zv8pwQFfoRlQ6sZedcl1RODdCQutwxtrS7MZRoqj4HgFHzexWR0MuSH1mRZg5
UivFjPtOHAH+BH9pisYKBET4wbYC/8HVUECE1RQyBMYorjEmXwEtU2jgxZx5f3B0wTAEh7KVvrRF
EZz2CQLQmLC01EwU0bJtMUpleKXCq0aGeBscMDpDusGR+fhkZva0fAzt084sKYwOekHkonGJM4It
cldJMIVURrKPvoJIgVkfm/T9uvR7cpdta9mTqXGkP/teOsqtgCAYv0blq1rcBznoyNpZU3vo2eF2
9vS1FZiwDbo4ieFhfCE/8+b5ozGQQlGIVl+OZ2ZvVJ1leilH0362hbspChJy/h1NUyuiVSv6KYVj
QZtyHaC4RlZ2Rgo1DYVfjbnVabY9vsSHDIJfeJP+CLvgtFKl84BM4RkGkTEwhQ4PeZVbg5rBoAXZ
/dRQDyz19OJ/C3S7Vs+lM8ofRdN96WxizHllKl1hoACRHyZaMdF8nrxXWU1vTuKfIX0xEtoQ70VJ
EB4yCw4PxW2q6/gbDeTNdjMXoNf6+a+r8CymHi4l+NWrtfOo8h8wXGLG1D+sbqs8diVYqjF94oSw
9oIZI7YrAa5GxMaSYWnM4IUlk8CoTLACS8ASc7Mb5VriVyMVW5OCQT52kvvxqyixZwtqY+Zpfk9J
Q7Nnl6zXUJFdsmYmGxxPKfgdKtjcpThQ6v+3rVW6vN/Bg+e6mMexZPn3Sec8zPrSxLYazBjrTjR0
xWQJF1ScJO0ZSZErOLdgft9VxeuSJQilWOjTo2HF2PZ+uFdtUgv4GLUjtzYyTn7GP+6ZW4ITa1tc
Q2ZZaV461GFHPtVIa6ETiUNou2hUnCxrAYhsDx8o5O5k4C9p5mAJnf3RtJubtsqJNoX4+y4VqMft
vDm0QNxRA2LDHCmN99deUH3OAboEuLFYo/yGyCAT73FuGfanUIgAx3xEyOx+TvO8q/lDOU5SI4Qp
5GVXnVEH1ZOar/vAMtG7obdGvaTvo9CIzhQFQzXPRDtUSx1JNKfHtRnxdMjFgYdpvO2lKnQTrvkd
rQpTZ0SAMF/0AMIuyc38qVact4KEDP5Fv506Ht6TcXCMjQp+7rGN5+lZItQnrIZ4hG47cC/aLYwa
QFCNHyTdjeSgv+y0EuJarmaz5YxG+l2mQt8U4S881FSRTt3esy3NnuFfgRFzL5YtNdhutK0WS3Kr
QgIcIvDdeOd1xcTcyTjWxdAgVh4xiepzSSxe8KvTiUIWm1vnLJ8OpjVQbRBzAkngw8YfIhYcMrkT
EMWvggE2EJuFIS37ywAY+rFo/slysaPFYYVsLChVm3PFcDZ7N7ZA4CV0OA6ft4rF2GyxPlvlpXJe
pmI6dnUkJN0EofUXusfY2Y7Mmz4V8XWD4+k96i3giY6klh7qfyvPwReKKCvaVOvfbu1UN5LwoaBq
+vlLK9UHkphOhq17piKyIEZKAjqT+sznbXEmM1NIq86JZa2Az4QbCHKx3qOO++6oGICpn9y40Lbt
TbpsBEtaQ9kaRPawoTnyyZLG0CY+81Ol6cl625CxAZsgFQrAlP9TrSRIIxrpsPB74JXpdgJG1fNe
sedF2aMZ55MY60AEpZPYUyvSJlDcBrxxVMwcNrgh2F2LKGXObnNAeDq5Ufq8CYpV7cON3z6Xhw81
zItomWd54e8Bt/YFtwbFIrll1Xz8HTocjWVT1J/S8w4VUmX/Ii1MiNQQVY26W7kv4cTL0oEuMswh
2xwyo1xaqH5pIt6NEylbpTBbox/cztI7URpqGAbcyAQ976fmoVBpX76PszoWgCkRtmtvIUHAGSe5
8pO84B+ZCwggBYqI0IrEilO6q2EmL5gmysv0Zk2PTtOAtpL996+cEo3qssMG4q5F6v/Ww4plu/3b
CtDWIgnLW/2P3/DBCzU7ygqkUhsHFPNmKhroehBcsfXvnMk7RRgNgAWv5TAKvYHo/tMx6McHC2vg
cIrWE0j+G8LLZhKuwZU8XCJu9t45XLvpYIBUrAR+8NTB4xb329zWw1/0oTcjS5eCau2Yjz7x3q33
nBMo2hoRrKcCUbZvuDv890vL42n7JPjlWovwaViG/mONbxeMZWrwkJcv3CrTHm3uBYJrpW4FLzpp
WIKJaUFuu8W9KNWijdWXkMs16c/Ez/tTdLskGHIk4ikko2opi44pW83yq1QPYqChDAGJ7+EVObFh
1gGfZoVJGD1rTCfIfNvFfnnj1VD2qIIaQ6Q+KLQOJJWGqsbaLlQ9x0FjI7twU/5z97MurIbgqkA+
GSRIFQpCD5th5Z/a5Qh1gQ0aHLfXa6vFA1FFTdkPlrfTI+Atk/WVWAEcMRXyMbed29izL09SFh9G
N1p6IgLTlVWShIJvyD3PktzvsoQzjL7NnoCJKYMJEvOsv0z9MrCcTyyCMmaf32NSFNZ6C2uo40Iz
UIS9wVcCOWavQb9l1+5kD0EhJMyUBfszl76gwvykKg3RYW5LGf5gBYV21an7P3fESEFk8YeFu3/J
z67tsWKs6O3DizISk8H+xTxPC62Xs8zdZUPiT37kL2p8nJ+ymCj1Rrg51jY+EMo4wAaQQz+2TOKq
380r/xBrL/ASrn6YRW38h3BOOdtkkI/fO0MwyKYzF+AZsEoS1CAsu53D7S3bOrV/BgVoCpajzFkN
fdUq0pXKTTiFbB60klWzdFdyQlIbTgUoprqtNP435L8JXqM1yiATTepgva6JYaGQyMClAwM59zyv
Eg8OKEsk/lzJ1nnytoopijLUIsRirHP9ZMRYnVlbtSWCdYD4MPswizeNUbIHmcnbOCgiIlhoJ8Fz
2HJ2lkuUGqGDsjRawld2W+HaKl7iC+0J11aZwjjEAx4bhmkI6bAjejrj9v86Egvoq+8bOWKN9ahM
J4vQ5mLdWNSAMgDStiC9fmlLujmsUpBpk5LzJ9saxvfx7ay+t1aweSTsQdUgL9k2hECl2oyylxbO
CGC4m1sdzR8TZmGuDRIGYRrVuX6B/Kkoj52F/4JOLHleCaVbsw61UFyQzdFUFDFqP4StxiDX1Ym7
hwBh7zIaVult3tIkbUw9RgnvcNzswQD36iW7Kk5lGBjXQaoeJhw0GNBbzDsqkP6cjpdsvjn4H54c
QX+/9xX/+L36FvLiTpREHLueEwtjUFJchwiq/ak9FWznZs8DwoFXUXpYNAZ7nn0t0Y6wG7xjkAxE
+q69K0NetfsQjfjpAOSw2vtLBrTIZVDsGrsnMTkurkGOkMPcMCGYVFJw68DRM18Fe7tbkUrbBtN7
6Cp/2tFdfvK7QDvaEgrEGlIp8e3wIOB6F2fW/kzZMjIkBlFKJ6XlneGLXTfh4PbNFL0UzK0g68bN
HzG+S3jNZuun8pc6dpNnBLCcxzuEVhOCngc9YjxnYcBnZw8FlVZ3ucwQSMlnk3gIBfudOP7A9EoJ
oUnDdrBK/E+oZqrwaC8S9kP1cYZyRM/7FR3TFfD4KCA7KclYDsfbAhMeZDbx9EdMo01Br5VjDnES
UDLyUCU61M8ct/jFoH7aPoHb0XzWbc2xMYVDdvtjUqSOk6ZzqAGHXt419Om/zX3pOedNt4kl+AUd
Qee3I4jtWBevSTV3rF9cFWO8nTEzMF+N+0el9keEix+2b37wdfCJGYe2v8HXPlZm1/ZwZpXBEi/l
/jEq4pbKnaTkO198gpjZX4+FTLz/9nerKWbK8MhHNay+p6KMWROGZosNm41Kqvk4uC3Y89Ope6Hh
ROk9mMxyt2pzAKDJxqeVX9JKKjJLcdN+TXdsseJ3DVtJTvsa9O85vUKva7z9XYxoYV6xLm/DH1kx
MqU3rZTRK7yE/dL9dESri+3hIzTpLljY1LyUBGuGRlQarC4vRLKAQWSVQ7RAIfeRIx7Yw3cYjDUM
ys5J8SKOH+gaAdVmV/QnVnQnuOucnimsBpd5v1U+OOp34SzwEx+qZGgEQvzSGQ/z9brXBzfIk1WC
K/g+ypD1sgGDX3Q/m7N4u5/SW013rE5ZpYRzm7ZU86vQnWOMdPG1QfheI2gojQHExbNxIqamAOD8
EZ/BBXlQt6ZkKZiL29pC7CIXhpOC17I7bDLH9t2y5LJ++8+kVlxH9nGU+30obVfiIL1CHH0U095a
yHBuhzJP7m23dLqrzvHLXQMrxqsbg2jZAfl8xI46DM4b3u4yHKiNVknGpBq+6mfU3dWSkqz40WsI
V/xjPPn7ONa5mdbikDilfDfXd9WW8PgLPZyNlT/dF947QAp9qxSfBKJmgjDO0ep2sC0iUAV+ayv1
S+HFF4ac2SPmqKXavq7Zv7h0GyaeUJGXgKNyekjmPvWRdclSEpFXwQPmJnusNDE/LYb660211Irn
18Hycu89VsHK62O71bcF15oKkDrsl2zQvN+f/J3fLhCTn9GYjeBmc3Z/0av1LD32wzF4M6hTTGSr
EmW7Wx+ZC0TCljA72LJaZZsLZxKIwxbNF1rE/EQOEx3sIuxeiGxcCBHo7zXf12sa9ToSNpYlWlMS
yvlVr4bBThRiOR5AcsNwwn5oYqBU00T2RoWmelONsFhx9LbaADKOERF0rPhAjp3ejKQmr7sRF/X6
btUnzurE0nUZFin8qAQppSPAGce0OpuW3ll4OC9YmZcdCf+M5DEe77LxcPKbOwZ78g9MDW0tXe4Y
unu6Asxbchl+R3kxRHHqtCSxDalhltz77xA5xDKR5J2A8Wqv7l7SfYbmdzmV9WWYXWYfC0ahPYZ1
8VP+YAzn8SO9FXrDC3qSSVMzHOwwpcIpv10/K4vZwI445yIUmGqDxL2Nb41MVWWQ2yD/lw9PqLfO
naE7bbn/wMjRmmdfpGYIDjkLxWSCghZM20UkmD7Sjdtx9YAiIKN7HMqiV+iTtFnkNjAM4qrHpAOe
J0UaRiptT74DI8PS+RlpMoAdxep/mV1Kd574RzbZDVr3+sWoEvA1O9guiXxv0uCPOuB7Za/bWvKH
4/Rl4P341mhtPOb5bBVhNbVQ7gxrHDOxE6efH/YMLEz0T0f4d+S/c+eODJAeMDQvIAyF3oSB9HsW
RsdraY+F2nq/B2P76x9Aa2mwLYeyzr/wLAQd7WTiDhMwOC1+BAkrfRRhcbx1nJnU0qW2bM7F7uB7
NfjbtgQ5IFTGBnHXOCI+t7hlOcXhHk/gwyd0a2t/N5kX8GwJNEOkZMFWERuPgAYSPpxlOov62F1h
d/QK9Tftk0tVnm8P31ypu45lRptYKP4rSt6Y5rqIi+gwPl5zvfvDkPzTr4gLc89Wao+SyhldBSau
TChsaoemxef+iFKyrh/U0AeWFYdwIqeHC8XUkH+Xt9s4FzWh1g+Ve2Abpv/Aft3zoPfbsNYAJ/Hg
Av8tBPWXjAzqo+suq5VZsqeTJodvSa5u2t0MQ29rC6kL6xJl3LaiO0a1b6VIxohguK3Jn3Zbb7bE
51jqLOXHCr71r4U01eQxG7dt3JUR+/D3QhTqD4zVbFz0M+nW7QCMxw/FARFQFWFmgwq3JsIUDMRQ
ArbGVVc16/0N094Xmid3+r6WwYRchSUfnE+fN2naHg9v8cMY0sMhjnDzPpXx6WpDWNnsKUVTC4gd
PGeRHOdk1WtFW9uvZzNoeUMgGkPWFLLd4W37yoZdXO1HdwWuAGEw/mWYMeix47G+TDgg4cQyyp6x
/daSk4ThOkjlRs4KktMDRkA9/ZAcnINwEoz5Pu+iDA1Hm+/dF2xKc1pTYT8b53TmydalmiBynTIs
ScdNfApX/qMuJ8pcF/OIiVducwj6fY4PgVnR74CeZfcr85mcJbNC6NToIluXGP9SB9ug54JFF7Ph
vCr1niO+WCG7N6j15FweyOQJgJAG8SiRix6cQ2Cnf7wUWsxVuTrHGA4GhEdOKAoC+7DS79wYktOG
Fy4UINNfcdUurRN4e4KkVwzkp4Nl2lTEMmhS/TIBEBkT0TvuTBowqGUxMU0F5ZHgNE2J6M38BivI
HXZdtnyrHgiUvifxN/8Zh4A6Ch8plX7putlzX/sPGcHuikwmxiIoYVwl7Gd6kBDtB1IDCAgIe7wP
aKv9NqblqBsM4JyfmPTBPbpUaFyr84ZLGr/wt14QaVvDRCsqCsApaV1qdm1wzk4uYmw29vJqr3aN
eJDnY0VPRZGGjCOJS7D9HH7B3MIY7S+ltAWIW1VrCoCvEx1SKcTBirKjw5i93FXkhXQddgOlO/2m
Kg+7eNXvk6lRZU38yHJTy1fpi7RezbOJwu+4NGcRDL+uEOfzzvm0h4bGtU1JuLGfSzqiZ9FNnp8O
elOrTi9uPyP7epYRMboK4OIafGJAo/c0Z0Sqd+jjzMNkKRQNf/eaqzcIJA0f9zoxKhPttrt8Q1Wt
ZM3btmEnP6qgxMlo0yUJfqoZTbqXeTMSzGJ4/TTPoorZwdxHmZD1Ii2YQO6cUfxn1ijPvr7GFlsF
4eHu83c/7AP1exE3z4vybipoLZ3OoBPzZ5sIwL4uTU7Z+wsF8THNtU+tVgax6Xh/SX7zl7gw65OH
ssbWfY/In6LQrPGVlSkYXonxpPeH5ljHc6Bq2gCdZhypY4GM+k4FDSDBaao7XDyx4T/MViVLz9Ko
PbS9Dt/ndzp0pcn3SwBBSOlnZAuOGgweRDYSoH+H4USgwMSDc+VsRiAGpx8FTSdc+vvXseayq18l
H2Rpxh1DDW3Pv5PQvbDXyvKfDloxYma+Jdhc9C3tktopWV7MRA5PqLQGGlcVhEr6/hvstWSXhyen
u8/MhRXvptsCl0kg6/BM9n9CT2yNjXnvZ5sC3hkTjNpbpkJ7r7Bhk6JzBU7PepqNYehU0cf+Lr2m
P74BFC7zHqavnV/+/Aymk7vXPecJDu6LbWZJCViAN9vTY+x8R88B4pUG0TZgQJrZzci6KC/RIDU9
WBxkGtS4KPe7zYOtoAx6z38m2wr6nFy3EM1qb/JB5QMe72W0dm1BqfzXma4blTmnMv5qpqUMZhA3
bEhyxsZkp19scXiHwTsI5VVscFH4URO/1n0vYNn0BIzFDkGtF2pGQc2uAsZmJj91HP0KyfB2D5aB
KVY3rM2znjqcKJwSyrjmUh/jzXrsU1C89FfYAqhB75JoJmK45haW1zaw7tHxNWSHvJZEESNhyNFd
x8ScoABSAAWG+s/A8DRuvBKe3++A/QBTWpjkDkMaaCBR6YUdZ3J5PZ++AMSJvk3Os5+AuHhRnCju
p8akyvFck8vTz7dTpe3Psk0HReKUQUdBKb0mBiqiJ3akRINZFYIKap71e0k+ywRfCvqUaupuGLF2
eZfk2FV6Thl5aazOSg61xr58xhl5g+iJalshdXOr1QTfcavGIG3rX8Y67QrVayS/w6IWgnq0K+/D
2lvPcNziKCwzyRO4JNZ/ENLGfufos2jMBPihXxDQFdYfuKkCyiuzy7O5+hfPXw6sL9fdY12pNASM
UGrT8Sv0qrYwgHKfEZYEH1YGIUBcUFzF8nyxNEnTWz6XsIgU0yxNkQ1VxCVaXAsta8tnYCSLF+9/
bnznaJP9Q3sJ7HV5JhcJ25pw1vWNWyeEpAmCuskNZ48c7Qc+bk8y16OjcQD7OmY9g4hxbCQ64i/8
+kY93hdI9AlecNLZMn+BjVRypUDvWQFOBIuahusfTijMIbVxMSc+a9eOPKEpi4q/p/dBrM1CeyAv
1WEiTQUY5TbIsaELjIIBWBKU4B6FWLZx9l99bzR3bkNxog4Rn4uQOeBTUfwCdWizPwxhom6/gUiz
z20VU3lxlmjQ7fM9rQUIOLjpkV1vtgy4DkVhXdigWCvEVbY6JCB+uBq9rAaZ9r53ZQfgGJ95G4cf
aJa89CtvXpnp4SaXuk7y3el1nS2CClk718KUjE4bgP64z2HTKOJLPaIwuaBWpGsBtZET4pIHZI6D
g5Kb8yhs4mHqx+PP6GvxFGVw6roLcJBR8CWLcS3VlXn6zGkzZFZAx2srs1/sIVqM5IUouRKXNorK
6YxxX7t5H2DP68V2cZMCYYqjErlrV4f1a13hRLQMmz9Eo0wHZ3nqSL3S+0RgSUrUSmiuVRcKxeBC
POHJ3ar5DCvafYRxn+Mu+F/pQ+d3gxRxxfyqNpvAGd/ZspBED7PUHIGToBhDU01VduGReK8oIRXx
8U0pmjNg3wnGemyEmVpaPEylETbhptt611RJJqG+S366xPgcJiZBJsTlvsiQXTs0eZihpvp06kQI
aDp+jyjK6/AXYda5SHGuS/30a0uuCEbpZpTs0HXpjnmPpIg39Zv/8Eygocy4d2Na47Uj2qCcb7bY
/lKjJ37KXosHeB+gEej8QTeMi9AsnXz92iKwiNmG2Qn2jKUf2g9MXY8ZmMcGRk678u6iSS5NWAcU
euMZ7rDltf3YiNkzVWcAvSDBmH2zeNTe60TUT+wRaRu0ST64CSdquRWvvXLw0mGxxIDyFFo3HJEj
msVpUMxgTsfku66vVjFo03DlGodeJNMpjo1A2IRhtdZ3u0bbwaebY5ovO+jMEbayBONCO1KB3038
S/kjkaixUXqCIvRkh1Ei9LgsIiVGoTgVCkaTGkRbV+OwTCoKJqIldf40VStZ3E/wV9y19xKERH1d
0njP1sC36+soukiT0QmNoAyRSz0BB10MdVpH21XkjlJpFthQQI0TODN9qyf5mJA2K6SfZaAQI4Tr
xK1tVpzTAyWjiyG4tDfwPMNGhH/QXE0pgPrUDZqCeBXgYTKVFmaV5FJI72dpn5898rPEgftpbic8
qYM56U2roDZxXu+kcpO4wKCVbDIzvgKHDfTWP3MAmqpJaGtdfoFrGVrc6Y0w7QBz0RvvILUosHW0
Te9xNQ5ofLYGL4xEm1McORBwd4zaLUVB3SO9+kZLwkXzHGTalYG2cZEAt+uIVODPkB5XNORAigXb
8Hhi8RK5HbXqTYIzJp1ZlvVBjpKgoqM6mFUdZjV4b+kDKbvPvR47AfRZf+gcuZK5WePsbcdmdMsV
3ewHeNaNNf/zQ7Tv5hkcYBcZfplMiuJhIDleBYPqj2wqVv0st7ONI/mPa9Bg/3JrdugNIQRRWZwa
0M6aJezfU+xbhfNacWyqmGEdiEgMxY1yPiT+MxITnX1SC6oe8Q77bEM22eVTiDbT37BUq+o33aa0
31MNayvDXJwTiHgOupOfQxEnHsajFzsKvpaHMGTwSmSVjdcFsWLgzzCpQNlk8D1/EY42u7jddDkR
x2AAyrsKYuSJBdNlQAzAMcPFhcXICkOoyEvx3UBoKaT0BJlUVHPCQTNK46iEqEAkXdMG+pNq69DR
ouCMZLgGoJbORGPf5vATS9Ql+TWsYy0UnfGhFQ3vkuSKv4B3YPZU4qwFAALnAqfDYwo5QkHkRkWc
s1vNywVD0DeOBPRXeRSCW/MxmbAKotu/d+w2zsb+dnT5oCpMTSsj1+8l7yPCUuwLJqd1sUFRTMu9
A7yHKWl5GhidDSBNJpYPvc5TnhLRAQoKCHPlQdo2gcSfcWBqqwGrmeBTyQ+0pFDxzRjEZP9usHos
ii16rZj6aP4vHKg1qRCajwODdR4A68V595AKZzfGySYHKlruOy9s/t4I0VTMlGxunRygzLnys8A+
cjBiAaz9NXl64karfCBpl7s6GdUUYWEMmPcuybw+Y+7mPCXsWPEAFgwSgxOXqrnvlTWblZ2puoa7
FpJaI95QnVtvZVoOeQYp8MWEZFMNKsBHvUK5jUaCcJlGCZjvqmPq7FhF2GX2egKzgbsYYFn4CMuw
iIkFyppQzJdfj26hPCWHkoqwHIcWBvuDbAXYQWLr4rBNJugtA798vFfXmmw1EhYw7FzbNn1iC25b
v3AtyGAzdYcC0c6GkCq11ZQbGqxkF21CSw27nvJ/K7CCjyWHf4fWOgDk4Sm5+VnkUEMB2CikKXmF
WO0bCaEbgJ4XjYf1lKc1fGLsWMU8uhdHEVQLRY5Cp5wz+6fBKrn66f+WcVcc7psdA5yg6E/qVhK+
20RgErwQGm25ksQ47B2prBOWuE5M3v/Nn85JzyWIIiKh7oM16BlGcCLfkybrrVlugyak8KVDVp/i
/dRwspeSLXDFkTJ0BlvTcsdslO4gtMdoUZeeHByuuOWPM4cP1XLXH4W+lUbnU6CizZBUmgU6y7uF
0DXxCakhrRwUR7/82nY/y06kXpjRYLXw3ABYbV0KVBoxd+8Jgsa0ZIk6RG1Wu8CbidfAAYyL8prO
7EUOpCSrIOPeDO15C/VBRqcXZJE4I5AcQCTkmvjsYKsNGwkBYGaBlfXOnueYcwF7gNVRvMrnC4jx
vMMbm8ZYzMcv8iP5pMbGMpMx3JlHuMAPH94tpInx8AxZz78nDwWXyWVEyrMr1l7m5IGNRf/Ccltz
MyCGZX1YMVgvNDfspY5CVwc9QlmqOl+cugNve/CwlLilG5obubw28ylmQ8BBn326oeqJPRwMNy5r
aOb1fjWXx/WPALC95fG2FHtb4CEDIJDDk7i8kKw7r4LldNCgs6rS7zfS0PYGkyaSocKsJAPrEUHS
Ls3fo5z+SPCa1fLA/9jcGvk+UIy+LEL/yLRGf90LjE0ZcDyAmHERSLXdYYjZQ+EcUcozJcukc3Ns
o4Jl1Lyjywk6vnqfni+qTjCMvudOXMKHXY/qpLj8kBP/0OPECRJvLGSIVZUr1A9y4nmE89V0cNhu
DUBFwjIOrtGY+m71tn+0dZHKYoDrcnTekUeH4bozKfQvhuru6TfQMYPFM67rDgGd4OqrFyj9dpgo
U0X2KRPJPAsCyzhUGJyyEpUis/CuRdOpFjuTu92TkW2HsvGm3V5Kqg/Ph46T2N7At1UtLgUL8vwt
iVvz/XdCjcg9RhBYCdVpoX865foBr7tNijz+bm2gZKOBGdxKWKZY9PiuO8f5Av0rrTRJOZ91I/Mo
jaIVGWXYyY3GkmVUy9uAytJQKujhRDDbRYlIS8jre7mYtgcbB5p8XHHUwg0CBHHmTGQODyTX51x0
5yGEZgsUM34YO5nqEvVoq0fOybvEX0hxPYT+9t5XaHzYRmI2xEy5o939k7+v7NZLzfdMkFQJOKEE
lnv2iVoBGbydqvtjekF1GuK5qAzrGe00DDv/qsxyN8ptQLLqPhxzDaIsGX1BYjyMUDQR2mF9JCkb
C39JOdsdErpcmVTEqbHjevzIeWI982U5KTNNIgQbq4bd/uoOzNn5+Czu4vJPJ6JxxUrx1yeTONEK
8ZwQovVizRl9f+oKrTNi9XR3TI+RhMsI63yi4rXm+LfLFC0bRLa2DCpjtxJLBTWpRc51ys7Nbyyb
oQLkHwyDo5AoTO33od2EHWUmMLXRXJP2luHBxJUpIwupprB5QWCNUXQu9ZsBEmi2Vh1RwHs5ingG
Z8Mtfu3YGVgKwvE+rmMUTAxXmSrRQHYl6vhWeswTt6XuU9kkhJSav9rkhJ1dEv6kVAwPW2yJoWAI
gPbQyTT/TTLWPKTAo8de9MQVJh3/8xM9mMLQ4ztw2Kxe/3zhciuSJ4Y69oe4rLy2+7q/JADdVZqF
XUkivr3HqILkAroZjf1u+n2qyR/dHSjjfGpdF8hjlzX6JMjjZj7FwF/934tA5oThl+GKsJoexDyZ
69X+YUsiwg5dXlTEgGOW1VrSKAVIeOGGOfRH5Q8Ls0vd6EgA/7tXBcddFoQhgMv8VW3QENdtm/Hy
yCWFXicgGp3jIwLylhmkEzzeiu16xnw4yHAeGZJv0ZmbTl/XnH3ZrgSwjreLwqCpJARF8BlfeigD
NZQX2fjh+B6DIJ9VCY03DPH78JFnIKD5xNVKn2zPYNzC5ZGCPZR/lvWwhZ1RI8Js0T03ysxEPxX9
HhAcNr2m+LQ7yOOlhGWtR761GDrDxdHAwtmBALS8MrXTujQwgIRw0sx9VsUay3o6OxZtrnsSFuut
h7cigbfDg5Lleq2r4bukL/gThnqtzdwdv5Hr0uuasFBrN+ge1bNCLP4/sV96Xjvlc3FFnhH4CZ3+
TwJeJqnj7IJXZgVX0Y+sZwHFaSBTCF/mkfraOCrhqxBxrhe4mkZlScnChu75TjsEJDloF9N1vbGJ
8EnhgSRLcPgXheTvjNy311uHlW3CdsRL40LfaxJ43AS3XuFazSKsYD5NyP0D5cmSUjn1okwdNq/e
HgOE00eRnJ4uaKBWmu6P3NEKhIO//m6Y91gdo7xZWtITC+qo1ekScU2oc705GsTVN/q3chrcEIcG
ErRG6uY6+7vRz5f0p60KP8RTBqeDCOkYCSxIghFRVw0XVPw/vL9L5ZI9ez0ReGEXksaRrClYXUd4
90mMvvkH1N9ii3tE2/9zWzHKy2WhlNGMg/DeioXKFCCO4+ggU79G2T014UehXSew0qQnKCHpJPL1
xLaq9U5e+l8YpbmcpeZm+YmmBYjosWstAyIe6Q2GDd7DO7O0hJL8AiTG9zPGedbI+trKac+JvO1r
53Tip6/LIrLn46hAFf4UBgb5ERYtvjgWfjCd28hWwj6BL25r3DQ6hF8FZyT7m5Z5pDqo3fL6idaK
VgtBf+1hdTecn5MzQa/1kcDWwHYB9hql0bhi8rDt3STbh1S0GrzNxPwX82bc6yhXpjxvyXHmPw4G
9/Mc6CGzzGRNrTiVu1llq5v4P/B1yaS3xupdJjkKCBKReIwcSNnlMl1dSJjesrpNGjeZqPevIFJh
FFrYiHUO7AuTu/0IytU6G64OZS3ojRvtfki55uoECY3MftDE5dsFtvDPB7OqqmvORg95cj0Iff8g
PUH1000gqvmW1tmvxbnCteecjzEpAhmA4GWdAbLNTOX9IG2/b1dOUEN42leysgLwXVz2e0q2HB28
LCF+JN7YKZtAFdNOhEaYa2QSIGlvvqatPAsJbF9dqSH8mv21MMwF7ii5vgl2HDCEgwhyYluTB1c5
88UcrmKgprmMKKDTTTeD1XEeZ+D/+LJ9mLfqoi3eJ4OlJnQw9gsgUe5yRp95Nb919zzOWyWHfh0r
mYGJNtt7FLdhI5h28BMLPKX3Sxo8SZ7a5Y4Xob5bHYVPSJ+M7OCvQFeZ8LeOpoHi9kF295GQsoVV
68HWtwZJkGbgHcn6XZ3PssqiRl8lX01UCRizniQWft5y23zkNxSCl9LI23j8NVDQCpNDu3TKWMSG
VXCXnrAxvBQJcyYikGUS7IUk1ucZKqYoni2A96pF7u70CMxoja/6g5E9ZLqjHyg6LVR48kFa80aR
5RMY2ScniQE+iSz3Pz0icFzgArBHLBYzsI/uMxZtiQe6Z62tK8u0s65UqDlxNP/4Bsw57o2UUObF
2K0pZmK0sWEBQCw0WAV/HGowMGy1y8ARQ+RR8GvuFls0rtr9iIfjDPEjcUF4WrTyyo0pBzVXDqMV
UIh2b9dfGhgzCk/+KI0NE6z2GZIAcTQbGvJsp2eoWx35qw3PXmJ2rsfGTFG6BqRzFu2zl75bQb6v
jjDshMSPSp2Kg/8p3Znd4PEcNGF6gihrKJzE10+k9KWgYzHxRWuoo6DWs2iV6yftaSbPfBoqg5Xo
OR0SscOVcixaEayO5Y4qs3KN8Vaom7B73DlfgwifneAn3C8SYBEVnYnmPk2qBSacHhsocD0zynD0
ZLhEfYN8YidLs04Bi9YB2TNbNLdeRWPIU/ds103aNVQI+l+jA8rD2h0qAfxvE0qua+oUATOK9MYg
bxH0j4GS7JoOXm1LKhmalbBrlkqXYRUrBiieLbYwgwT87ubuzYwF74tS5moZzucKxZizaWpnVERN
++qeY0BmztE+/GosoHJzEN4mpR9h8kAD0ntIeNOfWlP2yy3xjO9Wmhy4pZkb5GAhRxemfQ31vDCy
FW41E0oEXIxCvjGRYed3Gf/s+lhRlGQlwVvST01TrdIskKfEsMsHM5tLby6OErZbozBiQNq82iJZ
7FqxA9iMqYVbUMlex+32jEkWEPw413VMZvO2sHfaTaqds6IXDsWO4hexQoYvk0aIn9JriC8u2IOr
2cbkfJ5vG7+uAjZ2jgKirmgT49QwHG2CLrHBuIgDXLBqkqHr8p4optQSKG+zVqiAQyjRrFxdjPFM
tCH292fs/JT4oDIO2KgTXF/DpLoKch/3pXVECFuBZjwM1eGutNEIjQt1N+x/FLlzoa/RLubqPLO8
4d4XXpC28pJhL6mKG3B2INwl4WG3bgwsG5QwK9nboXrk/S+x2tfyUXHZTpRGH2LXsWegKvIcf3EY
wHMHXHcsMncnN5mgqmWUh9Jg161Ck+ONMisE2Pz6+iTVqqwuF/sYHIPurwZ8FafK3lOjKmXRjZEb
QuFbzQXrlgEmKdokK3YPY9hLoiDu7D1qV28Sscbj39cTneFfVmRfjAsBBhh+qzZ4e1pf+I2BaE8w
3O+cK8JgTxKBSbCe5V6h0yCzo3QvUU+ocuBjcgBRK39DHj+W2W2GftzDq8DOtp/L1CSkL/IoL0SA
SRTC860qMsHqVSMKBsEyrnWC8GxpPAWkQjs892HbrKvy1MQgrjKYjNie+ylNYlDzRm+o60PKALg1
GGlMWdzyXcWHSDs/s9Aj4Q5ixODIVw1da8rIWDB+C6Hnrtt7+Y2id+iK/Pd4TRspzMAVN9GGu/Cn
hacUReTZAxUq6aXomyDegnO/a8ZtRMcJXr3FDkeJSJ2cDr3ed5fqpsec3LTl+JZj24IGVGYajvA6
D8oPqAIFtLAsOqTTTyTiM+xWC0T9wKs5SjrVXinxQOaSB2iPL1Xo0+5/tdKJ0hfVuq+3lPG3X4jj
FAD1a0ALlbSSyh9qFfbPkCpA9mzywXrTMCSTMn2uuq5wKdelLSI2tVniWNCv5XYDQhk4RSROSjWK
pUFAhjx73erImM0BHbODYPRWhiz3yZqzWnD2koj28ZYbGm6O5r3/hYstKvB0K0k6U6VeHik4Mj7r
0ninUbGz0XCSB8vjAnChECKNmYFePD99swPx5PegLdWYWoX9e+ClnWoJVZhmo8ssP5WXm1W/u5DC
EmlnIkIfpX0ih78arLbB5dYcqW38T0uGHWmrxS24RETgfcnbRcLBz7uJjeRkGUS2S1mZmdI1CGaE
//NzfwjlumPC0UsjltJsfYy36jUCpteWxVWHGFm4UMqh2nAS0hjbKKWbg/ZVtMan6yj+lxR/zOQw
DOb5ERssXw0l+90tO9jmkrX3RhAc2c5yqWVtNiblFXPh/reurBWIvG66XHOTqPE2c6tZiM8UmKO8
Qga7PPLsZn/hy+YQIAEiyOxQSxFZ/AeERy77tjk/0vCz/yixtnfp17YCDhk6uOJxueYml1nP6Noh
XFXugLlFuBeFpUxPNWcnVghuUEQ0fNeLZ5qQJM/1e66njr73VnDpbX1Is6yjcuCXKW7i9kgnnun+
hYVK2xxdZ2r5JGhc+X1tlYrQ80LU9kCe1hWgxZNAKWMMlfd274lZw9GOxWA2gs+3UJLuwDzSWhVt
L9g3aQ4ZU1S0uCUaCbRCisFweqXx4Ngpxgb2HCCv3kZiQlTK+fsaN0Uzq1tGNQ7zaiyFqvZoiWz4
JprhQm/zazoVvE+wegxC7oi/6KIwxyPa3jKiQnpApf2iyYewEug7b+n6HXlrFUtXYQtYXel0klnE
b9M4+SmgWEqyYhKbKQzBfHuY1UQixzQhVmkBVppLNHgp01va/kaYxrZfQn9iIcyeEDJmdldBCWyb
ZfoR6joX6wPzHjG6D5XCz6x8hXVQBisd+zKhT6iIbBdskAzw4zl7BWRp7zkzoS2uFOnFyfrjxleG
ynkYqYuidEVSAmTwu78p4SjNdYTiyjcsFP/AmPbY03pwou+I/35WahKRzkW+LkL4Q8y0i34Q1yA9
MXHjL9FwVbsIRS4wS6qMwOY4QSdq6/n3aEwzbuWS9UWEwPNTbrjBANuOeVheLbI6ze8s0xXc7AkN
eRRPhlTe/omZG8wExT7ZQUqVhvlWZYYrJUOoF7GktcG8iuoQmhNgRoOkftEXfBiZxai9UPikfHim
gY8+6AaF6zMrdk4es04z6h9fp19HCtJzJ6TlGl/91fXBeqYD3nYo2nfse9u/0TXpHfaWnV3drtRh
yV5RblTenoWbev3wOIs2ysA84Am4GW/2SHorB/Ulim/mcFGcFERoF1AD4hmjvgL7JB07j38eVH14
vL6jn1Lm8kfycyEebwR8X33TLuRSlZgEPy7z3Kaohk0kFgfBCtXA5x2TByehOC5r39vzIZChBcLa
xxBt0VfNGkF/iwTyIKQRl0QUjZh7LgFsCZ86iDvCZV5jGCqmYG5ro5Y+jH1S1KNcV4Zw6pnVbZhb
+WQPn0VWyk+DLCFxlGiRK1gIGk2n7c6i+xznIed2TYiMTNMltO665rl65Z8uDazn8rMn3XD/oD+x
qLCfZcyE6zncP0s51/+ph9o04qPw9aX6t+1/0WXFPwMvZHNUjWD3q5I6w3W374KRurds7CM8I2kM
HqPiWmIbT0QhD/63N/5CQGm04KGBzW/anXGeCwkiU5gcys+lY7ynUDuAubvyqVlth8zc90LT+Vtp
OoZiA4w2wOe90WK7aXY6/PS7BBBGDcmLY+jRwRK2rzizuFg7AfwCuhY33s4Z/RAVIHFOUHy6Hqcq
iRcQ04XGxvnsYulOKsn/crdABwl5WekByouG6KeMP2mJ1Wtsdc+RQW/cgW6f/poMJQuQOGzqS5Pg
3NpRsBrqgyvck1eLD85Jw12qjbACcVbM5g215Ilawjm3Zt2jkra1lNERm/jYfwv1PZJft9Dkcx3C
/g+K/jWWXt+RrqMgKkVlXwYrDk4ePjQKK3pE3HvyeRQfBoY1obTxFBpLICM0m/qMPFFU5qRgz4Bc
jWRI8Kd2XeHaJO9NWzuN4Kf6xaG3vG8ZjMf+ovW9DCS8Xr88u76v2k4L3csDmGWYwRGcHESxZmJN
loCgA37d86tDyWcPbY0KTxHlaULn96puU/u3k6GDjWn/XE+CD/tZ92AiIivLabQhtaJwzB/9vYxs
wJqHqzT4YyuJLUtOW8gD9fkhheHq+yw0VVTrJzVPrwIPgDzQNolMy3+Kqf6Qi7AW3V3ciK/Z1ra2
4jzA2LVmBVFw11n0s3UvSG/J/a5H9D+5ynxjrEkHh71vadKPdLhX5a7wqS5UX3K+xS+GLzhA/GYy
AZ4ctvjPKC6bc/jNeRQZpAvFV1/7OWiEbWB36UhSfFP817liPzNw5Czb77j3mG5JbZkrYy1BDlDj
oCQJnB/hpj2WPLQr87t70e/+tvsqT2gIjG9haivJsNqZG4u6Njxkeo9CZMjGbbUuoSXfkKTkvU1X
n+CvuRhLbt1nV7dbwr6XwSePAeQm/fUi8xVZuRYfW5Hzdtu5LLLmbyaUNfMPDC1wyE916iaBhmcv
kiOd0yAr/QjlTirm9MYLpqXT2IGRdl0dcngp9hogl7wAPkw8oQyVbxHnsMJ2nvzazo0mpqePhe6t
8JR6JboM+HCdMHZn/wUf7IbWu164dealx7kPqQnHTcoOHh0M8wSIU4gtd3FqMqCCH+qwC4iim8A5
uOhMmtYQ+V7EA+pViD1WhGvWdix/+31oeEWshzip/aMxp6795BnAflCZ8kdQ9hXkQM90YjXcTy52
Tkx7itqbO0AN6QcETeRgPS2e8fb2FVKA7ZBc3JvuB5p5Xyp0tkwethVqkkofBy50hh1gPBppFrox
rMdDE2J3J8C6UxiB0XfXw8z9Eb2LtyWHISCBgy3gDP1YauLrK0Cc0XaUvOQRZ0/+4G8HbZppqVUO
9HrwD/AcJBe47a5jGC6KPjySGuHKxK+BilM0dpV6jH/5HH+40GB8Qcx2cvl+2TV+LeBu0wURBvjQ
gaqNF0MGT4iHuVanPrnLgo+e3ru0aNnIvCKFty1A5Rinjq9CKplTAWIHMMEmymh4mFmCjrUL0tlp
DzkUN4EVtYPBnK6Ff/AuyDigGf4g2GCyknpC980tEnqQQtH4cX1eJgTMiI8NcsdHseUkj1QrKmpT
GD9G+AEIdW4NtqmxW2lgZCLDjQn5SsXUR3opZJoXVdEO66DxVkJrRcpbstqcwpPGKmoPv8plK+ru
4WKfNYetA51izsHYrk9kV88k4wcgcZU8TMP3Ln3hlAXzRBCeCrPUGMk38KXRjak/oigGOkIcZndX
aF7FfR1YRN7veKK8iX8S6usty4UpNgtCW3R1fYllzKBj3+tbAHIkh7xqaGKqmgh4dxKN9LSCJbi+
hHcw80u9AakPUihtEWNgNBvrGxecZaUE4TZ/PJT+6txsFTUmsF1omvt7n8o2hiyruWkbsYVwcN1w
cSZrshSuVVxp1jbkBgczX8dW8kzugMzqVpn4NdCwvn58gQ6GCRfq4ghER57SjO465HKmST1dYIPh
IA85kvkMvQmgOFd/p+7K/pHNnVgcfpl3nbMBbm+FjFgjccf4L7+dxN3wyK4JXZU6uoR4xuI+ZyeR
BKugg+BHLW44OE4uT3JKzxDQWWoTLhScGogiPNice4DRzRfGCPyfkHil2jQTAjCARvlCtQgqi6Ij
7sAfYlnb1lI9+HG17RFJ6zjISBAZny5M+wbdSRwYgFTFN4gIytuZT8YckotCyTp2Bu1gl8Ia9d4o
zS6mflBGKl4ofoxr4AXUdjke5QuHWTltTf6elZ+dA2pE1GOK9uj7N/77/MApG3I0vrHdYD5ubvBU
RO/aSFbmJiEg50uzzdICj8WoB6rxLK1a+KY6QYdeo3AUM5sDMCo5T16++E5O1vNUCh8VF5bLflwl
WU4/9Wvh582K67ZREXx9OSabTOZbSZp/QB0T4iaATI6lKeRtQSiIZKVMfNiibaP0H3iGZroNadKk
Z/4h1tzjX+BsyFEStQGMbHVDhDUyAKhaAk/sS2mqzpgsKCsZTdJPzkosInYIPJ8ZTx39jgcRCoJX
2P8tGwFt/FdcvWzmGb+QyeHtYxeq6r+tRVbXO8+h3QWTpZPm5SLmd2mvKzwUB7/H9oAJKWd1kDJn
13u2uq626RYLKixr51j6ze0ZzLSSNl+lQ01asBChc55/2bQUsktvMWkXpw05fsdDfpS3w5PZIsFy
wcfi70V7GMG4BQ+VwIkKtgx/40eHetzDu+jjOHV4egh9LZ6hthXC8SBYRAjgNnlHw2RaGuswwYDw
F5pRi2ggeVicxT15zuBmv/e+YzBaI89QrqlQ72PUs+dF41U/mMp2mcwlg7p/LWlg9L65xgUX7Isu
flVjm1+4Nn6KkqAazrLh0WHoUIRo4x7ZdnM3YJvRf4oEh+7ucqOvMD4gMPxr57aEOaNjOSLCvJbR
rxTSmC0qcj+zsp2eB/msd40o5eQ+WRsNrouAVWOGGdRcbXMZIsVriGLjLnRosFzR9bNlC3rVO3MN
qp0sUtj8o0wA+mTmsn7pjZ82HqgbJzS8KmCdlDH2SJnSdA56cVD42nSpCcXVi8F/8VDRxYUJkRSb
lAB1ejHvXw4oYyvRlOlEypommYr5H5h1cXLJH1xqawpU0TQ+7XIjtMre013GxIdG9Aj5FCpmuOd9
/cnd/FMC+J8oL3xsv49BTOq35gFVl8ZIi2WHDTCf2LACtvA9W/cpV5ocR6jBdinePlEb1/BgyI1O
LGh3U+vfAa/vtTjlQZH+yDSejjzFhVHvy4SEqS2AQoV4Gd00RNEWZ1YzKA7Y8FNG787xdnGChYWD
sqkwHEdVC5tprPdyRjRQHPBdsy237IPtG1y7KuqwMeq85OQ6gldQp3XCtVGamXcaOQSqj8qd2MC7
15/czLdrVWVmI+W++4bf8CONLOrPuguhS6fKbnQ+ScM/nBtR7mdRItgKJ+HRI6lw/6VOhHAsf83S
JPVNpkL7XzMvVB02Yqc41r2hHjhFlxcW+BrKyPH9VcThrQm+3owaps+J12D1Q8sjHvk6Xk4RqUSu
pZ4D77BXeFc8XiLySl10x8En8xserRwMDlBIBLwLVTVIUKlbW40qWpe0/kTs/94SE1vmjEybYIZ9
Iejfdqgf6LcTQFM6la7FGH5crM6GY2wuxnxNAIMpGkfKAkWaTodNZaDEjOMeXIJCF/gDd1XgHJ2k
RIeGI3S2MOHI7YC5b8fWCupNjSbVmugNXgJLc4N3KGH6LMl1Poy84MZToCnW5AaQsyStm9lU8QFY
eNPBXmvqbUrQZKMj16PMsEW5jRty9EhviUPjGwwUKLyzHRS0zPqZkSLhuhvKJ99b7CZnRgQYnPOJ
Fwv3jbCQGAqmfGO2f+z9PIEKQC2Z6Q4oPtCt5Dz/9+YInvR3+2TGgruAM8f7t+bOAORBUt/eTXqn
komPKhBA18KU5Mrz3vEMP1jL6TszPLt07um1EqR74u9eBR3wKmlxxdi4s5N2b1p9f7THOPa8q2sS
asLTiE7rEaKozCn+RTHbh9w3VD6jiPTxuIZGVsKhlcMBXQOP7Ism80j3YW6kFkWJRgyiHKAagmm2
pX4V3J3da2Z1pyD2awGBqln1U3cJu0uZ95Zipo90q1SUiUBHSdDuNh8E8DYUorH6rfa3bd5JrOfQ
l9O2ms/S+nmT/ZoP2nXuLJ4u+PmWpo/Lf+hRnZmywitXF3tt9LmlB3nuQpFQZ0au8wJvKwdXnx5R
WgH6mseCoMLT7NwNKnRFHnxPXVkWsGMRuN7Sd1qKpFmX3TqMaOKBFrjbr+Cj8OCvTGsAqaGJxR3C
wVlgt+0Tv6LEml9e9+LHr4GqqLBUpoEk+uXXRbIJipJ3cTYASQtD3c5m0WQSpjJJgbBl72VS3FrC
qu+XOayhdUPg78S/Jjbim+71KiALX1EN1gqoP0ihB4XRIjQrfsO11pBR/SxHh++FNSWlG9F7S2aZ
sebxcZAE8We9pCI6nPHj5Ushhq3NH4gY7355xAyhS7jgIJpvz8tK8yGmfU3cgFAzu8CX1j6/Tqtn
NpNXQAch9PFut7h8Uuw3ZPcKrEWRxWvfQgMDIPpBG8tBAm/1jNIvsJMVfkOwWer5OBSsiLL0KKOh
wBTmDT0ixiE2qcNjWeXGXh3OzSSCQ0rpc5UA6/6Tx5f89aNVJNyBDkwFI9hjSJZYbnP9BRFX9seg
BltEOHgE2XOlw8GWKjpCKZ6PLWXpndJ2Mb+SY1mkRmdA0XJMDPsaZbmyMYpGrQqytnqpyUdg9G0o
ZbTbxVQdEk5Mxu25AKhfS3egoRiDCAd3JeTPDb1SyV0YE+qWRwm7HZQ1eddmifXa30IIau+Z7UyO
fKOVtWFBd8hsa+4kRNRL/X0s5E2DvHbipLoA9bMAJsBesmN4uB5thyv8BN2hJcuYRHdYYgh4b9CG
2SMJOs9Q8At/uYAmfWSyH08cKNogQFEjgH2HVeMqIvjVNzbYkDX/xWy4R5xWOrRJSP1OMgPAokrm
7dtMQw7cDnO8Ctfxd5o9qwvlweFb5sSyKxg1Y1WxLflR9siTA6x8A5LVlkcLUXgY+520FDBoiOU7
x5pQo4MnBdWVq5zs+ru0hq4zpPsql4DbDWbadq+ztanMRlZlgdeJRJlLHIumk9SCnJC/eM7uReBT
mS4tQyofppoGqsHZTtmT+UkAMS8Kpn0HgVwtkXKW7DMjKC/jaHfdLepJNQXkyN+J/uGZN+SmUHub
Jfa9FYb1iFfrSOB6pdocchaOiN8aobdISvcYAmlpBpzmAiOv1biG9nrrCWWa2b1TsGRoG2Lx47rw
swwehmlH3HWMDeOxYqvjwUZEy8RblEUmD0NvHVmA82Ng1q4NVEEgZqorXlNmZkfkPy6bUM5RJfpb
POQH9djgTYt9ad4OgpsBjoIC9ZsYBCaC/81Je2UaasMDCBvBiM1Jthi5ESA8sG67xfoHKoTnX853
4BxsDHYdiUn8zd1hAEbX8PreJyHHRwLcrqEK3oRjuVzBkLoeXTfI5vOyBlNB2QWOFnPFsXnD3g+f
U3b/VgVAYL1xUeZlGHDjLchWMFtFVmDLjp7DsA6Bx4pfpbc1bb6HesF15VSHCaFG5vNfeElyOSOH
V0fHMQDRxlhTkO28RGQKLS6m03gF6EKDmS7WPMWsB29Lp1HqngOWh7hY+FKHguhsRi9rtwuAZ0it
gErT1VkuvbfPuV6aW4VY7XRVo2wyzra1FxjZmC82o9sfRnm2Tjqzf4tgQ+2cOANto+mmzKq522Z9
NdWdw7tYIzPtoXepzZ7R1WJFB7OTSmzyh1Um2Dw2ElmRN3RYyebyVsaTe7kT5dUuM5YW80/zqsy4
x9xDh3DPdCQshieS2x32IqMhRb61GzZlp2mCb6kl3zTt46byRtL571XI7T9YkmGledUL+cr/9MPb
wtxZ7XYf1NzKT1FeEtt9x1qmRMevKJwPXVWSKUFVbbtGG30KYoTQpTTXO8+xaXFT80A9aXg/Q8fB
K0mur6BAK6trycskdo3VJydyIbAYSBC4MAsvSWrwvU09TN12RqYq13sX6bz/nA3PXQmSXemq3iwJ
1v7AGbTHWqROc82E08/o3mRfQrzoeSjxxeVeCRKqnUohFP2MGp7a634lyW5J+V80oelO1aBe6jvb
LuMCXePB1LTAkR8Qy1F7qrqW7qgaOj5cv6gqv483SNy2oZd7niJn2Eoxw7LilxZzLXWhDQsXGKR7
kjIhWpdqi06Sn6RtuAm9OY8eFCra9M7Y/g684CDodTnD8cPD3nsjpKIT3kARgt6jsVA7rHNhxMbE
DXp1ohEozpSFElwC1vI1AMNQ2X1it+7ZnLi93lKBb2gXo9Bzm1rl1cYDrdmEpvkumxrSMdo0aW7c
r3n+v9x8HlqZRZHryRMHmmgdDMKI9ZrkIJmolZzseSWYnXAqniXhEt4U/xayoGBfJ+RVcOJklAfI
4vFqJrndWLjUOtP0WcLuMBNjvk+25cZ1loG5YDRutZXQRKt6a/i5sw5jmpscWvcGI+SyZwUbRp73
4zE+XYtJWZSUDmbjMEE+WHRtHT35PK7ZSrw5OdHhNXEXKudk3//Tr/lVXR3cpJscOGq1HhMMXJRG
4iZ4AXVknsjresthpD0y16nV0rfbMdwfgNSzKq8dYHg/UOuoA7XjERDRNsFI2SBdxhCFjENAo+8x
tAro9ZZ8zuomZMpRA/Ub+ydx4LmudFafjv8Sf7wCN7kvjve2EUVCbBHyjlzGRGFsDNwId5o21RZJ
Z1Y1dEeG+D0DQdGauxGZ54O+ks8cZvLF1wGPjbkY8h1AwXoP3F8gu67iwg58xnhK1wE0whwflgN1
Axldn1RmrvpBXt52ZVCF8spcEk1hqOpm+e6jQ6exCiEPiQbyPKQqhxgcC28wUfysQJcaffHX89c8
KMW5cIOt77ilboiMuOagV5JHPkYbsvrw63aUuLRtYfCwBCyVrP4o6//A+B9CPacXMISHVvjtj46l
SEKL81+xAwSgtprKCO00jQ8oqVzXSn02Zb2zJE0pR7SQuA93WLzuzkurlfojiSu7LrxuLVjKt2S5
+y1d0c7CqvgCmKxAudjzEze7ogGAtSFN0jHEDIv4asrBEmUu/JllIzMfCSDqW4FMEBVpIj6ELoSS
7H5evcc55DmMcxSWpUMuNZ1fmfCL4j/jmJh+Lee8SQVkGW4a0FPsidlP8qxIg3AgjdMNFVCdav/p
TB2ERhuAQudpXRAEMo/WtcqgJoDyR+Ek+KWIg3fVY+sTuHzpAkBmDSZ7ssyK8Szajm51ax7SmewD
C0evoLkC3YFupoqqiAaG3Ad6bmNQWvhii/qUE4LqaQ3sd72rNeUXGwaa1qFDHqXge8ckWrmYFcma
qGm+FNa53of7MyG8CAr/8Zwhbf2svm3gyC1D7zciK9tF757twyEFC32N6ZiGBcDDbvI5FJjnJGKS
UR07qkR6HbI/6qWx8ThyeOt08hlWNmKsbSmY15YV8/dzrolUKwT4LrmMlTqRELisvG2dnDf9L/g7
QOZauY3jnadU75SFKb2eWaY0GrSzZ/CutOXh3ErKW8vMtQxx6iORItpGLmEb4RYpbTwJUf9RNyhB
lhRp+W09yu4UZsHMdm9euPbzpc8jkRJR/MMEUonVgNiVjxkHMr8jNsnk07NFO7PoSkricQ9mICJl
jLGszNz8qtafS8HTmRUKWnzjlLxm0G2ZOUU+ztT9f//wXrh+qVClGWQgyClwkTzBmECKC6/O1A6B
qtXOCuiZ+6KTZoryAI+9RLIJfTUdEPMfJ/yialSc3iAlet5p3VFl+ymGKwwZUCj86gSqw/2g2bd6
zQGm3gIEeDIXHfKhov7u2xaoVwSbOWA/y2Ue33ifnPILbK0Z9YDR4snJqwhR3/JbFPz5sD+hIiLp
PMGvF76fhJhsgdz59ZmFYNoqImpeFKcU+N3/S3pUAKl2YHxYpWDnyLa8nfUtoMfB1VxlF2+FfAHi
rTyjT/pEPd0UH5koAwWzcCQ5/taB0jnDObfwKkVbpvT+O7IAIdY4Ov3UpcL0BL9LqV0oUcwNF8Ok
URyWEYvAFnf2ZXNABPbdY3/pupJ9TzylrjtHiLd++t0OJijiwCuJDvo5oTLsKEpJOfwavrMZZmph
T6uKbIske2hzcdHVF1JLhvVwpzhVoCF6JVI9WkAnv8ql1oU+WMlEKjXA0Da2piNOKCTj9zeBbfUd
xJShzn4M4KI6Bw7bYekojgIYSR1uFWUH4Iyr41MPD6opToDNqTjph/L76jsvK9SsiwaXjwPafezP
CZA1riZyFB7TYnk21rUWr6h7Cv/y5d1+Gcm7YP/TN1PbcdvB21nxBIXEXQeBzNEs8sKuI87v4SS8
rRyZthibry7k+ow+AXLYmiEL5FAvGikQQlSk2eAR/YcTcrWog45agR2CdaKl5+ZMRQ3WONnaWITy
6qBbE4I1oI+LxfrpRSa5k7IRQQ9x8kXWj3pHb3mU21/NONk/EC11bUI4VW10f+owHQmvTenExxIs
3ew8Ym2GYF1o0nRrp5rbRk6Y2qm156Enl3CYeRzNv37pi9uBjoCtosoIkC7Mo6AqaedjUMxBg06u
vp07f01q/T3cc7KRUzAHFDeNRcvMFBDSDAlrTd0qZimAN7LNbQlNPjCVH7/E+yKze+uPEUAjNixa
ft0Q8k0Nl4JCJ9A++dRy8Gksdw+rd8B4GJJAlNYw84/s2QVsObyF9zXyIo8OeExrtSljGNQDroUT
MrEY2yvym/Na5gse2G+APFdbRjvWY2aOPA3hh40gTEl49uaNJOxb2ZDFwH5020G3988rhBytGG/5
u+7GJAs5uYuudww1vGAB4CLZozpd91k8nEgTY6I7wH8yxTGoS1UdMNRQjDZO7jU99M54kYO8XUVz
ZqsMgZL2r+Wt3skt96jK4W3zVME/qgC2+S4YZZdRaesVh2oYl+wX1stdefrZE9F1feov2M49Yh+S
BNM2CDh4xfgcwxl8O0IN0hSRJ67VvzhzlxjhXoV6GZm+IpL3iV/MiTUboDQD+/fXuZj/7T3eiVV+
vsAovgnhA9Y9kvJKSwdf24Ed90yR3jhRBser0pVFfvY75BQAog/2USRqSydFV4dulXt0NyuECXy4
A2g1ufUJslC0GIXC0ge/Jl3fMrUGwwNpYqv2S1nkm3ezHs1o+0e6yNYfS2UXuq5rIOpUCrhoupmo
6Er0lxVrYe164dYjsgZ36emDG0feuDLajYbiO52rqMZXXE4DymXtG0lhyvOElPbmxLj1jFsek8Xg
vaMLaI2iOBOri+XZLOI6y4bT1JLjao8HrTiMH7nfxJI/QEpv9ZWBcSBcEPWAdL8FAE3CZTTesG0m
GMMthyg3L5HUqDi+t1qKDPqSXR5XFnsSZYSkMUBbAS6PrDgapAnhgOEiRR9IzQJoGr2OtbN6hpEy
3sBQ9K1Ysb593pN2FebpMZbZJWi90cUVJn43vRiRlEDnKjbu4SndK5QrQTfolHE4SNOIJJPkWYC5
3j4VRUcSUZrjcYKxiS5LmtFDIS7vDmKQLQgCKq7FsjH0ivTQswxfOthMFflJw1xgwTSebLLbfH+k
bx+gEaIjJ4PH+7Z1hLFz5W27CrWlck+Hmax6bdzj8sknK2akQ23rjjsmeOqRkGdCg0Vx5zoviXD1
ZODG2Ky8asjo06QJ+pvwqx5jvsSoy/9svojARz1kNu1iepW7SPPObx8aotzjjzxaukV/GiLZfwSF
3m59TrraKB+jIjzdjWRqVHrT6Hu+9MDOLFv4cpeN6sQS/6olWafnsKCaOg3Q82EYwUjAGdaI2xZp
JKvnLVwN8WuNvI8ntkWcSejCfVINomSSJkYhP+DxTmRzfXfD6Un24Se2QKnPOpGmPkrNgsbIp6kp
eE0R4oU5rPklGruI+1pW0hL9v7jWNLYtsA8qv3+sFwu/TTg6g/UDn6DyF9bjUX4T2pmAsUi208cp
20IX4zieKCBaY98zo4oAT08WNMZuKMb33HgJx+UTgSw0QpmXnq0Ha2lZQohP+2+VtHamHDIunRjW
VTdATl8sMMyDxz83+zpXVk3GV+PkloT19V3zaUZC2yCrPsyfLQGX0dIBMwstM1Ndh0NXnf+FUyL3
eaPn35wVeBz198d+7kbLLA+x/kwDzQObOjuvAg+G9eTi5EJCp/ubAUv3q+yWLtuLDle5ULo+GEb5
SysFdalRQRr/DVhxc8Td4J8dfM7gDvo8/UEo1hw2Y1No4Cn/fHYMq60kzq8tnP0MOniZJ47xWpgk
dNDkNcRhr2pHv1iyCeI1TLUBunabFb8UwtNrlqKvmX2q6X5tX+E5eutAHS5JA5CbZkHP0BTkVnz3
u2U0pbSgoDmW0y55S/Jbm14ZLJ2uDl9XhC3Awj82xJvQdne3Lby5277XcIXdaKtxZQA0ma8faGjS
rXnlx2eXtPY4QRbxOQV+y9cIoGrFhQoZ4TAniI2XDTFxP7qvonrn2aJvp67Z+0EQpNXq8SKvgsLh
c314+jO/boQF4Y2uMl2SrzNUo1LDj08ZPYZp3VVuTMJsozJmtsmIJ8lhrlpB+7DQ7OAWdNouCBok
3oTIZAJeD2yR3HwTD2GN/Kyyzk3CfMqBhDotybTRCT3T2X1UXY2DxlL0JlDx5RYDtRph9T1ElIAl
KaCovlYOFvh2xDwsu0I8eYQUbyah9Wvy0Ad4IJFVRXnR/UMFvfU+0/v2MJMJeviZozkl2aGQY1i3
p25CDlFUSUcL/Ls22CVgP4eqxO7qXlF7S+pjJtX+B/y1xqGwpALAAhbrPCpmBvs7oKFlj0Z8oAmg
M0RZ1X1BM0SyLAlzX3Bdn8tacrBTg6hBX6L6rnLjBIbGlReV/0eyD1ZxKOFpFxiXwyn9PxO2+NXL
WziWTnhRC9yD3q6TqBLmYrU1iJ6H564dSqYI34XR+CYu4UDsPXhVx2SYUDz/MsCG2C9EMO712UOD
9wsxetrqRZhY7dIf1+3IK4lKHdRy53jnWwuChvwOs0ixx+P/RhwJ9jpoDv2W6w992osSntMNHaKb
Pdu8KLKvYOLpHRspW6Lt0X7b+wzOOEp0ZTiMAN2LN2tyeNIKsv/RH5JtIf/i7526Cmii7eSMdllM
1MgzdAumhdaq3XL7Aue+GmPbgpF3KTa93A2PbRx1QL1IGkY3NhycbCq6Sje5msmCCSzqaKWC5yoC
a7hRoiK0R/eNZgKqZkq/aYVT7mMMb9p7nOXhCOoc9tUdCQYWD6HBtwz6xd367VSzapgJSGOoryNd
QUPEteufvpAULzSYYR/dHsYH2nnh2fg8/ik06PeijxDOJ+b3CJ/nvStpnK5x+ZhCg2RvG9ezA1SI
3HKI61XBCBKEBWvAj3N630LmLrfuKFyVwQ/jkdKUiSgUCiysUMvypLgxGLGx+iEi/F8YZRU0YxdE
h5msdmiI1ZiET5kchVGAzGFJ5jBFoMEWKRuJFgib4ndOWcoaA8m7nJigonDMo4/O9zv6VsVjz8YP
W/XPWulyEhEgIY4HKo2WSmcyHL2W29+u5UioKjuPtYqrOMSuzijth97Y2d5jY89OJyS30D9P8Vsa
P7g5179TtyOd1EItqZXU+33YY3kJcfKdPXx8Sg0/5i0kQ07I9Up4pZZzR7s78QCdC4A6i6KG/jdH
CTDFRr5sUUNk16j8l8VdICI9uax8ph+Hl+/I9CmN1D4k9FnWkX1tr8DUxQQQ4n0BJJ6yp2wtU9Eq
6Fm6GZUZA0FTTBD6zPQauxAysnOqhz5ZQ8eNnv/n1u0TmCXsJBF0QF9WhhMLPdBlu3FiUY0QZEsI
KutaP1m9A4yF/K/4nEvcePwvZurACcs/rhxQuwj6oLz+f6wKQjxysmta4rMsb/Ecl2V9cwU+XzCJ
xPDxa8EoFpIytJaq1pma/lTSW0uCVNZiS9FNh3awqgqevjepNbLmDDxsQnBwZBjh7E2CGkOIsZp4
dB4vZzE18TvK4K6QYuPu0G5noGagHrhIZ7iJx6mKA50ZRfIVmIxSdkgF1IdHmTB+VBvYMT8TifoQ
MfFicVskkXMDfVSzp6KZsdKhZRIhEG4bBLOx8kcsVLSPhlLGY7lDBKuyripj8nakDPCbppdHtm6j
ozqYpiArZsDMVTv1alZ+PZwgk+WVu1oVUpAOZJRkYI6B3j/NXsbWm6r2RCflNHGFGGV17jVj1sdr
1Sd+wQHmAEj7yGxI8XXf4hip5dWV1DqTpKoNUONEOOG7wz5Rwdj4g7DRtqpVemZzLd2sA0yG4JGn
6DqAfqDErJM0CvXTuRioTZz9WV2UyGX+noZE6ccBUbG5brjFkYecNbjfK+g5ot3GtD3qBs+OFCVy
jXIP7M2Qmf6OGA7E8RFnVzMf+LY5JxxuQhIeppqP46LHyeijaf+TG5lpg8qgI4Qb6plcz4Hb1SkZ
pjylukH5RuWOc4xc8oAdRmeKnngIPMQ4RMweSyG17j0sJ0xF5opqUl3to7PB9hCS+HSj942OZuxp
x267xezZINWA6B88twl26BcMEMYV9d7EA9VV02/XdbYjmhwQz1KkBSr378W91rW/aPswPUSMSzBe
dR0JyiuIcy9BtIK0fY+Lii5WphJqwxcdYnrh8xSQKtDsL8qT1kpD4YqXzlDA1LYJuONeklsYmQvr
ZE+16JUmU0IiPxcv67V+cOXodG6hI4qBrw7naqcRSJWa7AdYRWCwFEIsrZy1tXgL2t0J043mJz7Z
lLDY9SmlpdrbM5/j7eQeXZwmlxm7fhgvfqVhzh1Eofa8IbHhmuPU1clNyuVy4FuyLRTLLKXzWVsU
xCI3fm8ezHldkJPDpUjgWEwc23WSyxaXtNMDbCZBoyaVDsXvKMyvrzHpXT0/KjJImcGU21e35DKy
/91bVNXh5lp1oOGHxnvqu5HLATBbEeiEo6zbOflI1k7OUJQCrCH7eSqQbqKIp8/DgTcD+7aR6EMz
rrL/FlOCrXGR6OaOSJ78ni7Ojk/2tIdNdt2zeVyIwXZiSMc7ZfFtZjIgNbdJ6QsvNmtRHRmVGGpe
hjDchHe6+LtsFrHO8SvPdd//qJYtFN3O+acCDXSjr7x5K3OZt9aF6YUDn/nRvzFoh1oKZBrrSMEd
wrViNlt3WjknzUOXyA81NJqMrE7RzrOowLkl76EIPPdq26ZFjsqq+v4ge/ae3VnCR9WSHBH8jlXk
mTe8qsbeAc1+HxCwWjhhGLvF81yD5mIKe1jd8t3oKnUj2mBlcaXp8cAaK3rSkfLsunoq6dFxLrb0
TDxPgex8Gt7EnBvSKGhX6YVO82OGAb/ZYCnwh7MDk5v6X1u9uaEGGZqj9japx32EK+/znYQ8O3a9
tFyxVvDDIHuLujggp4RRRUaGh4UnZxsjSmL2MozhFtIaTviy+DnJFe5BDvX3GcX7fn8GWEJ+qCGG
wjWeQTSLGN53kYikkZi3mtj+wsRXZNWmdIhE7IXftL3l84ob7evH6pjTz4DMqhy8dNw+SL8TOqMS
PMuNedzcYQRWcXPQm3devehNvl4ycJUMvsDInguvev6p+bHPuwstHRwW9eRSoRJAUe4qPf1ssuNZ
IufBswltUkEU77zzD0lbnLV6ukA4vfwmmAXLiw2K0vyzLZi2QMs/iVQ+LJTRIzilTJ+IZ4h248gf
+2+TiP6rF3+6XCRZbIYCF/lsjQQqY1VKrmhE6ofOtVuAsh5YKow7kfseZ/mwxYJBWVJju67zjRkk
pd81SrlBdMKDbUoUEg3mv4tdZhRzrfOClEUgw2xRrxx/b3m8t6FT8PPHE7KwssBtX8PWU56idWGf
KaubQHEzbgzqmzTbu9GbsEheh5Rouksf3RtAqUbZ4/d+rDkNGiXdUV7j937jrP10kDL10+DFt2+b
1XtXcAeVo5k7GFw9lThIj6VofWWacJeuvLfCj6l+pfeIgeRCuAuwsKU4qHJcOJx11YyxP82iVucF
StrKtgFyUKbiB4qiAaRwjZSuaaqo0mJSp+GSItooo2vxYiqRPUpAJMQa24sgZ4t8dFBbnhfPS22k
WKmYBiaVWF1nWF45W59YWibz8gH3HjUO2gnAFru89OCTdS+Hp3wL9Tr+gopguI5v7EPIgin8UMls
RS/52M/3v1Kp9IfwNQsUHNe2/shak9Tvm49sMHMadVU0Mv1Na7c10GZKSgXVieK4i5cwLLfTdDRL
kIxHuC4TK05XN2mTeH1oBRKMsOcPgq4bMKHyINHurXr7tHJlyENup+WMT7HAckFT9tbc1rPQgUof
FuG3AMSRZVBIJZ68Z3BMXl3DqBIzcX1Pvp9tMGNh/rCvX2GllxHwu0zvfLb/ToYx4oeSMvlDhhDE
hGqQQMreDFo1ah4Raw+qmKNKbKCwN6YbagkqyCrh5SelVfoCmZ+P9JbBDoVgQyc9U7m9fQ1BIvcI
Ipzd6dsARC66vzjLtA/vDz6Z3z/GLXRwX9eKTcKppTssuGV+//lI/3ZqhBfjm91N2xfHsnQQM5rJ
3VMJsxl4w9lm2clpYPFDrt+RD3zjs6qqx2RT+RVlZOxwGVjwzDgIigYGiuhfhGxZbppDMH56aIwO
o1YhGhSnpAUAolAb85wnMspJQYH+yIlIn+Z8dgAdtXJnr1hw5629dyb35H9IMJP9NEIeoQmXFgzE
SZe8Yi67Fg2Glr1YWp1LsaGaDmvWmj8eWdrs9siAJ2JnWnDFvMKDBQYpViqFA57G+grLRzxqYHjZ
MHWxooGneun3clThQxlmRz9E4jS1AvX4A7qkRngvTaHJoog8Sn98ZHnUFGdrqKsKMg4P5EvYzwQM
ziDNz5iirzylcNyLSodV+JHnNVjlhB8PMlLR7ldT01+9CsSbqoS4dd30Js7ZHHzq+6OQVS81YRI8
nS59lATwcOY9VSjfngmhJS4n+IUvXi3yx9gI5tEKiXOcEO7SKiJceHD8/sxHxiU4ly4H+j0THOgj
9hemG4mKpSiaqLZO/T4zlz61fznO43A0a9b+C6eH9nO1Z3NRS5vyaMzLKIgftdjh5kAGqy2qZnFa
ZrdERSXwEwI6EvYsjcdpJJMhaMF2q0O8UU2rmgOGUjwBe8s+/MmSW4kbjhisACAMBUyVk5hoC97/
+kY+gQvUELRjxux4u6kXbbduDGa/JCYyyaUEBdETnw84NwaHs/KtNrIkX/6wt7fC6xT383Aa6eGv
sgdk+cPA6w9XhQ+r6jBOiZLH22Kt/fTnKhuUg6qL3fwUBPEt+pQdtz/VIfV6MdygIIQKlMtBikNa
L8HUGXBgPzEzepuufhysbIKm5qz3EGHwCPm3a+5U31nyaus+bitunTz++Qa7zcgxxI1bo7dS37cK
P2aUcXTiK9rAiRF0V8tn2qQDGWJqyVW8JcMWJ1kZeJdP3p4D06GGW2KGW4nzKXCW0P5b6nkoh1a2
DZYeovCeggGNZIL4WL95LoAAxeITGHkVa634AAR4Nz0aD4/dkD2vvGtTV2b3FJm3P7gEkwVjV2A6
Rr+/jfDAqrf/aNUsNkCyAjVaZldA6T0DbRre+7zCKGXpCjtnNjuQvDkxkVh3zBPpYcor+gsVqwLW
X3T+3XcWZxV9/Wkq4AIhEgmeMzN5Q4925Gh2hoXCiXmaXN+9QLEXJsDtULhRDWSOp0eBRouPbeyg
93qGGEXMQM1KdABo2m3Zkcz/BXzYsCATiOFack5Fiyfk4P7xm+oVGqxNZo8Ne79Qk9yZq/wKbiSd
kl6eSm0qq6lALaRmgBUF17t2951caIC0oH98L1xRv9WXG74QOCE7R/AMTS+s0GstYVlcT1M/5Am+
3ilPpxXCy3qxYMEVPE8VWhcqGMzJXH8u3j/YDBagVVjEeSNe+NcyAK1tJUfsLHMyIw10x/VgSJjq
G8WHW1VtKH/XiAv9Tv2H392Qn2Eyr8xtWlg3+9dWw7kI4zl40cDX4SS8e6encfv2s5rZaZpla9Vk
8yFpgm96q2tbIQsjjK+muMPXnRw4V/4FyhXuIbvWBykbgKANn2JjEn7pJnPYzkD22m63/f7KXzUl
v9q9vaUNyUiWbXCkSxfS/1rr0TRF8V4cb3MI9sZ8Z1e/3j1Oe1zESLr5S94V/WZiHK+jMIz5KqEK
gHga2V3hNyfggi9GaWRv7qm+kntb+lQZSkiMA6pujXWGYnDm5obMUYoUOCWkFBviIKyxXeBEfrqv
ELugPCvxdD/9yh9Fsm9UCj3Ille6rxVuITLFg5af5K80LGRMNSg7yBYOzgbmiMdnpARRmqf+blRF
t42WyNzNNHCgjGCZ+2mA1FIpNqkBLuieZgF5OtuI5pMPlhwbMm7IYTscYgLovMm/HqvLuDqZdFI5
FDqfJ5sW+MjDmCVjjbSix5hYvdylqiRuhFt0CIiF/V60Ua4p38ayyGIeu4Dwvyn/odLvPC75Pk1C
bLiPmOsRlrKohbAJLtwGAeVdy9MGpqM/2CGF5yUXKEY3rfxQoo2lvJjSzlHUPMTFSkGohRuMZY82
FFcjBqlmkGbB7ADlas1wQKFDRQMZNB0djUeHx3n9j3CdNt3D9mcRFo5762T8kDvrJhs85TaH0XxI
FVaxRayFHomhxp9AAtQqZIgl659f/qtJkmYZtB4/DuHZyT/G/Jis7AMbd6IOWDwOEBkN0Sg6FT56
v1ghmjJ6KO2AwHsG2mTSqpANKfSqppueIey9DQsfAhP2OHFSnW8XNKIFUfWcm8InzzimcJ08uJiK
Oivab2EIbOccYuUdZ4oBiYtNqksatp7H5YtHp9fRiQRfXHj000ek+uW1eJKtFe+Pn26vioDBSX7K
Nk9gM84TXa1QyGjZb4fXyxHEYCi/FmklriRjPKgAz5gTSvspwM6a1yco2bUf1+rl77rXm7uua1N0
7c/mOdvspP8HPIpR0A0orowagLkLmxbcvsuoLdl2t0N8X7YSNd29KoQ3vobl72n9iwtFVwG7JdC9
pZpuOyMhJf3p467LN0F0wXPIKfqxyvJ7OR2KeoHx0B85YtODiEt4E3FXrFsTGw3zlyidgID4NrPU
+HBHXPB9vGIXv4SlDfpDGjq8WrOZ9uIfzJYsAT/aynXogfNxbjWRnOf4dpxoQhhMIj8ZmUaHpoQO
WHI4L0uJFan4kg2kBfV0YK2tXomuIeWA115q5hb8RaSRa21ROMSuxtYWivGXhJyGGyLHBAUES+Cz
74IZL/i8H7YytSC9iZndomqCene1vpDShacR10pR8lTLhdQkUPjNaWaOQI7einK+twDA9s8qk5zS
ay32Dm/yUkrzvZwGQ/16ie8CTY+sXJM+vVltvXtpKIMELiiBd5tQJA1FK9w3gJtSIX0WPRdZwMR0
fLO4Lwnr7JjrpNp7//8ctv+kL6V7v6cIkyBzH95gyp17oKgBW8/NjRCclcqw42D7vorr+6vBdcWk
ARotriXLxUSa9id6SbW5aWH2rq+S1aw3F9UhpZkqQQvHGKv4hGgf0EzJn4P1MUKIG7VDfI6vybXG
Xag7vcqcYU6GqBytpvPZO2MYuDrbV/eNkHrZKTt3+DjXhu74NWqvfqT3YIDgAv2U5dPiIv1RDmxZ
y1PyDSiADLDqJraBH6kYAlkBCBEyvKkWl3xKrJUznivHL8ffh6kn1Gx5Ey9c73XYULV7Y7EfFxI4
2FNaLYD8Rk6ADqeWCzCxQowXukzELnADEZPh5D7xnslBO3Sm4LwTU94a9/syJ6Si+yTJwaxQgFj1
Qn/PrI4aFDPP8d48BbrJoksrJboLXtMtc6aTNKBv6GQsnj3++YnfCSBjL55sRb7RNtn9X3TLaF+S
lBB9IpP9A7VrkI9wmI2BFhWRM5BsgvVBZPb69O/gMQdOLSU7/VvteZxxuywd8IdGW7Irf2vznikd
yudbSmlQfNus0mQj6QEASzfehjj2GOaX7sijYbHAfNF479SJ0UaNXnm/i3/ad7qR5MvC3uTNZohR
2qOnbCEycrB+lebW5sEHJmC12y1P5Af3gOYYee3v4W80d7AIq4GXATSjrYNfXlSClp8tAbb1BgqP
CEX7NRXDS9fyb/ASR8egvrzvJv3TtRFfPUSVJEy+u/dr8K53yUjLxjYxAg+p0y33jRn670u88PBe
yDjT2MAD9+n4Hk2LelyoSwEo2RAgEwVRbZjsLwTG/bkbnVTcfvzIEfcnxszgYjIBmymE4ArdmIgp
TA+PRiw8pAzfICo4sioXMUspEsW33TKd02kD2CnvqpZGDdlMLfBeKS3WXsXTzVQITiojDXm3efwt
U0Cqndsflw6QMYh6ss6qje4olR8rptL5FCEkCJi9khLU0xR2xGv7yo3TOm/y5rxuEV0HGvIZHxrv
o2pK/REehkyVi6F7PA7iVIfQVTxivDpqP2Cwq7Fa+opB9QZS/qSKW+YuZwx9No6RLyi4jH2ELygx
PGrJSAuz3Ne2ZxiltXwqczZ3a02HbO3smu3n2Itlf1eiuETC7k/6qC9nne3NBq7YSphXaFaz20Na
076M8tbkZyV0X8K0DCuCLGRQjSeg4iVn3i3amFtDX1GMYOiE4HEWAOEQ1aP8AXhzjcgeYANiP5mP
l24uxu9tWN3Tu40CSanv1UDKuP1o0gq7mPM9xTy1l0cEjroEVq399HyIvdi9MUWudp2f3O6Zyoka
YNGWOFLyNfxwWe37g1lcC3DTMy/pj0hXEiSag162jhBfKoonZhnWMWMn2vPobofFfK/r0BPH7Sfl
2F8DFaeWyXPjYahTH5l1/T43XyJcGYC6L/+Hmm/it87puFFzXemZMg6N/G7JWJHrbSQpgY270hDX
4CO+7Qt5eQTB3/R/jonXfqblUvkpAigtw3W0u+1S3LCZw8quvU5UeMAomQ5mdKet/8XE/rbwLp1V
KY1T4vB4/adWHSyiaETbjVsfyi2oBRPaaZEgvN6uw06LDLU8A2HQNufDS3+DphdZ2IrHy1cBntgz
ij5YDUq8LXjiz2W205FbOKSPqjLPGznIysNEdtIO/OqdUTIaKTN7toEsQB2JZQ5xW5bi4XfoebEY
EHXiEaJf85dkevgoXbXcNhh2+LKPQwW9eEIntv8Egm3/vfJHOW0fVCSVWYF4pqNTsOAVtFSuwOnf
bc1mr+3H6XjDyJyto76isqr+ZPKyVJpCXyzy/4i70svsK6kjGLC+wvfDie7lVwE5QyuzaSd49yVb
mRi/BifgvWD4opRnjnrrTl3bLd/Orb+v2+bG4vv0UilMHwz2YfwWgVRp1Vf/hZqR7AApLEMeJ7Wn
tfAgRj+tkGpSjYyGmVb5VtaiovIuZwwTBmfhfuGePCet5gGOgc2byWeoCwXgCTooqvIfFPO6iFWg
aLn+fVSqtzEmAGSKa3m0k4xEDGoqV/4fjF8zjnCx3oe/jnUh0NHuIVgi/1adk42fVnSu2irXrM/b
aqZWx1+K92kSlbSy5OfbTh5ZlzP+tYh3ikBmrM4Ort5/3Q2FQfVkg/dOc1VQ9Og2uDGF/JQAnuMP
2088BmhfOl/9+V1TIB1d1wUy/W01H94op5PnxejrvRN1Gccvb+KRzicTvP/8q0fr5F5vmh+43/wR
wmnkaM/Vn8VVqW8PQ/88GgeFwxIScVD6gWy1cPikQp5nzu/fX7ZTjcf+jwz3ZvV6yxvxgGNDwnRb
jw0SSz1p9JUzrF0ES2Owmco/7FLDhRI8a+7H6ov1DaUYYnoM4nYZi4pq2uQ28PkQiLdnTxiYbJJ7
mgXaksWrzmIu5dGCEAOCm55Be4sZpzHvZfDw1nXPTN7FXXmvK79OaxtKy0FYR2bqI6rlvwFQQ1GN
d4tPVIGFotwPy7tA2+AVAc0YwYrSPyBka/vqJm/e74yMaJ/Ig7jkiKG2ck13D5PQUCs2mz3S5YJ7
YREalFVj29sX+apvlp9xekeUsMRHmlb5oWl7d7V6u+H6u0Dfg/otUzydPZSnPZgPoQCk6NRakGqd
mLHSCddZ3qV0Uvc4O0ggsw/hHUwlP4RaLekRoHSEz4+26bOqeRvkVxUZD/PjgR9F+Sv7xlZkDmK4
H1nEj1aP32GUIdLpkt+5KakccDbLtJnEvt34V9y6Dt7k8OrQblUdQmhfWPyCj/8K3rTiG47MTh8g
vG0+/Ydt7NhIpu96wh8ZWJ8583sqH2T9NpIERliQ5/SppAToJZJHf0DF3EINgCOQbg/sV01C+9I+
Z0AIds0X+HzNpEK0pyKhVYLCJ/fwZ0VN3NE6ZaSiiOZjDJGwlxDFNczStRZF+wGv4X1pQpjaoDKp
UzHzqwcECpYOs2RkLH8TnisaGz1X2284Ng8kpqfnfwkoQ3EO3lrt0WSo+GMYeSjMEoDbObcdy7Mg
l6lV5N6CY3fTniMl5eVd9gjzUR8mfWGmoQeCwwxs+y60hK1Hdff7BCIVASCmnReCMYCx37drTOCa
zcZMWT7UHfReFFc8EWDs1D/k9cYnV4yYMNgMLGiIr4DsEYU5EcfXbSHCwA310QYcZUW1MVM4FgAp
74jaMeqt6N1KIz1MfDBNyQRlSAgxe8tNdR6t/jLae/de/vdpPQVaOhtihE6Q007OY8nuskVEwREf
XVtGFWYkexSL5cDM/Gx0wqZnr4IwpooZVIC5LsQfG4u8uFqVuNOFk/fxwNVo7+534r5zqreKUEDm
aX341DkhBAWyusfBwQNEGmXg0ZfR3P+n6TN8rKpF02h9Q59VXthSOe9UZ1WDfdWV6R6hACPcVtXX
PZZoubfjzNzaGd3+OQLVIE6lkEGrGaOPlOluktep1hanzSyqZhHqBgOcu+mAh5JxpLzZnOd0TzA2
JUgRZtDd7VqlLTxt2MorIPlWWmidtm7nV4ikIloPxhzFi0dgdS59Z81/SEHUt38RUlST3cnDlIq9
39vyhxv5aM1P8j6OiS2jUCUitl4iFBY2t3KS+ObbF+ZZQtsLUCCABFJE40FU34l7H9GlX8MNkIb/
3ZFn1ovbrXn409CZ2+U7XgldI9SfWmpMac4tYRwMBHsutlPh9fQPcsC5XyZorMtHzO3pZh24bQ6B
xey67dj3oaiowEz+87riSaeBOWHbUpBViYm3jfpnFHtTMO/FclAmSlJuEk9RlfRxCQBnBng9RLHv
mIlEwgrGcFGlnF6/wgSZ0PoFhbUjpGR3hicSOh9zlKCMnFKj6YqSrLiQCh4TKHJCrxse47Ux9IBt
tCgV7iuD0teMENOOrypjiWuZZrV/nz5gZqEjsC2DmNAF5TUUF3wn/DdXDIQ4iDCeWZJKrjo+5K1e
tt6hNwHhla9se3uNciEvBcV+4oirD6LByHp+n60Ql81btuNC9X4zHp+rL02HPn/iwismdAOgVTmM
ZjePwxnihQTE8XJQCbeamQ40LTb5ovb70UXT9EpZaAboEcNqCoxP9ll5pQMig6IblaEaJgYPXBdK
JP9HyQ2zsEm9nkxo9R/ibYhWqozWt2HxbB78YACFogLvSu/yVwLIYJ/Qy/rRmjggfR76V/sk5JWW
pGPlIuTYWTQmPogbJ4me7lNEzNZA3JU+6alEE8jHEMMTpFAMyzlaEkDmvjKHYfPonWGSCYl65yWJ
0paAXgtHnElPtAbOgqm9J6ModuK3nBtHeXlXb7zHg7OTLMjESd6rqJEp6jgQ2IAk8fjYKJ5q6Hcu
mhX0dIKxs1ETkQo83ZkGH9XXqNlTjQeTDNH0l05Ik1ozeLy2dcLzA4W581UOfhGgPP2719GVpQ8w
4a+NjXWXq/UINtGbpwNKiW5fLogLKTJWPPlp1cBWy7LLICLxnG75MQza27OJNqClFkCb9FBsK/S6
w32I9yblvmJE48EaLJvKEPA9YJQGVoJOYQ52P2DfbdoNsXV7Ba7dfi45daqBwwgU51KVOGzG8eD/
yZ9jQdmTqVHZKkUHqTvjMfZRnvEcTGy3F2HaeJbDUrTkrxASV4iIpKLj1MrDysUW+xAZe/tHlbjf
hfyDM4bUvb5rn4LJToLQ1BpuCPlXm4om0QSX3NoSxXyVl9QeLSQsd3CaScyntTYF9ShSDdc/2Kau
EVnAO3VSDEWPkVSgUd8J6hQKVD/4l5vaMbrLk/uxWbOYtiU2W2a3WtdZZzoBgrYs04cVSw1qPbUR
z4YaIap8C+f/gJbPR6czXL5/Dyicj8rYO2UTsbiHVkPsCgCoF25qJz8t6PBwWRDh+uZJhGwmwGM8
VhldIANTREeEizXww4MQ3vQch3tTQHdidHSaeSCYDFO4TnZhIShO7WwtnCWAE1lHvdFT9V36OEy+
Mtrudzww8oBO+j0jaslirQ7QeFIM0lYCL6d2c+KFnlVvFIlIPLjkcWWENnXwxtxcz5QOBRaF2kzJ
I6nOvz3dBRo6rUmSXsQvtxNNGte9glqnzCT05lwA6dLBc1no6x2YH1OCsoN/n1lKbD8/CckRlDSw
qaeR4GwgnvHarCzj2g1roTVaQyAZMBpOzEtUPymtlmhMGAFlbXCWb5W7XDMZLNS8MZSzb4ivMhp/
yrU8NFfe23SIlPAHg7mzazQQ9SJjSsd9ERRAz7XU62v9FZkStPkKqMh+IJkf8DTNLp35CEo18vki
Tv9j3igBd2S04j7EwCKLKUjnE77/D94q3zIQNXfLcgG2B85pR3XsBQ5ubOa7Ka/r84bPz0Bpr9AN
4OqyKKLryrAmENH/+qBoj/uXYivV2qexLuXqSN58tp5qkjeHgneaLLBjJURIFkU3SzaL6it+Op7d
9T2lE2FkJkgzfIVLGWrkq7k2qSsAdzDQBD7t30jX0FOU7wWeLIBpZ7w1bjjiekSdvpOzGO8kh5gF
avYSfoMdwABza0+ZKuOcEKq7vVLJnwfrr9K+dxTgypUqo2kEJo3dAPwtqEkBVSDHkv5SUf6z7n3F
Cfg/jQz07tDWGbGXIJbfQv3vlGuTwWS2DQu8CSBl2sH7kzQ+nkPCEQ5dR1dIygMbikyPlRTdaZfP
LbKuCsBwmzVFvKYNO5BaCdnokT+ug7OFcYgXM9EB09Pq1wc31qTvIyFCpdz+/XvkTVtfyMqtXgUh
cy1355xtoBvOAPxeuWE8qWGkL2+16YH4b+DtYrbJLL3BoKh7Ccn00OJhJ0zgwD/qUExfo/3b4DOT
eQpNG3dxKdHvqmZyiDRBBnbnkEEzVXIuoK9qLsnQU9IiUirzbuV4Ou2IQ3iAZcSsXn6+f6gPcieG
uptr8gUl5w/t2dSUZgymHVcO/tvPKE84fNJMoMspDxCaqSgolp8HFem3r2YxGlbDREomSPo01jPQ
9Gl01FoDr3UovelXeAGzJKupYFKsccdyqVE0aYt5/Fsp8bPQZFV1oFfFu4BmdrWdyTO+DtjOz+EU
l8zXVjVvTXPE8exfrp1PrwJy6nlt9XNxvR0AvVhTWK1eHh/VzBeQbnLrk4nOX+zsnv1X/Z1el4v2
m3fB1qkJQtnewHaKpbUrtF1PJ02GcIFccQhSp5N+V2KltLRXgaj6JS9Gp7tdJ4wEqxY+KvBiBKWB
Wqz9EPlly+KX5nm4EwI1i4+pdSHzEKqfEKRveD9KyVpIyevwGmXkGtTHb5HyHeZrhc5b0L2nVTpd
mzvlNDEAfBYRnjG4SvUkCKWwmDkEgxXpkG88zDnK1dm8RN41goyRuTJCRlX5jdvpkRrpfavpUWsT
sE7gymhjieSkUOOVIFCD0FsMk5vrQVCaaO0B27WqbkhHxgwDNgrnhxaj9DMrkj7wz03Dgqn3UZsP
dg/vQLlwmdcMnzgq4/zZen5o68HfrJSlayLc0M1EdyUwLASFMgzxU6MJYVjXKFB7gbj4kRoAfO/F
E4e7JO2hFoYLmtMphL7Sjktz353ucwW+Qhy5eUgemk4rNPg8yAva0hQMOIok3wKl6xLTeYG0xlH3
EcTo6t63IKaBG+ihx+M502E498L73vl810cnR3ekK+GV0CCJIkljPGtkmJRHscdNP9R9V7mDejVF
hfBCiL6yzzVSXAbFuX7Aox8huKiUm04ZxaNjI7mcsvAs+gpONAP1y9DxLBvtbucGq4ABdS2d0mn8
iTum90qwnPZgtlf5gAjkuKJan62fE0JkbMX0RiEl6bSvr76RXXrinuWyAwjXwhLp29l1tuuwofRb
UPTxeiS3SGVSseV6/+WhzgTOLnYWqdhauA+Zi7CzKQfTxueD5TNLcQSLjRX232TsE8b9j5b08KgT
6Lv34Q55ycPk7cAbndSerK/LPAQ2oWoVyQQMN+uTP0XhUwpLi9R9Blq4GQNuWh1PgI3U4zHpF5lL
SdpM+jgWZ3yhfnApkv2sYTQKjkv5OjPUoZwS4MLtasva100bozeXrawYm2qNp6gUptYqe8ZM+JUx
ngio0+Es8LzZbL4KScMfN29eCDXFrKrO2TlJSeM54pCNDg8LzGsreLv2wfOeXnD8+JzJIrB3VVIc
rLrmuyotX6kF5kn9+ME5u4FWb+bmOagfgDR6tNkOPe1pxmHACn8SfiMfFq1iiKYmyzTK46OakJI6
f4ReCTSwLWRvmjjGKULk+Btp+8VfpdLqnBL8Nn0z2QOh5sGSIswqIIweWR37R++t7gyQ5sCLEaB9
M9Gq58H+cbu4x5dvWePCOaf9znmOUwW6pe2X3ljHDDAqmx62ro5BcPw8chvjXxMLGgXKKP+U0utr
Uo+1UAHSufvIFTnYK2s2iQLAzwAHXUT4O0sbEAq+v8JFGYqk1pJLfRan+rHCbJymOzXCsijxXCvC
8OFn/GMnZPkA+NxXg+6msiUKq0WmsqMDcps+mKZqGpr3yeRjJZttFzIhuGr98w+/t6FaxzvIEJpE
YLw7dQwnd/AqZhBhgh3GW1az3dVX0nH8qoBzWbYBasg2bwCuEZji33k8OQmTEqk7GNOoy934wXtu
BlSzEjLyKT7cwcs9FpyFpV1U9+wZTtr61Eg30ebXktf5NLe4cPPjIjSG5qWp1QSAFNVXfOhqrDho
Q8rLfuvv6RNzxLGDTwx3Xq0ph/h65EF+6q2mHgtF2wA1fnoOZFedQIMrZ8+A/08rM+jF3O4zRhPa
Uzalh2VNc6OplKiFihJvGbdFf2ar839qlOJBQnATsBcopHKsGMevAsa0aPQQMFhGZi8WAywG7EWV
gYfsgb++DtkMj07vpNNm/5+pvOclDHobZ40mmLLja3rpuzsnq1LidceLVUrBFlzjfyPheN9cD3t0
DzFAG+fGTsAlAABMai3HgUbPcto8jVxY4vaaONjjmV1OcNmAYOI7KIKuWYuEAW81dqdBS30SoAjn
TzFaPSJjBe9V5GchLRYsBxcyTp1uWWfaPomecFMxNE00r9qGFl72C6AUMNXbhGcT2Z1Sf7KlgGzy
BhiqDxmFc5hpaejAWV+Va4+WEoZ545GMxZy6EVemNe5bFdtZGcOpA5JOhOM3Ga+m+RVD5hIwmxg8
HKWB8F1pvnImEVw3Il0PkRMDTiqRL7GDDw9tb/LK6UwzvLTzlSsKKcT3LI7bx0jk0s3HQxkxxCOH
FzkPwKZWUc1ZGZr9iqlpbAUWTbXx46NivmdAc61xKI0HdX72KaCI64KAMfP8CCCgn8xIKkBmv+aF
YOHAQmEQIy9G/tbeNU4rN+8FuPJAuBZLc5ZXdfrRdfv6F5USdtR2N9zF9izLNR/lZY/F8O34oKqm
+A+vezn8Yt6x4ZzkwrS8g1Y+lH6l/R5JMSZ4a8/ksKVKNwRwlbWGvsI2a+hOOqwyEqEagYJ7xTjm
FMRFa9xGr4jyumJhbOCaToImt1pV4qL6nMTbsp1JqxzHH6oEATtLrsmvCtpTnLldH+JzsghNPDCO
NXNuJ1xEX2hRCqDZzZ2LKOUVlz8FojCCpxlhBUT37JSP9v1batnEq8Lbege1GQp7C5wMq3aTfLI9
JQ+340252BOB4aF7L2pFHrpHc/yPTKKID6r4bPO4Y+a7LnoXlOBM2BL8WCeAKER52GW7XMGVcD4D
p0g0zwB2ZFa1qP3i9q76Xr897UhVOIGBccg34c59/QKrCptmLLBI33sKtdP/R07hJ9cMUbWZuZTC
y49a8b98qX+W9y6z3KQpFuFiAwpePbgrt2jh+0jYw5CH2mKnfZG6WN0tcRhRo7R1N32Wgk0GgSs8
orwVHTfum+zeCdyxWWYAIxk5dRraST5vtO9l5pHVIu/07nTkkTs4RcD0jhLBqsAoybLuoIJGdZo+
IAG3dnR3tOHRCdsG4mVJjX+HVWnk5orTPkskg64z1C0CJ+u+x0Pw1VqBNuNFeFpub6gTGlOV6yvi
X2bs0GrvaUTUs/Yy4arQMwmP1P54PgIwlWiUtsYdNYTTFoLB6BjUkMfID1YoDQpl5fop0OiAB29R
E/39h0f2HA42DrkZlPda9hot7T4KfJrZbEq/sd0gkg+OsjRUu+lj1X6Sbza5y0nfWLLs/auZCM9W
IXzOQk++TObhAO9dedUaC+xpDLJAkGfzYdszbjo3pqzW3fftAt6KZmcTYel+Kif2oUHL9VdUqoVk
gzw1gqDixXdQNrEomPQ820X5U1DlGf4NvfCdRzE2IM7OZI777bpr727ehHXhhHYIvIl5UT3ZQHgx
VY9TCMw7gORGz4B+bkLWAZX8Mb1uZSm03v22z3hdR8Nz4m96yztCSSYi5b7n3gi+4DH8qid/owSI
YrziagJJ+w0OUmnOddwrpmiAsPBsCqsZZbnKvQGQmeBHQ6UJ8CtICym2QEJNw7apFJ+mY9Okx4Yf
iaAX7XWO1R/YftBsK/yvUc0SOeWZ7eEqNhClF6O/E7DAVPuGmHol52I3zMPxFUd1JPa0V4LtAa9X
r11KRHE1ctBOC3w6Vvj4vFHdO51ug0qtsTZkZd79dpvQzEI0lA5JQJ7Ah7XZWsXBoXxNTqz1DCO0
SfysiTc9o0jHh0GA3fssIFdmibfPtcksK9GogiDUVvc8jE/7VISyUBGwaXYDiQS/6q4fR6tw3Vf6
yuVOA2OrrXso7hfo7c3GrD26oB9JQE+BSSp7H/kaX89fo1i2oo+Q0576wx5MW7JqGMviT1zyLkvd
qaM7ck8uMxoj+hYHnqMg4vxzZp/AGsTX1B7kcePOymMkqgT1ZUWKs2749EUZTQ/axEQQ2QNv2/8Q
apJeYabWVfQE1oA7ok9DCcfK/iKTZ15QPh6C844QC/9iuTP3Faq2K7afa+J8c/th5x/X/YDAtgKp
xBhCT2visMfIuZsyug7S6/h85RTYAvSapbeUf3L6SmQorP94dWnsKTYQ2HDMZcXCthQodvKDp2v1
vrP6hHlsX2CZxUSjniUFe3H+EVyZtE7tFVmxzo1bCvI5YzMBRO1OwaaaWgwNjU50b5z53jq5jNWy
owCSzBG+uqXbe0dvlLH5Xutx2Zl98fVbHC9BfphuizIH3r8OFYcFmNRQV5G2HKURJBf1MUM6u9Nk
edNCEX/AKi/IcOFY/JjwU2jQqLYjgcIDdH1cdgRwubH1aTgLaysIVOkd5GeR3lyhzuEIA6ouidqW
VCMsDJcWAzvfxQ+ZGp+JD3U3csuCiGRy0KGmk6jri063A0yFKHcovZR82aVBwKJbsgPC+ilRZnIC
M0/z0v2XUMT+PgTZbR7BMAwAszumPbHsjptn5MO9TLDimFRVP0wQs6mUk4J/im1w5ENVXvkCwLc+
rZ/tVZouSiEXmGSz28PcbqAQFKbUg4i3NblGlorw1jxUQo/33Wf8x6EiuDHWoZwC45Yvr6gD5Ygb
kt5ybfJ8WLq4wz9s2tn9Rlz5D3OC7gr3ArnhDuN2iPcTrhJq61qfj27OCmw5y3Q81V7mDlIHahgp
zx+bbX89PPzDNlUMIpbW9l4PLFEUcz2/MU7LEXMn7IUx3QDka+XPIdM7HkNVxmQ4fLegGcFqxsJg
3QSuTIUIMM1KhMdgsyyRRk2LgpGekZa4HCnjmjh1ZtWOVpeKRNh4rlJwS2+Rb2Q/g6mjnmZfFU4/
XB1E50aE8v30/fVshGAHOEZTMEyt1gfKo663VHtP47wN+4motbTQhhohyR5AaFcGynNiF7PpWIm/
GV8JdTUpZpV91EAyhS+eIBsEopKXeT5isPzRlmOCtg4S9Y/mQTgYkZHB5W06aY4BXeSKJHDXagnu
Dg67OOq/DMmK6ThNStFA3PhJ78TgKSyu7xUoGqqi9s8PtYK87hCvauFDnbRz691Ge9SCNcmL2nHC
x6gbICt2LraY1Ag7qmlAPOANP2XWCm4lJQ1b7wgcoW37DA5GHhwgoBRBG21pocKZZu3iSh7jvjgm
RtAQT7SW9PdRvCFveo3OSf9h0nqObLhk8E0/Yie6oQSLiHm+/DuZ3csqcFJuXinK8tiTKUmPbiey
9I6BdOAE/7NtWRAXW3msyIDm1fC+Q3F89oDPYcvgp/a35PYBjSm4zs/vBWcO9pQnIrqx63jZqMRK
8/XirdwhYDEkV3vzzo57RWyh+DXSy9xASDlB20vOru7oS94qqnVDx7E2wkpYVmG3zrwZw2iVwpBb
2ZU9g4ENEKPmMiXo+jMmlpap0Rs4QjPIJe+dIp8wA0/fmb8IoVrNDZLgf1US5nAeCr4PORTkZbgJ
jBCdf4tqAcBlYD3+VwOosaVfL2yIwQUXvzCL+wp397qedJ6fHSwOtuhXKNIYpx8EP25iMfKYXnvm
g6V1xTMkddbqhsNvN7KNKR/c+btA+UYsSGM2SAGgV7d27Kiu6FEtkZK+HzqlMkX3EEqx8ub0W6uA
PojQX1kf2xzt/od4HV7dBiKtx62LhXypKYXXh1vfU0AI4gYc3Ryf2nwZLt1l56zfS03Ftxkx01RA
wl5PAaGWi/D8rvM1Ohz0Vqm9mqqQzuDUUUyaxIFO0WgfiznwYq0MIP9yJG98AFqEvMgkbStAItYj
7pOqQrM1JZjm/f1SaKOx99S35iauu3HtiO5Z5k+aPR/UaEnGTOfjyoqP6dz6FfFnLPMALlI8ajKx
aALNbb4XHgyCub+jaX7wanwjfJnY71s/yCYZEbgqpclmfc8zMdWf2fVJKSWLhs18rxSBDNP/F/Cx
SR4gO8l3lA1cj8DjwO1h6jLx6wRlA6zuk8d69EsKJXqIbM+QTvDlkO8j+iSCG545bm2kLEYrrnS8
Xlc20vwpnrJk+DUZ8MHzQ4pws8cCwHBZ+E82rkCbMAIb4vevvL01w6gOWi9sMsv1YwOFBakUXvnu
lIxlvb0tS/CCE2iXqbh2O9XyBJPn1cninEaAOb94lS/s+xRBNIM2vsbZrcMJ7yVpKY796yMfjkYT
rDyTapfRZVPUGH62JqhUrFmmtdezaEnIJ2/PGD83psh2t2Qdr3LwsDonV6PvIcfdMoF4r0iIcclC
fKjmWyrhVBnkdH76FRXOL/ki9m6dp56vTntqBuunsSQnwoLTDAK7EZbLDA7Mzn0ZFIJ3F5OBsvKt
IECvVQIo9mhzUmFOLkq+NVF9kisdm0k4TptN2s6Rd11eGaFeI3tmuoyuwC6niupqp+6cM1GqfYO3
SpzJB0ss8JygnmIJfJuYbyvFMgYkA3xMHqebak8yrz1z5qH61EF7hpiLo8ccYRVPXuB/7xRN11cs
1H00LRTkbgpnA0dlT7dX9lu30/U9gc7PzKCgUuUkMWroti6m7izQHwOlFb+d58I9hsgD+mDHqeUJ
/KoU42FQ4jrQzA0NtItQDjdc35jvCPqUeD2AGTqiCiokTGA7xcb7DH5fPoWWJlVLY97yvOvsQGCm
PJiXcNAIZ/WLUjd4pEwgdyuNNeBc0pjqKJgnnSFxnJStgYmacxvT6HXuMdEyorr9P3uTL9Kr9Nl7
4oFhHzfYAxdZafRyOkEbv7KeF+7yMHUDt7mfLUT626FOl1X/RC2vVie3l5s1KSRdkN2FnaRh+07B
QRjY4cbgM1tS2fy/wVX6u7Z6s921zTyEsuPgxovqEtHZ+1JV7Nz3MOvA5OVXik5LcewQOluk5n4r
zgeEgtatvKwMfktxu+Csgl3NwSo4Yp20PNwtBvWshAYJI5sGj73XYMDr/vJ+pJeCGylKmufSDRWc
3I83uKjkvQdB9sd8sc38E2vl2iLkvgjqMq/uaG6kJssrvNQl9j96FSl6danGjj0Ofssg4rZ00Hrg
ol3mPAgUx8y8/VmUOVbDhClBCPlD2KDdzIsYR6HHYAtb3No9tFP1mV+KAg9gTsczmXhex95KY5cF
foT1eAStzyaRvzk+kkf9oTK3QZADVgulq192buJ+WXJptkqa3nPLF+bvB1ACMQfUU/Hi6tf/8Dbe
iTeqiR+kXv8AwLuExqA6xlZu65ddXVBS2d/atCOIsHOF6arK7FPZsfkxfQ4UQIIDB+Pht+f5rIjm
bX7mEuWyw3vkwRhZ+uggPbKYF1zbrlvs+CfvwCUf2eGI3gTppla/kl5wM8p8JCNPmkGAh3t/C2G8
3f11JICD90WNjIyWypXMbaZUathX9vs59HzV5o4CHOmMibagWGLyR5J4Kz594lGGbJdtbGiMyR7a
hPRGpzfQ6s4twdAzVKp/4HeIIGffkpQC3lp7BtI+fkNX/0PBslFEkVT/13TAs45kuduu9ripbgNe
hL1QnGi9EZMdXKsDBsrNzplHoPjLTobajvXZz2Iu/zBHsbZTHLqppIWnv/yphGj4ipltCai70LLp
cUAwSCiYMId1Pzr4QM4kYzs0zcbpatKHO/1w3T/FcDJ9BRf6E9otSYnqU+KxeX8cjY1AbrJ7tEgX
XnT4cMBcNMuO+cngVgtoJDDnN/NO49zdo2cokPdzYCfyPqdlXOyGJReazr83PEPKTYeOEy8CUQpN
voYzuvoualFPS9uvG/mtRmQgBTxh7AfbXrwtFL36zYVoe9Tqwq05IhDEoVfKaRajE7KodvLQP8iJ
b9UYG9DE0Ngg/x4G9MPClSfIvK8EXGE9K1JsM86dq+4F+9659S9amPW3+A/2stREZQKweXGpxOek
U/E7IULmj4nGK/5q+0v2BquJr1ygPI13n52auVnHZnQx/A7CLpALLWufA15bJVnyLbdOI4VKDHVL
S6pJaEfwAFU9mitNliQK0vfj1esxAU2QffaIsxVUZEXkmnpVic6zODzxzANOdUn4elQQqN1fOK5P
E4Zqn5ZThZVhuHaILARAZvR/fxSeIIF446KD2PbwFOCCgaOFOdwo0/2TNKxN9mZlZyAavF3ZZKH4
19+DnnZg5B9shCKKb0qkoR0xAsW7BaazxCYCbT9pfbExArTCAd9IxAnaeomiEqTUrOA5a7yJjryq
+nTIw5rmdM3Rt9CQiqY3QK1GOeIe6Fsn+5qCUeTP4nlfpfLeMCStMtmqLM/vSYqBt+wxFVUoChAo
mXAiJlq8xa5klkoF4kcZHogyRZFYqujTOpvi+YqJcAPB6XZbk870qMjGbgtjgc1zelL6qmccTiK2
LPZmONP9+qQInZvdBQ5AXoLF42UnK6fA81rWoQ39khoCkxQVh+d0KOlTnBEM9dwvZ3lrYluYKjJe
vBd/jtCjw6kSQHBF6oVZVleeZdlGCIPehIGrMWT3cvLu88zpwsReauOqpaXftjepmrWLN88gDkLR
hLJ+xU4RTEDccCtyaVs/bHXx5mZ3B2EKLSDFDvmq1QArI67pB3B1wg8oUj0Eeqx3aNWr+yanAXg7
yemeH+NWExM5FAf1CYlABYsIJ3j6cRnNXzfTN2C71q4wTni9topJx1hyL0bNwcj1gKSRf3lREub9
vndNX702Opwv0e1QYWuCPuxt7rE7xurxNP68WKRR9NyshoPyefvqjufvCSM4xND/fmS7OxKMLz7e
gmVotvAaD8HuOe58c8YoCYkg14Xmf80W0KvvTo0GaN884p3ex5H0NbKjzGzZBZUpQQ+ZqMqdKHPA
WWh6c+ZC0wIYmRunY9XTiGPqFLxpdvIlLlxKSCOF/CC7hh/PISG2HRNTVcYTsjw51H/qcpqJqFbw
6rXs5Yg6rQK/pXEyzXYEf21obNhxJxxuTFyQoQp+PYBaaHHLRbANtn7PHe2wAiHfmlM7MNyeQTkp
7RodfuoqkVFWn27eBWpUY9efN18CAteljfp02VM8/Mpax1syw1DriLpzX0C1Jup/PqN0gv5xPbrJ
22MME+fT/yGMo6/qVZuKQIyHH5hjbsRk+Fsv4hNl9dLEXYoT9Tdib95hNn4gmEDaM6/SS3C0ER6I
yJWa6IAptva1SfKBCvQBNMpvTYNA3PFx9fSudsVPZd4EtZDfZfl/4oo1ll2v4WhLhH3kiADlE+ZQ
meMw8/PwsiFYk6DMEmSUdO/3GGFALyzmX+EANrxOa0mhwXPvMA0KCfN95OEEcWusydc2pQXQ+bWs
nwKezEZhWEBEUTkaItMLmE1jYhjI90WgC++UbrIn8BVVwJYb/KTUjyLc7+tk59idajkUw/yYquGQ
mmTblKkULpolKSsDWs0YQcrcuWyfxzAxYcDUa36DXC1s5Jd9HV9uidMRSBnU5+2yB1Ads1Dz8OQV
omngvyPOcIiz/EdzzQnCIGIuN92LfJXb1FKROTebPWdKILqgKTRuhiPknJk70TbtQCmangd7rncF
z3o2OM8lXwWVyEFaxJ7qsbUhHQknnZsEK/Ji++2SlX6HnpSGhtUcsPbTV9JdbwzimhIs1588Av1p
BeoEO9rj6V9KtsR2BGIt01bcWmaQ1jsc8kYFxDB5TDGXkxX2rxNPbNfCs5f0OvvxhuwOQVlqwBjM
BWx3YMiAmBkwES76RdR/sh4CKf01RjhPRmxTM5uMrTMmLiGOWf3nGcyTT2/tMweGIJ4x0o0XV/nx
PId91EJ09d/FAvYS/PW6eAn920iNR/OwVNqpsf4FgLd/VPzhbsY57O81XcFOi6Lx00YDIwbn9e/j
gcFTSMBYCZhIKruIGSehWfoBbD6XOL93hjno3zKcIUw6+zp1Xt+sGFcsabgL6vc1fjmWbkORsGKD
wk3c0X7TO/GeRLgTSNtdanENv7oNW5chBgO9K4jxke2kxeg2ggsVhvtw6Wu5vbBrYVHXwAepsDN4
V+kJfXv94nKi9+/QMRgMPJqABuSVcKRf6kIKdQn7JDWz7uWe6G4EUQKNn4PmBC3QZcO5qJBlhldd
laXESv0Ata86bZ3A8JdI9Yu43yQuTyWuW5nVf67oXFTa+xsHSbsktjeZCUu+omUIdBaOp+rdcAMx
LmNQy8sxEtvjiPao5IjSIAssuE8fyPOBzKuodWhzKzsnWqYTsibJ+yL3RnY2gG5cftEkbvk3jox0
MSB6QWgvHXessxxayl93BAetIOMqUfNekpefUBeFqXPl2dasHtCGnoWXpZbhstuifKHwEjJgwUE7
Akes+wO4SGrl99aGtZnF8S/r9C4S2iOcj3bDnNDcOEdT3l3YKqsxI6ipFGwgrAx1LpOWvijF6a5P
ydEYW18CeC8Alr36HCgAYgoYVJd7kOdDX4GjQpAX52BlitPap4H/7UmAa8yckVCAOAsHN7XlOvFL
OtgDMJpn90UfNr4ABlFfgdw2UJ1K/TrkSPgsqLlrdaB1stCsRmi+Haw1ZTOTjzWSzgKbZveg60FN
Nt1XgEr+a4YjAFMrzLzIBRLrwHX9Voxo4k9l2wFNNQun9XQj0kcG9Q3e5ogLa1fnhmY05daz7KY4
pNFOKR+vgojBPBOlalNAzYJipNuf3Dry1qeTXU0t/vh9I9FCWfG/40znIoLNvnHJfUeOhUWTUyQu
R5nklgX9P7idwkb8xa0H9zEO/8zGm/tYhx1H6Xs1ok4RUq4P3Gt5w+S6TkX2mef8frfH38nwSIE+
AWaFAy+oXXS5cwfz5VXaKrFOgomzz1zx+2ZJhUvQRbJagNns19DnqAOiV7hIehrmLJm3/vcDTmcB
kKQWhXqjFf9X7EF/7J3ZecUDilDSYvJpTyf79hC0CwaHbMjuvEF7J2igX++daTc/fYiLa6WLqcBP
hjTWScYD5BzkKYBnevqsmkt47+EUOTkkKlfEf3J8zGIl/NUnKf1R285G91BgxP43DjoKDg52OSDE
9tTm4wTn4sMW65UXMHyL1FZ5UGZwbZN2GiAeisxfQtX9xSSYNOO4F7503piC/duY2ddkQypNy+PB
CMRS8BXdCq5zexjT83i9n61dfC2XC9q2CGGLDmPc7dX4EXCewi96S5Q1M2ApMx0y/a9tjqhx02Bo
ALTlaoLmVEG/b8VgiWCRmwUc2XOWoE3K0WHxcrcJJNgomrlqE8zrV2Cb9BtqVvLIG56I7dpeLh0z
EC/3S9V0I++ND+Riru/efn56NpDRd81kFHAJ5YHliHudu5r/Q24dl7XPcGyvNTdbDHBD7XO4L9cZ
l1S9tehMXXTiViHnqI3vHFHfZO8J7yx2N2DHhaYB8J2JoQKIBTR940wBCo8avss9EC/GZwme+trW
I2GmGTn4NxbYGRYqNEL5f0KE3FsljeB020a7oUw/DSwbM2tr7oa/jyV227ZEgCm/DNxiy42QP0na
q5Mr4uOlRGkp6yeE06Zoc7fSdsJS3Dtdghe3ZpSp2Bwyu6JdkbIlZNQ08GKSDxWtDqgnwdM/5BoF
qWyFMxRYLt01K8qhPyyW57thE7ya4pDKqiGkVYRGOgim5Vj21dJi46/m5nPWBcxFjF/RPMmnNJZP
gYqDFkSwONYmchsb8bGFrEghbUVHrQ6KGYL1btFthcLRE9hNYibqoYR2ICZXz6W+lbVdVcRH6X5A
bdcSKAGJ/TUe8+afdCA+iWZYGWNitn0MLFDjF5R0AKDeN9mIMDFIiLGnK5Z6ktRkTPx0BjpjtSz0
YvD2ROmD1A8TdtECcyrn8/QXDBKv18Wbk3map3tmRc/pd1GQKhzEXfEd/AraGLL0tjRFJBjZEPen
fE5iELiJH/XmTFEqYHP3agEdLMXJKQCS5064a1gW7aXPcY6pjW+GqhUz24H3Wek2/CszQ16P0As7
5O8KBIzX36moM15cCpVdM19izW7Ea0b+gC2hoBA2DfGi/tm7Fmflw8/ea4rOsObHpTthGZ5q+x2e
eLaalVOTnpZJ7NaxL7T4UI0Z5K4gyRF83JNelAHUHfD6i9AvaBVG0Zs4pE/8KDD0j/jPS5V/hxtb
a9NTKk9qYxbGqCjMJ9WI7gm2curYIbaxQVYbIaoCEAtUmpZAlw37KV6zeL34PFJk1IW2LonKZSXB
JXFQD4ui5jnAPYfIRDJsw6QDKsup4rutt/JnNdat7eVjsU/hMX54esGZPNXv+yl42YmLbu5h5Gyh
VXmRBru6Bh4Q27Be4WiFZeiWqXdybUzTgv7fgzA6jgqP8fcJb7dZnbjGyo6Q12nY0XuJn0TeAgKe
bGm8vYJEu1VCA+0Br4mI3zCcQgHdJWiif4hkgb+Z59CmAShKdTAUwVhTWdWw2bK7QxvY8YeotGxr
+kDIGuGyJ1oLiFpw4XydyDI3ZPlq23uegNMV4WVbEfn94ChSjzlFNqxfR0Ce4xXhJlDxm8C8VB5w
E2ARQLA9F/faaD9Zgq1Sqf1YU/BKGq0s4OA69SJ8dA5tUBXcHrWnbBdBP0Obbl993bNjQAtPYJ9u
pUkLLY1qmamkqb/LYNhPKuk03TmgIG3g3RG0YYNnIIL/+5K3qZZCiylvVzOcEteBb1tmwvC/5a+G
8yj1U8Md5gLMM4MBKwoUlO/K4BashPYnRqAENJiH0RKIaeaDz1zqEU8bMZgGyu5nZQZMsnNhJr6/
f3hjUSM7WbU9w1KWkHxlQSN5vkKGiOc/uO3Fgcyf70bxI9FEgH1JXrkSS7EKBNtVQ0eTT8gCYj/8
5wkhm+moeu4+DB+WiykUcG6HUBTIKbHvyA7z5pZpQWejdbNgEDq9OYJVOM2ZTfg+zuIE2NESrZjn
AilY5gC12LcWJ+sBUhHsnDOARb250g8U2fMuztceR4IDGXvWCahInllLkVf5xMTrOVjLnmhz/hZX
2GCf67NquKcgD4eElHuTwyBtopQP1RIEVHvw9yyCI9JKAqjgdJgRbBitufLydzTuf2qOdUrWrrm1
0e+wgv1nojCuuP81hxEjOAGU3NqeN/6TrtI4KKWwfPbzNUGzrW31574RwWRLc80ZDfbw3Gw7ih7A
tDqQbw11Y4EkQhReIbtHU+76njk9HHeQIRcAOegeXtk7OvxKVwwPIsfmiW9TKDEQHdbl0s4n4P2W
KppvhNxtaVtihLLaM098qRi1NYhS/aw3TmSSPKJzCDKaKdgT5lquwOkIT+Jj1xhuOJQvf6j9Zkpv
V42JMLpk+2OH0IoU9LElCOalTQZMgLlGpeSbgTci4BURzQ3E4zzuLE4g+x3ZZJ/7FcsL0JIeRoQo
K84z4An34NCUwMcclY4C4DsTE5FgdQo9UEKF3650uk7JK38nk6vwthlV0DfCDsr6+QK7TR58r0V8
UFmpI6+EUEtDlgKGoUX433RmQII2YV1gGt4hR1aSNkdWGlkfylTW0k3JVuZ9ydZpNlq0Eoh2StKB
AI/+juNWzDLo1wrvzavPO12P6CoAvBgT2gSJ9NbNYK7AYVkm+6elNPMMI4/47besDjntaQO+GInY
soQoExs7fjTJ+tLfGHMbMo6UouxtaHDX9USbj1Vl5Q1MKVo3lpJpR5zU9+pazi3GXmTYCasbLwru
FmqCOMF+I8MsRrQdq04cMuBvhZ/J+Px2GvkP5dh7Voa2EmZNLnsQmc4RmKwHg/c7Ej/eR/ItYnwa
2Z+O1C7brYskNMCwbjlm8KZPRiQjfT8xnN2E1MeYKQktzknpEWUBS01LNiCxvxZBnwX26mClQWd4
G0AxVtIgWLISPV+0pLRKgd+ru8JXA4wB/3QSV1lYu11tclRycD1/K3sU9of9brXE7HwTy8sdF4V3
9dlKdk0uvG8uRC9ED4UTJO+ccTCJqDVq6HPPYAPWr5Rj2yLjfC/r9DMhJ8CpPgdUkZza8JiVNBWK
FSzwDX/8joPE683IrYShtGhy0WM3cKs5gX5CokWzHc9czQ+UWv/IofKhnCEpUt3zr0tv+g9jI6Eo
b9NXC5HjTkNEwFo+gyoBuJZgKHW+o0cXqWZM52RquZdxCKYUFb1Uc53lURYPjVQxSD5/fp3KPNcH
x2lXPuKhJ6JYJ83uG6Lpf/p5y7u4gBfKCkvJB4tJ5eXT/w6gqohAP8l+QNFwS22fkOvAComQ9fO4
WkPMduhZWRCjZ51shwViQ9lFxqecbrvvNhwC7uVh+vhuckFAQQyuAR8dgPxwgDqOcVP6T0PgRsMQ
D3dfQwQJ1U9GcpncDt5bt7glZaet9EcAmu+yHuDsIC/qRV1CZPgh8XhOfxNV71TXWe06XCSdK1I6
eZOGcevFIU1BUL3g93Yz9pjd5F0R+MlyPAK5TByQ9HfdL6su2JTDFTt1yo6TYDl2a5l+qCA8FEwT
q6moR3uVOMKlmbj/UVKF6B5aLvVPwdo5elF3ToVbSNDyTugasfdAyqhLJmTNkTcq2fJ2EAXlZsDx
R+iYG3uInQUhl9QSEZy1K5rlSwsZzPKA41vIJ6SkY8B3jhjTuDyFfaewqnjK1yRUmPXjWSdxHV0K
84p27AtUrBalsEvVkCGwNoH2mDNanqb8+bz6kHVFnNN7uS7gpfFu309JErYLltLowQ39aJauKCnU
zi2AcbXpNUV6eM+rGzEKhIhgExsx5/wf/YBczfE+2Ax6pB7/DxpG9fFEGfhX+eKANdPQU5bwLdiU
XiaD9TNPgfDD8X4Gg7Rya37StzGcCRADUewTvO6yzkJVs9mLOxj6cxMFLzD9lXHb+mr30kvn38b9
IcQicq0Y1ydUvSadt8dWPMvANwB4pkqoPZvs2jsDaXbmyIx68kUt85y4xAp4xEoh2EtoPbuR/LDM
IIMFK88pQ/Ma5rHlUeq/EYQ9QUmAHAcUW2y4wgD/MgsNKnJC2Mly6xcNcoK40gmbsPogenToTqLk
QVQnvnE0N5XPnKimFbEIOrqsk00bR6o2moUXYmY4CBWAJ1JYZSkyJdKQN9+fvnYxF5uJqaiNjjaL
sr043UNMo4c/MdVBuzwD2XJUnjc6kwMq0etgWjndUffJgyifx0Ksh/IFZNNIJ1tIltr0cWDXnpS1
6Op3DzNZQ6oECt69SkcmxDjNa/9apaFMXQHDCsACyzFR9guz5CLxSvPiGq/lCDwFWYh0i55eBKXf
OvOkHs1FAi8NlfC/XHvSFEJsmPAXIlQsyt5FGbu4wq1lFljzTidHeu8spiSHEgohfdTZU7mWsFo8
Odcz8LfVHSq3I5E4Um6cbbs4Sx7BbtAgfNjHTmBxyogvUKZwmeIX/iOLal2K9LZ4WM9+tv7hN3ra
iBdCTnB0z4jPZkr/zB8IAxNE9nsyfp0bpcJuip3ZZmqcrEJR49atUgjIUE2ffKgdRejB1JhIO55x
Zv8Wd+RJdISz+e/MSFbzeBW/E3mdndLhzg4UMIzYk0MOyovGmPiyS/PkHnniL7QXgMlADSGqtusH
PKZVefAzEyS9Vj8nPAG7IpEkbcnedS2Q5DyJOnPPYZPVrS1LBUP1hNNtGUThom3wXP9HYbHE+ERO
HMGT6ZH6lVc/6Vy4PXewmg3hAGhVvWNkUmJ4Ar0Ze5Telj99UgZsMM9Jd5iL1YGQFLHhv19prXkF
5/L/nuipYBfkIrMqLx0i+SZnGiZQzxfQv5XZqOalGzv/y6BLIkI3RpaoYb1qc6PIxdtmeFU713v/
3GKPYmTcM7ORri81OBzNp4Lcbwgin3R04JFZIPwAxOjWPxf0c7t0kHAUjx2gu+DEpxJd8xXok3aP
d8Lmmoz5AC4gs2qKm34NSx1fBvkZ/XFl7UX8kuFkam0tdSyTW9QBCDNPGZBNEqTFGtEcs3oSBP7q
OLrioJri9HubqTBO8EL7VyPCp83O6TEA3Ab8gXEBy55dFmZfP6rsRPw6w+fZas4MzLpeguN6SERV
uRduIRGsTkYwUVd5dvvNnMVXc2Hy/kKXfaDw844ynKjWk+szO9Zhn4E0L/mGRJvHTzDeWQnbJ+ix
YBdSdDV8Z0j0aS+8dRHZp1kQbWTPoLM9Ca0PMnSX0/bjng6AZ5LhoZYYExLoyUun4zancfE9KoI5
QGFUAs9ctjcjjRH9JfGkO/8DQFCLr672lS3wpv3BgrYsoXSIdZyMa95Vh9Bsma13vSyv5f5xlncv
/2Tx67d191ZtYNzK2+T83UYR6Q/3qO1hgLPXU7yo/RPY5UmWa8bhXNqaVbP75SAVsr9lirOUAtaz
myTXIsH9OmDF/yd0b7G25LBInFnyKy/hzXqHebH/zGZDuLITTjbVNAt6Bz7kCkw2HSm+uxxog9CG
KcjWlVnYuQvCYqTmI79A/w0YiWocc2hv/hyAtV+7pzUSqknDAsSqA3ZeCzKZRYL2UPNjWTjMlHWr
fexbki1fXtsS6qjkoYoe6MGIZ02L/q8+Ktei/Z9ulseBEzMmugH1BWdzdlixUp0bUCcfF898qh0r
eFhskGy/RRVooAYTyIonE6C9df2KGe4Zy6dVZ0tjuNMDXYgsgQggMK2EIOFYhKL/S5MLpda7Ckxb
LMkcnjDJP079d5O7Wwd7KBe1WYlFCAdTv8cDvDkxPF+R8FxOnUpYvSSgUdfeJM9gdgIYFwpsU5ZT
7LCWbYbl21ZBfz1EiFPx+3aAqoqI6BOrajb3CAtQk3l6QgwLFTVf9hvBYc0mtz/DtdFvMvNIxrP9
B4F/xqzqCbixB7IIpi17uhIt+3hR9XSvMX5qBvtTAsph1kaEsaTKobzI/i5L2/tPeRjOy/HsRTcu
bfK7CZuAvBVMmsaYz5F1pu6GDftJyeNITmkKix96opQcj05sZt0Dn0xqf8Hu1TlVugYX2hZE0waG
AClSHNsNpU2bTJ6GCoFVvHge81/hffIu8hjrsmawja/zCAYX/I9OY9egcByi7fvltwFeCRiIm3Ms
to28684eXLXq95sH1QuP1mK7mkhykGt/EGUaXR5GxeX0508WGzzc4yjdHgjcM0q03mibrU+/LDZA
rPX6NeT3WMpkg8PcNe/zGMkIoiwjKLjslzlSHGUyuRjY8FGrXS2B4SbVTDTQO15xlO6gCaQ1q+N+
7qH0J9NxiJAoc9GEwXM7Ey1mrZp4nVtaK1CvwOoJZO2vKy0F0/QnV/KSHOuTbYeZQubPPujKGJ0f
YZRglNUXqZbHSU53818qqZ4rrANpVZoUUS4q8mxjB0/5zIQ/+QVIWx1AOAKJUIKUidHVpP51MVTz
VE18ueiQQjlkClI9RmfvjbgL1ck6qXdjSp40FzmH5GxdmsYEsPKsEdMFyHZueffhLb6gmTvRncAU
VR0jaJ8i7+59dSmPnW/2gE8OsPDYSvCAHfYlHSHZnVA95kQFxa14g3B+gsh+OCGjkwfanYB++HdM
A0Fd3YfugkqsYIJThxgxBbGtqgk9fpdyLhjeLuv5W514AeaNbqX2W9nURhefpB0+ka6n0UpNAKFY
XSNfhMTloNDH1p+gGXASJC1IZiRX66POpmoHTTRPOF/Hdc2DsH16T2dXGIIIDBvcMwOE6nSpeu/r
4QXFoJmmaEDVDRDWMSTGFGo97ZahfuBxShvkd39Uifc+UVEZjJEEhHhTGVj6OGRlSgD3tWx6dWTf
ZpnH2wyimTYT+A/IF/VFFM+zbXKIE/uN5r+QZ2e9hpLKrWH9Phv0/TtSxDgutcDKy+dgimLW4K5U
uRV+bxp22hA8vziLJlZ8b6Hx0IxLyVvVhurJRHMePvnmWgY25XdgBa+VhFAyT35Dd7saS0sxNf6k
FQwROhfgC9VFUHRrj9BwuTovgPAO76ZlBdPAPrfV1m/jsYb5UwdxJcxr6/whiLfSpaw9c25oGbFD
IedBLd5gQ3JXx9FVen7X2g4QHtdu9sQowYjvL142pdqrr1aC76w+Kv7zZWrohGgVz2T2yd6/PVcA
z0xJrdhobqnxvBv3bzLgdmpoh7GFDHORH0xe+pk9hG1mq6t9yege9KFXeNBfACpAwwNGqiDQp+EU
QXrrFpQAtPJtKD7zeBrImhtXPTSccRll5yYmPB0jLyeKHVwKWXOMVWTCEbGlYGyTvmdFxg2WthoR
489CBTeMMA0cbvaDKiS2sFYN5eVf/lFVGXdltnzed71K6ypMNOJ5B2tfC10+F7bgsJ+voxAOwDoC
HT+nEYnToQGFYoMGjhGovO4NRb4euDTpDhp0WtH8docxop7eOCh/+JT2AWP33XOmC6vJqtGdvGo3
TnUqiVan6RwQQnqn8aY2xs9gA9yoz+ecxGsXwm9pe9o2FaEZOg3nHc9FoJO9Euoai9JpWZqamyIN
++F8JqgnQVwZh8ZzXp+nlhZ2Ql8mZ4+4wi+zNAVEYUmI45D6bSFud4jJ+FzPSXdppz/O3v+QTzWQ
CFtAobk61kiM/VidGnucEBqO09Mfj9rMnRppn+o9T+F5bHUpPDdftjT/7qJ0Qadf6vZ37j/z9Yhm
CsrEzQkH8wpKDwEhNXRANmLun27GMWvain7AbpfikIX7vubVJF8c/+aJgsFi3oe+e6GnkkfJIgzM
VqnFbyfSvLwvBfEXVNP1sRJI8ucUZ+3Ku3isj+6O2Jy8LiYH33s/Hoh8/F6sx15J1N/iKV57cYyf
xJ9sP+vxDPdf0Pz5yxXIAUAsRzv8VTioO8aXyMFHWcHyfcYJ4dldIn3exHvaU/IVn5p3JMVlA1I2
c8jPa4AOujxf/wxiNsHTq64x8/pX5RFTPWbn/8v1xQ8CrKE36sBtHc2qoKwbQDigqc9hbvs1TWVK
4qoRNHJlxQkmNSPLvAVK1PSdqDGO2Odho1CssL7kzF3Y648Tq+vp+3eJohV0ybD5f+nSDKpSXvLJ
OgZdpMY1BU15+xMrbaRY/1R4LW+xXQTB/GPNZSzldED8g+rEhpzXa2rDcj5OFJvqiuxcj27PPdA/
Ka44NrZ/nrxQMHetGHkoLbw5v+/1dOyIeXs+vnGPnQCY0d4KYrVDns9OvS1m/iLHqscsuLMUG5eX
Lp8KumyvMCUQ8wxf7VPlCY/E+zVdE5YySg1F4saHqhw0NVfWCK1SUibBbF5OwzBtvQTXFwTxCNIs
6T2hOPxjz6ecmR9fW6Gtf1VHVwESmneORGlGZkKfGkXk8Wvsi9ULhVhvhXSWmedmA640uJ5T5oZy
SqERg1bWbGWWPLC+RcREnGPJtrtW0GermtGTKBQXyLF7u55z5JHuDfppl0i3ODg+jBSdCEgIuLs4
OLxwNDKo8ZXllg/bDP8aisID+5xULABcBt3LZ4O4B1QlwXpNGXmULSqztgtRVIfoKoVMl18WUzrz
TRfLAbpjUJnMsmyQXn9464UxWlmpJT9UR7h91wvLPKWCt6T1cFN+Vx1XM0H/TZYQbOU9cNGSKg6s
8IGw5ujoJ2qsUn6gCNMFhejdMMjSdNxwp3uOemBWTobFkTlP65rz1AvdSiwkxu8bcirUw9Y0IGsS
nsk2wOVByZYFGI7ovmS4pgu3Gf6POOBCuwO1+Eer3SM0nQfuMZ7Ta8GENiekepHYJzp2Uv/L+NIK
N3ZCz+zRJl3ZPTEW06Ojbvj+MFbs3aLeDeWBUv32OKZdzaCgVwQegyJD2HGTUNutya2FX6IJ3vt9
9g4jtVX9INmL3SR7uHT6F8HqlOI0fryUKfxlgG5RBzvvVpoShvlsd/7kIIHoyW949efNOFPXGV+y
asiXp3LAxDQBiG6t63tK8m8zBj0TuSGXS0o+bcAliXI2EopMfIVDxvGsrCL0Q2Cpg0GhuyWOKAKk
4Llo+YK0rVVPjLwN0qreO0f+8l54XSaZZzHlh/XyTsGfLnxoTnxnStotorBv/No8VJSBplDKxBqU
L+HvjW5mEVzECf/uorrVXQ85rWX4Fh26QcZc0X4biUj5/46OKpHU0/X9jilEZpOccHZcMw7KTARQ
iAgkyAB42bn9ZO9nGHXA+cHGy3xlAYUOGG0xMhZxpOajMfXJXeD/CzO7ir0OD+hxmeYrjh/n02W8
UW7Ec76iVDyY0pGRYrrcwViMhKi0wr52feu5ZuNtyDCVhub+Hfnvxqyanvsvrnpsld0ybam8Vapj
lxQLbdnuXdVjF5vpqBFVGxYAi+zNq6pOEt+xPkleSRL5/eSV6Quk0TpMzvP570MIspP34k8oxCyL
Z7kd5xcFcL1/O+7VNm4WEogXRJ3Akxl9CdMAp1ZLvZoE/YHU4aYmlHp+kUcehPi236z4iwM/sAP+
GYT1Kvl5WzzwhSbzk3TqhAcofJV/CxnPfzfGKB2wCDPmJD/J+Nt1Z8A00a3FQgtcwd+YOhz9JluJ
2ZWnYLpKzynB51aQWWv37AEoT1ZHVX9XJhvuDqvU5MbkHb68LBvQ2NJVUqfKoYoj5XQM/Xf3odWz
kwJYFo3Nyt9dhfhUMvRMeeJwrqfoxZvaCjRL1IULPuuC5ctBWI2ISg91iSFUvPHWa2RfimT3sUVk
1il6jd/vs6ezixZhFbvDKM0PqUkYGqQMvoMBcTR8hPdcDw3YM2jwfG1N2IWt4Nv5Hdq9V753LFsb
5kFW5sjvhsgLblBrYcNILe01YMKRLWw63vyp65q0izCVez8NcR90QCN6zBD4pPKNbzevg0vkpF+s
wCXWNw9SF/p91Fk1Qsy8ROk3uTIRV/BCGeGR3N/aHOuKSf7ftBXkisoJ4cMtuEv3cABwIxzy34xg
iKRbK5SSnXJFGPlyR7aJNyyWvLSe8m5a9b3d7fDL1xibtvvntTqtd6Qcq36GPMdVxkZ170UFDCWW
TyfTKfTeVs5HjYy7kSOwIQI0RCUCLyPWRrG690LhBI6r+vsa61P/yPGz6nlHOwxfyHixEJdkvxGX
8TL1NN1vocYkWeQQPWEVXajptstNBINHEs2q4lW43rUxEraexggPwH4aHsAu7GWoCB5pUcXt1U/B
vSFMpFAucBdPV/KZRs0P1tL/i5WOzMLbg2r6qPdTlQZOOGylL5qM3SOim6ETRsNNP8P921P6aD4Q
ervsxJS/PUIzudIUXh97zcSJ6+JV1bXzQWsELTnyDUxh8T4LdoeeqWRYZmYqa05t54EyXU9Wl1rs
22Wb/41Hxh+Tpm0JUYYoZVWJYyfkWAGyXEF/l6nBQjq9ootP6QtRfebKKwSq/YvqIEmWCqmUuuo2
jBLGWkLEiFqjLb8mpS56asDfAvVI2f0s8us7wSLkr1Qr4gWoNHA/qdcf0XuSsq3RoBxg91sDaBHx
C5SSX90lDpzZKGyIngu33LgHehCtU7/PrNzCi7yXA+X1ntC/FErML/lf2isBEDCc6btbfO+vxMlV
tmfncVFcJy4u21Bc/MJ5w7ZPVY2RSXf7QrZB+8IbxtRdOvBiECpZlfXYFbnPeSN1aesrZ1WyzaEd
B7aFH3RCYdlXZMh6RAbdGAJQoibQgkS4oXwN5GYJF3o/Zu8gwjSHxYl5+BqFbOxgnqRKps17d6I3
ZNx41A9BquH5z0kzH1yA0G/v3y41wAUjoUoQDMRso7kGoDJ1kMLNV9v4efNEMROhHIM70dipEeC9
7CVcw8R4zNC1S0HqhTSjvdowpTNjRt+6bd/MjqebnXW9H6ZMzQQhUGKFI9UH2J40yHYCKYMZYHZa
v0qcZPvWaVMpY8gXPH3C/zRzfp8wJHNc919XWf2UH+R20PczLoXh+p40UuciqS5f+2BlHbjy6tS2
bWsmvHSQEnP/HrfkKAcv28n9a0T7vY728JsW36r/HHJkvQ/VKxxtniP3hvqyaMq5wWAGPQ/rPZ7l
ow14nJ9YNqRVQB5FIbatrdoqVvwxLOPyLk3CylNabvnZsWtBoqRjiRw29ZR5lV8QibVU+wnBh0Td
8csl9iZV/NSE8H1JkCeTIsWFXd35OjSQcmu+qkjpGoU3lXjWPHkAjssYRzTyeyBxGcGLdP9ev4gx
PZ58awNRHstFep/JrvDmptZYNSTl7MdLcDPn+zVm2zMVF+j6fVqcqXsqb5W3uOFCjmJNFdmzCQGc
CINjioaV9+v2zFayysRSJe6yaIX9+W6zft2xivdL+SvJk62bu1Z7LZC6NYnj3/pzRxKPTQZbxbCR
oKEURAIGCvvGpaJpt4nx30CMzAVYoa4KKxPdL2MTkGAI5jMhryd/F7GSrTesjoPzx4yvo5I7L2aY
MhlZecFP4rEuUegyG5giJ0NbYXiG9L8f26FYm5IL7TbGHwPv6BWANO+Z5iqUmQpzWUhOgCrvUB11
RJEuPdoDjXNvQnRga44HSDWxO1gILr4lVdUsC9xMp0rWITsIRAHxOyjUXduvHu+7EzivOwnWbX4s
t0JWagzLbNQPCLBM8u/So9mDgAWoB7jCHOKWy6kOPIyXOEVwXx98CVyNP1M6QDBjinQAbOnvEAzG
fYUm7gUIwIGA8nWeC5gkCEMdjlLqepbXezChyqYfnkYvRgj/1DEWwRmFU43lxVdqnDpdxUUDjSTN
QzXJSFSDCrH2LRcRs7g4ksOioEaKIiCjS2NYxKkDxoKV8BejgauAPWanr+Akufd7yJA3KNlJ9WLD
OKQJH8S7BUXkwIOt9NOCTj+UW1R5LU92E3VMTw71j7CeG6r+oSI1h6gY8LtXh9WsoiydPc9YmTMY
EoFeXuNZaCaWrijpLUlWq0grbfWyAxG/Kz0VrLB/hcjNt4ZtpTIw9vfk4BKLfCdnAUcSRYZo8Azr
53pABYRjw+8iyIaZryQgx6/OIJtaccKs3zMe8l1B0VKmTQGGKIbwgvlhV0kXYVEpdN4Xxdh8nbkS
l8U6nOIXqLRa2vwUj/G9vFy2U1YuJx+APwgWRP/THi0aW/HM9vuWqZ1fukCrrersP9jlzQvz0iOY
FDWRDuD23W/4YhxITfCIL2VpjXZEfsNHlAJbUUe18MVtd1u7RPi+PMsgcIBrSzGoXzIQBnvgHfaL
tUUFn7prpaUIsbwjW8a7QxLovp51TQaWNwNsvtvX7CW9XNSIKt6B9r1gISk/hjQgA7RPPiLSVGFL
iLicoofhMhQqPD8/G3YurnMsVMLht0ipfCTtLLm7a13QAB0kmN65EmG7E9F7+k66N/sjodzFxmAh
ST2WnZE2j9bVVttfrXjm/02Ntte7HaSpm3F1UKkmCWEZQO0DUQhBT7ptCOeswOV6OHFS0XL7Gn0V
KCACK+XYj5S/TUWT6uBvGW+LxHbi3YGR4YwH4E6GlLGIe9vcMgfVnJsOpSniY/8mAmunNZfhV3Rt
HmEvr6EBZGTHzuwPpylD4nJimCo063gr2Gr5ksBHZetgQRF+/E6EAr8tNjswbODgXLW5dgWe+SUl
clfsSf6UziSDXT9FuYLPxRNdjLkLbBOkAHe49D7ViAZx/x8B9bkL8IMUnZlrGhPn6T63OaLImnFH
7sV5qGOsxucQw8sbEGEVc23HdWVAI/I0mhWm28NHckFmZ9H9sUA3Ltc+x2OjL6XSozY2wPNTBPe5
7pY7+MjHNJA/yHf3kZi7g5Z/w5G50TDgO6nwTbL8HVdJOK+c15bLDxE7Fq+pjE6KTA1RrKZ6tV2Z
ZbCJmI3uhFog7TUTbdVKcxdgtpfQDAIMkvlxynd5/JvAbYu0gAvGT54qpld6YqREcDwkPaRqK0Zh
ACJ2+f0tI3zsUYrfu5cEKf3wUvuZvaHYpOxJyvIDaPGHQQ1wMv57wojS+cS744A7a7ysrYjGsc2v
2FhJvCItCE6Xj1b7V1hApYY/CYQ1pqaMQlj9c1oGTu9VahX961+KfsItdgrB1tQBAwGNKvcnr9kP
wWHhoEAbxWjd4lUNQdL+hNSBX7r9CbMJ/1V6OByo77mxFLmcwRUDyvGSGBqwjLb/hQQmc5UzAtAJ
61AeqxT6q5iePzSllYlUTfEFzOzoRQyo1/nxFBcP4uqkzDhL+u06gqWScD+WkXazQWJZJqTAO2AC
c9EP4gtq4ejV3gxXIu6cyxjLXLSbQCoHYbN5DDl1UGZ4w/SJHgkoRewYAVNFVzujWYdIMx4iVRWT
EB3EK7e2+Qg8e+WgkqHZbRJUqknZy9uAqsdDyFzv38aHZ0gihfOFn62bz9EeHcRkKfobvviYCi8k
kjumpwSMhjg3g+CvOLd8qJJdgz92LURWQsXj+Rv6siuRpA6Ecc731af6nNa99etslDiHRDQsMUQ1
geTPcg3XBJuYMzquLkmkgIObwsSQ4Kpp3bEjvFchiF49LObipKQM0A5ch3glzUaGaGpyT6FqIJqS
mpighxW036NkDWunK6UHl0k/yZ6UKXy6zLTfbgtp3BwzgNJnCBQhTUwesCXqjsBDmibxTH7fF9u0
gyt4HqM4rbECV0N4ITq/ao8W1nqKy524NWHo9QhwnQjgCal6lOI6M9WlrWX5eN70e2Z3XNGYI2oK
pwUphayYqHOVWyguprxRhkhGJJkdbGI4DUEWHFNtu+TFyz0HfS9yc+YnDbZj9DTjlzJ1EuL3jtFt
gtJQqldAtgExUo3734q5GEi7ToTC+78sG9KtCGwv4rmTmvDWlVCiP+NGOsRbPN+BtjWNZ0hGnSq3
vLI6jlceYc0J7AS24mUUp1kzjs79XJXGo6Jn0DdF+cN04Wm/l2ngUyqoWcZMKNDxN8A+6/1jb+AK
loBzLflf+RAkRBPekkhjC9NNn8ny820nNr/8/vxqmGXxyj00dW6byyQ9J/ZLkiYqMJZvaIJLUz0Q
+tn67a4EUkUZetL4dS4Oc9DTif31r4kfrnRoMldVkYEFKnUvVaKxAY7YxhQBjWYq9/3lYRY9gEeJ
Qz3RLmzeSD1WLSFBDTnR4XvGvS2xfU3ndewXAJgV0xLnLhGx3WO2RfaRSWZ+THFRKJ13BvSm5x2S
WK1tZcgOnYXvhlaL4C0hWE9dUCvREeR8nQkQSkduJDtFGT5fgpYr8c0YQojLqNHrZ6nF4RCJPjJj
I+GbOgK3wXV3n7p8REH2qIWD/9xQooEaVPG7czwIVPt/oGjcZc79bKmWkzi7w8HunPRDVVdMnQ2g
yqizrIRTEdjCeiM3OYR2feqYre4vcABV9wYjmPFEZ77j7ehncGGfqAbJdbzuqXuAxQ7zsLSfnU8E
6qC3u1+fors8v6een0i/f1x2HqTgVAi8uAJW9iU8EO5ZVD/S/V/vAylsQGSNZ0Fmaitotc0S79lT
1XjVg1wg71+CVuDowx1LnvKDtoMVLzCV943ld+8AMj4HBps4lx2IJ5Wo8t/e66g83K442q/kmRJ8
IXFZm7r+vWjNW+N3EV4ARd2N6RmdNF12/7v6ZwxM7w0uVtPNhPpdfTquqFroMgEr2uhBxgDlkDBF
C4bBlbMjPGlzqrxp6t1w1O4LzjMMBvrw0nZhiG3ZYdPDEVw08WRuyQdb/DciTB9/dMprh4zaKjiN
Yi+3VxXk2BGAVSbsCGfVWfx5iIqjCDnMyQpG7FILIC6JLUh+O9SH9nK9PGvW2MGvtK5PS+1NVGwC
m9jTWR0jIoWXxRHJDIuyAUfiXUtset7VmJdvyU1LGVoFSxQ1lXieVbFgRZSVwebQRZrRhK2HMiZt
jPDUUpjUU5qGB3Fhm8IIDD9NsPXD6vf56XkldiogkK4dO9LjnKIzAz9syWWVLVcnLoEwanbNYY5N
V6eIITJ4M9zLrmTQX97+5CEPC43YsAv7qVKuj8kh/7EdXQxrdXLmhFGNCP1mMYRsXG/4hcOI5Zu4
hwGPyoShP/y/HpnFAk6sVamfYmZy1vWjm5vr4K68tn+67lTaWo/Ee4hHufj/m0qfPrh9tLa5cB19
EElp0rCgbMO01VCVDkaBQh0XZ6lURnMYswy9R2644hpvSIGYnQ1Q/2Qaltv8uOQd0zDvMMnxNs9k
mLJU2AQt0JvCyvzbECU26wZAUb6eipnTuxT4OzNM+Iob9fHtIcwbd4x+RkLe2w3PEASPtRNgs/In
FQ3QG+1pC863kQZcVzTbzvDRv6i5li/4Egd4RKm4QaaMloQGn5GcB7dD0Y0ry/1CN4vQ2JoN4n8u
5ufE31YnFJJE4Ft5lhX5wUse+gTBIySdwUZaN80FrupVlOA2WGfqyr0TnWPNHoG5Nccdc2nPio+L
XEDmOKFBX6V2xpMkk4TrWm3VjBJ9iHQotwwZEZGPmE5wQgFshznxbgFRXcd//PIONeYvA6wOoj9v
AXYKu46q8cqkyBpCtW7pvo7rkp0BHPxXgYfTzaBcNclEPNOWRLaE5YBegkuUvuJ3n2Jn2cVpPLNR
PPQ5Ooa50WsZQhrA6LhenwXZFUQ/X2q+F/GtS8lo0c5zJSihjN9bXJH4ZuXH7kasuAQH+HxRZ8U8
vwQYRetivPwRPYSJdsJw+uNmLtxXYS5Lc9EkrMvxdvhC8ZNWp3R4DT+ReInSr1ZVE8Bpt39wQd9V
Qu2DkAXq1W+LuJ8TNcsG+5aQvli9ubDYUypD45cmUozAvMGlobuqC2naMrDNtWxWWW/nmGA6iqWu
QM8s7/t1/qOhLx4V/PsUkMHtJqklPb6l3NvYXSQmLLkqaiV1miZb41/WzKF95PRRWAH6Qm8/dWPn
lxVQ8I+3qfoSxoMQnLNU9c8oXoO3XE35RAtVl0qdoycoqbeR5fuEuo/F6MVelznNbOpspJyb0yvG
VxqhCkvMebKCK5UM6XKLfNZhDZoe9L48Q69ohM9fMw0e8FFmiX8F5WMwY/8vAvONSdBO2qIsYKOo
8TT8HnJSH+na1kLM8kz04WQZ//wv8eronhKMyo5I2jcFQ8cdP7KQnUflaNwAnVBDJz4sN3Oaejs5
YfHcfIAckTxTspQCp9bNIJA6eeH0qAQBxhRWhA12YCNMx/KFFdf7QO/l7WRVrqt/4Qo3wx59kVq+
R5LIXFeKZ9EPTDT4FvFOmq5zasgeFzvgUjd/dDidJYxZzYGWcWXV8pJ4utjsjG5Rc9MonorYvWz+
kwXjkQ4igyuwZeJF0Ap2Hg5CsIiN615Zx3vvX4bcBIuLQwHQyVUpngCASRlX6CYLCJIvZDacDH4W
Pn3peHTdrnGVG63h8q4J+7jT9qbEFJO/tLrtLaG/81CqYHynjILfTMPACUf6KXKPpKq/qKFN5OF1
BZ5gPHsL1mR7w6YfS7QXoJ/bkim1S+l/J69TkiZ6LyUrDHGhP/6XzmjQ/TnEg78PfukrtKKXai8P
cmPYYmNX9bx1D5jUPeN/FwxwtgvLn7/P5RJ16XR6Bd+HusKM3n4LhzyClwRKDG0sik1cUqxhWJa1
HtfkpO2v2XZ7wucmZN+vxtQktaazSXSnMb5/y5beFhMgROq5K72XfJ1VTc+91qTcsIsWR+yDSOTs
FloWQINFSNQYI5AdvEBqBw4xWs2oOHIOJ+qdmCt7IdR5V38EgU66TsaHp8rkAL5BavQpSQ7Yhuf8
EeLQrwvGkGyU27uLLJvwcsFXqEE0voVXt5bUH6tDBsgrpHjM9PqKO61N5RgGIK6MhWYCfYgxPDM5
3wFXu2b3bNKG8RtwZte0LdOgg4KJDHaIyncKQrMJhH0gHv/zthKqgj2ya+rQ1r6h7BUEbh7bdjXN
nlKirvCWHvPW0fD3BVq9N70OQSmVzof3JOeVquKpeWpTLEF6pO2DSnoQgnJnqW9DayOusY4l/Euc
g7NnlCgu/1H6PJQinGIXBgQuDrJUmHF07iQzM/NvzxWW0Pm8ACfuJ5kn+sywuR/MTikHWaUC/75v
JPq9bTpL9DzHooCpUuY2xSZa2GTYcXLVYQ+oIKmplN5POtO2UasakSjzINi0Sd73wnyGcWLIVzXR
/QpRTMTGuIJ5+cP4EWxA3iFIRMGFlqGcLGKdM50dCZ6wUTsZUV5v+tWHNzQHgr6/2FOsJ6iQ6csE
Vjwvqu/TxxCXUhHMatWZA9IueoKQgY+Cf3SaeVd2u3cHlSImurvVVRNxtUZyzamKxYIekbnXBEK3
/ci6DcdcxZWUYfqe60CsW64fFnE2ECdl5slVpTdrugT+HJzivx32tw23niEfdFeJQ4oZAJlPyjOU
VHrwTi018RzT8dJyXYzgNP4iGHqSjUcWVyqPBTEm+IJx2KnodSoK2Mf54srnzciOqtGKCJ/YXAkA
cLUUqLyrWK2DxzXZIecyhVTxm85rJStcJ7s2+5ZduFvGbfada7dTNDGtJ5be2a24pdn09Lj5muPn
3Kr8o/q6L3iEkAqkUL8TjFr2l2z67dOlHKMlwV6Z49j0AZJRiT1/mEf1k+5t+NbPPIHu/s7gF90b
kPsbYmCl55LQjIAvhX6jDtsGAqfkFlYxW3WMeZl1nQ4k8kk6etbcM4xQx64oMWtmWIkqkTe2fTZ9
GYmpnsUk0SZUMFLwN9um6SQNQotKKd9CoJgzojCUsiesOBcMNIWx5lvgGbyjNjstVYpnuiqM/MQI
CYr2B9L0aijxbblOrrNZrIbraEB6KUiwalxvrZgfni0Av5d3gfSRJ25prw3SKk/O8HER6EpRX6tg
ezU09T5P++rv5AsLg+rMd2aUnQwJA97O64NcXFUOmvxba5irjn8HkxT0xSFLAHS27GPtPc92nqux
o7Gape5RkT9qMTgZ0xIJ7mFDlifEsLgMRH3LT9V2z+PvQL+mJL2Ucj/GG9kBGvRLKGLSSBtmsOGe
UfGoIc1GsaaZFnQGl7kP5SYAJbKcEzNB1Ueq8dogwnhXrtSTERHNVXreL/BdibdXMZUEiiTp3L7Y
wI/6jLucMb1Q1YsqHrTZ9IBCkVVSFDlc8MLBIdI1xhTMiRZbLlY1CMdtHh4g+stpI4jfCdcFNtoa
FF3e9u7iKM7DKbtHVe7LUK69qnO3ZF920ytbD2H9oQveuXaksFDq36nU1f32P6sacI8BuhZPIxzZ
FbHij0SKzwAn6M2XGhR7wakrhWq4fKwp0Q/Qq44rUK072T2hWup/41GQU+d+v/2pl6ISrPwhxwqi
UxQH4IBoiM7vFVqvIMvFKp+UQj/qTnHraENdu0nxrYUKq/XNNsBeKTy1CmxwjXpE2ec6Uav+maLG
BW5I0m3pYc4qVM/BIVBrM8y3imwKQfAtVDvOBXt2KbZFLEhQkafFntsOz1S19mo97eIP3+uq1kPx
hSv/lO9i6jpILNaMY0RS8rXOH06Fz6c3sdnggxvrqrZurJhueX+PTqYgv0KbB5vkYV+2KNzDftXq
ToYMO1JbnI+qXcLSlm9hSytw9C3hRnIThvQXNTI5NgxfWDSwVHNikL08i4NRe9xj3xVHPQhiVijf
tRm31PKZ9hUf739opZT5XaR2CRu6wcZ6sDd+4hA+kUsA4dH39acmyG65eJda/a5UCbCTdYyLHJyi
mXT0n8Q8lW3naEIF3Y/bplXlmDaoh9hNQWdbipcYqq4H9L3jXBj+uVyueOWYd1GKdOrRxYP7cu86
eisygBiFw/Ulhod13fXBbseL5MYdhXNRb5++zybzqntzDeuUFqIZJf4MB3U5LtJChCpP0IS4otID
nbMAnG7OvoO3fyV6lCuanD5YxzB8XDRYYFpjLkSUtUJj+GV66IwyKrtDGPkPtHL46OwUe+T55Ro1
00Pk/8+akURm8vsPO2kPjdppC+BexlGcjNBImeIhyKSNskk1ZgqjLhBXvrtzeDJpSFWrkEqCIAmn
W4+LAZQRbZ9TupP4IW0SIf2kOFqrgxoeZyDGbpAWNBfWiEYLilDRnThvytL+YyRMkjH6q7EuzeZk
6mcOp6dXmZooVeYHkoX6QtyrHDvxmimtZwqSCMUrZR+SCwRTZuD6VtWjCbm7+k/QAc+jU6IQHF8X
2iu+vEwD+0a4l5v55lMyVDY+WbFpwljDoV8TaI8iSXLR2UhycsWSVHxl7/TcNPFN6u0J+MrL7QoV
mRUCRnZvM6JCA6ZaTb7G5OZ/3b1oeeJA5GB5jZH6MHEt4xumU+iPuZQlee99gfeBDc9zF6abySGw
8ZuqkXgD+ydS03VI/e++o+GzkguySlqesigfJAdABAZK+HOJCHMhwnNNfa9SK1yANAvyMMfzXxMG
kFaXOsAtcobY+SFHcxjMrHSalEv3dW0CD8AyyCOuvFfCwo8Q/ao+zDCwZGbZG+UMPC9GVhm84Rg7
VozRJSLJ3PjPnr0OMKvzIAafB5NdnAPIHysWXz4h7itZWen1xDuBnDq69JC95KfyOIkzYVmL0irZ
hbEqdvzpJpo6krlfL1sjfsLrq1FEb7JaJCd3PJJRP1ZVGqABLdOFKqItKrAJ7URs3EYy0VsF1RWb
7lv2EPJd4YmpktijVyzCVP5003fM/SzYfK2rfHEp1qZ059MpPfdRqaDc+6WrtYfvrxwF9RA5KIqx
USo0Agja7Y8uzT1im9LwbK64VurNBf6XId1OT62+Zl7D7+K2Eowg8M2wDyeoedKBYcVp+GCaHTTn
BKIismKBV+ytzRNQivP5Oq3CVpiKE5K7UusaNc8W8h0Ew6PU/ORUQ8s7f7sZVju0HwEIMLLe5GrA
ZXoJX+bet/f6M6OsHJOyhKEoizM7jIaoX3enX5lQ1J02huE2fLZALdMWh3bf8iPxS4+fP9PrIypc
us5g/X/9OF+fw4Abo3bVuWZQEyqpKhFol2Guu4CRUUprdE5rWU8ab67+EUsraX0fVKo3xJWvbIt8
ZFD4wIE81N758Mg3HLi6uRkPZrGGaIZcHqW0Asrn2rmi9ffY7sFofVPAa7TVIfj/fZz8VNBOlauJ
Q0RFKeV1c4a6A1gDjuhdNbVQKAyp33VVkpbBF4l7EsMbNexH3O4DSvVZfcqxQaWyNXUi7k2cY4XQ
hmlr/8cOsqbs0a/kA2GAO1dSOUFv+evTAwo42q9FMHyzfoAdED9Y602erfu6OwOY33I8jzdK0Xg0
VYA13+eHnKypLku3RrBnyvo2HvBmFhhuAqEcRbpTi8x8GfVan/AwwvljKDX/rxUpx9/w2QLJ4cDM
WT0J+BXj25ChNe+sujxUvEBAgiHUsLfdniqctGgYxNP4vdvM5WBJsl/TNAfFsiw78k2GGo3bZKfi
0XcODMMgDj/HnOQmemtGnIuRM6pnUMU0QV9Eui4xxhOvhzO93U6tY6IzF6CcIaiDsVNeLi5IzoTk
5K1+YlPDAVd8ec7ZkuWVUQUce42HzUrf+m03jrQ9Eu37Uvc1oMmpuVBQX1d+ZpoRYxSF2BHgxJ6g
R0y0CVjj99XapeuSxaJMv7w9RnxTQZej2DD3nyBZoiPvn3/y9ibKhbtijR8u791C3/1Hi0I2uIZE
O9zMACcFa3LUa4gbfYP+bRxVmJcXkvU/D3+9X4xcYK4w20H0Bima2UqOgWJaviOglYqwUWPIihxW
/ZMP7CpHQ7rFTftyKwRaWhJlhOqRRO36MTh/a/nh42cPeCLOaMrpAGmFs044k0Nh0ueunNeqWBbm
VSu9mTQpUCAPvAoP0bEcmnnb9ROYMMhd7YddR39d9Nq6/3EVzBviF6oiyuIHqAeDBYaTDPaIfctR
EAW7GuBd4kDxU995Hcdzpnnh52vAZpMqpExWXtcraXaCWbCtcBIJUxZfvYIDaBEb7MJpN7skXPSR
z/bJpuCwscOl9Hb6fSW88zkFJYGn3kOdl9SOkx4Q4J8F6Ds0CTAGtUNeG5aZk7nOhNasY85GmNd6
ig9/TrZfmUtciHTeJfQ5v9l1PUa6vyhcpOKxAMzhrfhqVnMQus0rAUT89BOKWSwMTaX5VymeJ7RR
TL0XzlHD3loh6sigMG7ZPZInm2LldRPp5gSyB7R3Jtq1AzqdJk234YXq7Mih18GjwoeebfkvkSPh
HobzXPxWakFvGGsIKva9NJYX/+bbZa8If3g3KBTi2Li+RWdZwdaNgRY5zLxTUNc/qw6urqY/BRRF
sVmspZwl3lAeQnZ7cAUGXEQqAd0Bf1MA3QVhDSq00ejzhax3gPo6THEn7sCrMhY+zi0EQ0ISidmX
8OIwLmVXpT5qFGNPAamUXHwdX3vh1X9f0d0j9c0H6F3nMGtJtdQxbOK5l3Ce6O8WtqshhzQiF31s
BfcEvKu3avIkxI4+wC4PM2+aJaZp2lA9nXFXfDxtN+bc6qoYOqq/nFMWoTxyLZRSictM/u+bhrK4
3tjJkK+ZkAPS0+SqH5xWcjPWhJ8bGX4SZZldkUWyYx8WEKuih/NhvMqmH6IlRhf8yncXrZxINnru
sAbyzVA/rGFy+jN2Ihfswhw+Bc6jIwFNHf32hbKZeV3R1yl579z/GmxYoEZOzq/Hinbz76lJrjsz
Y66ECnBzUUAmM3Lr9k8V0QeZ9f2gODEDq8QTJEJOgeC+hMK/dLjwJOrbm+jI0OlTRyYgnfRcDIwC
sJBtztqWEj7fJyLiKuJTF9dqW+KFU6qCsV4xTMB/Eq2wCv0nhi3FQ/1ZxSg/kRVbqdkAQJM+B8pK
a+dC+A2FpStCJ/EOAriS4QqH/zD6C9SReEx8H7iCh/yiC5iR1/AouoPIUg6A5JEMuw94XTtdFbW2
aIU/d4rvWsACoFC9bYo4DbCgIfewSHq+KcExYOBNaLMGXRjhNya87rIfeArI6XuHlYaBDiQ13awa
AEiwt1Y1q9q9+vrZ5fowzdhZZVh4dk2Y5nA5gBDR94VRxQpa5ifqNgCfscRlV7WrQMYAYkrhGxva
tlX9VBI55c+BjyzrJjF4cGbPe2ElvaOSd7biPZKjzWVIRfBxmObohDcvtrqfXLTh2i8FcpiL5uhb
8/gY1EbIQFmsFJDyzobtXjO0M+xhkl9/cGCm8tAQKlGiZUL9IocomKVf+UZfJbviQg5MriVpvg5J
iskrhUBFT9JC7LZChrjU1MNN4TcXdjN8bZt+DyON1zMhklVP/lyLNDcjZsHaGwq2V14U+jbFnOWv
aexq8T91Lnssr069W97/xFoE/4EqIkJugZNZKrIt3Z3GrtkNX46HBvjgpAQRKAdMzjz84HUb2ZWC
Sb9xamRmjkKuR/ywVbEG2lIdDSUMZh8QbTN6+ng4IjqaLRmXAobAjokHy6fNKMy3IcVHHEBPHgvR
hu0tfjgMqo91+AgmcHOPAAEutEw9qDTOu8HqGXXm1QJeU3+aEoZ3CWs0QUMfMtEPn1zoLgk17WHV
JaWadHJeRgsy/wLgTXBRUHxs7oFXz2bKlDgwRUBiaT74wxwG2+QMZhyE147/Djsk/OKTFgROhPxu
edChWdrczacMuK5onkEFGigqyfXAuELijo59xqjOf96XakzcSSTu/PPuE7v7HCShoiSgYjIamfJp
bWTbZa/oIDhpqHxuAD5WBn3RJ7/oZ8foK1vJLdPu80fBYUf4+zDguqwS3VC2JN7dl0DROQuzyCUi
uBI1Y5Vn6VLb+F7/bSfnlPMkTwNMWG3BeEz/VJt3s3/p6t+BMTjW733WG2PbH1tB1XaubweqJtLr
1LaE07HHmnNHKRQacIF5D3x3xrEuggdOUjl9zXqgJuHNx6iA/LjbwyTaTM4tKYF8A80maFBaify7
gV2WcYdcFDHH0uEgz7r7ecdHtTVxeVo5Ygy+4SDutLKZMM5+/eML/8mGJrzkBJFRnFdWlz+pjxWe
LZzb1ESefD30gF5i+aHDlFeULIbLJIK6TgrvCc47ODKBxrynFD+/KuMs0Jzz63EKOSEKUr0VFkqz
lyEeGIDRGzE+oCQkOCgfxFBm13gfI3L0t1tBv5mvPOHmMgI9Jdidr92yyFXZKvWoKPK8+FjGAeDC
h///SGHlHwEkon8G9azCAXEPwuTiWhKI6C4wS9T4xL7SSBFdppybmrenxG533S+IjwXMMmflMNud
yM8ZBPSflMemxYuubEypyGaNLcnrB0kffvkyt+FPJhy5RswUQ0SYd0IYBkXAPKV70d9N3tXCASdP
DanALBkpOoPAXBe4zpbdnJUBN/e8jSbbzJIXFXy2fi5etZEreJl+KWnHR8u1lZ0Qxo0jlkx6dyaH
KQ183MyVjdFRVV+zI73tUDhI4sxGWnM1eP4DpZr1PSQUmLL7XadElHtxA+Mogbk0hu2lf7rKZHil
FICzGq4RSSZVommD+HrMg9Ll2qcEtRS8jpG+tRlP8abbiOpwFUJkZOoPoCD0bXv5FTy6jJzArD13
eHvZJESM/FrqtctKZOaq6+09yvQVsPPMvqCCh84u76gpUy4Q7zEsZCh+8EBGVfG3nPFvJn3AH6P/
K4W65Hqwp0CfuiS1ccUvU6iA41+r7wJ5EoK/Z0tNloiKZONxgPQYrMwcgf8XM0ShdMfXkqkou7sx
d4X+04u6kmRUu9eGmZo3ZdTGyf9i0LfCZyzvTgXJDg8wCFId7spJMIQO+Dl5jz2DogJPyQhOh5NW
vKLqxCAfp//dT60KidBD5IXC3GO0pvNKUiqBycmHKfTw7340TtOWCKOcJh8OBLtiPzrkffxmfNTm
xl6AKxb59saT6u/LFgzD2JuoShr5xXI3g2lgZ31J0C6FCJ6F/ZcKnZyvJaFp07b7PgY2bhV5Gne2
7FV43bgqA4+wyVF09dVbgqqTaYWhwkbv5k4RbstFQPIJrHteVMoW39/nOUrQNGIgDL1Q6O3zMUkB
vR13Lr0Q0sIIR2yRXVSW2ufW96Kz62yYo9mz2brUQmOMh6f7MylUUC/x4XOqMc/Y0O/QCoNyCYHH
4vetTCme4zm02iQER/HPabhMhYn5OrSJSiRxcIawdd/7q87Yt/i3v1UGXI46VFHDqI+i8SmV3zMb
p3Kq2x5YT0TJC0nOtxw7jNrAYGOPQ9WYCkx35fbcUTwJ+UdInC+Ybe6iLog/rFsqnqMBFFJUFme5
A8q5SEeqO28U2WRPSpBKvUbZnGXkIBWPrP7w7dxH5hudtbjzZOfo/Yx/Ud8qBXs23ty/M87Lz4EL
yGOAmhy9qGAg4o9DKxGnwSp+o8lkS+jfRRVImjChfSTT7VAo5PyUcsvlrbGlGvatoJx3dB3I6WW2
ISDXFSxqzehyJeYwHwn421KBE+tluiOeCVksv33wDo+AbEbm107XjZCYKDT+jp04DwrqvD+mBzxy
W5sV870Vq5vT18lAI5kLoHXnV3JRVUTO6YMCA1xtoGrE7sLP07tHwFcB6yvsDSG/1jkjGXnhuKup
ST+UIG0S9MnLYCn9LQ6ZX0LP6R/78Q+oqQpuMiFXIJQyHEKbAJDSVGon+W7XY2BAvoGCAKoZCfjl
AnZf+AhKr/sTjmQkqBvbp8/WJxlvcplklDtN/zR1WpMmO0YklyUjp5+rVITdcy+q3XcYNVSO3a6d
R65N0NgCfHdpMAAcBka65FSo6Vc6spuHkTTZvLq3nNdOn+wzzEuddA984Osi/ieiYYdl1MF8OfDk
Hq4J3Ug7B+MV3qC5Exi19pqKDKefutIrcFHuhIP4eMSO4ljL7fPtvpfjk93I3cvPq2CfPBquRNwJ
HVkrr1vxVBufRZKK/7NwWMtAlax03Gk8VCx3CZawiXwKHcQSKleihKTHXfNM9r9l58IVBIgPzfpF
DEpdQwgrZxb+2UmRgkB5lAmBFhL9HT6V5FerAQtiRcPag8fL+XSgjAk7uMAeS2gpYv/QzxhENCBO
DEOt2LiL6St3V7SOmKOVU/fyjBqsvHVYhSU5a07UL5ZnHw6xVBm6eBveogF6/vzm8W9zNGsi6aRA
jY1cFg5JyYxaCBQiWNlJkUfdK05FwZ1A1Z1SYgcZEyba2tXcjzmvtDqyDwuhPgDaxv2O7EVaKHzM
lQFQOAX0xLf8ejba9W1MuAYzOusvEAxr22y9qbSTFA55DPHpSeST9nXPq9EL9J3tHgtRnyUbwFaL
SIu3o3tni7cm9jg2dQdWdsXP4/RrKOzPZUt5E4jy+Oaxk+tzvzkT3+mkEd/hCGG/R5ZkTPBVzFTx
u3eaf7jI/GBFoJ+r8VojM+af+YpxWed0G5dMSKpLi+d5JClTMcAkwsyKQ7buixY8N+x1wYXShMlA
fc+EHAUEYjHVsUqbqTqg4tKfYEAiTFlfhXw4buD/NHC9dnxsVyeaHZuYdwNkhHKgP7w50+Ar6j47
PDymgGoDqMg/y6mSmGsnZHCQ5n2fBvq/JA5c7QaS6dGCRcBrcysy6VqVcwr/qkjWv3OM3grZNaSo
9G3kHPXzF4NnO5Gm0/Ylrn12hRPV2dec8LVRgu1939OM3yEQcTQTDI5zKo7ARFohjrTX4tdJ7Mml
LJOxbbQ6VDgRJZp/SvUDFVOOdPN6DBi4EEHVrBvDRsvLhGG5yZXJ8LiR8K5nsTRvxj8WGtciZ46e
FteoEWkjDVoXfBy+vmPxfi4cgUw3ss2j8xzb8jGiDZNUdWNKI+4Ev7pfpBepcOWLit/8Q8z4vPVB
ONWgZMZeEFDTWzeMO1gR4BGfzX7JLutG3/moeHSDgEx3v0ZavjrMmW4qf6oh8pyedh/3tiCpnj/u
A1bQ5+QCV1nm4c5GCuhm1cwJ0/swpMTQmD7k02kURwFZVHfiSoMQww89SlHrZEdGzJ4+7matc200
PXFpnDqSVvpC6GKmN1RWeKmg/9Z+SG+cGk96CtumnSDCBuPgAFfkeHCbVdBvSo3CHDx4+77RlCqG
caY8N5VsZHyPuvIpfWzMX/RwxxRuth2dXAaF91Y1spjDnFUjr+33HB7ofX1U51fATm0hMWUYqjHK
uVbq371d9ItsYKcvTdrCqU+EptwJVawQU8+IbVB3DDQPRWd3BarS4iwbmxo8IRvDglHFSRO56qg/
mJvfuf05HqoBN8BQKBclRE/oXcS2a3IEQpyLa89M/MEAaWdSOEuQGJGiJRN/0KevzO6LNAd6za5N
l4fhZ/ZeUtewY6ZrbVfHoT0tJOw6vU9XWnvk5fJL5naK9Yo0Fgok0trZdxwlafZrvMACAEyLsjPr
whZJokJpFsqQxBizTHVdUh9MUB342bbECotZk/ILCsQ+M/zTBpjX8+m8FtLMVDfEY7BcoT5OugqA
nuZqrml17mskRDLS5p6E67r5PMkf9xDRHJrt0uOGwLpemNZgTcyl9mR/6yyVO8+eS4MXqjXJZlE/
jkT2iO9psyAV/e1u4fXoJukgH+uk1m9tpD5wYqj7gcKOKrtJywG3dUUiUxUsP445WZRXh1KGvdGW
GnAaBt5uc+aaqiSsqO5QZL91jeFyO4BLm6V2/Bn0ws4sOZa7kDgfiaVsH1N2vaKUa8ibDhY7Har2
g9BoGiQIQJDyJ/NiOa7osd8vClXM4uuUG09knmDCC8tZu8/LzJaidniuerJ2tS5zKM6Qzzaq3C4T
/3FrNcYeKZz20XJrxl9QLmPLKcRD8Q0yxMYwRIej6SS80DRtMx4TpGB1sYj7Vzv8dPCbajiFKGmr
AsO5p/2d2RPFUElzmfcDCW6kLY0jr7aKn37TmMzk4asv3WwBxMbCkmpca7/z/AWMKwdDP2cCoa05
E6Yf58P8cj9RbkEKaBiQimyswDDT0ClEl5ihmgiFcIWB6bDmdQCGMh+zZQ5Dy7asuetIRAxt7C9o
khOxJQCUhq8whMYGPNBsJmfvpqCDg1ku/xGWBk8kEZapJjdBd76+mGRhB9pgj9+k5NXmY9xSly7o
pBJO/thMQwtGuJaPJVtYIcJrcg8NfjYJMOnPxvZc70rEB3nsEnNwHuBe6dgkx3DeqM5L0vArtfLp
5cSQH+XVssKTL+4xU+dogFY5hYykjTyRHiqwN3OtUkOqqXGt9j/22UkKcXIf+GEwuY07HaHhDffo
A3FpKqcNueq18oiCpiprSj6Gv0mcrMpb5o3Eq6C7cy10jVKt46FygkfxpojD9FrGMWh6CzAjpUBb
POJ+od5uJpTBGbL9+4ejeaQAKgHr4q7YnLQ++YApDDVub/FH8qbkGSTdFuL8375m0cISptSsmXBu
1Y5KSaQ2kb+u4PXID4F+3vbAMqE0dV0IZIKQqu7E9aUD45d/maZ2el1DTUScd1w0Ksggeg0EbQko
LjhspIZWkUT9HVZZZjbsKhA5NVS5lCcqa74Eza6kiZR/7f2ogkNPFrumjGXsC2rLmuSmnxIHsTdL
SRs8e/If4lQlsaoGlDlWooNenk/tbw/wbsggjE552lYzZwlaF9TQXF2aP7kp/nPCRM0F/kMkdWVV
M+Fjq4UGhu98g9uRpZysUiWuJusy1ztl9yBVuA+v7Rcvo7pDd+x0JiD+HyByHbsoZ/VYvBzYaq9x
Nkv0J6eBKZN3CnnBr1rpCBWyCGPd5SW7MAAROyFIeDtHAjRTwzQCiW7WhWQkw74pFqxgkUF6gAxb
QIEQ6bmjLiX7bGgOZUHI4ZEhfW9KgqRa4JNb8jg1rX/aVcBXz8CB1LuGI31yNWikdYg5YA6V8c4o
eriixE9/yxfDbTeLD/8czGHpOkpDKlrg15QvjWt0NFY+i1sC/vkTIVbZCVrwL194tlh+dsr82QJp
POTxUEN6HtO2VQAEfhQpcRS4UqierMjPVIYDzsgqVLyFVFOdvMzq0Zi6TrCpQLBNNZBoPlXWMSK1
KGk9zKTUNl5gaY/lo6w26y9HHFq0gWCiP72btP1QQTd64wgLbI7Ctm1UaYCb7bSdiB5eMl/y5lHR
ADcVybHizikI4KSulGbt/EJltGVBobllGAJf2E8KPGW7u00MncmUFVEwcJaeu4ktg9YPMGrmaUBX
ZhoRgQVH0P2Fse6fey6mPmgZvgO7rs0NpEefogIu6F3xBACxIgX2HO65urNSs5vn2MfKoZ/HIWUE
UMBijvZwEv7+TPGdGAePB5pCkixGkNhBcFTNT6TNAAoKdSv9NKmZLdQ/kJrR0xJp8+68v56LoirT
w6vHPaIZcyt9+Dis7S2b0LOU0MW4zuCkJSdjFERRb4UjEFfpsRvXagm7ioOZ3l/NKBD4gJ7fFlxs
jBdbdvZJ7X+jR81oPiVRTevYUDNZ5QCPNPh1b1gpUnLSfITlQum8ynnEG7qelhe1u1tLGyBx8pP6
qRejMwh3J0aVrYS2shhpsM9X4oUmNY1DJZ8LSQlhOakwFNxjuRRCYvcW0mLYTZ1uPjF2LVgThg6E
j9Hsw6HDGHfWEkU5XDn6dzcFjllTiPWoRdWlz4XJi/6zsXhBBqMQoDOF5fiAbVd4m+Se/M56fq3/
kP9cOHPQfFU3Jj8/RNWwrs3lboJ7zBXzDg7CmZFYJ/Tg/zTudrpdiFn0akei96e6hlaAuejlTxDS
sHLRSdJ7H9Iff+XV+k/nAYv3LqfQhMqlTgiLJdbiqphhg4J+8TY1Phuhp75kyRPvymqekkVg7KEw
6d6ctaTd24YDAyx2VNXo7+argWRSiRflZ24tezYWPN3gBC3qmH1apQQopCXJ4BPd4bY5kLvSiboX
PrQ0wCcMjEqFqa3Lg/r1RSNU7IaxXCh+h/lCrKH7e/jlFw0pST7rNOx+g0uECJgKr4fln9T/v1oT
WuLUXE48nwi65B+SIEbE6ew/H8IYyeZRWTXA6yAswD6u7Map7VKIoPG2lJ2ZWvl2kHsU8aiDrQyu
RilCdlQGiD6R4uY+6HT1K0eSDSQ4maJw7Cu2HjkICm/33DSiiFe0Jr3H4yfS4FpfffPnddBRMlFp
F136/Ehj4Gx/TF9uaZRTQgyFF4DMGUkMfIg8GWFw3sj5Ynd5KgkA/w8gommQ4kIxU6KR6LiU0Blx
w0cUiYaXkhS5YevOQ9X3g8EkiIcBpdjY9669lKg/5J/QNmsm8wORTXkm+2OsKdgp2wA72gg5oIFw
9xyIEwaTBhoBf6BqpJpYgU7wHllIxh839nGern/yrHxGARVw+/AKj2rixCJ2JDSmxS5Q8F3HN8Dy
0KAshP5hOFNVbAg1t1A9qsqhs9FgAlwQgBZecTnKbkpQTNobpb9AI2QTSPcGZGrKuib6ado/f0xb
+O8+uTKpeKdLq/zZE6208QhWId4ZL3KGXYwuF0/IsTiBFUuuIEX7+UMZLDwmxENvXHXwClYL1/s7
ZqKfGZbUyibbs3Ezxr9JT41AE+TxqW+wjsTmJ9Sc+yRdbiryPlPV/Mvp7RxS44+IEUTGLgh+2pl5
8rj3qOLDAz3s1+Xv/fUBtrmTQ1lW2urGSml1I0a5vYa9xdH3cPM5MWfvFLJQbTX+Gl6TUokUexVT
2f2uUjhhmd/S0bs9Txrv54ta+rusl3hcLfPAGWbjAc20/3fJ84gYJqa5LbkoWmwwU/3NYvjCAxiV
t6xR734AxjuoDN8e77PNvAa6OytUNBwnHg7pZhHIeNY9WHLR8Gr7xuWXjfaoIjlFK6xFR++rN0It
4aE4YauGQ4PqBsetW9CAVvKeCMVE0mH7CUrhDfZD7z0tC0gkgg5gRjLw9uQT8Bn60rjkVzyqSp4E
XP/3n2mgKibAdzIW99qC1Hv7204+B9PXqg5gcGFtPkhhzZujcwzue2HjKvAr22Npf9yN3CSxIuHc
QQprQmoqQfefZ/9rAmV5LlPpG03UnO32QSwIIvGZGF6NJxGY+MgxpbykrODVwEypXeZIGwxrqcMm
x7/ZCcev2XgOSNwLWxY5G/sPlsOVMgoG5Y43x5H2fTX1T13qNMggPro1HX8Q3QfioeM2H558DaTs
xp+i9DMKiLguH5/crIfdwdeqdxBLK1xW9x2kpMn9Y8AZ2KtoL94W6jSrpi7e2UKY2lkpU/9qYk0A
kAftbDlyHMjb0l5VTPOHqRvCmPuoPBKeVNFcn2LChmeSnhUBcOhYWW81hImC7TIrMUaxOzboPOWr
bYTvX+IBEbMNMPKGKrJEScRuEY19skshmt9+bbuH12XRCKXRvnZ/Z1NmdY01qxh/jpARQgWxCl2U
dTuESYt4xnK5FP6tPL0Kr2GKD+4UH3UuG13fGL7FYRO9RsA2GtCmN+kBTtPKVDxdCXH0xbJHd09G
R98DtBJ60Lyr9uZds6vWBzeGCm0QJQK2/hugkVqLDAwRyHmLDHT4G9ChBYoe2nH4eQMHhQXk4Bpi
5quC6HNdjbASrc60GkyIomwHv+czKmRYNmS71EM8dtVcogW2OlFRVRfPu0lOua851L/ob2fA7mZZ
6IU25eBlVcEsbSdoUHGpfs49ZzxyV33hYlqwNxbHVXoeDBoMg4RhChgpoSen82A4cnjE5BEFQdqH
FtFrSB/mTjy3RTqGuRZAz8RQ/QuYQ7Jc8Fuz7Xx1NM9d28xZ4YK0XeSXaj4WsrVmL+/YxAPT5gHI
SIkce8ea/gi547ZZepwCLEFTRDXlqtnWhBtdrNsUtw1LRSB8QPB8EBr4ZsIhU5w+Odn0MMoKBgoE
Epea+mpDdlLd6ePCHSpLNW5JoMNM+Sl+negIakmCMKEdIK+xE+SGZ/EnZciQBnVUv54rkYQb8OtN
5V50IgeYFVX47hU5CqI/2jkcqtATvDkLXFyAgQ0d3bGrBELqJho6lQwTd75ainbWbysz3EFD3S/d
j7BO4DdvNvPpGiYmOtEZnGP2wkQdHrGit4Qz0+u88b2Hw1gmeQc8jFRNiPtqFT8/9/bU0lDRvICc
SmiM7PqfDzvFpo8jR98UJm17spgAR6ouMuLa+wyfFwyhEmNH2KnWORfQ/Ub/ry57fD9VHsrMuFZx
ZoAilQMd8CSUGjrBNR7Iq0WhL7WSO3q5+MRgKTrzfr5UTaBZXqoLJjmmWJO7t4qzjKArj/5bfhoz
bUXaL2I0msRf4UJPWAtcZil3qgS0xK89O0qYd615DVURvpyopDNBuGJHRqXbJIzhYJNXVjl0KF1n
YLtK/zXK0kk8EDavlTk5sB4vmeM+6i7XY1Cxc6NMmJH27BZeSeFI/5BvwyiXKTCzFVGu+u5NqS2C
BCsfYqoevCyzxJmhoAQ6sVwmJvwIP1M/XbIiuQNcmhLG72Pskv/R9GjWIQsPELUxR1tcDPLy1tbg
J/qt3KQQqO+1Of42oynbMexz4/+2ULvs91k4jOXyjLrThjsCOhiE2+IempfcSB7Om1heFRd9iZ43
7EF/HH7PUeDgPjD8QbKQojuEieIT+LQW1qhUw0hsTty0BpErBhJdvHss1U1ENdtQGrH+/TjWwyEp
eC+2wazjib5fQoS6eWh8W5APl4LcS6Ggz7cdyH1C4BgpBM7KM/1AwUqt+j6zjPwBvuyQmSl4QD0/
degS7hJ0c1yq4wX89xPJPJBlHUrSJ1VE3jK9vYEStZjl3BWqGpXCEmonueXKv9D5U+z9whhJsOTd
Q1Acn59Iclpd3ild+JV/D+N1bH6quzLcGh6KTcgpU6JV31jXlQwP43JO8rMjDBFhRdHu4jKneu0C
huRX1IgBuHDIaCsiRDsEfIR7WDnExeFHFKICe81hyd5peGnEC5MbRUITWxxUGglGeLvt5JB5Yxkh
HLEiAY+pmSvIa2fym5kBbr/96d0yitzZK8Zyc0Ea8Du4VIgm+k8pTgY+LY+2ULWvZ9Vf6ReuIfHS
Nl5mN4eKttJitJstaSIXX2U1FAUMDbtwAebZshm3huLRT4DU9vE1hu7MwVYBYSXvmMUnXpfFORj0
rWSHo02wCu97tvVk+msdXYnc5PgCbG4lEYTeaEHhBri3GX8qVvvjfkE/Oh7zln+M02KSOmdo8Yn7
ZG4QR14Bwenw+vdROErnzXQAgawJcrlc5e68cl56meeeaCUoFG0+n+aON3AH7kjl5cZVV6Tq03nt
rwYD9A1w1AIqnsVAeaIpE7QUeQ0wyv04RVHF+nfYEbITJlEqXgFtzYtL4/nonhKhIkgdZMM+EQZW
juyj/GxMNaqCdy7wLllX9WDaWkso/hIjsS7wBffB44Fa/fL8Vs69mbq2VG/fayC/QCjqkDzRmH7F
4s8YVPBw571nbC8Sm0SH8clCW/EP7dQKuWd7sWE9ETzVj8TVQmJwoPViFWDAzzixgWbE25Tb2D0S
olnVseLmARi9OROpZLYgYz7gK06zR3/itahuGvuCZmWXL00u56dEeE2t0Fx9zxyxjyF7LU37wfLu
K7GSFa5Pjw2l5yiWfq2g6Y6QMR8K+Q8q1vwRFNRmbxEHe1MGxSHk5N+/1mojmXHquheN6/yPJjkv
IYSbee+i9COvBRNViAukQMy81oW2Qzo8lV48ZO5wHmKHyKoaFSEFNAnhHQUMgKqxXOkxp3qmpSJV
nhbvePFSq0cs7yTCJVL3rFyERVNJ6vfq1CrZ+kGMTyiCH2OICQNLBUdlX0VpLJbyoPRSp6/8p2Wy
FpDkQPYLQyeru2x6dos2N8VuwKCxGtyNs0w8+APAfdIk3LWj2oMMaQTCjC5HhGyZPdRqgAnB2/Dr
RrVHdG1A6Us0E98Y7kHtkwVOywqzw5yRmkDdZLxyM5+a8nfsHiavDpzxNCT9KWuXalOjWAQ4ID9s
S/1nsio0oB1GNG0PDsFyYT9Hfb/S2Hzj4A0Dw3LOAI3kEIXku8AZlLLGY+PyMaBcSbH13ezRRLGm
9O4krwXDFL1quVNQ48zXh5CxEBR/+8IMTDZ5ww9OUOpPtbXDY6ZzogXra+TN8H3eD/yOEeGNBOdK
SABrdbn83ZU1Qkd6Hoi6okYiSszjEKyMoWTlEhQedIPjPa9okt/BEN4t7Eb0BbP2ONUttt4u7TUy
dM2l4m342m3iGeNxfIz9wt06dtW8hsK2FxhcJnBy9kQ8yBgxpnfrEdMB37SfxRUVtAA6PUTLaYvu
X92hWiKKtt2r92Ti2mVFh7jPH/9eX6Vx2yKnALXJ09ZBQD4tuxsGryzgxCPft6sSC2FkVgyIeUSE
3QK1b27Fj1e0CmyEn5ziDWJ95buvdVC+OI8Y/a1hsr7BXa5qlkiY7var00QXAuO8qZvP2SrzBDnM
Z1hmUbcOYbOCAFxTu1X3cDfn/HbifuVK7PWwnYwC3BwbrkKjuKy9Qx4fSU1I4EqHfrxJ9fVzp60i
/lEkp+iD4hq9lqS8j1ikrhmKltKhVX4eGKDEQUajtVSoC8YdCAe+i56crYZwVBwAN926fvhbg6vC
+UpYVrM1Px8xXEuCl6L5pbo5GHo2fDqxmmq4hIEM356CnB01sLrYNelpYkfzZy3Un+BjTGFeXUPb
hWNR5iQxI3vw7J/7sDBqJ+/ChgiUSWjPQNfZWAQzT5j0BSpHg6I40ZhNEk7X233f6p/+77M/wL/p
BvQTwrKURs2PuOFPcADZSk1BH9YgjeossXhWmDtIe8BSzFM24BDZ0v+qBvycykjMsDzQMGLMxANX
lMZQ5EFtaqk6n9hK+5vqVC13O5uX3KXFjW4HTrikf+eNYoTEynVtyvTfqEHAmgEGPk0xkuyYZIK8
0dbbBYqVch40Nsq6RgIgo9HXT1I1p5JTLFW/iE3zlRfqlNbBolyqaOROCC3m6iW7oshOoCUReHg0
LvHtNDX58B00Mcj510x8HcH+jV0bY3squsyxOBjM+ZHAyh0dBIOxI36CMmNUWF8pNrn7vdiY7t2s
9wn1PlIPdCNHvk5lTS5g4ZprnP20kvtwTfdqRcXVsOEwMAQX06ciX8nbAUtQUrrAP2X/X1I4lo0v
gmYiIs7r42FpFGVEaa8cmUtOo8Kmi83QtvlYR8//TKX6xOrF1Nfui0RtfFMFO0QsHLhLrfxYx0z4
Z/LWbPPjL1EeqGuW1Nczkhpwou3lNm0LilHFdZRUT5a26hzoDdXz7wESxmm6K7cbhmEDHcsSBOwW
nGQZ9NQxst3vmpF1l50SF1PSXhHMjGtyZYouvrpDuXeTcyk1NkLQ1sKoU9igf1AYVWO7o7BL9wk+
Ucs7XjRCl1ZLUQnhMlm8XpMYJlQX9j7jpPfWNy7+9kuyvfzh33imlaxeomIniWY2AffgT03IVuVJ
wIYdj/tyPkU7xvy0ZCeZ62aj1Crx0eAWSmySfwkGE/fQM6/c0yGCNwvq6Ez+bLBx6IHKeH0lLT0R
1yCCBuh+0Rk1+aUjxpjhBEcYq12E11U9yRmX0OeLvy7g8b0WfiL2vzbkZZFtyKU/gr/SjpspIqXL
9rVwcZt8fX8zSr2OhLaOaZeb2ZRtEq26oQse2E0f1i/9OOvMI2VRz66x6GJhehEcKzpoLSzDeSZH
PV7bVgv9A07XSfxi1vpnxVvMgYfJOktyRNYTbrvKdXRYRIMWDGv7Id2HJfSBwNmxKyNPk1zZq568
KRR9vKcFZEo9SW0/RSf55R0196OwpXaigkQ0md0Fo0pyu8zbF2FKVwZl6/Mw9+uMucThlQk0+w6l
deERNwbNpbn4BBr7K6Jmd2Soov5+a8Ypx9+USSGsAcDonOVQJg9iWc1fVAPJhiVF/tbXsQ+Zg2o+
1Hae+IZP2mIYT7f3jzdrVLfjzZsHR4ttgrziGDWjkMNP2iBGWxY0E3tJ4v8jF4/XmVDXBIkN7mOT
vWaWY5qV+BNDf3ln98QbF7WtWkRlUnC2FX/zqjUtrD/o5gFHh0AXGWatAdx6U3zYZdNJuIhUUey/
YtC6966bcrY+dg+hW2XWaXrU485qCrJLuy46V+QWX2cZL6CB6zsKF5hI2FP/IL3doWEMS7ep8vQ9
BHfSn2YRlaecMHNK1ybrt615uKAaHMHQRCmqotEbmjxJvAqyJMS3+wfJxWRyRftJ0aoTI8pYSIzh
YeODuy0TC/x3sOg8GTtJWJT9MnHvtfQONYbLfJzSQPtkFK4JUTe+V35o8vd0zv0hov2jUCRbK/mv
IRFKl2PuaKvoaMfSELopaos+IX7M5QEsbxlJuZWHjSHNneeZYA3/HP+/aE/BZtP3GXQMWKi+RApZ
nQJVIVxjley/LwVcAi3ET4GBX6jTnJC/oyIqR0dgN4OrDBbBN5R5VEAJccpYeBioVB3ldklT/R9z
eDlYLAKOJuMikzrxGIdWgErTjd+TiQDbUbJzW5jYOZ8Sjbedl1x0bRfkzkTC4suEUoP9LXOS5LqC
vfbw2EfqLgvezYIYJaIzK+mwVr7D+t1XLJwOfDKyEl4eLzAWq/SbRCIhYKc9cGifxQFbEnEOApfe
sSZDllr15GpkVUQq/AGEEovYYJB5hJfYzbYa4AXDtHy/ShOxIWRjndPPdHxqX5yBzlyL2nH4qw10
K/PCFqpXwJFLk2L4tkTj4Lrc83G7AMqP05e86zkErcX9mpuMnpmSbWC7M5lE0t2FtaPd5FEbIUUm
haEF39lnCGeQttUqmk3m9xLLIVSJ6NgLhZ+EiAqGM1rkb3WNHwjQeHC49WzWmWsBbKuTqQAPmGTi
BmZsi0ke2KsXSx4QkcigEexm88UEAfVfJJ93ztVicuTPveLLqGau/xtAdgMxZJKyJV2mEwC6ExeO
FBdU+4b4TlVVrKWVMlUvYBomjf5Nu8u4BfsIHB4PR01uIHRXwBZ1XIj6vC2qvKnZXrwb295ytzCH
O6tPjDomnl3R3d8grMhO3rB63KuJIDW+rZJWQCnAR/o2fXtWiVDZkgoZ+p5tjDrQI3JUQe3ZvQzq
tNEskCOdRwfIEkFlIwhmKH3P6s1aVPXvSbntQQH9I7KjoKZOO8TnN6csR/aHy6Ueyf4FOEAEjbI6
9nl5ujEtWWpaAgpCi9MtcN83G7Q7t+yrOVttUgxmEAa6JmYfv+jRetPkS+B62FGOMdbPK1CwO1bl
RsMeNcOM1i3jsaxdhocEh6+zqBMC8i3NMcaZ6+Qb8R0J+DZ7ztItWDyD1vMKMLri+wT8cK/1vAnb
4YProOHKPqeHKmtdHphahS2tc11y+5dU7lZbwiJDfExFCzUAO4tPEwNetQadH8Rt6ZDxoo59j544
Sx4VVM0ZzIm+y6whnt5Svwc6I1RYpieK7le8xLCBOmh5cfW0Y4ts2JFKNIT2LLUJzoCEz4S0kt3K
WSFoZZjvZXS5w2wVAAi9xy3vLpXvULApbAlDyQEDdjrCTxC2qCglbx8vtYOQzC/2PNOeZirjDtb3
HtbbpQ3XmAYjp88OrtoH/GxAmVWBnNz1IdwwO1seelZO2yAi6M0DLyP1C3O2pbTXJ2i//f4Tf99i
X8jZrNIHX68r9aphQazyfENKdhts6fntXlvGSrOSBdrGRNgghwuICET6ugmEvM12Dc5rIRZS0nAK
WdAiV7rqN3wgOiJadDMwbUmg+0JjbXh5Zvj9SxZEDPFgNeqfJz8RCNFvrsWXW4L7tBT+xQCwMbMC
WeCT/3iyFxq6HPs7D2mTs4BqRWe6SqevZqqKq+onyafeK3inv7h6yOgWIqxXTJ3bI2lOrMVv6sik
p1tQK/uDtuqGtCRZATaRGSyyGlq3GOBo1Jx5fkyXYvDvcHn8AU4zzLSXDmcGbXbyFZZtbBnaHwCR
b0ItdbvuKmiNNH0uTxowGEZUPS25M2fQJh7fMrfW+qeYkDKJTl4h8eWkdz99G6aYkhAzWPZahzG0
+l5k1hm+p04K10Wa09FhiVTjVuNm3UB2Og3NzN+3VPO3qoIVmTgu4T1uhXgyu4acFA+9yoTjD4JO
9uwKqI3VMgbzxb16toqEMKTveWdAXbTwkAiT7/xXc5k92079pi0KA6pWxpo+DSfHrKS8xN5suDfR
ER3RT/xZDzbDeQHXwZtCF6SUm17mP+NEEziS/av3LQgRp976zMSU38SQ10sgHsXSfn+KIMdN9Ps2
zVN2ev2OvyvnJkrtVyamYMpuhJlYg5AINR4MWHfM6oAmLEN/hNGBkFCW5NBb5UDdIAoMrmZY/zxk
m1PlYdtRwuYGD+DAstpewZ5ehUejxRYETDxDRHHWDFNgcZjvnLFGevvI/MNq/eVobskEbwOxbNCr
ZokeTeF6qR9OItOUVQQq7DwxTkX2pqG4a7m/OzBXVo/WF96HFqqrpKTE1eggM7po97pE7g3w60Jo
68VX4c+Q6fAl9NRoYG97ydMtEJKeOcsMkYzTtQOhtmhQp79SymslJcXqJtlP4UpIT/45KpXazb29
pvFOoJVxttAxCBdqIY/ZE8MjPKtZfeaRTRlEjv8RGtGEhXRUypP5vu1Lnw3JxYtwDpJbgNCVO1tt
UnVYUArVmNkZAWKBfNsFsPek9dIedZczGn9W04kAG6/iUHEo+T7hF4i0ntePhfsApK7QrmgLlOz7
UisflMnoE7al+KCML6ulRN9mTpnPWrpmVsFGWEYX9XmYX61klNzGpvVMgRdBxwAbfFOUHpdNy4jc
HA1oBDKrOp4gKdRrkcRPJzKGWoHmtCLP+Dh7jtzjPyKL+UIB6ha6jR1+6rVwpdJzNlqtwWCqM7CF
lNHxr/qxyJt97krIu8Mp5jnKPWQf9rWLeF3R5wx2pVHs80Q7+mvQaMpKiQjvBstwPzvlkcK3336t
KqmS8nJNh74b4uGdB7RatSVpYG471bm/C/jCs3KJR77ssWd8ZfXOrcM2vCRwpxd6Vp63hr+lgyls
yOejxBDY1daHfa16UkRb8w9tgMHvkPhzUICLbsUKM3MZqmCPLTZqyIeeRwACk/jAcd3ADltXVAkz
AR0yKvla5ZaxQIACbRZz+WRMae42yvIPBNoxa6M+OBqIGYAHGylxwuyO3uxbjllGQ+8Olt9150OB
osctoUWTXQ8VFgI85OGAm3213goDdoFCUBpUUluDFEDdD991gJfpnU2msknE8a+toYl1rcD+Yw2C
jdQocYyKzpRMqw7W2F2H0RY4Py/joQEY3OmxKPHdIGmQUvl6ixc4f0eLQ0GiRRTh2YCpweZPWYgO
EAzVZoraZWY0cV8KLqkudwTD6hIGYSbeevDIDBuuZJBU9x4v/sPx/yCYgHr6i5ibGrCD0lngCuPm
OzPQeiNx/aNDS9iHesiyzVCH4kYtQ9WEUDSvjAIwZGf4ZGJEkAkFgNX5yWJ4RTY6/AxHbbXSLnN3
f99pGBYyLfcAdmzZwmDfmUibHZ5GAZTTYNiQU5Fan4uojCm8VIGMAYe42IFIuGadl7trFYHI8nSW
HDY8SKf9q7AJ47owr/l/JvDk3+QzxpLrbYNf1CveS4d+oQvDAl69kXU4dcusmYklElx2+BeAvqx4
iByKnn1wRVmQckvzh38CUwepbHD2EeNBbkYHJOU0lbj6E6VxTch0935x+TlMkAFPEQRCXZgdDzmA
QyIWJKyFXULsYft3NQ4iXEmLKplaqxj/wH0DI/OVe3hPOvA5/QsYyYNbjLTW+/SiW6e/Mif8H3AW
MFFm1jRe42IfVMV7Rb9w40BOEVlQzNlD3pGtUIFi9A9EY6YKmIeYitzOdBBCECrRg5zeclX93EYy
4cj+9US+0T2rd1+zfUiH9UpSGyHlBkjQUUIMizFhd1WrtNbnSIQGwahdoIu1tTLnPpicJkALa9P5
P2cEqgtEJguln81f/v5AZHv0Q3Ij3/SMVSygN9vF/jLp9Uwj+GxIuVbuBB9HwmKW0J2RMiZTJcNb
rCpiHQ+xzZse3s6OqkuO/eLalt6iHrpyUp3KlKFD53x+nOU9U17xxqt7kd5XeuZVzByU4hiNNs+j
roC7VfAGnJsBkc17NhHKQidc6IqQqpTNCAgpYL1MC2TDF4in1eIINbG8cLPXDzR8zcemdgvdrv2d
elmDn2oykasR2AjmNhk7mOP7NFLnQyONLgbiBwirQ3a0EJ2WAGXEbpVIcev+zEZxXs2g+8qeHxXt
28Hu26jC/FChax40I1ubAEo/66v5wQS51A9i06ake7KE2EPMb/X16sET3d2S9/L/NWeBjJTDA8xr
V+m88tMRuG4zAggT4oJWxykqYTHO0uA/9zs3YffC68f2yscOq/ZJcILrY9dcKNrxkqEbLAYjgE2Y
My7aVzSUSxZD0cl+FPdNHRcixBTuYlM9bSCze4zwHJY0nyVfLVW6RGpcirnepoozeKfhbRxcCHPZ
r3fSGVZj3ex/3AlvEbTiSq6BEdPi7cQ/Exe0BQerV4KZ9fkuyG0OD1V1YHQ95DAc+E2wWonpVhpm
ustzT4mYqDHxSUQcThDGlG6VnYSSRNxS5Aom1G8q07ouXKscvCg7FQ400ZY85al3Q7isyaeKaPDD
r2D9L1IiEOOWsjBy/yHPF+U9zGhQpREj2rfzZ4fEhBdZDHw0SQwD6eF3fDvYJunnj1UocmqvTOij
+4lMp1kWilvPbTRBLqfRshWYyXqx+Aqsrk29dJyQ76XUi/1evJXDkFiP4dbgI2EQG2wW0t1VL7jf
QMY9nvRMP1dwdfTV3nXGqCK08HrlscUCP0ROeskeoDBoC6aqiKYzI52H0RWh4RngervSLntHoDWJ
I64PBS2TZQ4kXMEJCUl6QfBdkue2wDbEKpmkfHf+C+P4hLS8QZ5oaRg4+m+SOgnoeRjiHihjFAr2
zwkeEr2UIn1ocLGihXgchwa0I2g3pMoF/bExiISuSkPclYDSsayrSgigBvEi0n1XD7cKFuVf4KfB
ZloxaqD/eg7xaZSvHLR576W8QQGl5SBtHV7qafFMj6AOx1XfDlEqFRL1TcCKpscNZTs3SuF2lHdG
P6p7T0n2GppCukYQj7cUcnmQMFntTKu4SovtMyJw+ViSnNDSo6rAKW57CgTI6/w+5joWEqgNlsSZ
5NB63DmQQozxByXOXE28rBWxUK59VR4Pn9CBWIU7RXxi76hrvfVyVRr9W1670H9hPKvdE5CSh9Vh
YG2LE6aLlwvBWl7BR/951H5AS3sKl0x1MFb0qKy5tcGi5CnbF8rdp16k5FwDX0vx3Q0G2408qisB
bwI+Wb5yEY53WBNo6h5IbhMvD0YO8v0K9xX83X+VVOZ4U34jw3fWWlGiSrUn8DJZk1VjUdn6PQus
W/Nq+3ivuLX9KTrQyg7KYKdmFsd18E4CUFKe6/XfOJxY4BOFmBD32i+xHp+xgMTy6ZSYxY6yooX5
/zBtNRYEtPLvh9UvAEPllqlntpDW/EqxCg6Hp3Hr133R2BKV2UsK2tPzAWbizJq3k/z50oRisfmT
DTheune4sVplzNv4rUWs/Y3FHUsakDQrB/dmlvJQraxh29OkgZ0eDmrL6j+yh5dVSLwu0NqvZjEv
g+SYN4rHQ9BbCDt29g1cYh9CpfDgZZkdyzU0yh79NVPPajRWNuwperlHCrAGRBkHLqvEeqN9FPZ8
zSorD6ONGP2liGfu1i7IDYbnrB5cf5LO4VcdePfA4uZt+9p6h3p/rbrfCLGv5Yfhiy9ytzvTIMsk
4UTXRFB4QAtpd8CrET/31JEQAPBCiyhb0mO11Bi+MBTlAWDw6OSop0EJXiLD1QayP+0yaqFWgDld
FD4lRrzb9uyx8/zjc6lT+hP7F4IX88ZtRiS+7qOyQ5glEdLk+G1zpMnyZUXXIriWZ/Zs2U8shrX4
Dkiwu3GmIQkW3N6zbQjysT/ywxDtVUt0GRdqjet/atlvyJNsFgNJe4HJpfYtshgzhcHHPVJhg6Wf
X/V/R8EdCFcjim4lSi17EvdBky4MZb5Ly4ogr0uEZcuKD088JeN1Gr7X61MTdPNht2Q+BO1IfioM
xTYQj1rGrdSXBHDPGcN15auU8vpWSKtWPcDK4PQi6rQv4Zosdq4+zTpyq/enI8zvMmlaUZ8i8pmi
GcOaamI1WWcwGnVLcsRE6TEtHUBrCN8O6/Pxnrar3Xp2+2Vw0TIBPThGLj0DBhkf1zOYVp2SrYNR
nDOoaLqxBDhJ+Lgv5cjDe2Tdxe22x3bg1VLvlP7l485q56FJhg5shC3b0dA7tthJ3mdnbB9ygPv6
0It7nHRZKXRdeogBrXeAYS3szHEdtSl6OobWrXnIIdwj+ZpX/GHauO2Ua1UsGtJD0e5XxwEpdaSm
QP46T+IYrWU80yQr7ykY2t+8GkDR54zArN6CUtzDO1bsmXX1dYOz3H/1LM3afXVnW0q3J9ilL1dM
8g1zc2fKwzd/RyGj8VDMcROv6UU7Ac+OYo9QjltriSdcsYuNdPehJDmXPfj9sSbhm2wy/A7jTYWR
Qz7jmmlIr+BcUStl1980aPtfGs0QxlTOntFryDFcWVUn3KPFKRFDSUPmcdKschg38vSa3e3Dx/ht
JVKvAq+tFiG7POPj+MY+95ugJTgA/aey9qFfdY1G3k1hxMak9bMq77INhxYT0yfi4lK7tdYO7EKG
49/jc7cm8AZkok6fFR4mgElo0LyeueyAArJe18ZfwJaoLJv+mN8H7ZF5OjAEaxptG7zKnNbgF6A8
B/hhgYdrgtSqnc22GPk+xvAy/0IEm/4khAptPd0Lfw61QZgzcyWsK3BsAu2uF1dxl/cf1Gg/0xli
bZpwNf0G0POssm6Az//o0B9hYCtAfYDFB9lwEnUSb8XrxuCCmFrfjKxaV+TPb2OLl3ZMJZpbIlZm
i/FpU286J4WHz4pgSZFdHE1y8seHGS8lprdCjgeCZm6qR9OYPfAJNIAo9kL3eG6O6s7UspIfibIH
UEGOQtJkjf7sO7yA3fpE+pgL79z1YWBMG2Ux1V7o7ryxKKIYNGLrsnZvMyBmTN1Di9hn+1gAF7Cq
1yhBbJZ03GauXPmdRiWxmfuzde5debcp+EivM+7l7Y0qwXBiZoHFyM1Bd2H1D1IlR4ioQB4Y/mCu
2sB1L1P3iY4GMC0sHjJWMLCj3DD9iWYqNgnA34Gp73EYm6lctfNvTqAAoGJ7HNYozr1dxjG6EJ4J
oAun9uX4eFyCRtBekSVgkjBHFTV+uz+mF0OSLbElfHAq3vAk77RFFWB42iX4lV/uozyfdjuvy0GR
yc5PtLYMIQIrcuwpsyETORFdyqZf4RavQLICdo56KD85gNhZ0EezKVdCQjipJfpFKHtfcXDHV3+h
7m1NZJFJB9fUKQMe+VLHWrRaeG3xELqAurkyxmxNpiSz0FDHTRakNQ5V6Fddyz0YY4DdiNlQPklf
wxZAyKckL4UUSIlEhVHrKusVV0VZIi3u1BxQGZ4v0GlgDBX7cgNyD+ZqdnBYmwznnOB+nBqtYP9W
ZMJ+5QN+smojwEKa7upSWKgkFW3P2CsViXZwwBt7jPDULohbFQw1of3qC8HvhwKwZCOOerwmmDyM
X62AZfPq0DhYo/3ctHn6kMJAceaOa0cqTETmH+RpoRzcLyjI6oibAO9T2vMhn60LQnyEMXYchdIC
rdxb3G4T5UypISd1JaeSW5B1JayBgZ794AZ9DkwPQWMC0V3Yc1UzZKCSDw39LojBjzimdDovNUSY
kGnLOE8DDK573L6Zx01DMHJH/l8Su69BRX7XKk67nysmbvnl/aA0gV8BQ9VDSlXXx2x/V/4M7BoA
t2yPS2et2I9rw2ZCa7droa5Kwjfgjhe4zPjWL/Gbe0ireSiwlzm8p1LDGqijiEKFRJo+vi8HPR2O
R8HuA+1As4EeBEgkjMmufrSAPjAX+yE84AdvlvLHqQBiO+R73d5bpxppmQJUrIYMql/eXD6KusQh
u9HkdRdONZUeH1GQ+0SS7W/Sf7q0txpYM5qfuZtEpCTrX2vC3ix+tPY/1dCDjbd2SnI9/XRqQ4DT
yELWUvad1CY+H+sQs+3OzH3ZF15rn4p9G+2hiI3JG72VUEM8irwL9cZM6RToPX0P4O0kmtrXaTe9
uLqKaCRAQbjE2y/px7jB3BfRig2onOF+nlHFRAYanDdA5AvYtksiBnyZz3oRs+K3UxzMD7w6apyF
mafi5l/eeIhHH7z02j6e3KUgW0Muun7OAJRyCGGMWNl2RZLUMzF+uonLQHHua1pspGwmC/RbEy8Z
Qe7Kg+p1/Z5Rv66JR9DR2mSkavu67BODLdM581WP99Vluf+44yYhMx1zqPYWnHjz3RvC5mun+vMO
iXlI2DpwgZkdPLEBFhB1/uwNiPHghr0yhy8ucwf7PC7g2Ybh/g4FBnFjXlX388G75+3NapFf63qX
NPetooE/Jaa8HT5KN3dkeRAZNfkDMG6pPYthf/V3gO91fGFmDuCFXQz/jjGhUII0yx5c8w0dYzV2
jvKbdEhlWeMGlFaBwSiUjpMaiQruPBByP3XwDjR9mIeQ3EEZJzgfFRWgR6OdVmJKIrP3XRvmN3lk
h+LJUn1lEx8kZka9K9sNFY85OwGBvD/FlfShuKLGiIgSk9nVowFsFhJONJt0gN+2luYljZdndSyD
lO+lZhTETIyaRAq5ByFe99nc/RV922cjB3WykwNtOFb97L5J2KnjLd0Flyj6bMiauKH1grQONCd/
lPU1nmowDvn0LTGonS/ex7eIayEcaKoVmUMz2xIq3N9Fv369kKN7m2N6vCu6Wpxb5FoqYNyMcwWt
zbZoL6UFvIVF50SXiYcOiSSxiSz1OlebdhJd7Gu9noxrGc45Xnuvy/j+fPX71NwRKfiNnqAlhvyb
ZLMUE40H9GQ53zdqO8cWwjMXGf3ov/n1YFw0+kLVdidR1RVWIMFO2V4eGzUj1T83W43CtX3H9rcL
ofPaLv6IztKTtNK/tJBCQ/EUqgRBIOoKmyDMeiuul97nZJQWeHVw1MiAj5fpW4CYiN7cD6zoPkfZ
YKG0TD3gsThJrxyHzxiNQrWdU7uc/kAtIudjRxxsnWu7Mv3HoXhVKq5HIdXDBT567ouPFXX5RIBF
LyqLonA6eC8xzP90M5Iic1iqcORHFuVB4GSFlQyPoN5Mk6QCWHHSJEEjOWfmPJZLUU7bjLIwQeXT
Soqq00j1pZc99nLA2dlCqLpBdgW+j0rrjHQ1XEhfIj2jZmNLbBuEX7pfCsRKb0+bUNBYSyMMl4QT
XZU0bMf7DeJxoVot84BiFdVUbS1vciQrZZSn6qIWG5lN5i9xYcujT2LjEf0I8oaiAm63UP2UVaYJ
YrZp5VOaVqA9T1zIXAeaO604R40yjO4L3m4zvjQ2LSIZTvscr1ITedLtv3W6WHkCpbMlYt7lJ6uO
H+2G0btwnhDNAm85WUexyflcbyDZpSTRqZ3D+EYxc+ew7kIzdxnWy6q3BaYxouFd5QbTVtGtQbzQ
ZRpnOuSDRqyVMICBczy/sXOuZYJ1AURKHe/AB5vjOY+Qxxsow3X8NUTYFZnn7eV+pwpoOQNwNAip
KY9YDn84NildsC2hFUJJaPhDwzEqKIhznYNMClYB8U//Q1S4wGmgtRorBhe60/wFgCbRgXvZitNT
YNZ0tax4JX8dFAVz9SZBTfZHV2HBByAT9/xkRnIH3DacCuagKAsps/xTug/vqgOOnAtArLiUnNd7
a7hLHm3G5IiUE3zAWaPNV8wBppJX1Ca1nn6R5HhTmUOdgan5SbG8ufWZ70cDeQXrOXsWDtQPWnAr
Af6nKCoxo2sdPqO5cXQLvy0vHizrtD1vcgHthBSfCauM5fCRKSwcrR6XQtrSNGiretsGODJbYYRk
EgixpRtpysdQR6Hn3vSWy/9g8OmY6p0h6dLZxSckhg+py1miD44c7L49sWcYDJ4OPgtrubxnFpd9
27nTxBV5lWp0tBSBEgM4WngRzCb5JVXRacaizhAirRy05/5AyFiiJyUEyBx2PzEUCiqcAGJd0tFo
7UeY6FzP5U0zqDGhUvpkJMcktEl4Ck5l+H2fYLroRLSn4JrmaSYkz+7Pi1Ff7T9iDFHHbq+i+EKH
49SooCur7oFVK2ipAYtVlikLVMr9yUpnU/RjCDQZudIQE1RH8M1b9e3ErQ9PbvNNqhbZPJjUalaH
AoYnN56CA4bn9BfrAxRGBcSw3fR60SusmqxxN4Yzx1D5X6oeOKspgNmk+v/A4MS3gvcgQiHLt2oS
M14WVOfQr1u61iFDle4My0ncMLO2ePRMI5tkXbkqk8toddutBEF2U5XpqEhI1BYpd3ZQa0wl6yEB
ikbDeDVXu5GJWkQHhhvn1HUovfWxCrhevid+ZMvUBTq94X3Fm6JDdmsz2YT69qww//ncT0apPcej
AddHdtVrLNL5FzKv633lfyFqZkSTzcoWV5J9r/Qw5cwrqVDbikOxwY+8ObnlDQ92R/Cjsuz2uYQH
23ldYHXDPNXE31Gd6bfdZSZL17es5+nt56uZ4hBllGuXYPFni2ph2URSrquYXIsL4pUdLEfPoewD
Zl2eYzoru8uKobHmndMvlN1C1mJi++cHo3ryYvktdK7ORrIf5S9R6xQtMnPrUOgEo0rEVBbBkiCz
8RB1D/5QqFcUvWjA/UUwfhcUA8r2eBkgfPhyhZmfJXYM0ueHSp2DiuVQ8kpgiIQdDBT/WYfxZOP2
iwVym0f0hSw4tbYuaqRunwdbTlJNjQxLUU9K674uHdFDueC2tkGTYuHvU3UkRcddFyPUzQgW1u5M
DaEJ1xgZIiq29jHc5OlWDYK+OfBd+/Wzab7DpDof3fljU+HXF4jz8hr0wqRmLvrc6cL22QEkATLl
4waEjojBMXTkF6epJ66pnX8Q4E6vtvWPn1VE/LDh6Xfy04xz4VMDliqmXmh6G806YQ3Nq3Wutf8d
OTmFtpTDdDfxM3eHprcSHpGO0CqIiRtd6UEWIh+tBYQodZca88/tlfHMx3klOi8RwwpCw2eTRvNt
sxiZ8kixNdWcJWNp5mFz44e2wUCOknrRev9gX7tZ6DF9Kh5J45EqT9PVNc+cmu0tvscACNUJ0y74
3sUW3H6pAiwBiskotIY0/ds4TVirSkJ5jlnAAIm+BF7Y8jpgyU6GKq+/X3b90Yk4JL7eoZDMTtGl
Yn3h1JzjUummr64Zo23Rnvl1UNsMeeviO2quViyVBPxM8C5aIZ/sBKZ/+RFccy+GsKAHATepyLp8
jxQ/b9YKI8T9EeFT7VIZlZ0HFNq5bYXtqmXdo3WYRKOGr3qH3JrK8KBuQRkmG6wp6PIp7ho7Mg0M
cybvGrz8gvlO7tM+xez97HXUYRsBQQdTGqYY9/Hd3EJPD17hvHU+0Icrfm3PMyOqRKE8K7z6Z9Eo
tbw3AfrCQhaXwRIprOY67ni9pAONrRhf7xANKvrFP7B/MGmwFDJ42IaH6OMgmBrt8b/x0OHohTiw
RY0o3Wv2Q5U5gbzgqzvByopkQr2wrqp22KcpR5wUfEgryNrg7qN0TaAtHB1+cudGHVwiC18zOZ1q
JENU6ffVFCyjuQEllNx5wYYfwCSFjUUPQmhqFb5eO1Q0LLKIAefcNledoeaEcQxL1WTLCfpcLday
K20GYGQTFKGCkerob+ucc9zpT8NOfM5NsYnfpiS0hD1RS6ok1M3bjH1Yjdbrt6FGYPkjPPNpbP3b
MpUhk46cvqr9SQezwT2qrThtKAktbVQhvtQi9niTUyeBJ4lBQvTA+f8EVciOFOsryFV1poQaWZIR
zUUt9QF+D8gc772y45MD27/gs3Z2pmvoY4/8t0W3FtY+FP/va3iikCFvMONZ2sAm0Xl+nI6m1ugA
xooSJCVDeqq6A+ojZsaVZu9W9qyuOe1I0IjRR0MpI0J7DZvAJ2ouGXxRuSt2IFhj97H/x5dhRO74
aDG/9NKjESCakUhzczsbnHvOE/QucLOAv4wwldlahWARurftMoJ+IGCXYLnNnt852rDdinh+VzWB
B7lfY1wA30SH9ApMzGsj5jp4Z3P2OzGsinScSJqCXhYpFpwOakpg9GARRh43imftuAnjpGe9v2Rc
wgS2XkOoukXhdTcLfCRCHvbSQWlvvwv0yffBsely7itZC41ThWkLTAb+ck71BJnfvYxrOv6UWxfB
uK+S/jOzgEUOBnGAAPwYo+Q4U/U9QZ9DeH16H1F0zH5bRfr43DdlteAENLpjMX267TgDNTR9p5l3
uK0HgaUi1f4Jh/LYN/7vOxYHUm7+kEkN2UczZ0s8e/yc8zOVYJW6JK5TYtu4PZHBuzXxA40EUKhf
YEzD7DlwKwhKV8gxpuA8FXSvwzA7RMpOzBKtTpmBX+VPyIEUK608Be0aPnTiIW6xY03iRy+F3tRw
W8meDiJK9Gn4+k1Vu5iKwovmvQ5BDMxvZib4Tlq0R2xah4gVyAEigzm2JpWH3WAEQ9gl/mAuYR2j
xyuXBkjvoOKqRVbEdCaDSnYYhycaCBv8h3KKy4DbltvEcAbC0UJtyWcjs6H7Ey5lStKmea//yxIu
x24oWjNVfKDNjHMuEVUEyOVJkHV9qB6jh+wyE5iQoo0g9Q/j8m1uZddKDu4TLW4eufFak5apeuHR
cRMhtmFR5e3qSnCR6jnK+DAJPjL7QSOsWYxEbEwqG2K+SjJJ9Ny7h9HJRTIhxKmhZqvwLQDsD7pI
FJLfwplr+5hZ69uunWC1X1R+ZvPZzGyeBUupGj8BzcbLzsxOymn2iBev34T7oXZYASqxT2lA+z4k
lf0SeYgSKSi2F9trCybAYXGuj+XO0xs3IsuVy4QqEx/N+YkH5nmX+ziW1EWroOLDcyonjNapyXLv
HSrrF7aLbleygqXV55AUnSaV03vYJiUb1Hpu071NDzgpMduJehfsOE6gfiznn5sS1KF/Wx9itH5y
LFRgCZU/na7tdGI0pC9DSO6rH3Fta4HHuweQzQoU4v9GYgmpTHV4ZIjDMFgcYuPFDt0xixH1Lhzo
rkgvKpZH2m5yM47N2fCCSgAj19JLA4zHzMm0B1QNKaXKuQ2hMVwZB4jsiUTi6q+wdffxbpzypgCq
gWyZ02i8VEyJm5EJfRfNfQ915pSeWNxg+eRkh1tsn36Qpm8wf8zM9z5s5YjkDnf5EMe1/hENQ8NE
7p90eQoonGzp3qzuAskOfML5UCThOZUCbInF/jcH6dkb7uMuwLFeBegi+u8WZpWoyf5TxP9T2XjS
d8IeQYrcX6DBWs7JHAPV8UTMzoU6SLl1wXOyrHGrIMi09wNDfRw1Rifd8439p78Go6CWyspulZyK
nrreuAvnwGikucUrElIPaQisJYA/u+Y664CyU48btdUEi2R7jm7PF9Ze5Er9DWgcgqtwEJQcVHOi
fhTGmpUeWDx+UKOWbKcbQtePYUrSS00l3bAtYWE7arwkQd1ErFaXr/kFFkdyvSi7wTSku114XmI2
nvMbGS0sqAhtPtqZFyRRscToruBikHdg0jEW/XMzksZc8F3rfpTE6WGTm6ODngcr7eSOVzBfa4G1
Xh+ligxEugbpyyonDZdJRqLqjf7mRYtV/3Zx2mywaZYaj4g49isKdNGJYDNFm4XYetSMeuZMjftF
dmhdzSOqWx+GQj6claApJnk4b9pYgiGXc5t4/ulpP4oedUaxNsBmGNqpPzFDfkWjZu7b5GoPAHOT
tAZrG/XMDnKC3m0G7SSZLW2svELte06Taxw4dXC33nHjN+ZJSmsuZ8MLl7GNGHYnIQ5g8BTNyKzJ
fqqwnHYEUF+NOWlrhLBNGCgwxQRjJvZkeuitwgHYwdp05Tw2kxJzCrbP6/WY/iRt/w6F6rSA0N1O
cjzM51cJf+bdAqeKF4vSYq7APJxpmsftk9jXZ+1oHPvLbNPlcP1q+X7nqdo0S2cgPTvO67pSAf0R
Y2h0mH83a6RAapAZrCzoOZCqwMElTPbEOsH9vr/nF3nlkdv5rvCNR5xYbgVUJMVs3BqJIknIYBBC
ariJzLA3Wd1QDkIwwXUV5FroSKhL+FQUxr8H4c7ex5GfD+xDbRHPIcegQnbbbPd+TSG1iiQhQF30
H4XX/sYG2F1ND1MT3e7/sKmzPAGX0g2apEoc0m3xtS2M26Ra4HrYaqIyr7Pc40jrPczpiWKmGgOJ
bHeruYX1ugwqXu51xNBuqymS4qrdP/ghDdeS2a8iKNB0vzW9K9+fvnguchQwPNzQoSGf7SleNhvC
kY5vnMcvtb0ZYpnuTxxsHE4METxEu43BHwriU2Pldnd9IEo0OLTUNg2fH5vTf48YTRdfU+f9JI2s
t3snCORXAlYQ42LPR5I2IFXv9MITT7+/MGJOk3atpFXNCAn2UvP0OeO3McF4JuMXyY1gNg0/PHXp
L7eEv9oNVtBM2dnTVgAI1/qobAj04I+VTNJrZu4Q4A6B6vyGJk65iz1LygdL5mrtXdAwyL8zahkR
PwZ38BHzyQE2GJOnPvK454Huo6QG5lXOBJER56uqfy1VfHaIm0FMRHb3TVjRz9vFLd+EB8glUb+2
H/4rZ3gL9fnr8Se9tFqJ89N9UMmZ9WYcXn2W3pQJGUFxy7wauH1IL5MtkSr+FR53F91X9DhR2eJo
9eCznSEbGBwA73CKG7kTrc1TdqWqUYRShOfo3MgEbuyUzZeXfKhKq0HlrVf9FOtltEUVFfnbdKgI
00SRBD0jWAS9qstfO/BjKJ/m0AIjENAqHCkct7InB8cF7FxZKa3GVJU25NcJtxDId+IUSZvJHIrF
85sbYEKEMvgjevftU8or66WDFv8pT0liJ3Dm7rxWNpeNJyaxktCaJHEGoT0LIOTC6D99WbAHEW2q
BLaGgZFVRLQA9IT3tOTR/+Qu15sqbq+XzJSat6NLdXk5MvGhYtaUHP5pwih8SttdKiKPQ1DSdGa/
dKgeoRG8O7nFhjEyTm8ZKkq3Lyt0GffioQMa9Tfhgf1C44A7e+KO6p3DcJMTosIaxTtJVp/IO3CL
8XxqF4OkM7G7wFHzuklSNAdsvl2dx0t96I6IpCmGJ5hLz4D21cxvG2WTdjA4KZx1F5c46IlgXw3G
MT9kAqtC+bMnnOpCGqTiPqMd6MHcN49N6Khllo3fPuJsu0B/BeM6YEVJA/BQdhrLYimEhtE1HZ5U
uhHebg4TgnuIhI0sKhPVD6XqgGWiJJkOBtGhXwmD/hOUY0pY5/o3F5UWK95P49JTTAQJbnRGjTmD
zApXBaIzyQqvug0FOm+PPTE9BhNOjQ0LirTGQNKSWUD3CD4iwQ8CTBJyyMnYvcsfOrlQW9rNn6E/
WQdoBCah78c/H4yUw0ZrUxbVxSL//w1lgpYrLnk75NhzkPOVd2g1TV6ZHP/XbE7kX9PC9TmEGTQ9
UKu/Mle0WaIgCrrE9+Zo7Je/nrTIKSUkZ5vgVFKWhkVzAHu41tCAtgVPIhqQhWDGmae/luDVMSc5
sLi3wqYXUdyTpXUBzpRtFpzwDFE5j+Ico3QmXRPsZwwXwDjJK9vAnW0ZcemgMwvgvMwqYvteHQVX
pACyu7IZqJSgdc0vsMeeRDBBt1uPl+SJZKvXRYE9WMqPRzELqDlton4fzhKOzPitKC6NyHFd/WmF
AFYkUOoMijdR+dzRnd8VhGpcgWXsK+rcYYQ7tkVk9TBuVVE6F83FxK2YEbrH/GRnrPCp0s0z/Zlq
6T+kgVJVnh/2G4NJtEbn2NvdkPMBklB9C91YIQjve6rCC3k8qw5QUlu9EGe+ih3iyaZj67rSuicy
8/pFhXdogRiQUH3EBe7I5PbfFtxHaMupFQhAwxtUvqr3KQrheOUfviATrO4RO1K27rijyOZ2n/eD
iEGS+wxeqpf4lTR9KbOfETpvtidtbfUSi5e2/uXloMkrt0JtzbKlN17yeWfpVnY+OG9lVU+6OY4H
APEtYBchmmJrgtEqEXfnVTQpIfaDC6Bekdm8Riz0autPEMDFf8zivY/gqM5BVhK4W19lweng9puV
xo7/XDm+koBpdgseb7qv532qKfHAk7JFC+JimNnBf7d0Mg2/cK4dDCZSItXHeYwChqOsK3LJLG1G
rRhch0ObC11FzfnwQV5vr8TBygvkLaBXTpvQca6wI4MhOiGAwtpPsVvmFjnTp6g3ImuHqT53Qka0
QIkBpviZWwteMhSUMOofuIo3LSZjyhY8aWrewIgDhTgEds3IhYZmf/xNto4KfPl3DdDJEqGlS91U
IcKaUC8OmdQLUrw7a2eXBOUABKV1l9o1mK7AkCF+O+M79Q8aPoBmoaCYr3Z4KyKoafElyi5zsaFp
7ZONSL3HkDHDDh5wCL1hKvun98nXeeFG9TgcbjCKZbYnQMveZ4GVgeZyoHkeZO5v1C1+Iz7SIGeu
X2lmD/ZdXsMhzm8IjAPt8o0Q1DUB9F0xhAcEYTJlSnrkLkiRw2pfhF+QRcwiRM8CeUncVlVYiAe3
VpZtZcwmRgtPdDsIrxDU5U98aQ4ucci393I38s0d+2cddMzX3smRq923S80D3Gxe1WnWQfZu+L/K
mKhNgyCqz+c21+25fNaTWj0fBNtfZs9+XrmSgSqGpWQwx+tbExlVwgO9cCyHE3/i1m3SXT/g0yxc
1bdn5z1JdShHPCIMzMujAeV7+tz+ulg/OmPo8+7DGKtgHPm6GprlDOjj3cym7Iv8gcM0mgIRBR6s
eWk5WZDrqmyrNbYNdKMfIPVlh8Xo1YrD/PNa2RebXMgGgN2z5aNc1bBlaDZtvc+6TClbfHcDA/O5
GkNZC9qbzKGVUlgvX+JnQR70tBw6joo6wOWIvQt4hb4g8CqVIUp95m/lrPbX33HPCuUPsL7AgRZp
LokrdFlb9D+58YIdHJUTQUv94+oOVVruhXXGqekn9ibhipPl6ikW8Eq+NAOxEmMpaE6e7DPaPQdM
thxgIQuFKKWSyguaHtLyNTY1qYrZzb/Mk45UF/UCWcyZDQ63yV6s8iXAul5bFXueUeNVoXlUKEYu
xYdg1uOBny0lKskPx8kddHYta4doQXdVhQy47f22fUjyyMp8T+UaMAV44eEJP4Q7oRyBcQZbJiOK
ISpi9jkuOLx6Q427q7vuTk9KJsoMt5PeRWS9WiwXUr6AObcsi6P/VDeuB6Gu6v2GwiBpRWkE8I0i
WLAZ7l6hZeaUEIpBA/kFJmfCnpD6tdxoduASgkCewTQdN/G9ScjAgKmPpbmKZ2ojkwuXS1e3DI/5
XzFABmgCDPIgr9+rDr/Qlcw2sGSf74rf1dWoHXwFvsZxQ1VpWO/xk1pG+cIqhTORP7TqD08ObC6A
L0g3V7n/lUUJcReI7uOku8WnJH8qALGupXc9/NDgcD2NopWQNnauWYH6HHrLz8YA+QjFoNYL8ag1
HnpXKSBKPQ5dkK58lWvdi5jmQn1oqgIkMTw1EI/9qZwlDozW+Fn5TBty2sMURTW3RsEj2zBvDGHK
dOrBq/OIiTkSp831Xphmm23473HciUejHgAaEZFc5yQFK2PK/GKwRf274cdhyJmvlzq/FASTyNUb
/zF0+t7ckjU80MMWOfVuZGWutSHmGWonwv4OXMqI172oX/27mAwCdR5vOe1TtoccLq45PXiRL1Bw
xp5PEJqQGFacW6RvVOUFIhsanpqUocvq39E5aOltxguWEpVWn9m6by7NcQORpJC5Vv0RLALBkGcu
D/6fv+WJiM3BJ2FjY1NdJURc2tC+j8+SFzvSZPDG9pdOciuRJn5ZEXkAd83pWacDEa1seuMpGI/L
1uyYkzBceE9cb/XL9W49K95phGrqSL57BIPu0r5gXoOPPrEj8sbjOkUhSl7m+AnWsZ5aA/zGfPjB
G+pW4iYYNBYOU8QU52f6BU1rFNcT+Ok45Foxe0b5vEGUM1XCGlKweeb9L3Enm1xyJdYNMKJiAbRb
lIL57s7KpZPVJuGHevyBdP31vOHD7z0lXnTx8KkV8/b39TU4BZLpPP7AoDk5sLfMmwJUwtl8WAh4
XCtItKN1OZa7RwlEM2PwnSRBIIWY2EMV85j3mkn3j1hmmxszGJdHtRvldNl/FCPlrJOt3rl2DElj
HN/vwUh+Qo49svKeyKm3kXV/tRjvL8PSqc9ptLumAIq2LA2WW01te9kYyX1vGePv5t+lGtqhFKLc
yEw6PIWnrbPRAW24pi6SvywY76jq1JkBW1PrwqoYH+1S0pP4NUfmvC+Ax+qf0Kt6oS2E1vP3lEuE
zi6YRz9r9fCLo84Lj2Vdo1VWwlL8xCUX/YYTZwsZ7nP7Fs3sTSw+K55ggcdJOEX06JFrUgKHF9Dw
/OPFUEMbctTD5L5BS7qpVwSzsj7pMs2KZSKtZc9nD7bjR7It+poiVRtRd5Sr/DxeHfZ9nSbSSa0y
c7BN8C1+RTt9lT25ytCaojRjqUpOAiuailpztEPq3EPIE2FmeGYZDdYJzxdk1TJIbZmsQJxfAkEU
dAXX4q/5DoJSr1o2b8SsizPVLte9aLIwoOwGImpbO5EUGOA8+4O54+b74qNNG9NLlskHCpPFLOI0
gMdowrQqZVRl4Sy2L6LWe76IfC2MEhvuz+YCioSaJE0CssiTe4cP0oQirvkEc+8rxloe1y8Q/JYj
o1PkG761qtYSTKpkfXhV/nUnQObQOs5N2uxhQ/UqAeCNTdeBBT5IJ1TCwjk1RCbNh5pTotYHtRtS
/15hCE7TuMQVKqJ92F5cVxTzQXG+DyN+tz+bLeTg1xD7rPhSJSybSSaKkAjrKVvDbDznnI5+8hu5
nZv+EMQxbX6Gkb1XMDh2L5OrhPK07UlllVQmyTFrHarqnDtEj7ekLtZhpidIsXKAOjRag02IyKn7
D7TXfPxD3LOfiz7R44LCVhHPaKEorVye8K4EQvPOcDB1lBGd73aLGFCcRymXGOjD5WRwcLya2yqr
cAJvsE8C8fKrkGieUn7AiiaATBVOjtPykU3/02YGsVOqJmTIxD7VIIWIhOAckUHXkhWCS+73qubz
SNVXm5JSUJOGK2i+RQMjjvWmQUlBtdAyr6hdHEpQd130t4ISCSkjNBtcg8KdyryPuh2XzWZP0o/0
Egl9yDRmTM8iB2O4FLlmH0DkIlSSsbsVyjywktRZNZel1c2EtJFjDYqT3aYrJeRlyRuv6st0th7C
FVk4w/QDIl/AfQZ57qKnWc+2pAeLsCi/kZk2w8/16/lkC/v49zzhIQ0NiVJXW2g7F5OMtdE69/N6
EvFA04MKn7EA+rmf60Dbi0Gpa/bSa9ZZREk9+nQlWarqjSbYNwIRzG98O9+xaZo8wdqIyiquS/AI
Ierpaks+jIEuiMFnNAXxH7Ke6tN4VLIxMH6E4QEpIeIRRgq+ZGyZVysmmp+S2sz5hq0/E28FPqLa
LnGpl3Sg3IZBWxsxpLOCt+WMUZ1zhTGV+qgyGul7VAUg7F3mAlJa3ocL1hjbj6ALNijQsKkFuAiB
lSgKwi5iG0S/VImpM/dg+zV1h61ejFcrEhYKGImlM5pLdIipS9/GGCThDU9QE8DXvjDOx+Ovoo1J
575/TLgJ1IZbhb6yINk3///0FfBZt5I2Dk117at5LKcXhtxCLlkvXGzwdp3tEP6P6vUEvXhRBLuc
lWG6hHgOfm3hpdCgffVVXYd9IIJ0RLJN/3H92omsS7K3DgjxaWgr9iv4JMpK61XuCFYBvulGqfOs
bEZqlbHufLH/bktlsyTUqlZrlEkpPH+BnquOXBbdTZVoJtqKRVY+ifW/k56/dHNeLWlWsWR+N3+w
ld1e5+ZyqvcTYmdKHBPEkpUX2GtilDHQiIZ2YxN2ba9gtI+YDrSCgpMErbv4+JKRQJLJ3z6QGVtD
QUkb73P6LNa1E2G1SRFWeQvE0MMoJWVQVPqTmFUQ+fnx51i1t2B+YLiA3o4cb3Lpz5bRQXpRb8Pk
bvCQAWc/3yXy/ZdA0AAVbKg6923lKUEP9/D3vpG6wVOh4OsyzHkO+YCacDUylvSErTuQDEEG4ZEJ
ey6BxY4Q7X1bV6l2+ihkLYVd3v9bXc6Z9/LYCsGT0ik/I4+BQLhMqJzQDfNe7+M6a6iVwmM7fh98
Zis2Bef7BeVM2Xet6TrPQ4/5Ev0huajWjIq5KDSDYR7pzqgu85xfmnfjOUkTKJxGWQI+2g9ByD0L
Gghle40zaoC2ac/0NBQkH2eU+1lnn+4YEQfzsYNJU+VktZPDaPYJITKpIkgM1RQrQviSCFpCy7lN
gB0mmDQrZGW7UQJBwQXuYFD9XSCG/ig1tgAe3322dliYOvC04gUyxeSBeasBORZwwb8DzxLywmQp
wu3msV3cCIfIDBkU7qCwy1D8DAGADS/CX86VwSn6Ie/3/a8Rb86E065ehpSrVZmoYX9E9iSb62Np
F6Jict81K8oKE1pn85hP/OTX9nYtTL91QNmqxSJo6aG/19mAKz5c0cGN3wamYxDBgH3KtHOhrZgA
n7aVu8x0aM/aHn0QO0ku3dB9GhlY+jL6qWrhZD3BR3XbQbdL+rPbrUuVYK3K5BK6ZAa2sOOQXUAq
rnXuOzofr1wGXB2/UPqXNep+WD8idbCFAvQ8rHeKirsQjI83xoPtkviSlrPKgb7/0f+IGXds/Xl4
/Ypt5r3Gfjer5C5tZt5dLiq8+FXePF2jfBIKYRvc16LpeCm8MDGdRlfrHgLgN0pcDeYKpHcAmqIo
Op60qpoH4ELjfT92xwv49AXYHK2a8wAQzRax7UUaGwor2zokd4L3kVNDX4mP4urr4xRYTVUyb8f/
IoJopFdeJ2pFjQ/esie7bkbid6Cf2a0K+d5rgSqMH5dexA/lQVYaZCKbBdbu9k1SoWwbWUs5rmbD
d/eWS66ZE6X0RLBk8D7uLxUMxN7UfvN+wX534TUmoxPREEaEXN4B4HzcJueQbo6yaC+tngJ8gdAu
6FGFcfTQcAbN2IW0FhE9GZ4pzvYT+oqkOnxLH9HfzCWXeSeNnlylaKNIkidp5en642TJ6qaBSIR5
mnPexNy1ClN4AKctTb/6ixUEKoLRajsCJmAYHkyyJo7/zdcTcKS0FLe8xHDBXeondSL8V9YuXqUZ
lempScASalSz7kz7Gi+eeHK8fGbCy0LJTFZlvJi8AzJhfdIRJwFtD9BEN/rTTkp8jhvhIfjBRzs6
rgcsYPSacIp5kFVqEdRLuMwSUJ/zyaEuJZy/MLwIP74kfALKs7xrVJVYrt40YPYwpp5DCnFE1RTP
y0lR5ld/EB0mkGvuTWfnQzC0y4GOVQPMzrM9IUc3IY2ieD+DjlDvOgsOl0Eze4qPgaySoXWMCdLe
BnRasqZG/d80109kXpA5Cwjdi4+CwLBVGTfBJg8RgXE7S611QTdOwbX2QeBFOAVE7TjFNz+aQDpv
M/kgUzo4oBzdZxdBEGraQY9fksEA7g5hYOpXFOo4E2N+Q9KpubOQ2q8GgsWXbGvqjfL9aUUY0fOL
OaRqfUFBHpZYfbFVPolJlsW/NfGmjl4RalwO0ByOb/pzlUJs/DOBwzDa0set2nUBdiZEVHOXUE2t
pPVCRB3JS2Y5ZGFJKl5raP0sVI/y4wcppk0rDMdiDNPSetLiizP7343H1xIVCOwOIH8lpHn2evbb
xs4XmiNSY/C/XTV+rvA+DFDIY/IHyVG0hPJCi4vtbwKgcEwO3nrYMHaGFJH5OD0ZMje6k31iL7z4
STguBqFcWluquSeqc1nEtn+ISYW8SFhZt3MBzBUslnq1aX6/LqckJb1x88dnTyexslEkuiH2aVoj
QNzBkDQV0p9InYLqyt9H034Q2jDa+enKmzBp7jVBHyTZr8dz+p0scUmB9khMAMcl7QFO6BY5gEE+
3I9J60VOLC44U9sTm5hEwa3Th/1hgvpLjwX70SBi6sVkipH0uMQI7RYxNnMnTzqI701QnIxXUG5t
wM8dix1TMOQPqjRyX8DG/oK7OoIqWCqYSWRYwmtk371cGxhb9hR3C2LzY5pT90WsoYAS9jJ/vTmC
pJp5fT+zkOQcjlJqJMEm9g1+UbC4lEupbF3nFVs1nxs+mMbqwXVBbXoS8Ty0NdROclo9qYx+sq48
1ZqYjIcNQYi+jIo3Sx1lsclp95v2AdzPgsiBXCdGnJmImGx5wikn+5BgTqUmVjUe5LBL4f+rwJkF
oasiN2yTVXGbrgkJ937cwAmeX97GwIbAoLJvEv2VX9TWdbLSINlbL6SvunmLV6Qw758RuCQ5121h
Bm9buJnoIF3JPH1e+x+tf3GCvrQJGN5N/8jY9Qkhat2kol/1rNFwHof8dIqir01xsnC1oLuFa2wF
6billPzqOF5qfMq4Ddxch2xzrcpvFDBZvPf/d8Y+PJSLSCLd4sOZ/54qCyqmEkSjgdni6XVbHk0A
lOXV2ZbnLbhpeGRuK4sXLibFoCFC+TBQIAwdA8+N5mKObBG5/8BtM25hgz5mmMDF+dzDouRLf0L/
UIgRytcy5CzyaBclIbutaNkR+W0ElkDUU44JTP/+pwOGB3T4zeLOeD2hUCqTApOr9BpInSLcdHnr
gLJSu0y9Oow+VOHhPvo3cNt5N+8k/yPHy55FTX2EqKVr6AXLfwRf8cpJNBA237pOB0SAuOR5MUS9
6dDBiCDN1NoNIi8r8l3q7WnVAl9DVz5bY+BquS9VgCsdUe0cnjyAH75+eiav35piJ99Q8s3BeM9Q
fxyRoQwa2d1V6+muiBKPMMP9xpJc0oZ/+e+diXUJcSugVIjLjs2FjLT2bu3JupIAeTLtCUR7plsZ
pSdhvKBB6HUvvkWXmOMzeCeFSzmRVmy7BxBUSNv4mBJZygvFwxZi3xzZrP0w/kwL/XYCCCnamk6t
HyYg+UWKH55St6FAsrXSEciMIEI3897hln90OECgWTpuCWZHX/58AScQSxL1l+eozEeAh/TnSTY/
dlU6uNIYqpByApQxnZ3emuzo8wFxd0DvC2sqTx5n6Uct7w+m1dQBu7d3VnGLNW8z1qKnEj8J3hkE
5hN1bk2JuTi/KlyvJwqw/A1dJAqSFF2p3tTBz82IgRHgLxFfXztzgiLEkw9YRzUVrR+dWsU7uEu7
TaLFEfYCAAVLHnFpPJFFOBSrUPmBknX2GvGwY6BfTo57rCp6/C6acgHh6g5+37clSVdDtZVKzpy9
NyCzBBKltxbtUgIw6rEz17YFJ0Nzy6TM5lnZsctR2+LXUcvcifyagSlDSR/ua0QKXCVT8NTfo7KK
RdZeJooYM2Oa5bGHPr+Q9BoGPC9JHrcd3TkRIjzWzIwuM38AJDgXg+cNE8zDlwEcRU156d7mos+V
Jvi9vsiQJvqKOvC1xis0MIbCg6oLtATDkETGjvQqznZCuI9kM2RluDBoSPfA9MK/bt2qG+/6hdX2
dMekt/rr6+CmHS8sOLajFPfGofKgFv5DY20wIUkdcxB4Z6b055wL963St94bp4OfZM4Sxpx8hyEk
4vHjHQVHWL1c8Coq25ubgkzR4y2VcK6UmwzG/nsXQyJiDFFTBEzaGUaclaiFfNAFvUlNd/Ulvmjc
CqHTgsENLiInI8Sj1xxKC51kGIswzqaNbg374FedHu72mfY7sE62GnxtHEGD7K4nDyvGpxwfsiGs
GaYPQaASF2mTsKJGYryXWNORsdw+rgnT5HGkWPRy5F7b8yDpPFo2EOPB6bl/9O6SSC8HTDcveN1N
govL7CXxDheO9JTcZ/r6Xr1g/XW0zlGf0IhBrJMBT8R7YH9o30NpRPNmsPhdJFKNVZ+gW37aRSrN
YWmoWZv8YwYmbN0PEgCox7mEXSFHhV+P9EVuT5jfVeVhJr3I8hqqprw23aXEboQtwL3zqFum1SsS
XKnbIK02Rn7fEsUXANDknjyvxDw3iQNt1dtrVJOy8EC3VW0uQ7KiI2iExFPLGsM/R7/lvl7SSfCB
eKOuiQJNsDZtZtm8eEuqMJ5QsqMOHFzT54/yWb8/ekUOZE0OCXhKVfTr5r+SEpUj/AUQpxR6Xktr
tWEIe0OLYhL9WzY1vU14kf6BRaL/+YNgcZk3Y5xwdWxhkFPzNwQluQf28LUzTgwkD1PG3ULajqke
M0uVl5v7YD++JR1/XwZTreqAHmqomkeFcZ1wmJ19a0vPIupUADzmVOseKvDVV86tAjkNCM1rEQUe
Om0LO0MW22H2Cnana75wJGN6EJ63N4HJoSWNvUorNV5nDCG98tVbm+UAGCFUb+T/oedUO2izq8YV
YWY6lBJL7JqP5wYeLcYiGiOmMcNtPQsTV8l+Z02iwEPr7iybfziSkAkrHbTYeSfT4zJw44jrABUG
cyPKSS1IZvHHyYuBJNI/TRUx7q8hRFq0cwaS2XiYphZVA6Ycm9ajE5vG8DR1auW6NSosZm5gT04m
5t0mg+sEVD3idZho75Kt2qDBap9FrTcmJw8nGnUKQPkd4y1473LqvSrBup4avtMS/+MpX/ZRBROj
gPJZgY7DAO1H5uW4EohQnmBWOR6bsIhsAgX05Fbj2LWvG+QVkge93gGxL/vCn6zB8lkHMnkS2Waq
fH4Mwhl+Y3hRBd47sXbHmo9VHRcHIiQ4VViG3kIv6LGIaMaNpPl3UkaczHStme3sPJqVTV6R/gHW
6blNQpdEMXXRRpOKNCG3wojqW5eGfMICVKST1Coq73SvhytpEFaXzp0reluiB1KZIKF244Z1Wu3S
QkmJeIBJVa7papWwLlh9MuDZ+0S0YU8rdLH/8c03u+e/ejnL0gK5EWgdtxk/k51xdq7VOHf6B+bS
4ZgVnFoFVjxG4pNqny3e81ghTbdJKsVjiAtqRL8W10Jfj65ggn+tpxnxza500xJ49yMY3AdWDqZ+
XSh+BSvAY8O+5I+aGiUSa+ONxxyQLlw+NAm8VIrL8Y6/T9dcnZ8TppvEbO7eMYguu9yIXcgQOtrv
/b7hLzpByXt3fSQa+9yj7EkgN3CBP83WA0gg75zIx7O78GiP6HMp+GNxfrE88lj9B1bfaiWp8zFX
qdLvWoGeBAQE6E+LUtrls/gkILz90d0JNIS5p0uRurtDVkfWoUn9a1avASx7+PgqbNhSUDR4S+1C
kMwCLLC/czvxeMy14N65oH2dR/+/fDbeRaAXuQVtb+UJ0rjfUG+3HnDNfdwa+1v+La2t4wj4rYoo
BQ0VIvleN54lDFJvgpSROu2Prqo7lDCVaV5xkeFJid6MMVL656HPZ4JR064EexpW5FZmoO5lA99V
3+YZ7Y0goXFKrIrRY/1ZYrNQQJlO6A9Hd3hNqFNYtKwEPDsvQwzQHfdBWJYwz5jOW4kKsiUwAad+
DJyrYR/34rBv3pBY70XFNvC50mEdVyQZ66wB3gyCiQMh/0hYzL5HhFVPaRVSvnTQRY8ZnLiUSob+
4tvR45ypN+FwpZtCJ1n4SCMmILF1iogQOfxJZnsytqe+zNUY5GPuaBDQoWA3E7dMVxgi5Kgq9B5Z
FQDJQHDdpWMdt4OrLtWRJfhHYM1KqkAd+Ih5yEc9pgGl+D1RoQDpWSSoh3i8DSC1mrs5eoOORbF7
FZkdRwBOKCHNaKB0NTFllbpwaWLV22vfvsWR5MWEO/wxtcrkP2Jl/91xRV0kuoblsNwtxH8D6FVh
uubNGsXWrhk0bKCkpsRaIWSbrV/Y/x3VARkEi2QrPsef7sO6/FqWhTMS87vzWsxmhS2gD8zAxjtz
94OE+spjVn9MWS1Xc5FgSDJ3XWuIGn2sEvKkhuv4PRe2jyqWVTNGNuavWD8s63XkwdaGdCXK925L
pVzne6Tril/BxKfmVsbczWILP4c9xIRjap//PKwXfjBYORTKDlY5NZ9RLOcC0pY9kkw7Mc4QuOjs
1IcTsVO/A2AAfjCLVKX3VmdiPjdfZGyh4sxebYfs3NUIYtrnIYFTfY81Yj41rUVfERx2qQTOraAf
uaJNXNbsZJdP1o2d2fEyKs213r+bAnJk1wCykP6WtHYGLOSB55PA7+JKAwC9eAeK11UU3rW2bmjk
qw3NUYklYm0IOgdW0CfFzGMhrtC+CQGiIFpFkBW9QzQ5LE7gc8irbTVO4qAhDGQaN9OxXzX2FEVZ
U5j93/paMMWb/NRVUuPWK0VoF0qKbh3KK4VFJUtfN5OdQigKzCYuTfrJSP57RcBVeGFYcpUvq1E5
UvXXIDhDL/5YZNa8LuDx/aYvX461SkSbrYUhsTInP+eZUJ8CzsNaCOxSSCku02xOBMbDBa+IrHkt
rBEZoqA4EJvrfOsOlfv2S4DSRMWnaB6EFQjDVFwe4rgPmuLN92Y+CYn1PbnOqt53nielF14efspw
1Sn9i407JYSu4lbifcwl2R87JIY3wyz0X8Zo1+ZjP3y4xz+U9iPd/YAJPx1zGqpWVYJoJ7g2jx25
9T4grP97/bTSN7c8ssuNzO7Us/J8UWgTS5O5HhrDZ9IQyXZifpYkfLhwO472ZEB4bL/u4aNcjP5g
L55wB86QoC9ImDqEd+mVtQnTBywsnOhlFubTLyf1D6VU/mhEuFIxFAHEVPqkVKI5v5Y5VOGNU2Z2
ZdPvZ/Og8ouVmaoiEHyFJw9Yz5pn+5Ic9fI3u6gDIDjNqCkdeVyElVPVBgnnDKLuNC4KzLvrfx25
t1AVEf7ehQ/fGY/fLUDvaT8E8nD6aScPc48htSGmqxnl5YTGizFykKdOJ6kakAWk5kifRMnDL6JI
qP+homPyBsFNvBw6b1ws34wDk+hO6Lx+U4ETZbp3bfPB+vDjUu21uzfjzT5PIzP5vYL4W3V8HnCa
oxTXsNRfQoJxy8GHPsE7SLD3jJ1aG2TpcfjchtQ/9VkT5zxrFsCQjzTO6ZUYGfPIx3SHz7zzSBoO
cZu9RlWDtjDjtN7gjKlZQod1IUCz39/n8OIFxXMPrizNBDPyEYsq9Lapk0G66tXNK7972mUI7o/c
3dTaJB4Fs/Zjdo2A0YPRSh+lWrCm5/9F4VQwBv99F6ADeUrbp2HLJrzPBJv0+4XT5U8mKx96s0um
/2sA5Uj8rzHIDfuGIC6QQMWpFIEiZJQAZeDRsAr9O2KvJBPfangFd1+UZMVTF6t7LXTFmeJuHDMw
KFPUvqLzxDrP18UbqLKT1nx48tTCcCNvCCVoE1kFMVA4bw+RyJh+cTNrLsBS5HPqe75cRDnJW3fl
D6P/5ozkcJdgjCqLS8G7erUFiDtRUZqEB+ofwlkIGWUEnWnC7Mdordxa/qzUczKctRF6ylj4dwDf
ZCG3xnMcNamrv+pAQjmUm/CP+Qm1ACa/wjZXr5OF3iv6GOobL8nBiWtRcDUgORTk4nOjrSUiWr1i
h2//Af5+RoJJSSsuDnJjWgz6vxFO8V7VBcFYVomRo0fp76Tk8weSdEpf4ZixFY72HO5NU2DNhgTC
xlRcTpPJoni0z48Q9O0Z0nLDzQTGZX7vuDGsIQjpguphbmtZnJCR48zBav0MrzIRqKxQ4NtotIce
on1DgPEzwq58xv8HAcwcWaIyv2t+zU6gM+OADFqEp/b3IdFvlodhEwG/kLMyhjJw9khuonY7oOgg
stBMZ8H9iU0AHtvZ5F2fhXYpGSMpfou5QfsS+TWPKVfFrWRwvVP088lVvuRGaB88aDkHf9jF0XES
6RDgxmAdQQTQWnTHmNEiAE1NifEyNQH1uqpghrKGFBeYNVM0/7vgYlxlHmOLzP1Mv06vQ6zZ6oxp
5fQnmrNnMwLmCKBdrc7syxQeItU1oePXAS8Qo5ZfY6SDP7FraUsRHMcblMvmC0SVZ+uP2Au9QezW
ahruxmSOS1/JF47SRP7fspEb73keF3DEGK5BsKElFaMEl2uMjsHnlU5b6UmnEZeMKO9sZ8JqBzlM
I5ZxT0u1df8Js6Y1rw/jX1dsfa3XVLTjFX2eIf7FZamUI8GoWcsf5aA2aQnZW87xmvWe4vrMsvkW
OsPi4obgVkh+q5lQIOuwPGGTBzcSD6Lb7vpBN28F3Cv3lqzS2mt19qr6Q2SHFwEG5d3vq8Vt2W7o
SKA8kLGLblsbCzgx7xTkelCPrOS1UOHZ5YQaxREySjZ+kc4mwZTXdL9hlKeGdXbTpYGFfnHmxKHK
YzUF0hDNdJSHaXzzDAvrodjN6WPDd7XBpR0z0OBrPGtXjZv5A055LcIjECT4+vk9hK7L118sfDOJ
p8BnR+VSZg4/r6QuMawXNZ3wqVmuwrI9f/TMRI3z6g2gNy+IpzNAXz1j776wRlIbiIT02g3NDHYc
USKnUXhS0xRzaREpEiZsMZaBgACIuDc58YbdVBsnGRrSBFC9hCb4dyZAcdS6Jqg8sDZHzX/5FVIq
edba54A5pfEnEHOzjJINn6j5bHmcEZqsyv78ndmW6VH2eHPRrOg9r3wYqBlhI3Ee1V/Vk5GySWmO
rGs39gk8z9mesVUVIP+gLYwq2l8n5vwFV0aP4AnxMaYtothwIgblceetGb8Engv8zoLj4SATNIGt
NE9l+JSNl8pkl70Q9lHkmeBmJEboeTa7pjUrcE24sVfMb2gf9tW0fIIEmMAuXSDBWmmgBE3WtPcZ
g842jkffp3Y0Qy3jPMEK/ve/xCMjcCU+QrLaKAf+lusNMnDsbvEeDhyyiPx+q5RoXCtxaP4zA8Uk
I7hU1CR7fWVh19Jq8HIO2p/xuOfT4fsUlFQjm8XZcUj0hT3gwj0vjhxXe7E50T0D1j1tVef3MvY4
O7ZHwGkd3PzT0eM1D9TpQod1Ef1Gm5D7iSgI2tjJMMTtKU30P9fz26LFbtQivL9H1xyVjS0FC9sh
SNHvmC1ljp/AF/T0jfLrIKAtqBgOwSDUbQ7dG8soHDJXpKcJuoG/x03yD8e4cUecqBN5sx/vqXwW
Fi1Hlv97zGxSxKyPA3BD7ag5Mg7c7AP5wUj8SE01TeihVEYZ2O+2IrO0h7HONlKBuQlu04Ld5YrQ
UF1Jy+Thw+C2IrZPJh2mx/62XE3B7XhVIEIqhqhymCVNQy+FYKzCIVP2xzIt90pUXI3bsctuSgCm
P864dmtpOogIcH8QLFn64exsT3ihjEQhiZPwsqnVndhC82mQFCD/Tf+hrqutL/OLHNQhtvmd7Yep
NNiCCY9bRlwnh0EUirz7C1pX6Ac6CiC8wTIGuluaET2Xjfkcw8kqiPFsg5LAz8exrjG8tdcIkCHI
c2TJPSJAZGjP1s+2bDrUiWKa+AX890k6wU7vKKceuWmjUdTpQ10ZgUktfAyxU1I/RcbIwNODx62o
39SKM1ahuPa+pHN2YtsCObP7vWORJ3MCABjkKDYno3mhY64QzDifKPJoyZsjqVgUktH7jJyphz4l
kgMwmyjRPqO+ud/ehc8zb7W0ozYlpSnbUwqzuZB/UDzjQGys+laH04U7LuG94K7G3XbH0bCfuTJc
gfYhLX/MnlbiBgw3yM3ZwHaR1OE2oCaM7BKOhGwgNT8BuakY3gDoyH1XwW7DftOVO0wNFDHc7CI8
ari8eMVMRx6RS5aCkxiwjpxo+LDzXczgLnGHJY2uWHsa/n3BPMcF40n+iGDIhvrNBUD0eAtJ9wPy
dVAdzMveJEdHCdRiLtSjZomzRKk7+6+ygmnOvvoWpoazFYXQlDzi6xIGzVqZFcSn4I9ZS4+PxOEB
j7zdDGf9Rm4f412IxacJql1863gq2mLADMKk96CICini/XYanwEpNHoFMz6KvSEZNTQT/mcoN+a4
T/gjj5I2DUf68pGL2jFNr/DT7hFEIUz/tf+K8txST3QB/iOLObRUIb5+db3p7A8Blx+nh96tLcTM
IghPRd1oYhdQjn0pF6ysrF05emIEGHpFThNf5URUPce9xq9VKJ3KQkFmRTzKNKdztirsxUPpLQzZ
dLc7g0f167kzQjleUYaq8pOYmPFqSihp7NxkfAaXKTGbCmmWh0cMPVy/ktaDIfPiwMiV3CTCMcPo
zHFAdE/pfVsKHfDuk9FY4tB1L+Xv6MqjaPJWxwWfPkLoUMIhEodfgpty0V8gOW7p+IBb9OPlKuj+
YCcVhRe7cYAWtzkUFhg3zwI3ibWnTZtnHToq4pnmXNIWZWYLXl4oHyl5BkBrCV1ANldsbD/N6aoo
L/twp9p/GbjZmoJCCfwI/AYcUmx08GYbhGCyWliapebZczL1A7KQWyP2mJqAEcRyHB3+EBwwXUDm
YD3YFb1Q6R4JRWCCqkJfPoCmazeMh6/zW8HNV6fXeseGY0nHZ8/WEVlSEz+LfNSWM8zDMf67NnSz
Am/CAfk0fkYrDAu1EmB+lxvfD6SIg7IBRxZ63w59pYYRxieHQ4VpoxF8FfNnrSrEnX/8ZApjWNB/
Qz+y8s8MtgH1JiQCD6vmYen3wkOlSAzhy2ySO55vv34KAanA3wlVG+Pj/npmkSJPD5Q6DA9boykX
ntKdNuPb7qf9zFeSg858BVbpZW8NXPAJ70DJMmTzajoI8O4W3qSPShsP+y0SS4qP7GtXy29VttGi
wyQ6++G95yJwrw8qqZUmu90zXsVgF4keKZV7srfJxPPZYnFUFK9grKpvvpb/jrbSxmAVp+JKRbHB
o7rRNkq0vQPE2+I2ER5A/GK05jCEf9rzVQ61GnfqaJ892SCesXPfgvvGhgxkYGUs4XSSuAAYIsmq
fVQ1FTIQnxkqHW38sbkwmNn7zaum/uS3rBuDAoFgowyVPrm1gCXLBirU3bP2+xwDrSWE3nFRi2GH
eg98O/iMxKClYZlpm0BRUJ02S6fnPsu3HHEEqelsiB3lJdBFd+K0RnNpXeZrX5/nlq4gYvnKwuAo
ePOTIPGCssqYmquojuVnP9aCsQOjqPHarER6d1S33Af+uEvyvf822TFviaFKAP2rpG6Uc6MUe10S
OFtD9gG67ipTWWFyPIRmwxgiLd130QblejHLeatNL8JWULj78MzWzdN26toRxbFUy0RPV22Vx33b
bX/8LTON7AaJNQdzV7iAZN5NKM0t8tETmdya4mUcyYjc1qmvtkCPv9beAi/+oDpity3Ro09Ql94v
blD+GxjkcjIqWfDohgLpzTuLnb3QR/aun1bhvOK/p4xIlojIKqAO/FRf9mYxZmNLGto8G3xvNDcP
6qvHfG2KhxANwmUgtinhr9xYi3LTXVjUe3wTZe/B39Y3rmRlwYik6pg5KaGW2F2Ed1whOu/0qSHr
69b+hm/dfgKsgo2ceGxzaOdtJKMMWambfeiz2tkY+xtD1M5gBj3di5P4gZxRQZKtM0cDMt5qdg82
CDAljcmK99bcP6EVJpKuPP3SngOqFMr2uX8LIAlTs42srUp7T3z1qAs0Ki18W7FMyGOav0kY3pSx
tWxhYnIk+ikZJHL6iNo1coId9tSN3XZExIrLbh2V7/lLuhZR+28PbBccmzLK6Hpn4OGy5k5h9r/Y
N9M7eVkGIdoUcp2wm5fBU9FtKcaFPlYT5ToEWr5PntBbwjiwan87HLe0ONquDnI7pt2bw4mV2Asl
kj7vLTzEOaf3ZSwOwHwR9xcTE+TmCk1CW7joTk6zNpmlPbbWYfd9CX9vqxZGIo/+6Kw3NTb4wfR7
YU35grXhH4HHmJOz5ugXB54aoYvWiEeN+Cfn/fYAP7fNeLgwvgCtomjQ/qGNVAgXY5Lg3a+6ZFOg
o9LdAJdt2VNfPWuQ/RlzFReX+SuFY9y/QytnC9vyOM3IvlhVORymVpedtTQUTif5wtzi/UywVYKz
AzOhzvw6ItF21cYi6wnY/cHSB60xaQy1XaIAMAsX5k7IMmlLnqzLOUDM/J9ckYXDlLCZ49Y1shfp
j0xNXdVr9IjCR+6xjJ2rFLSCSZFvPLkhLGztom1HeLZr9s6JgRQla+/4RAfGNnF+79n9WSyjEpOc
l/EsLBFxX46HSdW93mIqhcSy0cqSg/V7KDWSR4kjyLVYeHIZEqcFUVSkrwnsuG3ssDS6WMBGONXa
1N07gxarIVWssZwvXjaM6yt3ubal3DfUh8INmbVvz17hoY8sbooV/QaFY+dxV/5ePHZgmsn9lK8g
J49fGukLLAAXXLratgrLuIXD8UJIcoJ7e58UlC9cV7ys/Sex5+tg5GO9E/EOm2o0LJd5gIJaIucf
vSBngxGZEGKFsklJBQiaLKGaFdehMQhrNq6MdhMbMaST5G8RGGctK57i7TmK9D6o5knLDWHjflE0
DocRE4Vhk5UFgRgTgtA3HOxhfkwOUb/xjsFTgS7nNsjRonbQwbP4mr5SeWmLk4zHFqzV2pkqYFHl
S9UqGV3jPKJAP35rYBEma/T0bBlUpDW5hhc8lHAJ6Y0Rx0tsm0qQa02oixRa8FMrvYrLVxKk2eY1
55nLU//0LXDOsA4j0M9pOOtZmOOcU3XxIu83G/XmlBO52r4xbIsmiWN1pUPlPP23XWHgT2rB3o3x
6sdmH905JBlcot1Sjb33J+HEQw+4tajGmhZQ1HdQFOdMJzzWtzLGadpctPvvQEJzMOaPY7U/Vbqo
kRYOwH2aMgvcMEibgps6Ak56Waepy2q3Kpdv4Oj4UjSLfHRhyyO2xk7ywBcsEBYcg25BXq+HgGC5
/ad2JwqYNk2K/d/w2Cf5LRJNneK8xNDX2I+cM5/6ZqXSf8SFHFOkf0XuGPXCFsfrQRinQ6RaLkst
0AU62vHIjDc7mlUYKMGWcaU9STLU9NdKlJ8/QXcZi4frb1AjzX2QIuCS1OF77r8LtinZKo1BVFT0
tGPeGqOWhDqpOTeptbJYzHeLAav+MFKaaVo8yDx+QDnjMGQPpFfinumvARsEDqtdbgJQ15DHcPFy
s5HD+gqkO6LyxB+qS775V6zcQwii6V/fLFmEyDuLJNcTvxJV0zZSVRV78Dl9cIcZs+noigpxuCbb
Bbdh+aYD2wNigov8ygCWZUAEkTRct6Mb23MwTRV475k0f5dhAqKCnE9lnNI9zVnGKeCSU1RbQ8z5
amzar7XDLQcV5wOUkkSqLSyEGWVWLStLf9qTHAHdAEoY5mYLPpryZBms0XbbPspqbGyGIgHLoy0t
xov9pZkpe6D8r6SDiAGce6IW6+dsJyr/H/6FW327BvbJCb5vtfTTlrauhNvVzLwD36L8e82g+R4w
Usvxn1+8NKwMJEPWhL9+ltoDCKP1s68//laiMIeSm+mUWg80ImMuBQEtQk+Xl6YjZboZZc+/fmgd
1bibrKOSZrFeDxRkfJ1FOsWf3RPifOXti7aOD+L5+Gq0WVFPf5IptxqcQQOIlEOzGLaLgmaolvWy
khex6T9ia0Ppnmyp2RiZyTu60nkikK7dg5yyspYxE0xiXi8Oyoifh0GO4NNn6r22504DwPFTvxI7
egbFixitKt4SKZcym89vcWKD8YRmXfzAz2Kx0yeJZM/Rjkw/nPrqtYt2FOxe2ZJEykMZzCyuLmvK
HssG6VuAcJxVsW7B08BMMQ0d8JC2M1a3YFYDg+Y+tCjvzc9otliwd3/W+H0BgDd/Ag9gthqlwOoU
QRNOwg/HOee0Triiea+leQRT+QdlstJsDarD+ahkCod+OOyfDgR3IJx0oZeBd7YlNCQkmCn4DsjO
Zx+7XWPvNXArTOsnit3QXfCNGoTUp5xIgeUTk66hX7he/e3jVzmh+f/+RZ8SUYEyozh7SNn5bUZB
WS+CqhqtRDEEnvuc1Kr+dGkT/g1oRGtbRHB/KUK+YEF2exSlZOZAlBdHSp8lgnMXX1jAYXiXYnPW
QQi/aro7OfbXVoV9YTRYPKLYbUE+8Rgm8DCaTzKQgMqMr+/dYFsMbyuQGMve3FrJta5x/KOEeK1S
9t46hY9/fQTUAdvdtH2eYO+dbybnzyZz4QqPWuY6bLlHBlDNA6hplzrNJZVh4l50vobxNMB+s4Z7
EkqlY7BwZR7vqktEixF0p5FGfbJjWAyISEoJTBd7IRkpjkSa5YABkva62df0RU5yh+exkCW+obeU
1p8XTGoL9aNpwTveH959M93sRonCaEnVK5G/vDSbt3t7r/8tEqgXoQG2fxFya1jvZB9W10NKpQ7B
9zHGCyynFpjemidEasc79z6UBHFgUcGsFosJCgeHMvkMsjcTkgXfOikakTnWDl5id8M2P+hy1q23
XfmxJM5UrKtUVAajJ4c5FYd6x62pg6FyQnpc2HldQ2rk+CsmUBKXFP4+no9WUGi9KexDz+RWx4hp
CfkAT90wgRlwM+UAuPTUVlWs9u3rsK2/P2aI0c4Vj9VNDlcR+EHUPyy5cpNhZXPDsiB/4DUsXzO1
h5eCYM/4vdneygd/ljNTOFvwB7EKS8w5NS4/xOlyXbhe33i4F4RPZKPUHp4uFnWZHz/vg1nmK84Y
LcI3CAlHkIlpAqWoIuVFTPGZ6Xrata2OGj57x8YFj0yZfO6hCqOVz9xIIc0x3J+n2ewWZR4hrPw2
OK+s6OsO+iZ0VG9QJi5qkV2Vl8uzxizwnRUDohiepie7If1UmgsXHka3Sha9HNTyEh4f+WCB048k
ppMc/azLhymnXUGWHQDM2oEUlG39TfU0uWXwA1aJa/rCZmkKmpdeJOSj6z2hnbJKwaEUWDI/BNI+
Epv1s6F63l0gnbHm0x0E0OMR9FiXrUIn7p5ZQPyTY2phSmw8wIfmQoCaZ8z0rjWiZ6PdFEjmhvyO
hJNbA9WtawvgwpjH50UgezklGgZhCioE9Zg0AiiH8apIs8tyjwpfqrzpKwnncYu4eDCSxIxzP6ps
itRyqi4fSJKElXn3le59fjARHzGWeJMpm0WasMtYNSP3edUEGE/V2nqYKZwy1+XdJMMqJkPfNjCg
GfAewUKZtTgODRB1juZuCcENTFqfNlcGFMLqxuPum03/+hHuBKjm6xk+QzE4NVesIvhSR70XDh1w
AYVuBMaI1qBcymVqX+3WhVs/5kMxmSdlJY88/HwBhIIosgafOprlndOJuX62p+kbX+7m+cyP4JI3
qQxLnT8rTJ6vJqrY0QGoroGOPbEuBlGEHEfy6jUQQSBwCnG7IbxRDnuJgIG9tjorOvNRb4MrEDUK
SQd+vStXslk33ln8S+iLYIMMOk6Aunnh0RCu34btzegJ0sFwksbGRL20zNYkJ9iASE1xvDmXmZeR
n3gNtXQGWU5ruM8ObyvejUw1xD1Q//j6DbRHCblNFR07LXKHtSCOeN1Gu3bgZWQS2vF3D/d1bry3
sp9OFrBw806Q5siLKEKNRNZdFYoaKYJ8M4Zv/rjpOjR3c9E84jhN0G4EjD7G/Ze6g7g9Kqs1TGdH
PLl/deDkScu8TTt8wpNHOh9Hao7a+0bVyNywBcjKa+Kjgk8wsA1FjPnUugUE7XsU3k50vZlsvVDe
pLyV0Qg36wro/eP4xxcnggJDzGbqXSu1rE1Sgc61dpBJz3OIpjhvQEkDRswUdoetMDxCtFP+to7Q
cCZFXt/OJH3GIQgYxX+PsWLEITigvIZJhF7FZ1QxhNfi1deQs7uurU8ry/ZNd77HXTtSOmQ7DWAi
0ZKIEuB6LJNI7bkDB2MffYo0WzshSDDP6U7K8Gtyq2iu/rBCGvC2xOuIBxIcnQVsFkigct5kx/hi
R7aUY2CMpkJz61YXFnN32nnoMOxxzXuUhVnVDIJtMb9V7e7zaqotb/8gaIgleVmZeWAQpfZwAnGU
kMK1WrpjpjwKCxEc4kjJTdrbY4waJ+znKmwJMHrXs3Jsf+AYjPdnU2ZPIV8Jtfr1GNVnUEL1IRyY
EjNq/8lLTzOmpvpNvuvBKQsz6DM6kg57kjPeju+L5XlsV9Gq7TTOWWtmwhl8vdgoTxMf54Mw1LLC
9i7H05GwoNrfbCYmvEoZlVoejGhOolfQs4LpNhsTZvAN9Zi2c49fGxvEn50dEbfexqqmv7U4Xm6F
66GWj4FS09Ph7rT85xkNeT14Ey1AnRrpSUjuAhL6E/0+XV3n0foj7gKpadCdwt78w7gJvjh4dtwT
0Yzc+wzgRiRIC2GcB8FoyXY2JbzCBetnfp/mNFCI6mTgFNVfq/aXM+HLFhKrBa/oYhqjc3JsCB1s
RroDZgUuo9lWW0RLeZ1EdkyPE07Q5HWR1difh2iiL0vWIFqTgzSxshu/PTzQ52O/pf7xLpRQ9KtI
H/qr+p14CwlmJkCslKojc+L1MShrmi1hiiyzVySoH8kcrMQu/w/cxV9+4JKFZ+Er/z/bHqNl+yB8
5UlLGn0FGUXcT/fpWlQYpGRJSRsxM++DmQEK2gh13PZfq6BPnWsIcqUjjzVqwUOn1ra/nBPWBR9O
3SBNCXiQK05/JI6G6FYd13jWyIvWHS4T1Hxff7iHY5PeYRKrEASV+qPTV8k1+WJ33Kk4eGdEgHj3
P0YuDGURweQxdIEN4mNglb6++lhGvK/z2zJflvV5TKQ7c2IWuy6AHLP3qjtUYnpPZqQx/Xand73r
yEw35whdRHsTWLbkbrXZJkxk+UXRt3TXt4c14Ud5FcY3IeT1HODzB/pmix6jXI8EN5Dg3avEjKQV
hBYkj1b0r/6ThtldbVG4VuF94fOX9pYPnwGr6i+rudsdDlJKaSN8s6JMeWjrb2RM7UbGTBphAHhn
eQUix6B7BzhU0HBag+NW+Jmbe9iXQ42j+cKz55TsqJu81lLiRrfKhgLiBAL+II/wGbRNavNXGpaX
caH+tiEj48kw8xuIR6Id5n+VTuyjf6o1GwOiWqqIWz/TDvgTQzFBKDPLoXyUncqwlyath11AF76H
nz01eoP/ykwrDMRPPkLwP22RIaTHeVQj5G4FECD11jtVB9XsH/FlF7/MKrWaWjPjQ7GXq0r69iv9
oL8MuniPCnhP+5sg2YuLVIJcRQ1PVpitFziSdN8R5Y52dorBfcR5N4q18I253CmdSNvQRdXX9o8Z
B5vW1MJHlNvfRdG60dQkoAYD19JJi1tfp+ZgUhtBkmgW+BnQ5ImQJ6HqG2t/MMYfai7Y5cbFOp0R
sZZQQyWDHcOFwSgns9NhxS1h+q2Ck8D3/XjcH3H3B2zQKOc0XBP9Vh0xVkYwguZmLZ/HB9ck1PP8
OEQQurHbKoc9VmWbSQ7tEmWfxObVkalNLRsxG7trNN1ob/7mwGjGjgtf+zaYC+hemneMEmuEpdm2
FGSJKKC6eiqxYunJ+ldeE+K8/wXPjAltc6CaeN7OUWvBtFV3JBN/xL5aDzCyblE7bJks/tdj7Svx
SKKpFW4g4hIO7ceh52/L3+DIxaIA1ENUquf5yjecQ3kChSOdbK/ogwvVBCPVCVMtSLyrBz6oiLrb
A0PtvN/RQbNaP9Rap4THBAT0PkOxiUvtjbQ+NYbC+rhK16IFGELvdin7N0k6nvmHvHCb8kAXU+5R
6WU3lB1Xe+eytDosxyWTRUp6iWXwTQJP5ee6mJ/VnEIkeZlJG/U5v+5SUMQcl5+oeL/W5MIznshj
jGKTH1z6E0kUOU/vKYnbpo4flVi5vAQmf9Q5S9Gh72zc6lREWY5B14qY0M7HHWvLY5tt1wuEjQSa
We0TwH5mSDGRVDF8/fEnx6iOiYWXNMTCtPftBetL7SeF+kvi2FkGuFbSdbKmdQFojqFOlt6cF/Sd
soS7y5HvBcxAQpdZkFNtiTgSNeoCIGpFNa8/NL+JJy6Bcu5x0KKJ/fC5kxqEqmtt5+iHkKr42Dzs
/zdbfLgYAE8hloLqu2aI13sDySlyVZxXUL99zRqDXQC4MeglVPdNUtlNFC5Cg3Opig98HFLCrZ9x
ykn0tRAEvzdmekXcGz2GqTmO6HDtvGg7ONgIFZswr5mO4OcojX89niDv+tClrU9+RS6h8QuFPYEM
uqpNylVyFBMUVaXDUvPArS+nopMxsfC/nma7LvqmIDGt29vF8L0gDben28PbiouvT6v7yzZrLyZl
e9LErHqJvBtClIWzmQPMSVJbWTuveusV1HZuueUl58zyl1DDihZwhloALfYN8D7MzNWGIphVST2C
GgPVT8J2vNffEqLKySdZ7FeNuE3orm6zn32rm//XTq3+xJkBrQ0kz1yA8Tf3I9cR0WU2XHjdvZ4Z
j2t/5XkWdhWQaiBFUPyGzMEOsdoHQpCRuOrPnmwD8jLQGEFlzhy7KHiwcc87kbFhZLWXWgbuFVKj
9TRwbh3biTDK0LEi1ci4072db7zun+r9OrvYuWxFSHRiM4DzFAs1VI8fsDcR5ckMiwyf4O8deYmn
LMUMXoc+O1/0v6nakscCbuDb3/t8u3rf9GNqY/TB2YWoAaibx26OvpinuAWamYXZyv1qSmetZE8m
6F5FRpzSVnRSbCECED94KN/K2/muhSsnjkJgR9+hY4zcbZrDoR9GZRh4hPdO3FUbTrJPUdds2Cy4
2i94zdaRMRvbBRpYoXU4HpwGcO3tPW4Gl0SGwahOIfLGC9RCFjRABrvHcERH+bBilXALEXF33uGK
PB8DQW+P0k7jxEZey8hTcvdCTuJJW+BPiFS+Bs7XAfRqrCw53mUK0hNW8Ud14wSDrJwnRTol9S3Y
O/iRiIvUIbFVo+ZIAWbCd2hMN+GYCdIsi1CbSuJQK5Ao+gwk3mUn4jfClv9askHPeLPsxLXeH69L
3bt6xETGUXRRLjEuZpdcBz/orlMi0z152CM6An7y3LTKcvq/DUF/12lV9sgrpOHigZhUyqw7pytF
N6n4lL5Gjlsuvr7e66d3nqBPZPgk9nbAZP8Bo7cH/7MsFbkZpCKSZtnyiVFlX8ArVuZEAwy4ENGH
5KBFrKiy1Etc+owQ+F0PYgeytFDFB6hsa+NGaefqM5+DXNyx+27XGs4ldYGdyzRV95K5OnAurEp8
OMMoKJfxfsvz/DP9FTUotXearFQjch+vtJHAbRos5imb/onXvnYl2poBy1fJeVSElhushW+1WjhI
i334Ylyrh0V2Ng18nBHc0e1NBbrRYkfoKBSVu4pAO8DMlbIku5y/Cf7gn76h3L4CcVT2tHDq2UEq
n/Ks8eE2VQmLvQpJEZSsjNd56N21YpRjDocGuewxodDesOk/JKf5HdWwlb/aD8jnqguYd3KTACQf
lPnTHOtQS9hSWLR55fzFTSXzU1zEKHlFtHa8FP2mP2EYfN5zJ2g9HcQzu0uMpX8kv8ue3VnsBW0W
I5RYAUmChmMy46ECws6yWjPYUQLyvAnJQ8+vuoL5oiVT95qai8fgYL7rsURbFeJsyGx7IVH3pVfj
Soe+F/wt3Dkpp/WjqNEJe+28vV2F3NpnVEGqm537Mfyazm3SqNYNtFKbUaw1Rv4xJZWvtSx1o/pw
7XE9Rtb1XBlmCtSlXZiPzaFl5Kaaqe+WsxfkghEW/vrO6pYEX7hN2iKgvSgRa/85ST0EQCfMat0D
6p9g+y2Ts1dJpnmFkz19YBxv0KskswDe2JXKQyIvlALhVkQR2h0T+d130anqcsulVXLu+rGcnOZE
Elu9t2zLGKTN4kWrD1gkBQ5OnsLaoORFKx3ecYCEVxBYkT5PztYBtYdrS7tO0vy7ckn276eHk4j6
oH2jp6NJnsPy/0tfjCZilfiKO1canIS2zbYQsc5+wp+fbqZ3qTgHUPds9yfSX1Roi/035Zl9jYc7
m4o5/BLFKAe44eft2Ssdz4R3vJjkuTZRkL4mFja/N2yKfrAar6fcHWjzFHSxU/kUB5vj+gfRgfQW
FBL/G6o7jC5dVSfAC0YvFmNVQ50BjeIpwxiazywgJur/0cHAuDlg9PDVfYN78I3BpZX727cAfUn+
fI8vVGA/nQiI44K8mfxCfxOZqDwL8gBPQ9ajUuaBuwqABg709HZkB+ejk4OCiREGnTLG/Q1GjjsC
iDXe+VogwSGlcMN3JlLUs/KXIwwjdFjQbUDm7p7GpTvpavIzgLLRYqtes0XiQmqyUv2zRJxo/XXs
jjc05uNqcRdbcg/Uj6BxwWHjId4sbw+ZxbgmK7We99Zf7FZ9fh/ZJW/fwSHc/jXZQfMjdpebq4M7
2JXg/NWEmJwT+/FVPZy4cApW5wdjmIg9OokQMaysuqdXPqD0YTjiTgrqZFBkTMbXZwxWgCuTBLh6
/RioRtb719wNeRZo3huhzdR9G9EIpkIDRUyEDircHlEJEX7iMwugWgoKQIGzU2YsMsBezu+rSB7P
mZYfS0U5fZSCXXUphVrKK5Wt9j3OT1T5HQsM0NxygcMT8+VhcDbb9MsFS6IRQTU/lnFQlkI7nZVE
2N+8gks/nKid3n/bRIbScOGkvHLS0T304rx6R4vxH6tZ+EpBqsAP3FacsQeBSvvrG1ziFqtM7QCI
rd5rQd9mnaUP4fKCowxKse54QOePZq3UPBw7U7yAsROdtG3Vc5y2Fur8f8uJ7/csn/VMM+pBape+
0BvOFfhrNLJW7rSJkSn5R3xrBA7/m1/HnzeG7JY2zNTL1PuVZCghvArDaXCAS/Hg+jLaIrgCQhbZ
8e5QFivMzja8A6euvIr6kWa6BLKRfC77PKIHwm+EZ2X9B+Qq+0k+0zSvDBl9hvmIwG2MduEniEQt
rsYgahnf4x2J+uf6Ve+xO0dj9idDFOn7AN6R974kEH05x0wE3N7PHL5x0gUQBjoj+A5XX23URc6D
YWm2QY9UYbgsCRLLZ8IdrbPI4WL1NqsBy+ih73iNdXYJ9u5vAOMJZPXJ0R5AzOWCouBzXReF5AgU
EFx4vVWHiKCcqt+3fcv5iWLoU6zamN9nmT5yPVvbAOsM6hvsS4MnlfaqqNarcmjKcY4eeux4Gm9C
YVBa4auS7KJ40JLyilSaXlp/dm2Rkyw/KdeQfLen4n91mgfNoN8VsRAx85iPTIQoYzCU3fkZ1VYs
cgd2hwazkQwLU4KjeS+Bh4kWDNYFgDRqFdd6ASAKVwB3ps5C4NZlcS5NilkCoFNXB2N16qT/Rb2c
9r9yDBQC59H0FpgbSoILa45ag+fLUeuZpCNKg1V9O1LXf0zeX7F95pv4ADcuczE/gGAaVee8bwOy
Momoiu3P+Ux3vNo1Fur4IHwCY3kbQ83rq2FuDuxAZZAa1XIit4y9vdhQNGZHdYuAydtaJVUYhPtr
R6zEAIdfd0Pix061AXWTf7OBhH+lGk9ZfvB8K1HllUQeD9MNUplDlM4szrjt3CRHglInUl2UDGki
IA216orrJL3vS0EJQ4ZI/y1cvMS+moYEt2PWexWSRkf9adXcaImYlZZaL/mGovZ0988MHoNMmNY0
7s3ig8c7RNeaX74BxprNwHJ/sJKIxiezRkb5gilpXIQK0FEWe5DbbzZ5YWP0L0hrcyrnPv8SJbrI
/gL9Ez+FUjan5L4bqPUP1QoUlnBoQ/4gzOmtIkUI9jimjykfsJIR8QnGF27Z+o+RDXZA1S0s8z/1
4TBAJoZqAnpcMbbpjlcr0FVs/tocSF+lB59b2PgguyUcYnQAJNRp3tH1XzOszUowNQZePSXgRGkI
lZuRUmGzZDhGYja4j48JW+hmbTK6oI0pS0+Alet2paEyDGGQZKW6Ec/pewCpg0LwBg+DzOpZXnli
wP/Bgf3ysEHcG3V00i/P7hS0vUarPKs+lLvsYY0PAraUzQf3tDQGHCtxRrtZ79Md+GitT47pGgyu
P3ITu6WYhS9Yb1uCYCmu3Su2LMYkwGkfkZizd09Y+I1BcxTFw68YD2rtWsE99PA7SZVrKv/AS98T
9nlu/fDBTjXbDavP3vU2HMtab6NofJ5l+Fy4RlCbZ9I+jr3sGWOH3JsZ3S5s83IIppu+juRDWjrC
brwD08tnkhM5NgWLNkxl50i0yF0C6hgK2WVc1z1rieMXC8gNuQxJxldBRD8qwwcvCaBs6Yk0sKLd
A6weLADDF203mtBKf6PHFStZgUW8DRQ1C6oq8E1myBKmY9kLl2Kw6cPL5qyPUBbaZ0S//wSUAqNX
vfYQZc4oV57IjMe3ugDrh81ZZyKwnlQ4wzIhJ68B3dxbj3oJADLhlrwevCII5tiOATxoJ7xHl5Kx
cLSDm9fJI/o9KEJoWZwkcHXLQWkgueGnl3S9cCpB6aQlyQSh3XFdPdP4bV+7x5ZqNlmOjW0v7+WD
QkRlg9SgawZFdlYp+reGgPIA09GC2i1YwksMs6aU+4vPsDycjQoOD3VmA/UrxMCX5JprTkvkY/lV
yoXgxXUA9yCl7M+E84YidJdjcGA0Uqq/tFBYuCUn77oz771LtXtBDu07+7JKqL4PGVMSViqDu9yv
dGURG3OPvhCUxQlpVzcZDhn8RFPeEL0/yVHSj+FuELERCvafD5KXKvObTnRhDermmhi/8iEZO1tZ
gbpAiHHtYd6URTzlRi1BddLKvUPYMVx1Q9t7SK3jgRiqYddt47Xk0C6nD7GjfDWWEjsYENyzqGjm
ei86boh4f+4rNXL3ZIV3apIfhBTxdoDDlUsZwDwu6pA0WMiMjX9mnVf7ZAfLfhm6coxzIRy13vQe
Ns29lLTpTWa+jJoWY9IzBBnRaokwboNAK/bRYJ4W46ebekxuiQA7OUk28ItDE9TW3bdEwxEwce4A
HFkTbM+DtdjtYanaBt7/KvYe6sXNhYSz02xT/PUlir4DwDD6MWOy8U60kWa5v6pfWdF/cA86QQcn
/BQZloMZUAn8y5oGv+LoKwlvKOJ3Ju+wM8f5+ZUYWctmiuNHZ4W0GvayG05tuTzWS/amqJGjvA2E
sb4ctjsBjm6g1bQHjTJwEr6fIFcqntByl0PtuTR2O0znpiTcFVXLxCC8vZNf3Knd3k8aJdmVNDDP
MEl7L+dZ0Ic9ZpT9gt1jVnQ/vC5QpPpCCxVsO3IT7w3DhjUVvGAw2PeTQAFwHxhRUxwTBh169zKF
3ZPvBOybVZTnXJkjbJGDCkyJyMS6Wtc4DEJZb4VEjioji8CmkpV5u/McIVwpdzu4aJ+HOgP4KWTo
Cl3AfjKxtRXlOMxoipbiXLcLZ+kCtLbi8mChEAhEY4YhiPVATcFDBcMJI7jR4vPOL/xrFi7be6+H
Jr64tWyWaB6osta5Jax2Ztvyb6vNCcsDUJ1HtOBL1cacZFTJl/ZBEeyfz1pQK3PCgObs6q+Mqi/x
p2YRxyHns0K/MPYzgxMsGc/e/nwOQQXQjj1O5uerDew6hk0FJ7NO2UiXGVroE9WpKgRYeWhy3jnv
+J5xLk6EFb4zAJ2GA3MfTwAuPGCrCy5nIImE+SyUo6YqEraKDK7Ea4WyXVmhBvltREL7HwyjDkz3
ibEwTjsvmV8YTisP0qEHBno0II2dzLx7ur/gGoIa+tMFimje5cOkfqFxQo/Nir7heaIj+RTNBq7u
HkjsPWs3O3QiaEhRvvpOc4Lu/6mdgnru8QpSpVGrFXhZJwAnsAPuI8/FqkgPsRKsdPL5lkJp2RpC
n9orQj0xzGHRyG/fSw0o7olaVmNCEsge6YIEMpfRx0AotXQQ0dzaAlUMJETbSDBY8QobP0GIuMgH
lm0OkuaI5m8bfp/zZ0CaDSARG/X2PRmjFh8muijIBPF2URLdIH9qaX6AbBWRozLZ5ne+7Er58gkf
GTGBoGUP9C9tbjcKeYKLs90+Bw9TXMLBfcwPTsYvJ9P0xPUqYKw4D3xqmgXuxPJyMDq3DpDhXb6j
Wd4rBODK4olW7T+o/dxlUXh50kwRUq9CM79Glqhqu6EO2F0tF3HMZLKHWscV2GfJpTj91E7EpgVo
sRCQIEsLRq8mfreSwjmIV0rnEw2tVeeNcikgxnLsAz2Yk3xnJ1UQnL2BkTlU5OsN7fA8W2ZyVqLM
tM4HggErCIYvyXO91/P5y0gusBoKhRi1nvBdWkd7yXYnwRJnYtCUx78RnFfKq/20O8lw49OdzICW
cF71h/4Wfi5l9jStBnbfdJOuLoi9RkvQ18XSLuHENaAzR+Gn6QZi/KyLqW7ZEMNy2IW20eKp3gSA
yOZ37+SzRRczEyft6eRfOwtGClo5ypb9VJCjk7H0SlA7BJX/pWVPZv4IduL4ZzYpR1R4KvyUBtQW
IaiYPWJYESwL2XUYSA9MImzrB/Afp2MTrWeATHUgDvGl8qXD8XQJBUhjE3BokJnluM3B/qnqBHYO
GevDYjyTx7SME8lozFXW3y+wjSkaFBnOo4b8qflGPMj9o1dNGG93hcXhjiaMlRYyDtwszfHd7XUM
L9pqDV+Q2T4Ka30/ZjqS9hRx6wsUnQf+g4wdBiopQxmZgCcRbfiGxsp+xGwAweERcj3Y5QfXlJFN
nRAKYtwQWPjWtn+WSe9EqWMeIsIvgp2+XWGT0YvpjlB6NmzrzL654AB3P8hf/JyP2EOAEJxKctYu
3iyOAgvmnWo9UXGvraVdty8+aiTSt1UG/19iK9QO94dOEytSg7d8R2Hx3oZI3tLypqmztoaqpwsN
XBHW4aSqziD0RKlGtHSq2MjzzzBbILFhRkL/xMZVcNtjiX+tELW9FVv8cHZsZr8l/8PKrgpG80eS
KpfkzU4ek8321uF7ZtJRPvZX5SjlxmllFCUWvefHxIfRdM5P7clw79X7/KNtQREtRr06ETarHEmt
GCGx39AseWvazGpg+vGoSuaLx8iyY07fearPUtleXulbncOPbyfKW1LaCvLReQd+oFdhUPCRonXM
Qn144oZb2PEW8WOkF3PBq/tcCChsvrUVJuLFqtMVE4aLlxT570S/kLgScmCGwZ6j5ufGnDZeMvSJ
g9PRmh1ZhmuSBqB8A1iRPvK8GiVGYHunwwvxTKNO1boceKH3Dchv1VWPCKJWBk9VdwKGf9vYWvr1
VP7pnrwB0sny5EkhQNotNisFrglRLbTDBDa6VyVPdxvYJlUu59aog2nK29nWqBPhkZWzJJKQkrKF
ZVn5qhcJlpAtKMwJObs7/291OQtZTwFzIiQ76x2JtRQ9RFCuXj0nJCxq//y1klZ4wHk7dFYnYTBQ
dP0Vc31sQtbBmxLg06mZfTdnemNDr4tff0CSWboM5qbL/9RozxzS0KVCHdIweTBPA3zZrYvgwazh
fL2eBS5yLNo3ZefQmTbEMQcN1XYUupll+jalstJYR+4N6ek1R4wqeuYBYIeWlmFnZC4fOpi9bkNh
3B5eVB9vqDhaR+zQ/+Gr5WWXDpdaMzfnjDyyYrhKmLv/cBHHjvP6d/XkSMuU6+kkPnUT6sCgmQLY
+3/d+dkH48dqblJx6idVhklwm02+pMH04ba6zMTqwn12QtKcxj8F5ODU/5/AGnIfalyC5Qb4cJSn
8lRnSimrwIjhWguNsLLpvTXkppFnQ4DluBnRl+K9UfLvJnKqZxg5QIXd3Xr2CQDyFHMshrVQcESr
HEnDL5ZIqTaRa2W6bhyzGMN/dubGtxWwCYVne0hUrhxhsPAwifmkw4ndHhnUbXrMor1qbffqDvQe
jReBwb7kfRiK/RNzq2ItLDgEW+ra/FWmlXZm9Vu4iKVK//yKx3GZbR1FDnzEKW3psz8pdMvpvpC7
2L9yIoAkRllgXbaRwvjKh0ylabng3RNaeNdh36/yw5YOGPflsotBl8Naga1ErultsibNnsTCibU5
FFZE80Pek/YAIAnRMKF9UFWDYVQ6hpxiA1BYIdOt/yTyONUl7SzIHICdMKSkrYDnar6xO7eDoSAq
7xMxKxkFmrpPipk/DaqxBlCIzbRaGb1bjePg3WGxvq5abBZfvREJoKQMek2pvSbV/fQ5jgb6+Atf
VRmRhvz3nQEBYP7uYF/48ZXLySMMbJjjaYFOIJrYJ4cW0zV/5i5VfPa1GUeEqUnUH+3e3qNRMiU1
oWELaGLM6GmR3eHer61I+7jLee5Oquy/Zm3QEormsfX5S+i/Tr0wJOuqXK4mUB/VCm6lasIoPg4D
ooQg1NGvP4kzhB3dW3fzDKUwKSN18L/UvX4sYEuYSYk/WDOomLPBVewJWYrspx9T1Kp2r3FblGq4
ZZ14b5xLut+Wmt+YNuKLvQQvZrjCUx4+nx6XR0VwRa2rVUBzhVl+HV3nkZ0NE/qHtulrXzhEz9cH
D5hiu7sTju94aUQ0cX3NB+R3NTHo9FjSPL/mpchJ3v6LaJOjukBa4WTCCn1sZ/1mux3jIlrw84MN
j8ylpI8PaK0cqQVUR/kBXmIuldslL41/rI6Hx2BWHJMpUxlTao8aC6euR8z4BnFPF6rHIsbeAwRD
onrUeVyNDCrHJl+Neb7ypsrumJ6Ir0cp4uvWdbebyUu4Ezez+tkpShl+SWW2E+80gla7NSewcfR2
XDyDXAO2RQ0WNnL9D4d+vuq193i35s48Y28hyR5RW0Nvn/XxTDkzonzLkoLvCC8sLNsVVz0gL7Wl
/vvtL6RsL2JfFf7JSuCjo11O2BsGK1HewtNvky4mxeoGzAYDdtFr2KugJ2Zh9yNWrLtpLRqIu/4G
n62TgGO5/P4a4C4BWguFex1RoXhV3iqfXy82MmjLt+gvyiOP46CigPHJjvyciq1QJzFov7jyJeep
sEOrr8s0KzEDZ3qxcZfbGOTzIYP2ihXsZfkq9Z0yf9gmdki/S8oTlv+w69/ToSJFc2F/nx9ZUoA3
pMfucXJKEKnGeIXh5JBZJ7pdkNa2vRxu3kRixZjSEBfKMBD3QtIarPW3TTRFlXPZfNszlozWfiQd
/1439aaLG0RTYfC4StswQeCQP1QLztU/H6HVXyYVaYoofeLkn0sQwxMnZTTb+NSb/R+5P0K8P+mD
LS5k3/a4T+/zdQr3hmT4zgB1Dxb+LJHECFgAvKim2I/SxukEFtUBEblHYafvEN6wkzgHI0MOousm
cuUxIhRR2CozFPcf5z+An5Gyt3jH0Q95HNspua2oYD4lmJ4Tf4sN3spzW5eIXrnI66UYm+qNLvjy
mvnLKjzETF48OjHD9PTeC1nVCvda+oau+W1ZKQKLQyglDUruYoNhxZ9HYjfUi3aeNmOzW7dr13qK
PIZjv8Bg8RVZnh20q57z4NeecJGxJ5lSoYF19CLFYEpj+NCSUoBj9MgOP55J6KbkXfLn7gnTa0Gv
tkWegrxsePFeL7a1wd7PdIz4ib5GawKEnQrh2nGkT1GzY+F//lY34tgdXkqyt1gKD6c48MSeZ4I6
9gIx+dtYwqn9Itx1v1iUL/NotlJZTbP5qRADMn9N8EibN7jB6U7Qry3Di9KqG0i7BiKQQKnGPayf
gV/vswZURVpBG31QUPFfdPFFt3aqFN2TE7gbbakcqU9LXMtOcNgWok9EuMwj8EQmwSybDzDlrNNt
nM1GXDIq0G9hT+O5sxU4PWqYf8ErACAU0Br1ltbedTJTPQbDKx/sfIOGvwoA2LrYr1vh4gqydzcF
858awByT6hFvwPYOyUZ0+ssIiWbxvS4Ay+KhKHbwxLOqxe49f9NjtLJfsYVrStYreXIe8DbzZYUy
zQeXYl1CGNyeLiW63zxXdZQ7YOHZwe9BdZbNuw5KiEglHQVxrJI71+h8fdrvw37tvWdXCixmnzRz
7Z4X0qsdW+4sbDrqb8jRRvDgABnNzFCeI3F95Efj8o48buocPYWI6MAf5bf+dLoQvjDlxhyFHXd1
2uELl4JXimgjVFzJ4i6s19mQZum1FsYJCZYuXshAqzwacZswqgvHhuVnlhEf9Is0HJiCCHuQmGEg
kfFWPJy0p4IXQDxOROILIo6f+ZaQzM43lpea9Ba0y/SGCjFGh7xMD/ZLpn7ucBpN3fhADhDlVHGO
T6pMsGgN3uIg4HGecqMkhwdAMb5ToRohbcyoOllKE1F/yniKHWvB5RPqfSwNKH53F+OfUYnNnufh
ALphRkG6IkC5jQOGDBeRN6UZY62Y+A7HL2IxjTezFZSd9GcYxC4ulWM+uqDyo60mELbHZ4EHhZGY
Zs6VnUimFXlsnvrkTbo2mpRKKrqvrCT8H9x0buhWR1F2x6FGZZj3vPm17ZmWJjCaQJveSAt5tpV+
lb5nogoai8Itx/Fv+n98gbZ0ACpYurHKDcXnl+6pofx0likHWMHnv/teMtyzAamgxrbAU912y9L/
+9E0mr2TjyULkv6zrCjctCWIJUGQ+DIXvLd3/yUQERpwc3IuD2SPJvsiPY+EIbWTqEypU+2WyhpO
REF36A6+ba5G029tzBFoFmUMFn8vkmwqoSmS9MRhk8acjTiCVMlJaGm7ocCCJ/A5tX9rb+OcZePA
gJ5/LLJ8RCOIeUPCPi5Puy7TJnxeHwzd937iuPzoKZxGSTQWdvYRZU3Zz7qNu3YNizW62f153u0f
9iNwSeNqwpRmXpfNnDs5PDRdfTc1/FPBxCbVRbn6rfL5z6sCYOmiWdmpxbZ1JsF1vKqr/MTor1yS
gmeNZs/WxC8ZL+Vg1cImQgsXtDkvXHR5xplsCQRlXk4SWkS8qYxuxwOOGNRG+659uqyV+vcaoX0D
en2lrhfq7uXPeGSBIiRyp4wqpa13Keyj4E5wOhUZbVNtZGC0CdyZK8tMaM6Xcpu4zOLubaEM+24p
QFFR54BAMPBmlgAVKPn/Po0/5p2mEox/2KlZxQvbnnDUBtfD3Rhp2T5d/rQd0bQhmzZNQWib//s8
XhCr28EYEWJ9bE1zSk/iDG3tg7yXh/aPZ9cGgvzFgiPaC64MJWdZHNgbsE0oIPeXczoVGX0fLzbv
P0NcB6Dj1oJ1QM55PubThyt+0ooD+HHrCtZAamAFF0SRfJ+LCnAYRhaK1BazrkT0nNjCoLR6976d
7Pc+x2qpWAAbMelHJpxn/Tw9829VhUQbEQqD3YJ0yS5+hcR1+kNT1TbNAnvKUtWU9aVRzmQqRhtP
x7RsT1kjK6bllPmVs1OkqnQSJmmZlV4Lvdp3HpWR63wOqQiJQxt2WDiIDAHnCaOhixoc0fbJuFSt
2FWt5OjbL12H1KUM1PpSXBhhupw609Fudmu3q0UrgyL6M0zrrm5ISMz3UK2x6Az32wE08q3neL8B
d1Ra1UhmwSsaW/t2US18Bkr6ae6ao7gdz7RZYv6t/AUXFqRVfWPqKqmA1LIZlOMXQiRyN39fZeg8
olx9LqRIEP5bmZuUQ1D1zcRTSrgYv9tXIsyfUqb5TvJd2aD3w2GCTvo6C5FZNOkfZAYnGcOk1D3P
FMiXNh3IE10GaQWf6GLgYV+1DiVGM550AmbYsz7d3wHg6y1f5LhuGzUFwvhutFLKipe4npzUic7W
NkGcdMW5n/taQXk9tcMW74i6RL9wBQYqdBIR0MGrV12WzuO73Xec9LZaGYOHwqveTwqAHnzINpyg
GNOqczQ8MT1QxZnrFFc0ia+zT5q1akfJhiIyjfaS+Z9JudKenydzGpufP+SN1SnFZu6+Cm7zeQYK
JmUcMaKLHXA+xlHGxRFxRtz6A/t7k2/uDXdhuky7zskj2JZeO6YmaF+2bbtUzIgwtij7rEtaMrEN
uoTw5XeWLQ80g7Sha1qzb+2C5FshIGpbE/4zBS0r0upfisR9ETcJf++CaGQilq9yCIvaPtFJb65n
n6/cPAxrql3A6gJNdY2EWHjFTl+mR56EjG6JswpgSbRD12YidbiBfiX3WyKbSLx0bL4hYStzI+k3
d18yjEwqFZjb2469KK95hDYCNhF1N+KcAVyU4r43NapReAg0/2fAdl/21sAdugFwe8TLz/x5nIuY
TfnfXsXhOakeYpTqZwMQnWYvcJW/7hYJfqhYpcJDAM1/pwFGhbgA4j+qOBD0bbSFMYqMDpwp2/ks
/7OZboO8ecwf1QTWY4c9ajDwMkKjPSOpFEbbjXY5q5NWoIpMGe8kEQ2gBVQQJECuE5vJTzkWhVMn
KM0BgCKP80RXkbpnGniB8mSpLPc1ayS142lk3Sls62ZfjzCNvgdt4u9+OuWRGW/tsL9qTufL2SA+
cYokxEpx0yTtOklKe43FzJKp0jyRSwedYT4+ko0/29DK+sTDbWopDMylLmKJ4lfDtoMoFs8Ehezr
XQxa/pZrzsL6rDyqdcsRNT6IVluXtU0bjzbeuU78ea6J/FTZk12VkQQdq46KaiVY4iZ3BDVsxMBT
Sv8m+ilca6/qd3bIC6csoY60p9aI03ZYTut1U4bVpSbn5WXrLL9NSwP5nr/TZ0jh9T0HXQKE/TOM
yj5EoG/Z2TgmslKqStrOaiX13n0vC9nkujHTbCaCyr1DPbM550uF0Hb6NvlCLpuuBcEsokpbVmaB
+0yYc7Te209i4WcqYW5JIn77hb6vLyXRKDaAMchdEI7gHFtvLr2LJb9kvwNPY/ORMg30IcTcpnbY
cjwpG5FjpKMLfX92DfsnbA9UZe5N1ZjIUXSBEDZTeDsHR4ckgJ6yEYzxaL4holqd9Rft3kjBXHTu
aWE0aNgM16Ybu2xophcEO+Dgl2reI0MWPITZMDScAxTOLC2psg+gjU4OI9AAcq5SSCUzsilFg/hR
ilGx8iZPuuyfSFOW3PEqfAHDFWkrDyKd4QG/Gi7GeHJEYySg5dIGjwNlTFtmLuDJbRI7axem4iDH
2MoUll58eLQoLqoI8YVcFYobrfYzupHqTon5nClZjQu0NxEXFLyx652hvbGkR2eoV1nk5myDuqVH
e4LNl+CEr8ELxRZjbrwzwSwxBZQMDALJ6gT4oNvXSdcJWcslk3NMY3HyJZ8W5Bi4jYwnYSDlgzcO
B2RgtqDN27fczk/XKy/vQEiX3vukQ4/rSxACVdMQIlQohbfONQPD9FDvY+UwdoEcaRag5oKcluLb
0ty5EQNtcA6dygzLfgUUfpFYCJ+Kq7xlzuE+2f4St31WZ+jk8DqD0r/jUKgXVECDhyh2BKkEWGu8
RmT9ZQ6/W0uB0gX7ORsSTifOxXc9Pw5gZQYKaeSUVMmT8eDsZtwQQYlxOiBJ3l2Mwog4oc35rHws
52NOUEBj9ECtgVr8CARYIKsWOu4FaedOkxxqwsEjv+CCEfhmc9S6FWoGgsQ1Hr57kzc08F3Ix80S
RMpoqcMYLTPBtWNEUuQwt/29Yb8aluZ1hs8lkGP5X/LIc9TjGzKbG7C7jibe6qDHJVNMunc/Cl/w
2c9Rmay1FPOYHCzd99C1ON5C/T9Y4lJab/ZHtMgigidfl7K2Z33pfNY6o/VxJAAcT6MdCc17R2xO
Fd6QfreAV9ZfbQmHrsPHSGBvezOuHeP0koFFqKk+TPa5GKAylyGths+CxAUxNhNP8ZapHWn/bLLb
+itbbbTJnV8cd0bIwNsxxHI4qw8K5HGvRe3BYP8S+xnrTjwYzLDDRFgpXHA9E8oohKR0RJMxKI5p
gjhl+eETMX3HBukRZoHOV9ZI6WG5tWfGZOu6Dn4tYiHvuUSD8niw9m6EwzxGj6YIXyfrkh+LK7Lk
c5D65AczBvt7/eyy9weqUgbSet6mTajKEJQ06wLpaqgTa2H/gVLj0MQAlBoKbvvwiiSv1ffP0QOP
ocQcLBWMmLFnjKMcqgm+J+wQmtnO3JJ0RQLQjzBz8GQBk+7kRxLvm901al9rCeKkC2K4Clp50OEh
4Gb+qQMKFkXkw2tA2DnbJFqonaw3WHp55umfaiD23Do3JfEEG0R8WnOf+14hnA9xu0yKXplcl2p4
d8WZuz/hvXtoKOov1cASF2sPIDeTSsyE4FGQVHwbmvxTWkjGgRpfBueD15cWJi7y3U3qQyaec97B
emIfy6Wj0wS45OmpwBeMFzPMLEJ2rS1bzZrkdW4plE5aUAhMdFJThK5IrWN+Ouw2k0fcVfwHIXOs
qm2O8RLO3PZHxPyXua6SHTnJjqlRTceywMM3GnP0nDS7qjIwW9YZmuCnHcpCz8qz5IwYRQiCZ1Md
amUbHrc8Jm81TJG8BBedJoW0apFHiXLdMXnAc1nNhm9yMfgsRW7us8NAq9HXwrY8dHWzqqb0YWbe
1Io2Tuz6soG+S+GzxBJYR8xcqB1gzr2VGq3oCN2+WGG7wOOuryf2OEsagzFyEI2sbyR03WCjYQsb
Gy6FnE1/7SAaYtiSsY+3W9BHZqYEWlfe9O4sTOHl4FjQGsENe/EpZpecf2Rzd0+BuAEjrs4ipQRX
IpEvmPF4+cgepe2GVPdZtEoyFuVQeR6E81nFPd1SwFFjAj4+3JKxBY5vsHFMiEAiCs28UtmCstyk
iSNOi/+8j7BuSIhdfDKeUNPEo5PCwtDRBD6sPSXn4CqPuaHx00NriZ55f2ZOKjzxBodMskL+YG2d
WW/rXfCFIn5ewYiE0ecuj+HStVZPNUkZiCK/E5gHwFU7i9UoqU3HQBYPY3we3dHQCcMZ6quLhuzp
c0s076XCMKdfkVRZJSS5MPACvJshSm68cwk9X05nB62Zh2xG3fIYnk3VoTPFC4Y/TrIGJZZlP20q
v0gxwDjJa905ojgPhEtDe4T26B9B0ICpQxvEtlZ46lnZWHV2mTMX+kgzsw3KvZHTBbme3JjToDfn
juTtyCPyYiuQeITvaE77C8ZEQXDY39HEVaHDU4FUttvl+p41eY2YMupyJ8rGF41ucewIPH2uENZQ
/XddYHzdQXBJgjfj5KpXrXzCQhzkiKLwyypbEf5uc/zKRY7XwE1gwJziGyNJIfs+AeAMFIqklunI
4rS0i1kep27ruAe4PzAnLn/a1P02ATnbxFTjfX8FfZnR1LuX2MDUvCkkPDDU1i4p9RCw+iX+j3En
eSwY9nGH6ge37ZH3CzXxNIfnCLoS3h4vMDQkvxss8ahxBavKSlR1zM509xMRC4SJRHhNKA3g5umq
Yc8LPU8HdCVK8MWBySX3eQt4kYnjzXEXvZgTtrFBQu7uCLjAYZHYNHfBTBoTOZTkZ0cxByO+uZS1
LtNU8zyrhlFXT6jpwL3z9c0sX9j6fB0C7eY6AFa/Scy4KvQFBFxjNiBajur2ADgjhN29RO1HFimd
ljNWv1IQcbXTUoyKiSJz+xwKEXRZxXbczoXORkhDMz9hLhtteoz5GPSSvaGbZGjGJ2doMQySj8x7
sB2X7bI5dtFqJ7bmmuoex2xTzVNms8KQOjdmf95t0AP3c58GSCXBRAdWqT9CCIEEMF0XLsuZDgcT
oDFL+2jbn+ZXqYSSFeRm700s5+8FG/XavqK3qbkawxXuwUgcya/GAPZU1ipStWvuuFlFnBB/wzlk
Caz0X/qiojPrpNIKYQloYNWCN5s9SVIp6B0mEtP4Bjw/tAVkIEFqq/hqahcBnds9j6e6SUYqXNaN
t79dgJYOzoffsSkY4Qx6M8WKwmqoFxJcOgl/2LIFoylPUtSHOMk1fYzCIU7tUaLAak0UBkT8QOpL
7Lpmz9usQfV93t4M+gwKHjNN1JC8J1iwYfBX1FzLtAlA2kGXWbFUpGWB5PXrnatJzhkJNLJUWogL
mQSW3SHp2PpyKKUd6ohpcjhSzM2IiBPZ04XrRyWyDbF2mlgSRSlDtN+6PwxRwQ0chYHvXGfs1DGG
gYjnJ+1yVn/w1VGu2FfyQOmgeoiANuH3z+LC+q2Rc4xZtKElpD2E/4FS9U+P3VPV6/OHngKeAVDy
mCltoJz4sUBpUQCryx7NTy9jEwgF6dHMb0PrUfVmmM7QcYs+MoPM7eV0tQocItrfqk0QkTQRG+5N
IyaohjtJejhUIJvm/keUByq3DP7FXnhulrKb0Tj7akiY1G9VrlMWCQzslfvR50GRKcbKkcERSGJQ
woTgvQjJixtJaMlqj4oVZfGNQRiELQ5wnrfJXfogOHIM4jSRSH4AQDTM1yN/E2bxryAOLUQPIUo7
cHc0SeDUmH7eUmMLBSNWHydhyTTAll3u7U/WvTz6U2/12lJbOmMjLo3uYmsIG0bkGaYD2ebqmD42
RZfC1VF+nMyBTi9vPCMvwPmcxt0+gYFdT5IoXz268RABZCt2jjvzUOdt3O5/k1V2SU245GqTHkLY
a/M6VNiWUm/8o3x43vMSG5G6pZHITd6huS0RgjEK5CPngFeIsXnfcn35JXbWzgjKvGPEoEg20qbD
0VzS9QT5fkGeSeecE+/8xWLc+siU0d9bQODKA1s79aBK21uFAiCXy/PuOYwf6L4fNQTd097Lrjsg
sxHemw98oyBb0Z26n6NtIjE+HxPdNymccv/Hsp/i/2nDAD0dC0DYTvAbz7I63G1YcRdKrx8J0DT6
x3EOhihJzva0iQj08TXuP4yG7jEGff+zPVjFBIWZMCJ1SCg5z/lCNkSxscvjCktKL56Zg2XM3HsO
JfTa/bQFV5D+46r4M43cM5M5maLJ6YdmJ+AahmPATM9mioyUFG72TzJFDL+sSIXN6NZTJ7f3D5cM
GqKnhR7dZkH64ZTO1KtLsqcEDjZ83RV20YLHmKGK1ZRZLQKnn5i3TCjZ74r0ai6TM9q9jY1TDSEH
jglxshxYG6SmBKW2dJbC0r3TFYOZC7bHL9HEP9ikQMu4u6oQF7GLI8nJdptaSeCy2+C6zw/mh8Xy
QPppLKaWktw8SAc/Vh91Pfd27sb+vahnxkrCXPCdr0tE/aKE7rDYNlkmcvqGCW9V4YSeK1kRw1//
OAI6mT/Jps30C9j4PW0cF+131THYSdDuDz0tB1zrswfnXvyeKMCkQKrm0do4nsfoavkQpizy9WLW
5RhijEFgfLpGjLJdky2R32tArPO93ZJTB84I4IlT3Ou1tnUBeYX7q/+w9BTthHVeYFynVgiFCgd2
Djh9vSLz6zl8KZh50zxCTlIH3nbz4r1eOfHUpKA4Mi5nVxaV/DbzgW2Is1IheuOPa7f1Hlx5b9DZ
JCa1SCr3vvbh/HqTmMVeo2C+E1kjTONECVo7fLcL1gPFqJfuWn1bpZHKi03Xj/NqKFu8z5qbLIwR
HSo1fTBRnyYW/XVMl/VviSJx9sF4Armeju4KLguKdT/TfNhoWZkjq0y0g/lA2NdvbSH0Onh3nXdy
Q0633K5yjbvUYS0J+Z9LM/iS0Yv0pj9yHjP6qiKyWDP0b09ClsHKG3qo8YS5GdI0yj1HuDI/Z3m4
m+OJg+PWWPz1G+0XUuPwD8hrUKdiCQ5tk6OrPm4rjGyjNABiE7Uw/eQtKKhVoeRk36PUJjEi+Wap
q98iiboEPMItJWNXdclxD+GcRVv6V5GKakT+/DWe28AI/DMhnQ1AzhB/pZwLLNwyP9lm4dRQS6uX
Q4yoNG1BmfjjeQgzHNk0yL+GLDz/mebgLjiDwo7TzdMBw+dbQB/gLHZfW6PdTXdkYFoxzcztvZoO
KauLllFYscRzUMrk582jYHML14QMFnQC2CC+6pEXuFNGV6NcNKfHF3OiqkTjBM1+4C9wJ3McUTtN
SZxPB7FlhSv+1DKO3Qe/0Pg5VMCv3q3wV53aDYwoVfzg4J42cvLZ55z1LhKw9AxBNHfzWZO5EFt8
dGGF8C1/wP0EKmJGU/QYuSkLJtBzvoQoJrROZkPsUyleQqcFnQfiGjMRt9vF1MFOT5zaJwEdDpDc
q2Bsnd4pIkbDxIv+CWaoDDFXBF9Omkux4JCbrE3Z4aHb9QdH0JcxlUkqyAdlRb5xSN4IonvqVmac
NDTOjGNFI8nVYmtHVFfsvxEQxQr+IYndg8I2lt+d48Y6fq+6OcF63jwojvwebdUjbCYnU8c+fF20
LE6Jdigf3PgxQLXtnpADeBqzcXUu/+23fnZ8sTn0KqeLnpXqVW6PM1fLoI063SY3yRTzFIjI2Ctq
52kCYw7/L+6ZMDb/L4MG5NUhC0eN4/irjgEegesgNdTCB6YNLW3RJuDfqB9JmZRjZKIDkfdTemVP
9Iw2hQCY4+4W66LUGZ82avMBk8TWls+8usJ0QeNS+eMiRS/aQbUV01e1iKzzz7wYOEz5EXFRMOWt
d7D4xOEPy6aZw8nU1iuIillu+SvOHD60PFEZxSQ2nuvTetum70D2gq4eS1eWZTwYcNukX37M/seT
cJ8LkmDwTHlQ4guYVsw5qu0LVTA9WdCQiYTcfP/ty+mh9+xH53GfE9yNJwozw7Ewt8N8+R3Yc4aL
mCURgW1LY8vdeAaoJ0jrB4qkIa1qI6l4/MZWzlYzecxEXOZ2FoaxEQ88hCstBHPnq/MdJSoSCvI8
UjbmN9NX2sR4PjKVDDq7GCXUp7QVl9fIo1rOIeB0IGGULqq3EdNOQ134L96H8ZyaRLq/ZR3ldhL4
VPYG9Y2hy3OaweGM5xyLbkZWN+ACsgpHnHAS7W4X1KKx9XMaKTkNWTSPpULfzjLo/QGdX4n5X0qh
Ax23B+kPyTa3+FRlDbDOfgKGmZe1q+oLFLPZWRTq/fri6VULlDRTDxC881wOQAWEwR6GRa1ZemlW
Q9+3qSl5lTQaqSitv0LRg9MUbowhnbLDLLNb1Embd4Xqq+Hal3BlFoYfSgVIQv4v0CzCIff/SIfX
40AL/HpN68YZcu5Zk/5vPsOdbZsE+2gqwKJm+B/mVGa6QKrgT85tzjMaGU+HyG0dV3abLqQh5bNO
CHauW51U3YAOOdd/uA+SUmYqRjw092xPyqnKCQH3kUM1j/v87SpUaIqU2UggZr0MugFPA4lNawd6
qVQ1my3r0+YzIeeUWllbRWEL4PLDvmg8yuYHhMMUBo5bTryO+93ueraz4L3lYnnVRB0fjnz4OhCM
clnE0fSKgg7NLsqqTdDcPmYRlVjSgA1j7gtKTiOwM0h8z//bHLK3m2vUjjP90KECZ7drrM05fpBl
ywS1MNci5v7GGAmp+9WzkdYlq7acp5/HQ8+bZnl237c9hLLnJL2diHkLOjKufs8WMAhFZ0GarouW
ke8CGmrz2e3+IsZZXAfW8Wcy803AomX1U5J5P7TjDupdJo2j2Lck0E/MbiFx4rcYbFz8zP0l9xlk
i7FEg3q3SUuGPhjIwuUI7fdSKX1T+HAYCepJjtZU/0Ez8opMAPEI0xSDhIcU3cGx1SrtA6I54hmA
xnFdJrBeb6KZ3dtSHk9PpYngGZcnLlebqIrNG4j/7wWH7Y12RScjw7WMpsKFScETvWhnn2/Tz2kE
LGxKDy1Kp/hJmJ/sHVn/XQzyhXheSsYcbEGLAEd85qzkexPmCI6vFVh+SS46G2O11gHb9vH8Apvs
gA72uv0aXLRfChxStHJEQ1bJJsNPD7TYoEQ5OvE7nbmC2fHzEqV7GLWmlce+rPq2AH8S6tV+NsCy
nkIAeca5jiwaBR05J0EwRK8Plv+8CLb9l8Ot0vcC0DBw19y1zvvPtKAFDm9CBGNFUCfGA2PWJXr2
Mm9Nj5kxgWJoorKbExZpF9FFhbULwjlaf3RrAqtPdq7NKufj0rgXuM43PHqRY4gm2nR3jewzM1UT
BZqvqCHnW1obyRRnOqrapjcLqMQaYaIMdqlDhmtNN7GBo0vIpHGnDjHma0W4Nx3dP2hOONLval0z
Z5FCby1y98+Xwoz5QeU+axVDzk754ZCBnR6Zs+Wjg2lvwB17pFV2rVY+KqFtm1Cliz0AURk4If6l
RAru2cS8VXlDPWFgM9/PZIOUrPvJuXBFd8MTzDPXuceKttCYMiaD3FYQeAOhR2k4vTHTaibFeGKu
M1/QpSSNBNS+LudEZ67sqWnlv1qidoR7Aaaw37kvIveQycVSn6ZLEJhEB3YgbuG0kgN/s7xbob7L
PiADnKEQiE0iR5LF4wdTUkDHyShQBfChtfBPKHoMJaqcXShp+fB8b3/k1RjqW4AB49hcGxXsC9YH
qwAe1FkZTy11exxgzDO1bw9b8XVwsTlAQLglP5C3DyVzY1v8srTo/C27hIFb+weY1V7Wb4C/8uiv
RjJ/zSINj7mYqxGoDqjq1iUZiEu095iBvAFKfVCnnzIyP8LXyRkJS10CckOPZiMebDeBSfDhUWdN
ssPI7Z4R2U4zIFxiEhhSsGTypvTGuu5nTx7SBBfyh2vbIN3M/ETyBUd9D09iQJFaMof+jx9eVauO
mnRtrUz/YQAhIaGVJ/QgptSz4oGa+QcTnHUk3Ju9ZH99qnr6R7fPX0GvX86GFHczzRZKN0wGItHI
ONQ/xk/8za4ws6qgU4JmkMx+I7t3WT0Eg/TTjMfkt+FMBX9wPlNfruT2sOmaETlUm3DMXRn8OQIP
e/CE5FJfEqiaWP17++GhT5QZ7s+oqZ1PrADgwpfEuCVLscNJI8QvUnqm5nC6d1pGgy84mDG+HSeu
swEtaSNczicDJufFPXUhEj+yJcI3y9Oyxhoo6gRkFqfwRN3Y+zxoB2+fjz1S/fpOqwNS4dWhIgf8
4PplS/ldem40rAocAdiFTr546CrWLsWqCsoC4l53io9pvaQa2E6ocg+56bRlRuHgU+804KdyLBhX
WCWYQcXilt0QadFnGXp1wypNZOcJW37OHdwJx8mN0YjaN+IDM4IVu17OBZVOIfBLr/xAFvQKt8m4
znN/9876Mizjf5i8shAn3z8/mMLCj7Y3LCrPJs37+QC6yJMd7ryqilj9JuNM1mpMeGxgorwrjv34
fXf2VIr3cNpsTD21atDP+BiIPWrUbfHkWKOzE8rGM5gZcFDACkE2wFDLxbOj0iVgO7IWADwty4JM
3TI5FZV0la9ZkxXMD9l3wgsEF8l2vC7jFAEVI1/jCvgda9Bdl1TTAWCpUV+BRAFO6CC17Kysdq3Y
16/+J3u+7V6ClLZxHq+n3u62zNXiYtAu/I8tgmJwom9Bwv5dsLHbQUQ0ftaz/yLnuK9IvJ4KgmP5
7TvxpZBQ519bNqYJSPP9F2VZ9S/b7JyEY2FJHoywv7fIt2nHkje4ZLAkfRbWNOFgmuSP0y8gLsUr
/xwWYpdnNFZkw/Ak54F3gSRP8TbfA8Bq040gM3MokhsK6CzreDSeC4auGJycI3G3OQhVPhtZ8mlz
wbiVlmtp9eAEkVVgU31lCYMyJRrTPuHhK0BhVcit8o00fJZ7Ds6BWeLefvMSPPbxyNMt8rukUVjx
X7FmzmuCmYsynSpXOPFnTEc6/7CScVK90FsarnKdXUOqau5GdkXP8mOatiZx8f5DjFSziBD/5gZW
ASp7HF+uVxQVep3UiZ6bRwpxKOMjDy1NyfKmBtMIQbqLSwLYCSG8cnG7qW3IaQK5tugqDljr6HeV
3svnGoRAxpdY3zRzwYJxpcE5EG3aBq5extHBgrecxTApGbdXDZbFfj66bTNftrGpPVBkdUeaUWRt
R0IzsR2xa+yko9o115JH9SSMXbX76EfD8QSAwLQYaOAqkLXtyIUhsJjLDtceFZZbm1b4Ttf8AyUW
nBQrXR8hVuV0u/gKi2fMIoQgEAKebqppvGJU4A60gPMuO+2xZDZzxTFd842DIG7ODSDrc05mjKej
0X5jjq8fb/g/iPYLmXovq+sckOt86WzBzmpdfNWUkGqYVyFpZYPfWs8xuc9wtBkDqNl0Ptq76EAF
kD0/TfbJT1oQpeez5buR2/Sf+BiogGUCgEFdWrIyKuhe/xcMua0A/3qhTNPK723q+dPLspdHzrjs
RtzlSZ9nYoflEAGSknxWiXFhIHLMPYWp2JOA3ARw92BVVOTgc+tr+M30s8r1WBN2N6W6Mijg6Fgq
Zz/E1lylxJvFIN9SdTUi1lrHcOlKxs3M4z/Ae8QXEga9fvfSQsT0hDj33KkPexlV9gmiD3m/VA09
l0/sN7UAj3vGto7ecM62Dl+Hh7O8HAzvhLh18wwioZchKYZV1K1IdIw3x6fXdKQBIhY4f7I+goCr
YCMu3xdtbJangivyCGX3qK4vqZkxre+/C2j+BNDvEyfJIynGu+x31R1EBXmCc6wLj5b2fXd7CVND
/uaAyCh5QXoIxsSo9s/LpD55NdSkt7Giu2fRSV5gYY8gNM6x34sq7/wgucSU45i0FfM/l4BMy2sa
uudOOWL8gqIW3I3kwXLC54HBVnHuzku9aKM2B/EDOmxhw3UlYyfkiVl/S9zPmhhaVBgrLjK8XU6+
DaH2BlaXGuDHBFOApr4qJbpukFj6jQFBNL71ZLM0CEvZkp8T4FUxjJ7sKvj5v5q6irDs13PR2ODj
4+oq58aiERXaNWWCwickEQy58r8tS+Ng5x+Q3obyEZV6x25dqqiohHLqfU5uoN7BuhGhtqeC6X4A
5n0xj29FcW0rQ4x4ntn86dvyAhQroRhTW0s6M5xuVvjoZfT8hBDFov7tgY9BaSRZsGbHDSPB/ymC
Ma0ITiIzd9D/JPEIQlIdLFk1/qzV2/RJecc9MzqPNRgnRcRdqJwbshcEyzJLJYUkf+PgbKbsnbCu
Dl2A4Druph2kyBPwmvVn5+Czv9fWRGthYDnu/hrPwjhBzinQc8ccX+nbPByFevkHMRkZrdJQHILz
Bfn0AQ0PSFmiyIkkahBtrysvs/QVttXfS5eXClhAyRPACI+yDJyyZEGed4cWGN05WWHs0N+JL9oh
4avYRAiUL6SBP7RlX4D2qd/tFxuZDJlh7Lytm29ScNKj8wG1RG0hEDB5RZIMph+pq6DuXvoSdKci
Mn7jxZ/QQRqFDx7kSyc6mrHifxJunvM1rJ+N/Fn5HtYPxqoFsF5fH9zVzTKyvU9CtusfWiP3hB7w
vlPBMNO0Cz4Wp+VDBB0KfjjpDmrUWFCtO10IxkoW0ogx2I8O8Om7ShK+DZvPORauIw2yJk9X+XB9
AgeWaZ5bPh9X4qQUy0WKPLnB63eHR2s5ygN/QihmwzpxGkAxljzjLZArU0bkrHsUZM5kf40EIt6A
f0hvlY6y9yxVlRy19A7p3mXWvmc/dsiZDksPPKeoZasADWtv4iVPyUGJENqSIIX9NSim9dEWZLwl
rSFmpKNcYP+1BPtaIjy76MJgPaAATLbG2LKWM0b6ADMnBnlqvn48ZH077FdwDUPvyYJkyNyvv83F
3dczK5Z1oPXFpvonsHTYDm9gjSfrNkYbNsMGFIzkobG5zK6J3T0oRJxqWQ7+e2I5L7qeXCLkMNYm
oNYeWrVOjshmOFHhY8ywxFd4LdlD/4WzN/PBoXEafVz0X4sfaMpNo1Bg7NPRl/K5YwTM0YtxeNxC
5aVyBvNhLYN6GLoK818dHmlVCEGl9/2zhrg+Qc3OM9LHMcixt75TNh5+eEzFRZDbu+1Xgprl3nBu
9g4yemDQsB8X7jo6zfRHCYBBB78sle/serdDuIf48hNn5DlWTEOqKPoKnmEjSUZl7JPwhVD5Dj+f
bp56BR9qQOTkZH6Q/it0u82XpSiUwhsRuyPzD3U9atrnXrwxITawrdTzTedYre6+gMvzBt1nSf7M
1dznRCwn+4UH68E6EJEmwwnTtArnE42AjaxhB+YZ9c0+LWllLIQBZxfvmewcTM+XLqPwMV6j7a+S
xvVsMMnRsfKWW5BbpyppXiLmGZvsvaeLZJweXlijxqBcy6Lfsl0V8FQUBvvJ8HiKi+NWXMOf1LjH
obC9CHlaS23sHJVCRHLrWK9wgbVNA9XXPbcrvjrFO1cj0PYVqpqpyKiDzO3FYLcVYyp97GqSUfEn
WuoO08eJh4pGujHfUmAAs78vk3EqbN5v3HrDDIgv3vMWqBY/JPeCPXbyUBbkLQaKVkAEBatpRHVC
dgtu10Ct/Pui5metL0hjvsQ9Gl0taT7cFza7d1hCwv+OdLuMfNjbcgi2/nOdU+LpMyBx2F9VZYWJ
K+hzIPCa2BDWjqWeKB+Vmd+wGOK9zXZ9d96R+K3rg8vvfkx5ThIBsVq3YD2Zi0K0DWM209kfRRzB
Mc3E6UZhDJMIJ/GemP7WBH5k1cQwLDRrKkL9OXzNrD4FAho4Ov4V4OGRcQ58vq9ENbtQxub8sGpm
KrKCwKK/0fUAeyg+4+AGOK6VQ7YFUJ337m1/gYQMJESBGuegqFcxLanoTHgC9XuODGola0Vpy8Fo
u+cFlLDo5csSfAJVCQJA6STB5vCsNfRPH5lMtoUxVxQQk/Is6JyecsYHavLZiDayZPZX1DFgQ8TH
ai3Mx1Ilo3JRjBa0ZQ3J6RseurWKgVN/RXRvEJOksuef9KOlu8d2q84bau7XJWlBG4TTxgXq+Xxn
nBLU0LZtlX52ZSnuHhETOBfMvjt7v0vYFCVtzh0HG+huat5BHwjKYkHX4gJWo8x25cnh/caiMAfx
JeWPem6nnIC01F4qXmrJbVVji6xM9D9nfAEjIYFP8ahz0YX9IWdPklBjac6zQia3rnCBad9Kj+Kq
Cx9WVVVCW/uwQhgIKr0WTsYUmwlL4UqYiBvA46HJ2tCzryMXOaP/8l3oKA+YxG5RGxX5dg3+y/N0
gLC7Jw2ndvYcugdSxqdrPKqMaoyPuCOwBkwEOaksa5SD2qvoU4WLNyVRYLXAnKXW/KRbDiZKrBsT
ShnzSEa2m0a414pLhFttwyy2YfOTcwjkvzsxI0yeZq4A9PrAgJ9u1zx9IL37KF7zbq/oSLwn/74w
Gw958BJnzIg81EpTqmjNljEauVhmPrCD1AZn+AtO835/TrPKV4Ngx/PIHUd06JLdGZ8DBuqCg8M0
hCkpbyUmw/KZbg0ytY0yM3JuWCQQa/JGNvbpyqGNk4nb0kLxGvRP3F60zpON3DF+WEYLhIxw+HMx
m0GdVY4nQRi0MeL4PXotkyYxjVab6iXGc8CYIB5voudn9UktCcQ/hchSiAOGu+OC3UfIFBEV3x7h
OEjkTCTlzeUYmveDXP5HZLtqE2dXCMQ1Fyqa31HVpkD895L/HfpSEbdWH0xDmiPbj30+D3Z04Pqo
ZWHRMGWfPLy9Gpl1Yk2H9cITUQ0Rf913hb4tqdXIJ4wJfV0xwnDxXsqb6uTnWTs4cAkyKEZHHEXH
QCl+3TykGSU8TvkCqjtbmMCszvleSatNcYop3MaaYMU5ldGWsLZ2ivPqPTSUiLyl47flLKFttF0q
D2mVjzSmmWzJ9gsmgT8IiXwB1jC6n2ZyfitBXDHfUdWI0O9uvaqMqKTFWDloEkmH4cPETx2tEvw7
KR/3/7q63H4uZvM2ENAmM6DVfiauikh2TznuiXglerKFBBBZghrKhD8/PI+Qi+ut6bpIIyuA9A08
+26l3uB2ukOtWG/khnU5/i4WpWk+TPtWrFVK6rKthHFuqC9iAw5H9R/R9Bao5Uigym6L1flqCzjf
wNxKFt79fct5uVfSFIQ3DNsi9YSovVQQoXypBg03j/lPBMB51QyTUh6IF2A4lSOlUPjooDRj+YFg
wyOYM/T1GUMLyCezwe7X3kDkDxe/NCb7FqKlHLMK38lG9aAB1UiR1gokHAgDSgap3Tyo6DnfFoEe
DT5FYZpl/cPDUct81nndfpbelTwFV7OX6d+O3b47EoCNrPPQXy8m2kibJJSDpe7BjR1Q3IrLPG8v
TR1xLtcAYh6vb/LOfPnQlxscPhiNC1zcG9tzURHlS1zBDXBsApI+lb/oj34x3QoaP/5Ba8wgjga9
eQZmpqhBucW2u+9rdiWyQ7lFi4P16gAcF22u0vpnGymikExxRRDYQvj5/DyQO/dl9IPtXkJpxNjR
ond8EELEcOXFdeDPcoiyN8siUt1lpJ3K9H0UDgEk5D8PIhF0QzBIunjqSARYX7fmHC1ylykVriiG
20rGTpSmQr+KmKAUF8lUZEZ1GCc+mESrmKa1t9i3zZpYed21J9mKuGeWWTtEFl3PzGnNtJxmL0Br
aUwhuE6216Tdx1bk4SSByi8+g7zYbCgIE6We2RDFCtvHUndnNdDTx202UXNj1WP8vK4k6O0rp4Xg
fUoiO/DYTwxJT0gbeOLZEinh29/owQ2ot1tILfmnLGCcg9OrHjy/meSnBQZ+6M7GscNzwo4tYlYb
SAhVhTdl+ADlulQde3T7+6N9QoYS0Z+ycGQUgCIuwzznSqB+6US3/GJHQxplpbAaE7s2/pbViwEk
s+1OCLPgI50hK0JNimukAWqnUOL9FNb5PYLvXh1hRHHWaONvKvdubz9JHFYLFhJ0AHpMjdVrO+8S
VhQaYKsABUZL5sBKxF85CAwbaG7vJLoJvQQRf/WvVaitFi9Idjjj6WW/H2g7TS8V0h/VybdOicXZ
/fTMFmbXho1d3DQAO4msaN7mieER/6/5lImnxBGEEt6V3139MvAC6sP7WcgWg2qC1If24cGrkss3
2i7Se/w/ZLOqhrE9UbUeQKR0WzpiofNDmTRDN/Of3JyCtmUYzPtny3hxMIZ376ZK83KFoAAEekz7
i1aLEqSD3Wpn5Aijmq2zwGs2DA0LeMHOU8YxDlFgPI+F4KOhWcpCM+Vd/WyRITTE1NrDZ2WpgQvJ
1VHd7bGXo3F1x+FVWD9Ve8aLEpQ1EkV2/M3U+Ttz9X2k0o8n1LKtRPhgZz73csUEIyo0cO2nxJKy
Mlx12c52gGKfmbf2jiOLTCL/70d7WQWDuHeOANdv/zsrAf8/nNIWm9MCIrrjvX6zxDTifdCXt5ah
jb109003ytdwX2xnZLVD2xbumKzfYRE24Wahyf5LtCOZpCZ0+SxmCmzNJl9MlBRkCaabcwojFsRn
vEL3p904rgJcOdmYqmzs6n+jBNW67i4FuTYs8dDJDSqaR4nTe1KdbmF6mCrZhBQoHrAWvFKr8tmb
9LAEq9S/ztUkhnB1GZjuq+XhT7qWi3yDLoKROkr/EDwQwW616DCLRt6HCv0wNyFCsn77RTy9/vUw
q2MuvFerD4JHcQAd6gIdQsfL58gpePxuldWBdTEwpxNcDb4SypRA6rAs5uWpyJKLG347QDh5uUx+
thY7HyJlQUewbbosGFPFhfvYWrfNC71Y5AU4d912zvCSVrbV8wfwPPKlHDOr712NBzVD0xTpN8YA
AQ5N8tnHy12CG9LslssjpTs01gjh9x2sBIq5D4SxnmT/rNhAjSHDY7SFN47Uof2gQumZ9x4DJLU2
Dfqh4ICIh/23b8DlABMQ3f2rF3pkjhjBka1jEda5n2FV8ildIbD89eTp/KvZpYvgnJT9p8DyBSR3
06Sm04hF6yeZxLsVYY4NDB/d30pXZI3548En7B7qZCod3JrtOYhNSxEoPmhx6HVkf6oBhHnQeMjs
5rRiC9KCZzM08Ov/t0hHaph/e21N/m1pAljEl9K3ekZUCf8dgagLVJ8Zm6kX8FZeE8h+HReSg7AA
Lj+lpAfptY3I0NOQib2KXqIWxjTQ8xCCvH4RQbF4rjUkmcYcUejd6lddeaE3t1oIoMhM2o4Wblf4
YvxQotXqGgcLqk7u1AhbKhUaZwv4f5ITvsvZB+zhF9AdGKc8sMY72TXHSiCA4SanyX39OIVxHoS+
FRofItNOS35cHuJmiwAckyV3Qq4ojBrhNbDAllt4xTT1UzmEr3pOgFzrfYd7Tf2FHYXF+wMeCSOk
RMtWq8hc85YXVek57MNzEdKtVFM7Sjz0n0kFQvBGFCaBRSXIg4TYMyxKmOHenBsoeMSM4hku2EJO
4sfUcE5Dd8QuLqLbss+Kzl6rMow1qkdgVNdr8nhdksIM5Omu36di+qRRENRU/TvwRPjTgFZqS4AE
XygkGPEd1UBzuj3MUadD6L0IOxOERkXJMrwpSd6TxZ6LBr7GLmu+w8aVjWp2XPVs81Z9zulZhQEv
dEyUN8RL+6gStnBHZXqZkG1/PosTYhvYvTdengc9fzGAbejmjEIt4fm+OWuYlyILpj4izmbehzJr
0GKWHjPVWj3lP7xipZ3XqIVQGJe03KAAS55s5HX2MfoqFp8UXQkhmME4KggHMmb+bk4mJ91cIDY8
i2nfMgaNURc5hGkK7ndXXaeDJKHG+vaAZfr+gL7fMxLdRLA/NLHYHb21M1c56z+Kw8mPR58uOROI
f95WH3TLcxZ9EpmtaEgg1ZHlwcm+YgNtT1Wx71DClaFZyL+jcddbid7IEFpu8BejwKNDHEdIDDVW
D0B7dH1KEvjeKBwiBFUMAUi/u2C6XeqDEe50dZJCtZVTZJdp8wtqaE3A70JQAnXZIYJPvZ0/wlv4
w1vsxkDTzo2//X7YALOaDFS3Ay8cWcE++/zsqndK0xA04Y094NUu66+qgofVqUSZ4yFoLjqb14Q0
ZXJSp925HEj74GpYFQFyGY3or8EA9qUhPJvMhh3Y8Xz24Wpe6QmnY+4zcofu7wKG+dFtVRrizMC5
DMtSd2PalHfOdQ6L4RNdvZkfzx9UN4Z3seg6euwSYF7bKfsD/yEUrKo8afeVkK4U+3SqxBAJaqa2
ER+vXfb7a5eAQwMwtA461ZbiSWvFbSFFU45YLTIdaxwrf7odrU/ENvb2mWXuiKrUiwaEwfSDXXFr
1tIXAq4XSz/LzR74CQAgB7fzz2OvoA3+KokzZTCdvV82OZ3e6Pz3eaLMSi5xfiopJ+o1glBDNts4
Ohb42sTlsLuKXHKpPvJglAuDOZU7/druOG9whHcYfCj7Ju8AIIFV6S4kslipzf1LgbubKxmiRm86
rDovLcbQKNRK6cghQCN2493hBPve+HBPjrS8PbAsmA/NRve1anfqHcpv1D/pgAV2288YLvWKEF8I
c01P0dPW5a9rQIFiTra2Ui9cJgAS3LRaE3ylIfeGLRl40fRY3QGkR6S+CDW7KCoovC2uy5LMG2UV
q+DeNjJIPKrIZFFdSJMrTKtDTtRthhpg/+3E4TbvjT1GDow1p0DmoKEk9T0pqc/kmlusX4QacXEG
hrQmulznAkWLYDKdUeVDoEsQX1IwpJVelPxvRfKNDJXi1+1ilIn/j2XR9reeqwRUUNHFswsp/LSf
rTp9BBkViX+qhkm3uzBVtz3vPrjMv6QTagLQigp2iANHuAWpMdJ9wHjOZiYBLdWHdMaiPL/zOd2U
X4ZjiYLpA4itiZwIdkzo/t56TsgkuOlP/S5+cCJpk84wlSbwvK3xVhdV155hKRHxOwiFf/mCdBjv
utw19SikRFVAzF3Qe5QlRVC7PNAln6zAbNQX5l+cZ453KmeC502QaRDfoik/UkLKjN3RvNu29vQB
6Qzhw4w3vhUo6rBTuIu8WyGxO/+mGx3jUVzese+rGth53YK3I5bIxi04SBv5KwKDG7dX2puNTt85
6ajBSwEo5dphoHkxg+5XZczHLiFyYfcONNHc9n6VppWRj/yjTViybVQ5QGS2h9ll68mn7MQYri0o
7w/otfycdfWm8TBeOyXcgQs5Zz/dETAZRVMJXXeVp2Q4CnDXRSL1iog56PIzHMFAwlh6TEiaDppo
NB71E7vwrXm5VtpmoTebV9arq6CA6+wPplsqA3MNOk/cNOrKAl2JrzejEkB6008oWtDHCC7WFcal
3FkqjGQd9wOeL44K55BIppa37wpIw/js9sqwsPE/y0MYm65jc2LASUSFkE0FLnyA7UUMYP+f8K29
EurLfZxX7UJXpZiryVzEw4KyzJuZxuywFL1886ivRfq05fvIdeuqTsA/WgVYIz4ataoD2m+olJzO
DmaVpPlf7/N/HiY0EnV4DKhMot0URncEQa4G3cUFIUBPSnQC1s9yaWdBdUuKgOhIFkZjSBh74KjO
qKJxMIVSDc8ykX4K9coqnX/XTz/0QMN+oo0BQwFLvtB+jciwpPv2Znb2oiE3Q53RGxaeBPRUDhc0
wmyj8cTnx2Dc2Z7nxQlTOtmUI4/JRWnnVL+sl7pwe0DxO5lO/uN+9IE2qg2sdTtJoMaovCIn2+H6
Z3jUKyzZnnDrgp/N10lsbo4KDrN2Z1G2IhpCvbSwPkudN3/d8Nkq4IBb50HG3oX/8wGDpaoOw0y1
9htpYAhkqwJWF7O7lkKqcmJF9/cqBj0oUrDoVpxf9y8cnTNMPWE5K2HoLGnf6fEwhV7EXE5UNF1q
E4YjSaCTWfVV7btU0g8vPACcz1YjatGN6EBRK7azrJpJy5vtqNKvhHaHNWbKlUyswObkGyO/bQbg
FpljY8HIXx0lc5VqJevY6mLVewnswBdMHJm5Vwp/4PWRAiTun157u7qRTRrqudGuLw3Bgi1z2NFa
Y4qcpl/s2YIdYcIEmqyKqLKiO7UAip6npphbfxTuQia4FdZ7iXY5VOeNhaCNwoGtoGevbOjsuIyM
wz1VAkLLZ+kD7/L7GFmn0WRu91S0QW4HC/mHboUY2ufjawz9ycaThjPkPTM2J6GTGgFFaWsQhtB8
bxTqYTP09uAKJhD+socOpcvs9q4w2ByLvxh+gA9X1fWiUtIs5kpzttr22/eoqhr41Q6fQOlGlzsy
v8p6fbiXG4fXv/Xr/+5fpV8M9yxi5SsugT6uikHpQ4qBP57HNVoqAGPGJ8cQ7Sjlxdk+puGqIN+j
Awv5tCVUI+geJH0hd3B4IHyLtX1MuSIH0qo1LRZjsC13TPBU9vtqG176U78TOhiTp27ZFUSxTUhJ
pt3H8OANyKp+EMvkhd8Lpha4x8RQkAdUPxXGuzQbGkBWjhNBl/LsFHsWtC538tQAKifceSTI6ml5
BgXGI6QXraDwS4MKuXdf9RtVAcyDR75VieGgEVIcJLVSRubUdnLw0GGIyBkcVOjCPpc1KV0oVTHf
jAdY/iN/To9eU0ZOGDaXO0MF+Nb48d+9T364hZkm/Vc/xF1Ht0TbstdZJY8Qpgq/lLny9s3UU0/t
VmemxwLfl3G7OdWJ6BHoLCb9KqptGIajkdtnlMr+qoPCOYK2hVgT2Q2OnX2bHnrn8Ox1G8hFXeSa
F7TV08yfDk7RrqRd7jZwNiWfvdsILKAt/K9C7rBuFLuaNNGdDALQvG203sgR2mT4zx6OqQkyAHpU
hguSW6yUwppBQ5sL2K3PQ0owo9LacSQ1zY6oYYy/xR4XVgNxom+aNcZdn3aw/zccMKNZpLiO2lDu
JOMOxpntpR04YGUb5JYL55vz9BlGjuuPYZSLaTAwgCCJJkgcKc6EKF4fVd5lU6+sKgcXH6R6UH+J
yw5QXfLico7G/9aZDiKHQd5IHvNQJs71QsNO/xSxsygT0DNbSTs8XeYSJ2r+SSs9Pwvbv2yAbnPA
mqr9RVsaEZhO5Ib9U+nNIvhmbEBhcz3wNwqW6j7BXEqvE0AWOmUHly9Kga9bwPr7wwS1/athjDzl
B5xmGlRWOMSC/BTyL6JZNVacgZZ53iQwwB3MwbyrQil/K0A+bLq68twCs7Q9oiIUW2CCCCu9R3GI
ABvKpW4lDTUK16UqqTANE612LmkJwOdR/dM2eUBpPYz66DguGRFTjsDyOyOXS597BpdYkpJdIEg7
m6Z020fBTZh5Vuls5Lh+7tMSXtr3fvrQXkEiiH7ITDo1Urcvt5R7F6x9pXMadbd3TaqHAkIs/eNV
ZJBX0bRqsuUL/CgtjKtZJti2GOzlUvXEe7dF1Ww0uOm5wGQAsPQXteSQmUSPviJm32VlvZJMnWVm
W0tZKK+sEAnutA2pRhSHZNRZuv57n9e64p3MVeA5MPNBH2p5R42J/t+CLBgaQOqmyn3Sdf4Gc27b
yPKusiGsx0vEgwJMxm7GxA/ZeYm/6DwiSk1zjefTpBqB2X4bt4uFTzFuqPp2p54ELPnESM6Bvhe/
lT/uz+84x3jg7GGmrfcyluGzyClJ8m30aUQYQDmeyKNK/agmrwFN+heslvduieQb7X0e1pqyJPXO
p73HNfqw2WblVBJGbK5JPqN/DFnUPlzEDTKlpgrpjiJNsIusR6GNemW6FXREkgkv0OzIuynEuMFU
Q9R9VPW++Zb3mBTRxlzmg74m+TcDpIaQ7fM1Q837AhnWKEg/f2iZgGdTpzBB7R1JIPrurm+oqeua
ZLXYLJqAZ7tnY7Ewz8hkOexi9Nr5jjwpGMN6boOO8kZuvn9gMgZNT/IfvJ33rG/hGU6dgVv4D3ox
zOIG8pYjrbXzwEm9mEC2vg0os6NxgmpiK4D1P2MTgapxjiYYGR1chURISUKHfdigVZD2NEP6EITB
ZgUrdU/oT44oc9uEKwycEj8sJqQ9m3+/VaRW349ToG5JjdfcqMT9tilhopQk4cF+4zqDlliI4jIu
xy7tVhpMQBmRWPqyO3KohMSPYuMscN185NY0VY0fEdhZORpnIyhTeXbFuV93oe65Kmpoa3sjuN1O
o03l/mv7ELqgffBxR58P35bfCVPVBRpAjcOH92JLUFJ5itQ5Pg7+yDM8YduPFvnsmc0KO8LmkU5p
yb/KD8bqvWDFDKJsCuPhrMORJhxQr1jjpYFz796k5aXQMuKcJud0G9VCDBlCu2gAjzbro/qjcU0d
ehY8A9ZvO9rIHNrsWgLsF5o/vzlapfPibRmYo/iZO2ModYgE51/Y1peyabxJWOUYN+cJLweaznpC
eZgCvjbmSC2LKOw1fSadxDz2M7fxlWNBsqLcWOfKvm7BMTNtn8eOO95qRE0aoVKxo1iK6+DBRHY2
CoFu/PSYBlAauw6F+CfXZ3Psp6RXoJ3XVD/QQdr7kB5g/cD6T5rlcEcF178Tt3JOumJ45T7ixkQn
fhbxitnzAUC1HFqHl0rLvGYQAeYza9uciLdavC+73LbA7Sv2/IiLOkmQV38xU9Cc+omfo1QyMNhW
/3JpB2La6G2QczDdVYfEp9bUz3OCMAIDDa5p5eRqBP3wpVOhMyrVtqtJ1JgGG9Nu6lFeNFNp4Vje
noxFydoZ3K2DuX7kLrJGwjPSdj1XalKGuuNmRNlL4dXoDYjroDOwX3Pxm5Mp77AQphACGGrvjByM
WW+eyejV265DdaLwZc1vfQRn4SXnCYTO0v9CIKqpmxMMdHYGczqdZBIZJ1sPHo5Y03o2kazOakUE
KtrrKNiaKg4Luq2QXrccLJuqG8mkdUrBoURl1c8KU0H/9tFw7PUcuaYCdPCRFGl7u8WCZo2LUk1o
6K9pQsMg37aU8Bpi8oY9xnqCjkELY7hMyB3cUgX1S0vsuqok9IzwLuQaWEgfZz2GYsVP5/nSfzgv
o5Lfzz46oouFqrjWYu3KSpuWc6BVvyc/taFx+PRtxNHuWPMeAHgmXZJX4mYD9W1cEXA+GW2JUUQc
vpxWM6W+Ct4+War3YmCsuzQwaP95Lt4Zq8xPY7lNTuqN9lEYOqQxs8H8jRmg518rn/bBtx2t1bPw
ah5Cjarv5K/j0bx9t+PQGUCGapw4B5X4F4vMHui/J3ELByHhP4YAe2MfvSxdrFOrjUv0d/6YHqDn
kKJrgfUPZedxvyvMKlZYsthqFv46UMJJmD6dmYiumxUV+wWxGJHyXHY+y/rirokkU9Vpmlsy3xvn
HiEk9wZuc+9hylzd3BklluW9WFfr6fqyQRSfF9qx6XSGNsYwBAilmG8VAyE/qvZHxEE+Lhqrive1
UuCTRXhX6AFBFG1ff71Z6dItjO4lBVmVEI0RDlQnhlR3Ra5Pov63AC+lgCQpNB68TmImnWRKVoIs
HpmoW/PS1vYk2NSOKvjB9gvAS2SXzegkqIgpokVDC1f172R9/KJDMYEuYpl2erYg9WE4y2cdi2yi
2fzyLnQqdda+x114USUPGdJmB+jVvu8M0RLddaY2fm9Wu5Scx7avoePn57jRhdV/lFjZSHgOPZDv
tqfX1Iz1wVNiMtmqZY8c4ef0qyGBrsI6UIk6Q4XcuHOjd2l9RFCXNqt8RKuS/jqTwArQfKxlE6VP
5p8KHCusRFLTLJg9DbDSokCK/QicssZDeW5LRo1uap07aVeDvj833qwK4NwOfvwy28bwhvfxdp6l
Lpt0dMwuTXRy5UaXJv/NEZfN4ul5gDtvUMLifiC6KkWTIv1Oq9RkMkbEItfyRsQU0gA9quWLHWVr
72PnW9v80BSl2R+ws4SjWBWRJ9AtxSlRllS/VwSMpulvAGhuH+9UrBcjaWmdRGzTQ6kAJj/6U7yA
seitgegXlME+s3cOlSJGZBe6RqkSKcdeHf2G4Et3gAQw3rbcQW3XoOdcHSiduQxqWf+JRlxp0SZM
CzujLSXSaW79Ig+WEeWke5s3+JpnTwO/dOMlV/AW0n/nyteHbF0qTM5Hd487SEUxudWdt8rOeJ1M
aMyhhzrZKuzkb3WFdY8KvOH8p6sMVFuEkJjCQyYl7DSWWKtI6SdUv8tXMG/YP72f75vqbG//4Hrc
hl0S4dLLqOLZUPDHsZp4fmkLZEdH6K860el/dHNgHv7GBQ1Q0jsFg+MMnRHLLj2HBLCLzqkOzzN4
qHSmJD0stAn0ZSqxdvevqrDKSqNk7d47Pecmd2wSpA685Ao0EhUE45A3wfUEkc+ITaDSJXkl52i+
VgS7pks6g3ueVMm4rS5UBciV7jZQf5BV+vIiAEZbMPTUHTH3u25Xle4AKzr650hbG2xL9dBZTBpC
lrMYXXn7F+q1Nhd6lub9Ad+c0ePoTgbkwTQSh3az8ah2WokvOqAPeCH1LBkJ28IWueLaEvvlM+hn
mxkDBAHIMUSYYtQm9OwJhipL2xweUlz+dYQoUXTcI6QnwNDhqwtQe62h5e/89qP+V0ISxplpQ0l2
VJ3V4YVHFH8HPHbiBzagy6k7+AUHgZZmkJVIygYpyrbpa2ni3eQZ2MgoRojU72y1PAjRDRLVDIES
Le9B5tSBE3W62CiPjU80JBQfCZnaU78VchcrwqoqjFxesjF20e+EDqRl7DCntn/tKg8uxgVwNeiz
Oh9uJhGp68rjRD0wO54B3yE0YjZh4TU/q7Qey+eph9g5PohefUdUOuMazpQoIlBBzQIHNaGVr3EN
P2ImWjkwL9QStYEDOUvJycOPZkMatsSFm+oA/xx2zFZ+CesjT6kuYh32vWmPjmJrae7sJSDjj6I3
K98z3WFa4XMZP1gL9pQDsvm/289nf14uCzgw6pF6c+We+sJ+ck1pegYV37VwMCSvDOe31idzIGuC
+xy5noxAWm+oWxg+sOFVEA43mPW/UYCyOJ3ZYBN2WBI1ZewVl0SibhO8R7ZE/zco95DKaT8cHA/y
5iLMxcmBbwBXfAYPHhyqnZibj/hrTv16s4RP3zI59V8zmJlV0TVKxoDRclY0M6ToHicbUglT9pNy
eO+5XlIxCT+fYPwFNkmpZa3qZ5FszWqxqsldzJytfwD6LTNC8svKVt3A9dc9NsLvkkhdWv5cnoOQ
zRXTEisUFuyc7aX0On/esXq8lRtdckBEoO3s9j8g3HTbdpvwPH1A9F8QsBaBb1rbDFFV9zxco1EH
TFnXmecresT3IkzlK/sQW3fyfpVd11hW0f7bUGlJiP961mlp03p5BDzWuD/T2H36DjCHiLFFkNL1
uVpkUzz8xG/FOqMy+zjmTtQDrzQwE5kqxWLJKZSxA45QCklZ5XAQOFi4m81g5SXmDOFYvxwSCn5+
m71z+5MW1KwOCfji2FtXVd6fSOsSDw3qWJ48Tp8vUuuXD1onkLeuSDfOfGukG/IM8v4yrwF490qn
boZgrU5v6z5EkJMu1G6OZoenohiuXzy5Uf4ZheVS8faq9FCVU6qh4exM0yUVO61dyLZm87SIBX0c
PKKJzcEc/EYjoH37bz7kE0jfI6SSTJetCzVut7JfDnN8i9u/zrBD5LXc1Ssoz2MbjiuVwpa7UtQO
maMrLrHpO8EzpfnFGAP0whDH5bZzyFFUGgdRPlV0EW+F2c7OdLHkolkFNXlNskFN7ypmNJ2sizeO
I09QgPXcpC2Zqzr2j98kUFbDiR7AkGlhlOTeu+uBYNwXmyry7jpeqF/rk3LxFzr7gIn0snBw/Cur
nJu18g8RTXGF5Jv7VYRofyxGQOM5wCDixdFsxqbKAl0UigR96bQjmelaX5Z8rTsSx6ef/UfZfYLz
mhe8tzssIHSBq3paDrW/FUrPUMWGSBJsemGWONoaP8Bv2gJy9KPVL72q82nvDIABB/vryFoxgvnA
huKD86PcdCoCjYwj3mWOsMlVUnFiDSqtXJxNBweSIiSgrvmSFoovFELlJM9M0pbZH4DgBBUaUtJK
WoWCH0qOkUYSd9kZ/CpZebMv/fMQgMXnHdAwR4lQXIBL3jrXrrh2QpTd+rfvHyj4+XZiBuWDEnGR
LR3y5GgwP4sO/wm64kOSqluF0VOJHcKCCxuR6iLBX3GRdgz9ezHwZkFMxgl1jYAFBme7GNRdUG23
QB0NN+VggvTuO3z7aEciwX4vHPUmuF/FdSiq03FzklEbzBYXxsrc3aXw5lBmTTdTlwQmcJgdqSI3
pJp7+Kd6bKRXUfAFNmxF4ogUFPxi3zblpBQkjrmwO6Ljp9M+BAQdK23IAd6Hr4h0BuT2aCS81G5g
dPLhIK1smZ9ABU0cc+ivGHlJDrqSKoaTclPiYRvSKwByO4Oe5EdFTKBYBDRaHJ7KDrRtf7MNfGzv
DDy+oZJb03L02wMw+NvO6bvRU12Klvfa5q7oP+Unc7BtkyjyoucMsz39JzihSrZ1r4q8wka6Nxtm
cuidjOm4PVBUwTamsPhirhBtzGJyeiDb8l/c6YqdSzEE1hvMk/R0vs3aGQ0EvU21IwImzzEcvV74
CSKhtLOxD2PjwkzMCAtETlbTWm2LQkNna3GDkSr+sQrf35CEDnWT5/WWQDbXh9mp3Tgy53Fe0pI6
2dJzz5thCeHhZA7Ao02wwJPoVCwLuBf7JaYsp2Csxks0uWOZP/WNSKNuPLJiyTvqFDvPWkmTvdAa
g/peN8MAR1X3WrGMANJ5Ldvji+h5v2MdOTMOk0co6GLK+CPKdQ+JmRpqkZZlvymcvBwsv+/rkFSN
l4no7Te1UffTLjAxid/+C5L4CdFg3rKh7GNc+qPvj/tthwQXF/P/5VqvwssLRhTeamw35z5t1IoT
dFwXbPcdBQ6LeN3eBeF5gbtwohMFm2uc3NtjfOINjhrwCp9gcS3QYE7mnY8LtC7N6T+MjfdleP6/
Ws7Hf/p/QkZaFJJq+9h83Q+qsbVoVVYx5/5Rrtmk/q6O9znnXwiX82Bd0R3NbFGUP3ZqduG398sH
0lpRbIxddql0pR+J0a/pCIsnvs8i8N8vUArweXkEwtOeQ9cKBErUceP2xH3TVrRdDc9XMNFt5rU4
2fTlQbpO0BwY1j00RHILtLEA/ZEVpiNLRQqoe6OXUEIVHfBtGQL5xl/COoOFUtzvr+X47dz222eg
RHsApesalhHA0Y8y2PMZNzyOmarktZKIhC0nlmBP79FIROiSB0HLvrIfN2o/hWs7zCfxLk44W7Tr
arLmTfKS8RqRk+G7RLxF78M6y2cZaPQNk271UW7h7KENwrGtkrgoA9IF/veNw8xOf59DXf8C69s6
/YltYfHhzCIzh8tbviB0mxRrAu/5i3/ANu+4RsnTbH3ltDo/A4Pkx/rYSwWykLNoYK5sOcXJFHym
brFAJArM9nSqiw4YmDJkk7HCNq6uFQjkicxokehIIwAQQOkgTCzZ0BEI/fyNF/zMarrzJkmiw/J7
E3femLVrNfeOw4Bt6f1aQqVjcGgDDnsGRO2F+3BhaFEOQYKBmaM56WFFm33ObxvU3I3tnI4pZPr0
F+IXFkx8Y4UozSZHLbQ11ZRav58N8iZRwFlsASruPCfEsB6R+hT5FTG1GyE5Df5CTh+hdfiIaUlL
Nwy2VOSyfAZ1THc1AHEj7zy8ON4vuJETeF3XYWhbirvMyWZqOk8pZwIbfyzBUIjSeQYNCxOJ7wJs
Ts3+cSH12JKAWPp1qSIbt8eSf35crFVuvfMiSawgdKlYYiwH5ud9BJmu0816mzWBheFrbtpW+7wj
ypjw9mUWHcPv7xZP/UqOdsjlny/coBM637S1Of0K9SZYJRDJinLapGExUglYKJMo9UGsL3GZ+lgN
pboqqDEHQ/sUVsk33qFbAKnyLC+GqFJIRv1USIXm68By0I3Z0SLye7o2LJmoyV524ujfv9nRvWjg
9+BFEvSYj5JTSWG4C+xeEtGLU2Ss6c+eEfXsExwEsvUYvLlPNY8ADV5uCv4hSzYUqkzZUEP1F114
DpeAxBOANkJOBBFN9SJ905yuv2YUO7lgRwLev2SlP+1tsEGdixEqBCv09P+x+5ZYCkwqdbOQsRTT
AUldBWDP6SsjvOYZ6yOkNd0C5GPHq3pK1wQZV2LYIx/W4q+acxDbXKCN+QVO/HV7j3ap+jz2/83z
RwKZ4yuBWiq+D8S1bV37eF7hEOTOZH95QhvQLCyJvHTlfyfzOW217v+Aq6P8y3V9/6fKO+R/K1Kh
M39KQxYsV+MoQxRoKh6eqiwHJWGm3TszjL/BwqW4IQ5XVuzrSLbhovURZnV9ySIkzC7DRCcpvEHF
mEMiY+ikvKCA0jeRMjotWRVF4n3J/d79JDctOcozGzQHzfEoGshhG9OJvMFadBN3dzC8EJPP+1OI
cVWAYIDnlCe3JQ4bXBJzczgOfXbvGIbhtHw4zui2ajWHIQLcRQucigC6W8FdEKgntgxyBwKiEOHr
hsR2fvHHqYBcZFS7Ie1c2DQoJrVhoiYVmAi7z91CJSH0vrMS3Bbz7ZzRkO7ht3mB/wgl/xxV1jQE
IhqlWHxHtszOvjinljcWdR81lEW3eZeQqPkEW8YVpVOovayaW7LaJ0njOgoQlX3xLK1/C3Ra35+t
WeYfqX3QqHSumwhqFFzYcqpRcMPAdtbIfV+iTH1FsaGR2jYumFzTSnuwEnKcbxel9MJCHKKwxKft
DtJ0H/HeI/k+CDK6ZIOAOE67HZlf9kIi2XKnfDxI8EeJJmElKvbSe40LYQ9ECkTihfGMvhm7Uf+Q
rT9uwEJG5UQ0m1yGjFnEC8UOES9iDc9igVunVaSZU/k3TwJvwITT3Gn1fnJUw0P/xJWzGyIwY7bR
AQYPZ+I3Uk7MXELe4qYE1R6o0oNaL2ObuwUnm/+FKhqnUF+3S3RxYzPxlWrDeyoDcNUcJ7WaXJg7
d9MqLYdjE2Wlahlqlu6tb/JIvBrdmmqnD/gZGsl9ivljSPT17ZZacMXdT6QDVtpSljuJF+Anwbck
Z+0CW80vfvyU0aQuW5QLHxVdQkJyPXc+YibcLp8e7tK5hgLMCujx8qx5A3+5MyqjlMCOyHROPzWj
JmtfLgkOL/SL728L2dr4oTh/eRPK8wkyplTpovAclBVyY3+kxUG4iYh65KiwX9nayp5ohOBge5go
TBpsUKMTYwrAhwBWwAG4diRTa6yi5aIL+dzqjQEsxWJPTM2A51o3DXxBZfRMUAINdYMto30G4aSO
xsYLFW2qrQOVD4cCIclCAFz+SIQdRqJBC9uxMiQVifHo/Peg+HWlT4YLrful84T6dnhz2CtXEfI2
QumPMhgXd6z9MXyzFTfviNtqGWAVQYK4bvX8oSB2oe9hsPiIH+v7w3ceJ5yJFCyezJbv1LnsPOIr
FwLqmODZlSSD5mFQpRkUwwanAN4S3h7LLfrP9q9UjylTsekTgKi62Ac3sy0ZQOUmAsIwCAYaNnSn
bLxwOVgrXrv0Ez6lhu3kEXagXnkKUUDsvfNwQADnUyDE6QXofPT7OBESD4nW8KofXVGDRluiR3zj
VkJymtMGC8D6iKXuucWeuoqrc47Wy99jOS8NwaMdukvRU0G22slO+G3vQEHzW/0Km6oN/8yvZsI5
wdL7iISD7PnwTB7aTu3F4Bg5jhe3hM3aWUQvSftwVbqpB5FBzwMQfCKwr1zuEtuD+7ch6ZAPLDkN
Erq7dOxQOylCoLcydCewkmuthrMuUW6yU16CTAvz2Em1HlQ8vxe7OEA2UKTDbyISvBqNCno/ZSN4
vtP2fDEBe+ZsJgo/9RrrA+eSaPYr5QWSwOsT2cCCMoITXOPo4D1yHSt9DjhhSUYjResQpjMQPW1Y
GXVUBDCff3LXkVu4wLod1sluUaDunuPZA/B3KrGSremvLgj2bXOlC9qSu+BaSUawi6Y/WxyGN78y
ivfqHAcnCn8Ll48weL1WU6XV1142GxWrGM2gFT1Qixhw3pmn7uj3bHf4fgnhwoW7cCWQllgR1E71
wvDwirzfsU41QzvxXv+1bg7lstR2HvbwYTBsobyXJVGRIsIYNQSbaKIPktbKGnyhNsTrTJY+tcfI
0azqewLrlKuOyTSH34uTi8D9M1ACewWwY6VskISncrGMVFAqZtvhPBxBsgZxzokOxLh+nmS7o6l5
KGhQWhqvGzjZobnW6pV7Ysmuc7xzl+2KnPE1MjXSRb2NMeDjhEbsN3jCVU4AE2qmTqaDi6Toq+Uq
+54OkxXVfUC0qz+ZwIfv12qx5HaWY85FA+qtToAHWmwRHckR817T/kAc3h9FhPQYYrGulnwMQESl
BmaHHSv1NRqgSV+QKRaO3TaYdeh87KXqyXbub8UQONhMcQNPjCfs/sE0OR3LInVKbLWBwwbzXcpI
UskedIy0Hpq0/UiVcUbEhh9XfqD58LBA4rdRuWng+zCNbMM/MLbH81rSitvksZ46Wk8ghv2JLRg1
I1Flt2N0hqROoIDDtXh2Im4Up+EjToywBJxpQre8sORzsd4JOlICAePuIg8dDncMgfCsCU8/YVLe
L/CRRlPxuPnRBq3lBzlBAD9dqSXd8ip6Oy3w5X58ynl9eK7xAhZq6Wl2YWvcheklawnFwmakgYHf
1/ewnHnO3QstQe6nVHkDDk7Wxh1RrC44aWTRuN3k5P6s4Cn56S05VevYBgL7B+MjDfQW4AcQp/8c
CRE/63qH0RcXGshIl6BThbQ/Ia+xJikqwxQSd6VKgbqletACbRkztu+J5qAgnZ67hlbG8V2FluwK
C188HcMmUanX63xuudN1dhLQSlAd12R+eNEsYrobStZ5M3YIsK2sWOXheGH2hXdbYWoJGwopmApi
TceHMiMq6D128Jui6b1GkCWrcO0p2LMdSyrnOuEpOh4ACfpadii1tubglJfScy9ZGd24gHSXlx5V
v2bSqMPwrJfghfsLPdyNCS5wk+NpTxQ7G3cho4Z621WdtMVlseQ/wRhYiI7hCCiZTPHu7n3lDVpk
rGMgcwAQTdIwuQ/tIo005d53HxWhU3J3sIQdxbHQ+IKerloF+rhyX9o43FFmFJTpUyP6rMKB4QNz
eHtG2pdvakErFw633ivf4QdtxoG8eSVJPx4MWXjt00FZt0iDNd7NQ/nYQ59ysMe6Eh+CFSeDM3lk
2L1z8m0/Xg1somfOEmT5gHczFS9aZ6mG602vyEfbqdEpbI9P9U1JZdZwmXgBPbEVOV4QlS2dKKsY
7CuRu8b+tf0VJff2IwebpK1pyAQs6NAzAhqP6T8qVeBruSKvySK0TeC6DJOLbRKnvFPabwAPOqTq
6cFWAGbapcIc+yNs+3SepXNvvkgZxeVGP6jjXL2TNj513fN3ASnqNgsRj512nxfSzDKSm+Py+/nZ
RG7OO9nSeB/qGvyB30aKpnekSAs2gnOFeXhSqaRjjZWD5yTZWyVQu81UWZ0fgcdZY9ke6my6aRl/
+VuDZYbcr2sCPkUe49ZOhUwhXLuIku4lHLEiKKWPdDyxnc5yCCB4h5SFObuHXDped47t/4wgDCDk
YfyGGfPs8XlbSMYyE7/yOKZ6Di0XpKrx8uxWG65AZFxByitf2yYIUQMtv4k/pKu6JG7mD/dGb2VO
uEXn/PT+yowHLIyAlOaZKZ9DUgrHIpdO+6erUm0Uiqj5Rzz1b5DfX6aM/PaV4FKgfn9GG+oKj87U
Fe8SZMyqfJGw+x7k+26oBYR/HrrMkjEQ1PhAOEC3LMpwIhz55yNFeCz+sH/Ne6E7TaBwwAfP0M3O
PvJM75HnaGjt43cxYSm+4WC8EKEZCEtj4DV3K1cfrLL5ju5SHWIiKWUQpr4EpEGRRd2VrT8dKjXD
wO0x3rNTLElL247IQmAQpVj0x0z1mLcgqE4LFhm/qtM9CfJyn+gdl+D/eYY5zDZ+ZaK3YEL/bU+7
U/S9QV+srnEnfhpyD8kQU5C/ulniag8vH4BIX9Dar0/ZJ3DxS3KLXJ8AWUPyeO5rcN8IW0lo2yps
DKx16QvankUFhuVzNCQhUqdoOSMnGx+N+vVUk2ppexAGIHLUEN9u3qU2/wC9YwFkrz/hDm+JRsdC
JvbRZffTXWfL/5kJeW6WrKIVvohY76BgPrBi3B9gmODBnjLAWvMAUOQVK96lJucUDS3i6OPE9Ott
xKQsXD2klc1MS1MdwMF69q9zC6wv/AR20+EqmThiBKDR3IVlYTpjXb9IEV+9eqYmeRNiRDy9BrDU
EZv9tEuxvagxSOpkGfjrTeo02VJ+UeQ3XfV3bC3gwU+Gt+uKqhI+P9CUkdinutiVoHBAAdIw4TqT
lk48ZhvzFWZzhXPlQJm5qqtMG4i26rIHAPM6HTvvrp8WwEPZKedhWtoVAgOj0cLNYqzp2Zx7WRuL
RvMgJVjpJQeSPJgZ+fDALpBUyL3VG2db28IQrYpG/4okSA1dOXoH36hZ63RL7VIGy9S3wNRqFioD
fXZNNw4WYkP0tvoluBrLUbTH7AFpgZBtHtDABIddNvp2hUHsOZCrrrLO8Zz2ZB4s/bVmAVIUIyAB
uut5YJREw5cBbnkuM+D1xh2xQmjNgfiIlQyLL8f6jrZ47Ua2/sJJG2MJX7LaGvtr+7UKMqZtZzpX
TJykSHxiSmECKKF0SfG3Cf/9XwxstvAX06nfZCJacdEvXUFJzK1ExlDLcSPb6MGenLSKaRNwMXEd
/wIZ4h17xjjT1V4hmK6IZ0gvAgA/w0h87Ryiw8E1w8x8Y0AHoKn7vhxQQgrd7i+0gnivcTLGq2l1
XZzCJmHD6TeUocAJwPM6Rh1M6pqqV7iKTRU+xRX78K8ts2ylLB6Do0YFmxNBT6ggIlVr6GdwLm8X
9J64zJ8ormxa1kCpnZH/4er34xWe8XIxUT2TM5iyhIa8yShBhRuIwQn9pBOHkofQlNLp8Qhio5Xu
1HUt382qQbNVYM9YOFzlZ6CQBUiv/FcWP4jeNm4SkWEOjeYwE5gzfZGzTRa95ZioLnUvP5Z64SGY
dYDE+egzJ9dtPCSh8IBgPRTJQMvcnvH4eazqIh7D38uPRY6nPcGnj+82WeU6mBJDWtjmLHYvl6CL
7VTupJWPrXNI/+R4xQJ8xtddbqjj4q8Yb32PxqhmFaHeisEEQvDC9ArnHsdL/Dxi6/9q7Q9C634W
7w3/HA/Rermj+nhK3aAggsIinSBeS5k1VE861nOB+vQj0LJyFOwj1zTgj/x3repPYuOeJpedD00u
A2mWEwivT4uCVke0tP65wu0kiNp4Rz+XwiWiipxggaXlsRIAXE6wyzrGtwrDcXVGMAdXrSopiBon
J+i8vqs73sYoWnKA880iS3PZW9rW68vlS6B76rTXEA8oHrGOuoVM+r9iX6vAzGYvYIGEylil+pXj
XR/QI+G4ELRcNEntbgJxLKvnsLBkkeeD0Tg6R+jWjPGJmZRCYqN7BGJI6mEYn/naVXrzObolWIzW
c7YxXN+yw7071O2LFNx4hi2I9iALUFDsk244F7ETyd4eD8nrDk7Jxd4NS8WxSoaV4wWVMfpdHH23
hGDj+fuiGSb9NaCwROIDcpuMsB2kyasA5QhPtYYpRYvl4DPjzqrvifRhAiYljl2vdFyDUoip09V3
l7b+C/YgSaAMUceFl9Jik9pxY4dUemlUySpxTcgqSuIcZi8sDjZt4DnaE5O1JTa2Pc8KFRik141W
hykfSCtGDv8CWwqpJesOjr0uU9VbUi2a9FyJ4UnKHN1lgXi0e0fDvfHLmNB1M5AnIiiyjDDrNMM6
sThFxEjZtY96z2swIpbd1dAnH/P6hQK4xnUb5r0iQiGcecWmCqCMYQnRN7LP7woO600dAwoY6to1
Hb3OhRefIFN1Kl3TqMx/FpIEb5FMK6B3Xsur2mIcRVCJSue8jPJgK5ElIhC6LVSMZ9qL91mwwCfu
vEq3aPaIln7ANrWuNbNZeQJxob1Nk+HJ94Ufa0Sk6r/NqMtL6ETd/72IDcdcN5lWF+jKGQJt6xaX
Td2N1LtRrelZKRbBSEkMPoiEClgzcGyX/wzEVxcXM29mwluT6cjg5mlvIxBVyhiaxpwdDHVKDGmY
fLeRWQlrbFxnZHU4YA/SH/8AR3VNnosvA6WoZjCelKhVyMSjcJu2JABh/KAaI3rEm2F4OKjVnbqf
msXAGUWAqLyRODv/vm8A2st9gqZLWHskGQwhGigPoHq3oyBAGkHMoLbARZylKsWbHsbJy4Im86rD
1emIr5xbNSfFjmV1PK2JOHQT368o51AVUrrPiz2wEfZ/9CPJqWsqbEtlobM1CiumMdpghfw7I273
W2v4BJtnF6/XUMZhTb+hUMio2VhsZpjrJcQQW14xGSXm7lwjEENHrA348hypRTDtS18ksCIERPsL
Jy2wbq1KoIY0ehV2JkFjOlBib6GhWD23+SaaObSZ2gqvjzet24dbUtWJOCphjM8qKI5PAonLA+m5
PAh+MSTCoZxXeBv3iI8Hshg9xjvdgzqnCottDB3Yr5/3K3EiyOOeEJ96/GrMeZ3KGOb69m3Tct17
eJFYbC/EmlCg/GKCRvYP7N8GSck0NVb4ciXmi2mfKK4BVyCo3dZ8pDJY2CN1eP8AVp8JBkOUMnEE
JviWmaKJfLJaW94+z83vencaLOZ0+ubSGTahQ44AoDIAcNlPKkST6U3MCsxXZCLzU06+uAtv00U0
LHM6pQtZVBPJn9xncCN2S4dV3QLkbuMD/o7pupqyYwntWqDpNz6x1w1jNUq8lEZ0a7QrRJ49ZnZV
9e2kmHbEYc7eiHDDu7w/XqhcUvIz6AHRfNUVrY5F1VXxXxWNF5qR7TbxBlm7GX3gaVk4O3fNRGv1
eoMlAbRIRxmYl8JiOJFT21NHksMfxUH3humjwGYziAE6nrHZRMHwKseUBu87QrYP0pL/jx1PmS0D
1qn8n203g7oLDtYko/Gsgv2e3ez0liUnPluY2nA4+GRNRVlIlgxSU+gRU43T+LhovxK6L8yJmKAt
YvV6kYtdLhiDe1LUuf70kaEvcYARS8nTzinwcLyfd8oI3BCKbTPsQ17Lxc4h+wJCqP8QjPdxKlLP
y7d/eAqGFv7J3LCp+0hJqc4FVHltQ5cRv0QS/CfsWwqeqDr5+b84ULqTFEhdvBSc3hHnUh18Cj1K
kDr3GjDH3MVBSTPryxw5RAiiTo61Pun6O/mh8iC6ZHkRJpc7+NRb6tzAHuPq81ku5R4/xmnUj17A
xjhju0rqkr6OkxMnPMOKaVVnRw/mH5M1XPyXKXiG68mHOyD49p2yBzhvY6zvk0r+QjPY2IGcwDU6
nlTrgHhPyycT8iZk2G+WM4tJEwV1Bx38DBmNV1OW8ZZ9neHKHag1QGC0QHfRiA7fmcFnWpwTuWtF
XKsrUC80XTVrTL+I3yJnjL0mlJm2k/od7jGf2J0VRNIAs7MbPwwBDrwNakUr07TgJ8uvWrHdoVW0
6osAKZIxXoBhOMmhfm7kLT8ayI5W4FLWY7Jqfp4fKTtlHbL2pz9MWOGrsMrIugRPvVf7rabYBL00
Xln03Edkr32XHeNbxjOmWKKHn8FGg0Bwc+E+uJRIDVCb1FDLTI0yvE5TgFyJew1ofabZNOmh1btc
tOGR2YKdaktOS+d3/UHgtGo3Z9CYZZDRZ+s3WbBORm/rMeD8OAeZfnJKtpJkebTUixwLEfaFSreW
oeV3jBDp91e30jiYM0x4ez90QfZaL2VYRgs4rhVWfzyrAxS/TBrqv2MDjyUZJhiHLY3zmlffc2i8
rhtR2DDTZgMFEnJCoi55SkQTrTK5eNtYqR8evPYNNpft9t33XbEkMGt8zXi8RUWg9PNQTMnND5dQ
fwhX02NSYanuL3XcMNSxlc1Vuwsbmkky70I1p/Ofb4VxDYBMfhb1kiu9qQzz9yB8TdghteTqAoZW
23vdU7gSKZRzCeVz8NX6SPmMTPPXADzoSKZD9tESi3wwTwNvGU3DtYlSgHBWvAao8HCXrTVCN+lB
LWKpe6Ov/UAMuhd4SOXbHxmmmWMWnYW/Cni5rVxpxWKnH7JIukbeSplcRJsPs12uPRa+XEnQumZ8
Lpu3Pbl61jLIeCKqEf/qvP1QZp3JcDR7CJzWC213C4u6m/92Tmzqm4cjQdgFEn7aDWewY7Q+m7aB
gMcRGDNAuWZl4QX7NcfThZXawyBp0i2tFgmTIbDATWZ+XI8WdfjtvrAAeuAo5Femza+jP+IYDTdL
jy3z4tHbg+/zyUZWgnYMNn45txlRvWM//t21QgXhYg8ui4h2wn8RuxS9/OgDP9jh6Yk5Ma8f7yKy
DdAKnyFNy8q9KS9Nx1CNX9aGJ8K0fyD4/VPxOn49/MHVlyor8GEBYkJ9+drcNpCe3g4+Z8IWdiSG
8RNAsAIq6okL+D0FdaiRVBMu+KX3C9w2krepma0MqTSndbS4OpXsszRNw6Keqd4R8RnfNYWY8TwG
1fjr8GvRNkcQ4cN90HfISgEx4hBFiqu5Z1KChKL2u9Yra8hH8y6rA4wZ/r5vf578BzFFQTLz3gt3
x8MYYA7uLdI2uBa3Ys1R5ln1RcI1/QxW5QZHT3kdmE2+hf84gyCuHSBkK4Fa24KefYqsNvhdtup+
YLMwAZZP4HLWHvFhqZt1hX1u+80MVZeoai5ERv2KqjGRmrnl87AKQsDupEGoeCrAKMxDxTo6Rw59
6GzPLAtevDnjkOPdYoSK8o4AH49sQ1qO4l0V07NzoFCdHvoRFLwn1bWln37O8fwFLDMSyk98Tu+z
wolsUfySNtjod9ARagZyZibyLQZXWbqnMljqY7uUgaPO5lVaXUn6mXS5BWeQgNk3f8P6dluD0y4r
+yOtzJtoAtkXTEhz3V5livl5kIgxVMwlAbf5LHexw9ScvCky3SCFahtRy1CnEJia++tI/USVjuGU
hiIjgTR5p8nq+YoP1/hlgAr0MSPvfGY3QWErPp55sLgpsKmPCFVcjx/+anN6qgmYuod03m79+JGo
rc3flOve0ue91S5gBSLi6KRclJIzoXXxZmLyyNUHO4iMo9jvU7yi/tA0/H8MUpu72I+l+bD/7gUm
ygYeqY0MIXa7rpa8rfB4FqhpcIWizuFPHEfEmYAeX1+5HgeJbkWBkkjtVaqcN6P3m+r3f4763EYl
DpRpTV5nSVG63lyuzT0cMZsZsExZ8IUAXS6Z1CRkCqWPs51/IP487ahQKGe+8pvf9TZ3MBm0ugTn
zCYQnGUQ7hrBjf/aQlZRXw0Fm+Jq9zr83doEA+umwyZQKeq+VtoP2BTIi26IbmMxvKHcH4uqYKXT
fyJOUelJU0PZFc23KWx/85MXPoDKLmcnNQJywkiCY/DOu5+jwRqv8r3JX/7UiNuH1f5IGnIGHxb4
YyXCg1IGOlWMOLQDOa2YZO/3Q1sT8jfvn0GbP/D12AmW/m669M4gWeMQF9VQKQBa1laiya5XqTCw
RPYl2SV4/Z0SgyVxkZwFLLZegDL7ymQ3RCz3Gy5RJxjVJEHjY8jPJKXnCiXObjdzy2004ky+VgQY
VX/yf4n8bmflAt3HqO3eGpEWYpV8zD26je3lFY2USxt305de2QWsWe6b9AezbXbT2PWOHHVk5RbI
bRiAhzNJr9e/LPMkWuwpcL30V4Bim9SycP/LyEW/w/GQ8x0Fx19v6HXOZgx2HqAs0+loMDlQKUIg
nYh+p/k+IS9IjpilLmz6XVdDNYrisDnW/nyNqvzOf6qTIemAD3c0fKFLr39Rs+KTgkSQgE26NM+k
6WOE6PI3lVF0ntKeGvMJIyMOxpwnqwTfAZ5PltJ4WEiFFxC6yYB+Aa8VQAkS6vN2PCyHJsOJ9D/p
UC/2I8I0oxAdyhXUX6rGxkanaKxOQRUdc1lWrKn5TGPjxRPYYrPhBJUIV6xWLnjdd7rEUtey7Tne
Y7pX7OqdSJcr3f1EXT68+CfaTHaMTEmQ5wPxvVQWUrDU4ZAyQT/nFjM7t7UTmTTtvMyTDnRaxWrd
uDrZPVh5YbTc6S6GwlzLk5OenJzGSQPjciCDRvbPkc2eqtW2SizZYf4k2Rn7YFCI7X29mbPIf9cf
iBg47aXvR6Ui7FI2UYhUfqRQDp0hOaKDFepS/hwY5WlgxBGuV/wU5ZwwDhdb9/pNFUP9vslEwFiU
gDXOTRxJcvBj6xwm/6GuqXf6lXm0Gdl/tTvPk39B4PIZq2kjlo9GrMewcG3ovKt2covihNS210qy
EI0s9YDVOUiSgy1Bj1OYRXmPvFYYVn4lKf94dgXOzcVDNn/bZICyqSbxsviNflDLtWezhVWBTAWp
zuufEnYvHmFjFpfNJVsFpBp7VORUclple7d3kNDo2BcPAtGbf+BaavAK/i78YvL3+lccwKNUuIiW
3h/16/gLSoZUsfiQF4ELd7O3Vrumalg1A04IS1jpAZZR4Wo66iT9fziVIqG0LmNDUgybi1cPhnci
3rRPdSxyUwZx5gmOQfp9ZAsQRGquD2g5s1OdzmXD6bGzk2KN4D+lLqNtkQP5lYsckml3FAmjc201
3y30RcbWFEZ5mZGga1eS2YxL9FtarkJ4iQPKaXN6oXRJxF2V40aNsA0unDF2WhffIXVSvIcrkkiQ
Nd+nzTpsM4ySo+gntSM42tC7NmVbG+tA4HgfuhlOWGabmhaNtl2nE7de0zrMfV8P4jSZXRsE2NOn
W4HuMFUTGL64dB4blhkmPtwd3OMeg1URaBGeYDetbTpGSjE1njrORclLOQDyXPrFnEt25vGvcWr2
/76d6JhOHb5EawUOAXNnZEOK871JeYZ/p9ufge1YnnxlqI2BL/RB/G8l7hO7AEz8wSnCytGQWupy
x4oT34BwbB0/A09N6a3akGr3VFxQIUdqmZYf7NK1fTKJa7rIPa9HbtZ5yuGQU6jTJ4Fd9PP+Ze2Z
Lnorxq0wfaOZy5q/caAEUEy1SI3X9W6H5RM1BTSFRiRnnwzduNY8OlApvtwKK/RS2meudda9VaBW
O+cmW4k5oBZpAXvfRAUv/st2QuIHP0NgUeAZNZWIkcfESTmMqqTcTtHD+LATv8R58p/SN5FNFLwT
9/pNtSnqQHw2KSBG/zHmwWmjcAnoEN4RfZQ5/G0pplXu0T5hf7/Cifv0bdP1xN+/lR9z75ErQJCc
8z3A/avG2S3palTlTOYVVr8n0ZdaQ+WcqLOiviT6bmgtziYuuwLb6QK015pogxjCrSGgtLHhnap+
wAREDPg0cMFR2u+s796TI1b5Meb7XgoPBYoO3P3QiQkAXVIF+2kpsWQbJ5L5fk7Z7A5kx+KVcTBV
+x4R+t4yajqiIbn3Hmmsaed43lrms1XpL3ccDooFqiyIF3dHPHtKt8oJ8ut4ZPBLJmqgxAY923y2
m2fcAxzHr7AuhxZSVIwPBUy9xP99FKvOioISjRaUc9CkchaYPbq/G+Rs3ZVLhS4s9gpDke3YR3rs
EecWoI6poAH8n98a/gpV4sI+gbXp25ppKnssie//R2A2HcnMEZBYstVEa+VxXdmzURbrfU3hq1/d
VWRpoLCGjM18K/tOm9rsW03nRGNEjXz3J9IDKSsS/Z+VtNKQuXo6Nb+MyccOWQT4udb8XotSdljk
tXJhvHHzRMCMMkjn/4h9h1r0ANMzGr0kp73Zsq+JQFvI8owlrB5llY31s2Y1HU3rcYHYbiHAEjbU
UdjsdPbTYJe9g0utL2R9M/U1bI9+byWvGs67yoXUb6BhRRAUALE5tn3acCpEVqkd85lDglN3k/A2
0PgIHkp+VOyuVpme3J4NN+MNMTI36BIZlwKysRQpEAGyULJt/HjhGAMF2D3rPu7z9JVHoQMK4/is
WHxE0cpYKW3MyYn3ezz1cvho6tenKprp2KCsb6zbBC1Iq3jgi2z1AdKDdwWN8fQeAArND4t8xtO5
VqA6saIQyHDqsd0+AktCAHsexfWfeESq3ZY+zlYCikQSK9VnkDHVAl8U2xxCnVF9AnmZV1ff8NAr
WIsHeKS0E5FA9G9yL5rufLWy3qYnQIYcEyMytK0tVBCtbAyPwuU81ui5sqrjOz3vfPQ6y7SjcR6W
a5eDizrUZqvvoN3QOx50j1YORLFxMt/LmHn0PSucIscVStfVmAi192deT4u7LgXipwUTStvkzb/P
/n4qTp0gxAQ26TkAPSZvWwZv3963QtMayc7x1FxpzHHZj5gzlYzQEkbZ/05npIszSUY5dYn/NyAp
aWYoaS3tGHPPIMCLDS3TI7zDxtnwVmKePbuFeDodOAc1M/uia+9iQG2xn3ZEXb4K6MVU2TfhA1JZ
v5JI3S5wkZoejz0pKTeW1gH5fgqd7zMiCoS7ZbUvr1WQp4JbI7lEwFf5L1lyL2Y2vKkyAi5qTFr7
WUh9QKzMsehUiCb195wN+J9mgE1QEx4Ekdmdo5ZpEdm0g/hqv+rGyVePnubG55ziflTdRar93Dps
EcIwWEyf0mBkJVUbqM8SNJowYC+9Gt4RpcEwvcuNONueDogG+cp45LaAilpkigLVArDP4CKw5Yjj
auNanD++/QsjM2QxV3Szw2lLwNPjIaSEdnb8SUf/gmaD4h9qlx1WanudJzd7C+JJKwaz+GfMY8NL
/taHGvopS13qW3azKg/I3/reBkvcVkrJFUuq1y/1/etq4zRpLhNIw1eMoanKsQEMJX/zJxnTEuLG
PGmqCl/A7I2/gy9AN2DpT9uHlsf2tTW3LL0pIA2Qh8/e9OuTAA+cafHWHXxURR0SNwvNsiOd9Fav
tpo9L5CULemAEyPI8+AiwjP+H5q8GIqLj29VLVtJEIPgoWPwGS0QJeYn81BZIJe+TcHq6XVnTdjK
3Yoxz/T6ItEzxQAK6iEGGuUThqZgVePNb9pNfG5z19Xi6Hx1Uglo+rCeGrTXuNXQ7xECyzl5fhi/
ydux5hAAgsr6YifK+rqfHurUlwecMXnUhdpzWZgGYnliYPRW0rHl8uolUoXJ93aCSTIROwI3rpZn
Zdjug43wyohmpQDCMKjLkT3M+ORQyPC/zfB8wItteJ6auOoIYkj8PhYiW6uVq/MXNs9reW2+CrLg
dpmIy6rRlS/2ra2BlVY3KEN+lfHXEW5xmEI7q/klLIOtAWVXubjUOL9P5ohscTZ0IffpwMv7P6yp
qOBh5wGJw3F8CXQuGA6yjkP7a4yqIhFF83oipuJxhhOdz6/tFe/vkB9rQqx9nVwolzSpTdppGd37
UC7Lre1SY6dbm5ePdOxHuAzkY0tnocuax0HLHEezjr+fity3Oz8pebrB9rQapXvr57rc5iqYyiuU
t2g8Mziwk81Vupbxm1zd4Tc7Em3f1YGmEY8kw0+3AZX2aaHG6wR+ypEc4t9176+m5SIX4HF4obSL
capLOi9EvrhhoZ2CHDNtLtN9o+fEaxMYxbzpkNVhab2ucOPmaCS74VWnU2na3vCXJzRvjW5PQWwV
/5C3MWKKWcZvKmySIlTce7EUdKXT0yLKlx9k5kYe9bK6MoFgrTbhAqd8iIZupy6fZumE1KvmWilb
JzRlP9WDjmfQHHH8NbRoT2ZMMRb7Gs2PzURJvc30AoUt2fYHyPuQ9ePyfIbWj2WpC1Blnez1ozhv
ilwVROOtyyDIiNwoc++GRB0jZWdGxTbc0gPkCwUXp5pZT3b8Q3S3En6+i11GfIh2tgkqKJ3DQpcT
a2+anXj9Bpnr60/Ib/DMFZ6uof0HYJsr+bTVHHTWohBreJa73o0ZKyLfixtQ2ZoCT8BuSxRQYMTF
SKHccLsdoyYMwFqoReM7nWbdz6wMIVptZUTwKoRkZ/E9W5X7JwXEU+jIgijRArvDg4j8UH3fA+wP
NS3u5pv4Ga3y02T5BVg0cTnchCRPjtdtVVn97IDDK2RzgipJYrZrdHcTuYRLMbXN0fXRnpEgNbEI
0O3zUjdMIDoVfI59as/Aobi3uY4Ade+USu0sOxsxIhhPzTskj+hfIvN18RcIcsIm6n4KKS6ZsbZl
UuCXcgkd8Zvj1w8bJjEBpqYUx2MVtwSnmgrEWr+MvVjEg9meDSby7rpJYJcESP8A2/VrhU9bsFXS
QeG3UWVRRQRTb2sVD0lnlkaDLpg69IrbBwqzbiFwoUafZ/xcKXJ6YQyhU8pGHaW0xkIykS/SBnMa
duXeNPs4TjLp3ONyRC1R7OJqqjOkta9921ekM+akwHVs9yd6xdp04FYBO1ZIj1G540pICYNc26e+
37Bwywdm6jG92GRgnn8tW7aLQxtsUtxahYsMzGUW9dwqPL1GN16/fhKfkasPLkjd2QTaWNACOaFf
oMwRADkaWjnTCqhdbo3GdWkn0SYhMOkVMJtprtUQEAgr1W3UTO9X9jg21ogRShzW3+mHe+x1Wqvm
SHgirgJhzHhpgoFKegbthzuda3ZHilxKGJ27eRxArYM3d1NEuB7zbHADUmg4RGXD5LercAk6rDVA
lssUKM0gbP9nCkY5AQlXpVIDPe6RDYTSEwehoXmjmdtiN/olhjiDhxtX5vvDMIOlVF0h8dKnMlIG
HpTRmIXPbipdqw6wsiUsZW0Q8YHRXyEoS8R2rS+zUlPzsjThicaXcV5CIih9cVGvGLkqbTYedV0c
KbAUcFup9+SbQ9OIYRECxOyNHSzvIYi5WWbXF4O1us9ZvzKvA/lni5F8Evnrozrb38rM07H/HQ9O
brvmo7MuXn6vWbPlSi7sImA0b4FXaLgtaOvV9H17Qv+PcQItBvze7ZY0yu8EjGMDlc/+OLz2rfWT
5gyQiEpUXN/59eN29N/XHHrDoJt+sQB2LqWWK/UVSoTbhqbw0534jUi+GqoC8aDXqxNcW9B7Zs0r
sGzG4cKm8CGd+f2Gi5CEBxywIEeW1vgYeb3bi0jrBGNN+ReA06syzZfGufCnYKnmFQdIzkn7wM70
i2rxYQdI8whwc7NuKf9EfHDRBjUvWILDMvwEQ51vfV/0QADjZ3IM45jKFrlWoSCxePOBb1NAvUSB
pxBEGQGH+EAAUgKtnn4nr/hHRjW7Nv6HBTWBTcXfVGGleuReiWJyZlr6UCl/4RlTjgUIs9Y1Tmxv
JwTsVxHLW6GsKuLZ4ls8v10yii5qqOOrLbrURN5XfHSg1YcdYwkvTM5aTCPOsdVZpsnc5U41xTeP
SRExUT2RD1fxxSKhUaZ7Lfh7Lt3XIopfPzxVl/nbTVxfmr3RpteKyG/DRJ/Jy1jmPKlZPJch7uVB
SnNNqnraLSDNwlsRqZsw1a/0/4B5xx3XM5DM2vojf/UQgBu/YcgyYUNSej0u4izAiwuLuOVFPzbq
YNxPCiBd5NPK/YfFOsn3mBvG/NlikLGXsk2n5m34oWzwkft9JcEazKhgzu/8nOH/XfVquwP8Ebkq
7t0LFrXum7sGsGc0LQWORSevmmPC5ld/SyHnEq4elLDI/6A6myNhBb+iNm6VYg1u3u6ol7mVvODs
2psDNNbBhwyAPmf7uXH83RU36P4ZANBnSiqanfQRx0B955/91C39FRm3Vj4XY7bB5um+YSEijLLD
Z3NfC+xemim//+tBNYtNIjTpjf/0sG+ytM/OngxnXv4AmwwX/RgbqA2kC1vUaAJEWFv3C4shOVoK
0fUNlx265/ybkrCJyxmogtv52L6xODRJxn1z7IyQQAERCxbjzM+q1B4zE+71cJVEI+iRADJel4lg
WEYSSEiZG4NHWIBp8Oj99SDdPkyDu/T/GuybzRzfwD9MUxndPYnSf68a/LL/Fu2X5FmrWSFu/k4q
QSFiGcs7ONNGATPepHmxJgjpQFfjEEqKC09ugIS6lSapKmNbQHgX6+zD7JbaRjP8MdCtb9UqPDQN
qwySPOayGAB/NLAfX9adg2Q5zTKfJeE3BOG+TbjuvddgUqPpCT/aRxYBRRHwhkcUFtxgUKaw4DnF
63y9Lrly6ypNEldxamRG/FsG6IqT5alzjNWty2AHzKFAF3sDZ7fKDIIoL24D3P6bClzRC7JD8yHL
7rLuH7BXkO8VUXvLiHdG7l9iaYzFoYU0teqRlgzYptOBwzNhqYoUhJsLU1C2UP1zNZ7+ls07jfeL
qzcl9v2cPzNFsMsrBUbXkVYTebM+srX1eMI5TLoQmI02CxH+K45MHzujgRyCdx43NS03CmXz7N0M
fqDRqvTRJt81TOEtHq2h5O4ajLr384W2bIe10v0aGZ7BC6lAj5JpJFxEU37OJLDseLzgOkWdkEO0
YH4ffNEkNHEi+rtYxdZYjQiamzN625S0R9D8Dgje9sotCu2yMTo/H8I0ZtKhuMlS3d7zt1iyt7J9
U9qNIx6MliXb4d43CfC6AmVfp3rbRahNZIYAha2Yz7tzEqEbGiMvSzCqei0F/kJ9Y0k7p3w9MZSZ
MBm19QPUyrGRG7asgpwAzjuFK3IulGqEMxsU6xjbUE6inXfvKb+3CZXUT6Omee9uozAcExbElas/
Ug6y/QdtGNi10/H+kQ3fJDaS5jTj+bSAPheKWfBbHr5tSaFjr7iOElvvR4t5F9/pj+f8He0y4/3p
5XzrUN5ju9L9tDNG3bqz+vdR3ZABmH90H2YsVO+TRvxy7E7+dog0Lgws+9IH776vlVL7ijpY9hFc
00S1tkrg/gJFVM/RMoVQPJoXCsdp06FiTK/FSAckcR8tBnfTd//+7l/blULLiJ92IRhmaLrv77QS
nMxu3G+k2o9EmSONObXPwvx7hegRl/fELzw5wxte8K9NZFfGvusmcn9quqJ1EV/PfMUFF0/PVtkQ
rsqCDjv5DC37MuwTqW97ZTG9b0BLvbdRJ6e2RsjkXhBjAZgYDRcwdbJTYOoAwmSSsmH3lk/+DbkT
bNwrI1iL8krBSokbsh/1JrHBbEAIh5xmPlm2z/H5CvEXipldsPuS6/EJBmF5Gi4zVWJww19DRlSS
14ULcSjylu9BcbBy4t81Nc0XH+vPqe1OoxWs+ldwauyALaMRztjLIu5lxRmWhOBDCFBbW59iQe4e
+tt9b7oo+EL5AUPwI8ErLf7HHw9V0xTt/BqR0AavTQGwcnlgqQyFJZ/46Z/0u1SibNM7F3h76pq1
6WcbVjXayeM5eSTAsX77Ey6l6mbEh28WEEwBswkCaBUnGkPiQN83ruj8HOkL+dpOvkeC1VYBV1KZ
0M6hWFfX0Uk8FKAjF/AdgyeVWxNggRmEXxEHBBx4by3tHbMbDiho6F6/WmW4de8pG5S3HH/VZpnI
cWytYFwqnEdMCCP89DhN7nlEDECwwttPBH41rKHcEpdjUeI8uSfKM1b7aLY88CILxUfyicbwxDAG
MRXDR3vLIDsmHkqDHhIo2/h4Rw79GQEll/+JAf89d19HE3GHkeEB/CeI0uI2qctIEqdhzvywjjV6
ll583ZwR0HL93JpRHwVzt5EOxK+ujjgC/ZV27LsXfO1PTToiSnFDlCGo+uYbqhtWHZIltqQjYnTr
cHTAFHHjbs4RvP+afcM+d+1zuIaBZFta7el2AoTKRZFizfhRUnOQ7AvHnqetTk3n8eKVREESbYF7
IZMDhJKsRj0jDRBwdGT3V8YhJusr1B2M6KWGQ8Bo2X/ZazTlatn1Fo1XsWJz4KsmLcwg+BMAtfuH
7/3vnAulo2m5DK1fCxO7DkExgKnzdlr3PqQqBswawL3Yv9Jzvx+uhnLpf1VgdwCgOMwV+90QZ9sM
W6hxLIUAP4btPAslXOT0WuCcJ1M4Y8dkfqI0dlj+vg2iDdkESGv7qog926YatfSLaQ/f6u4nfyq8
CaB+PwQ40hY5EPXG8ri2xdO/TWQnyJEtVwl15/25P7aKvIl4EV/JWd2YyW/NoNJR0V3IVfEPZO6h
18mtSMy6JHxIDH9ggxbd/3lbrXyqbNAN0Ko8eyL+DiW897R21TNJnwiN2OYj1gO9yJrJT6o1Q9Om
OvAyqRunz1TGwiWMZXZ+KU9v/8UTO2Y4gXYRSenvz0pqjS33ZO41CXj3T1cLmlrIr+fHhA2XZ70p
zmKdKIqbeguHs25bw/8Y1FoG+PcKLc0MT9B283FQqbGJm0RQFmYh6DBkmUcCHnEgaY0/KzKuuyOQ
R0QA7OczYnwvslqFivxRhb4+yH+Bw3uXr8iaTsTkDx1MGSP98VTNiQv0DjdvEJ7WJvyY6GhoAcN0
vpqzPKag+3UN+Cj1z/RDPGVS92Z308S38UYXrZxxLrD1jqxts1RVI7Yo5NJBGeaKF6MjlujCPtif
tIhGMFqdS7beL34MgK7eZHwlUC3KCGNJObKTLwpTqbtqjJTLoGWrYgewAVSN2u1OI5kS0KCRZ9ki
jSmup9AVaNHgbnY46YhzIb4Q03z/ZMWTsSOqJFt5CDzSTFz7FntTIRjRVFsLFA7fwSehzqj0XWaV
+Y/tEs7qp4PSC9OW3mrtMffDnukg5LN8ZLA9PkD+cK5dxGm6FmfS5vHp/icehgB4iSM9UHrgscAK
N+K3x8F/wNi6BEJGxPR0U/bDAS8s5V+kpTLxxYFHPEPRPS5zuOdrM8kuucFDVhB3S7O2SCf0MEys
uNHKhQPwVUXxejxJugeKg5+M+WuRfq4qGchDQsgUD18sNU/4BCSJoWtLXqdZWcuEufY2nRuO6fkb
yUgRTS29rnzYEsJyPzcoEwYYpnfIdtOIy8IrA7NgBxNIDCuRQTFyFj4JJK4CjXu8NIpWH8xtoMg0
cj2a3fdSqG9kHBLK5N+uQaeayylxMB5Hy4bsT4zBhGFpmEauII5qiU6HypORqP8a/KY+X3tdLHJP
4phvQlhmleXgE9TWLRP4MvPEVOGg8ZZKGXDoJQD6rHyS+TprCWXAkyTchr+NSzmdVaoF22x8PuFa
1R0F/7DE1Wg30ZRPZozFvAstYKovnphuwh7XCem1dyQek5z9oD3xrqFWA6sT5/F94R91x5cdBS2F
1Ie4HFPwt+b30IFvDql/+ew+i4o+tN5WVAhZMe9KWdnrVsrBjqm+UNW1P5ObqawcOvj4oZblhg+n
xXaf3mbzbSRK+P64o9evYrnjcsDMcg5BE7TVcZPHAhnT2PxThohq+aGwBW8ka3VmiaekBl6BvVlu
9ev9KZSZujzu6mziHWKH+v0P+W/cFv9EQ4CEGkSvnSG0HFa7wJj1+1FrmDmh50UNOHzALoVjoemP
eVEk7jUeTJTJn8k6eC+/RjdVRJQfMtI+6UiVHsmbUEjKYr+Elzd6bjZEfDX3Dpfpg7HrvtCttNDI
2vw31yxkHlbVduQJdPKVIcGIcc06YJ7Q2oFAaY0/dEkgqd/TEERsk7iuGdWttaIZrNV+fza1E0Pn
ELgC28whG1I6QbTSzXgjN7PFDnm7LRs9KNN9oVG0ykAwmF6WXXWbRmi/nZGoDqlw3m8PcWOHrCNW
BxFvO1XK8rjuS4mIJtfT0JXbF1lAEpr4WqgMWsggdMZXO6s/4vIFCoR5Kxvz/jNC6dgkIsN9X26M
QUCKFM0Y+Kpwtbd5ZoU6wEaI68M3vyI8P3d2+qIcHMZv0YDG9OCsg7xKaJbUpe9yUzImlxM6Hv5e
RtT4M88/i627jn61DfwqJCBoGM6ePMqu5Nln3z+Zi4PfSyN0JRwYgkwIIhIsv79LB5Dgs4bDYT0n
mGMAWHD4YYG+CXLXA+iRvCnd0JBPTiN7uFjoSAOj8Jm8TJjUkffJaA2+7p4Txu5K3tHsB/xbgI/2
8Nuj38Q2pdlSkRsbtsI9s/uYsBv+y1e7H10NJjmjFq7Xakdz3Gj7xTCGMxZi3gduOn89nd2B72oe
r9p2zCJSAxQOnZcrXWqYtj73xflMBcodLTiq4skQUPBJJn88qoconLQI/SrbU39gXegpPVzw5vo6
6rz4j1qxT+zV7LQWSyl98bjb4ob28yy+FI4d2rMkXQ1+l/5mbi+ohjFSVCFxyfaXx7Zt+iodUb01
X6Dg6+8xaPbG2RGurH++zPhdfctChu6oxuFLXFEAOVoz7h2+kVunj6jt7zDyhBJKNlxFnPAGYoQB
FFssVEWniBYqjhjGnl2SHK2xqanIeSed51ZtyqX8l/ER10XwbFZrklcsnyeMBisVb2paFd3PUKTZ
Kt7cyXOxZ4zxWkZ5wY4IugpsC/vccBImJJzrufNM9Nylhkz2d0w0vwqeMhNieJYPqJlEn+O2x24O
b8pI7J9ePqYuP9DmqerThVGQfIqeIRwCKoxAu1uLo6jl/ZU0437OItUPyg4RkF4BNeUMeRZg6fCh
Ra2zA9mvzHLUs3Wsu2BAW46rHihnvv9gtDZ8g9nVLmaYOZO/c2OMgsu6DgFr1bSnfAltiixMlgEV
uV1DPErHKf4keYO5nwSwRH7Tp+vc9vB92nEHCBHpFM0TSrfdP1dnrO9TyL7tdIOqnZbFQjCDVN4T
yR7vxQ5SPgkpyrUsf+/5Zut576X8xCGfWqH9kPh6RjGfBePuhDUz2AMtqqoHd92ESdGg1IEMKmot
729cQUBMNxG9ug+hBy5FI4LThqtsSiQoGwcsI9J5FS51K21Xr4xS9j79NwOreH5dNpciL78Y9J+/
P/cqmNLjS6/0N3e+7QabQ9IoHSMloC3JQd8uv7lWaFtAdrqBZveKVrU8O+FTkEowxW6OvOytn/NF
eTz1bGF1BTBtUu6kA9w+0ZbwmhwAPdk0PS4FMVPsfLnejje1ka+660mygkJjI1CUL5Kh2Ks+1I4O
dxWvypNctAbr4n3vHJEZ37sJMbn8NEV7x0hWmcZyAgOMHiGFYkgeseYtafXr0dxQBJbZqDcNXBQQ
eSXqcAQ8VBebXPXmGrUNLCGOAmpUfjgdhkZaUO8RMtZhKQDS9hUQripxmBEgs+6SAmXtpeVWpl3x
B9JIMFH0wwfrPpt2/TNi3IovDXsYZ8KQRDunSFh9qPjR10m6G/7NP03N5AjbCHiBoLpnKimN30ka
LOuD/VZUPFvyA29pz8w8osVj72HD/+73XQryZF7cMuBfgJsxKPtX44TWSK7da1dhv5iOfhL2vxGd
7LI9XcUVionznxTI6rmaqw2dHSIull6Ksgyv3nMB3BCfBvpKv4w0nH6B4bKh1rh7HXNPv+jj/daY
x5eL1BDu76c3ScgYLnJp+HtJh8IqBdQVvp1Q6eJAbPgyNCbsa/x1QedoTCvLpKMfpNxaQUOnSg7y
vUmZ3Fzl/ul3aH77XMTulvs9+mgy7zX0cTJBwZeXJrKicH9F89nYVZraCJ/zIoZd93zQILgwCppI
e/WMlHFLoOxBz3CG/6/VqwdTV1MvWInhKUmIPqN5fJRzaovhz+AnD9unOo+esGpK34CTa8JxnCWf
PgBZCGsuolx9DqIByUHMDcj43OEm5J3dF2Rlp19aB+NzwFvLaGZ48FTE9oqc+zoiB535E0mQegsl
Hp8DrSjJWnGrSniyiLla838yhBE0byA/V3fpp9NPtDF6gJ9tF+U/yqk6RtAOstvZ1ldsSYXTlt+e
dvVoPjQMWuyQGL8uULcydq871Jysuoi3tylccd/ClVDWRYZ7H3nqiQ6i8LBbntxADOlbIUYEHaml
S7uKl0KAqnsXgrGibkB/F2h+sWpSmjlYDQoxKM5zGdN68Z5ksQaUscXaS/V6TZSn9xJJUNyoUORj
dk7qHqUiVm3qpqrhOxKtge8T4en6HQvnW0vmHoeNuxQLr0dimzOcwOoyUlqfEpznM0iw9rCs+3Jy
Xyu/w7cfBDtHLDd8Q6vCpIWdnIqIXCmGHE0jev0qoed7MFStW6ADR5Oo8ZOPWGaTuXqH19YolIUN
lCR4momJudCJyzHQADIbIs5rLXPU1PoXbyOMKSk3MiEWs9eJ4jL8kodZJtSk8JEcSqwY4Q3y9ZOc
taeqWa7cEhKyBTegfexGIPxuWxw3V0sxzEOBWjiu7gqWZQSek/d2Wr2jxyMlUqX1LWVzSfhaUZ21
lLL4YWkxvTspmJsVMwKswebUH/Vkn67w2VpDBICMzDtcZg4oXio8cnL2taGlI/MxdvgRsysYX+By
P9dRXrN1BfYgdJ6BeEUeNhB7t/FZTcdOaAMBChPPhaes/5aHfAR9dRNwo5ffGP8L58C9gAR/GLu7
cStD6ZpVb6sqV4VX96QBPh8gXFo6iFzjutEU/6HwuH7IRHNoAda7ATXoPCB4LFy4gC9JyOmjYk/2
+IPVptqbxHkhIGRPmLW+SB3BPV5bwHvPy9X9ky1ktxEGH80X6uFpfxE+XW19hr/S5ipPuSmo1S2C
nDIvMic67Ik4r+5I8d8cp7g6jZlQUnBsS8zWy1I6OHwI2p+JJaLlXzrO8p67EhvUR+JAHrlboDll
yLm/hy1qnvHVAVBWcSLujvvDUGdKMkjYY+tyLCRpfByavkpydUwTmMI4YdSuexA1q2turKfd9NAA
RY9uTZTfP/hs2YPxH0/xxtjtoe9vZ4OQ7oNeHmDhxc37hUf+AuKhNDdbGELfIrK3/b/7GQ2c66G/
zH8Z04WbbN5BTeTVWOl7wxna0HwWYmDd9lFnaTtGUss6k/1Xlp/Ww9bUADmoFlxc1KQRzQSHCqkE
ZZGSItwD0Ov16OFZN535/5HyO3J0g/hclCMyMarHbfHSUY+DE2f2kN9sFw1OHvHkhkUyYchtRj3e
bT7Gj4Moxc0JP0/7l9nV+tHOma4v5i7dnxt8TZ4LXk92PLHR9GymOLbMTzCgTylSZzPkM3OWWPgB
6G6C/wv+JBd9bG7NQI4s5xvI4iUzVrQs1xgnz6acYqeCdaG07Mk9WTsSuj+Dw1MD/VyEy268hL5n
DaczIwvB0cM8ufFL4WQ5G3uBJ6u5fPNa7IQslF0bsmUYMzebQUnDLJVWTQ10qmHIP/ab86FeJJkW
OmHDeBV21Ig+A3vRC+CPwinLR49i4H4CwHMIdqzSse55yjzVcuP2bUhRp4AH1HMsZbMd2mJE1GmG
gIw5azoEm4Sa6Bx/0VB21WFy7y58DhXHybZvaV5lIp9ZzRdV0xY7E1nRea4yw1ZlejRt0IUsYo1j
kG39wlC3FWHYHYQrMoVJW40tfCjH10ejrYRZNTzqE15T8esbwN1q3UnLiO2nAyeRMZz40IN0UG9P
vqPNVyvy6/uERXaz3hlrYGyIJibqsjlpq5HPOynecL+gzijffowVZqHjTmoxhCJX1BRSn4y+K9yJ
0q8otqGsNnChdrnW/02nJ8cB4Cnf5EfxD5cKZBysjoMMCMxpdBE2uG0cc6kU4ZWid98jd3ix5InJ
cM45E3ms3qK8KPu7ZOCuQQASwW4nj/u5nlSqE14eFdeGuaKngVg7GcoQMJxotUifyYS/mtEgz6p7
cm/iSPCu9hqtN56bpToljVL4ZdchOjlzm7cJzf7GDOs7uW/7j7hWPJisUkhYlo5Oh2TwSU+vr4oW
3n6iwr1q4MfmXTkSsYo0iRCtUI1WJ9n9GBtSMEfQiV7JaRI2oGpR7LVRmZOzQzLgD4azv9wxgx4B
DzoAbyeRc7hOVndW48yyDLJ98cFOMff/nsEZVKFlk9Mq7KlZXFTNXK+utDjUrRjlNUVuyNLcKlEo
vHIkmqv64XYXLDgGP4LfByvqU04iGyoVxVtmxYE5ovHytACcCK0bIxMzjv/LEL0f7XWI0lUgAjeS
F+iPV9wPK25aoNV3Uy5CGC2dgcyRc9ZSWzE0J/FLNoEgGzAnXcngODBH75wHIul5GiugWP/z3n5H
8zN1ePF0eKUcq5atnk/Rtwcw3N7to68rQdUB0/MVfA3dsWs+gv+PiNpDI7gu6wMBiumM2haSOamL
4vxFDgbUhax0BEtZLROQIr8Bl7zyvDjCVyDZ9wkExHPsEoDz8zFFW+lybRphrxf8ApUmCFTPLS0M
eImAEymRWVbnki2cbgSQViK5ez/RmZEj550aV6omDsmNGQPutTykHgaEhGq6SM3Bq/KH9ymToEtg
JUibG4F2YUotbS0OjEI3ilz6sb42ReAQNOthpwxLVi0fndCnsx5oVFubMy8vttioZf9lF0fqe5LM
gjOHDmCE1XwzBtACGvgQGhRAM2RB0RiqoolB2PDLz6F/AOmdEJaotkAzbdg5NWklQXpnOJFLfuJe
n0eK/mR0bsDRt4EWK8/D+i9J0V7zqCoHVewYq1Mrvny+vBl9QKcj75gmZz20j6oZZHAsYjk1qCFR
sog0jPtVbOC8swDMtmrT0la9At2u4HV4fGZBofzW56sLgfn9GC6skGkcK6xeM+nQZB11wipZnWc1
EnFI/8pj5HbGhc7byxRaKl/xrTHk5ry/4heX404hy7u12VytwDigeQ+Rdd2KU4xvADOBdD0iO7yH
Di1yLzLNwocnARbYpDFp9ScPdqtuQL/JE9tNbV6mGrfBLLYmEs1n2Aur6BqgolKfmEy4DbbknR0p
zJjUZX+DWrJrXygOhBGsJhnjOrmolR1hrTm25L86lVQ4qV3z7Pv3+p6ID0g1C8gpSwelfmvSdZIR
iUU5xrJ8WIKj3jaqlCNE3e6aJFrSU8pApVaVWinsbyXLDVWn2vtU1yaMa7wKPY0pGxZ8l6nRXwci
QxDgrZVvLWUR5Gg/tkWSh7Suj/9+IsSButYNvZKod8A5v38E7mCraj1LCQ+f3laOAm3BssTFXEoT
N1Y8eK19Bfqo8W5Ouwq9Crq66v0cjo2M8urcEW0UNUQeANHAsDz2SC2AfGhOp9yNP1aEnctQcuhK
jQkYphc8A0E4f7Mhh7rrzEpEz2RHnjgSCqxDeMr/HvhyWkXJs/ZwJFaTpSkVQ41xRnT897zygITr
v1RxVfWDtF1a0OG5pidr2XrvN02bzhJgugyh4uUOYom6scmuOrD5ADUpKnvjqwLVXxjOAFvaQ7US
vXQqyVYnKZRvp5aMC2+Dlq4hzO3QAfKyk0JkrafEz8qrOdEiebkio24GhqmLbsw6T33/uk1bpuI/
jJsfy6JqeH+HiIhji/HyhxkB6wZqYU93dBqoThxROumhG0q6u0Noe4yB4AhyB77vUVrcga3peLIs
hiKWBjMPm2i34QNEl5z1vl78+vDu87lmhWUDXASGmgEBvuRThM9tiwAg+mdGrb7Kns/VawWo1Y48
iPRep5MJ2wfnhi1iK8B3F1QzOc0ChV1Uigp+LwvlaFM4XqiIw+nWdNgsUfLE4LCinF5iCVCim/WD
euWAFZ/wyMlNFYytm/WO1LNwrZs3S5PVk/MVCgpbfr0EaTHK6eNRQp8wC/AUkZUGYAkFYWWhDByh
zsqdWeW4M8jRsrAeRJnfZZ/+uyELmNUXbiTBHHWlVqZPTW5kdwRWKyYpeaRwwAdEDcmCoHtjHclj
ozYT5RH4mrtq4pVu2zyTsRzL6xNt9hWc4Uk2Ax8msg0UTDK6brOeYOY15Z54ckphM/MJMNpqReN3
WxZKJHttUrv7cCnR8iwnVCQtiQdQSINnJMeF0sHyMVR95mzmBor6RYRZKv+C5qtcp5XG9jzyxzlo
Mo2alk55xAshHNM2PWvL82i/eKDdMliByXgDJEYpxh++vwhDkMRPM3yecgG3qGO64t0I4/lReb5p
tHERUFi7vicWVaYRRNP04HGwoBsiSaYl8++uM6M9q/8vxcvjELGfoC4VyKXXfVGUNRPhbELC0mTA
TyPUZRnBD30MZG25V4wjwcMdbGGxz36xPZ9whWptqI6phrWZtadp+h9D3KdTReasXO/WGoKpUOKM
L71tWgjKInKQU6CES8zzF9TxxxynugmrSso0E//n9zkyZ8FPdncQicl9yyQCPRJVAVYtDuWXiDRI
DHqLFcsNiLs1AhhBQvouEYpBkAj77cbTK6qeYrn3ICUuMEy2CZXsBU8p08mx7if5Lfk4FBkjmlVO
twMTjg0hC+Q2izJ9IFmN8JmvdNc6zU1pVmf8yUu0bXHp8Yx8LSltyVk60DXx9dcyB4yHf2U0pWII
XARoELYbn3d/cFp7tZQLSqYtCzJwKtPSD0DdfPjLNIp/Fmzde1eaekzP+jCdgRU/Gee8fAuLuzFL
fgCsaO80kjS2vZBt9EgDnSK+nBRBSMuF/xxjk4UenmmDNUX9/xAiTM8R5NhWjL3MKk48VHkJhYN1
qlRqGymJd5lkywSpaWZLPWblC+t5bt2plV6oIuyMZFcZNdbnQuZK3m/2Qvlx3TOb0ZkoNg82NQOF
KuIoJz8CE8CDD4gQWUBEVftORaWCHcsbTfC0Kx1GYo3evruN/7ZBrF4wpmyvDFc55vqJlmmsi5Ed
9hGJbjQPtcxBYdAyT1RbPpFcg/kjlxJxC6UAfqczYQm++CBd+QjLO+5rWXw4LXOcb6/kOI2qbhmq
zK0dx6nnYqwxwwH1/fWIrUacxU8X3eMan2gmJLbJgkuzGbHFCdcpAD55qOdRKQyqs2VyyfKBJn/L
yHkz4au1mUiNGe8Q5uZ7vI75pF/ebrZWQMqt2F/E40EEaqcgNyh9YyHcqfdBQwomieIQhJvccHwZ
sJm6fN1PBeAH039SHRH6d0aVAVtUe2xWfxz84YhPq/ENzAUhWDC9lMOWKiWjvxPjA2rKDqGNIFas
RE1PdyE1yU2t9YimHNPamjIgvMVSixACHhWnV1/pf/D8EVi+jDooyszCrp7xH4pTQ3e55LszQj9U
uQAm9EFZNU8ALd71zwGWnb3qxsgNhw9AoZyPjR4CUUfXyY0NV3L4JKXTAGy4+Qi9z1pqgSQosRLo
Fy8ryNYH3u1gMtCs0UlptnGI/Hnaonbi/3A4T3Oz42MyxwNYWhwWiftmxnoFj8SNl7y5zydmguOp
JH6IWgaowJ8nE04LTAhdLFM7cOVdYOwNcD2WjaeFeFK9iKe/+EycGxX70Q7J34wLev9E0zcUWr1V
A58Huh83F7iam+O5bPaX4sIwDIIRUtvhsYgCV750V8uSmDIfka4/f88AArN1odk03tEDlRafR8LY
t8RiDHE9/EIOnjZuj6fPn9Yg8Va87vcOWwwapQylWSAnrPvtgw4HgiSbvCZrwVQu8dD/P6xQAc8g
rOgUSrK7NNWjIhk+4TEQbBHcDwHjXHMWBEonEGdrC3wSOa5zRSMrJwAF6Bs9jkJXHiutQDWq5uw4
04HFv6wOYxHRqC6fp1iiWrFbuP3mlYJajhiyBLIycei7IsB6tKk33jEEKpxfQCUiuxIIXhsLiKsl
rT89FdzqAC2aCIU9pUUzDEHzy4NZ8MtFl7iah7lA26grCFfQCKwrbEWNVUOVdZVoAQDICM8hitVm
3rE0x3gkz3Vm9HSl1o/mYF+S+SKH5jCSVt4xHKjq3S4YNRNP2fkmnyJZ5RndIYxQU70Lg3F1OzHK
aZznmdf4wsDbxOhSNVh+XbTg5Z51Tm9EACs8tIHVOdZRqZjFD0e7ameP6Z6Rw3LNbHMDOkDdij9q
2RGiScctu74YUDAdCcAIEtkUpmnYCc/I/5g5B832B7EsVfayLe8kKU3pfzyI1uA72eRy++hvhrUr
pLGuQJGvIQ0Kp9mcy51qZ/e/KQ2TlztMmkMC2wjAI4OJ4hJ3YyLhYMiWI/WdwT7p3HT44IIGFe3j
g5GT0witcRvGEXSTnomCrvinN1Us8PwZFvhWwH/vGolzJQSV6jaG4WHBzNFUFPbM5cITsu0qi9D5
yzBGkZkpza6acP9QbFqZPP6a3bAummtb7uzJ0mM+SVmPaheErTFk5Y1+stOs5okmOemkiB9ERN0V
zrRfTQVFGQSH0efuGwQk6taadeWO7g4VFChjFulU3s7KS4rOShaz1YuKUFaExUwsFlTP3mm+Ecra
iDaTGgL4ot2d3g0iZYwtrJWArMn3y5sjhrOC/dQNmNaLWXzOkCdLxQIufb2AU+q2QdJ777FjV7qa
cbJW9TwSxjSVibsOmVYlYFrz17e2JWxE320OXvEkBamlfvcJ5JtNAWF1gS09bkf4h29iTC68gyc3
piagDI1y4laGQY0Bqhu7JwSElQhEB1ep/CYjszGh8LsarUTiZ4ejJOukzgcOOOLY0WMxrjXh+GYx
DTx6M+lOgM1RqXWVQAt9Ec9w6c+Cgyd62hy3mY3dNHgfVogVjJEcgyTljCNQKB9j2rCnx5LpX1LX
daY1XDl8/Uz1xwpmbyfsXzfCGuCXmXxypJRsTHM4GKnGPIC9+L03rjqv/OMyDeTtueW2qF+m4VX0
W52dEFGRK1qwwsXy2WVUU/vlaGIe4O3v52Dr52KibWwUFUWL/MkQupvE9YD9Gmi7/dhV1g5HqN7v
uhi563fQH6QFfMkJC4AE4YiqJf4KCfMsjR03ITyowlPCHPFPzuJeN4atL83iwUuVYXSJ3N7CFdx2
bVLLTc88lvn5R8nWAt56aRO67ahCJBN/yIfBMYYHTzsES9X0h8ZPzV+4ga0eza6NBhHuwUS0tG61
aTtauW+pWPSoJfRpYzTldOxsKUE65wJI9aylsZgd/fR0qoqogakcQbjghVNyD6CmD7/wzCeLuBP4
8XzzyS8DadABLyMgDh7IwyAk4D5DzAv5oduo2c4AqNckAs3r7hcZRSfRdn15shJ3+7etZZ9yOD1u
rcqOLdVsBUPQNnJQoOGWdeLrbhrtzbbT0MjTzyTh9G8V7OOF9SHvZ/saHhGNSeyt10bX/argBM4H
Xfk5xq0+WBvTZxSV1bPl1Ky9CcGEnDeyJ7rNwLb8a75JbHGbHWZH1UTkp//JOvzm9qE34wMtuBeW
UswRH0iVNJu//akmPMh4MAXM9qzRDn0mR9mQmskyWX+W7GMB7yT35uUdpR6fNhIb0vx696YuIGVA
MhtOkc4IOuPlybBOlkue8u0I3wURcIqfVu3N2i4FpkMpxInH5rbQxDGhR0pDTgmnG4Uy67s2eo7g
V39+nlbjV2xs13LrCHP6BvV8uMAq5psFPIGmU7jP9CBK5j3BMAmPkxCnMHy86oSGdACpn314gZEg
5Gbhxw+2ZQqw9Gnk475d+4PT5xuYygf7mUdYPcfID7DNgIH1rLQ5GlMFQneWQm/yj0YVrVU9AnRg
yF7vhHg39vek0gGM9pZgYoUCk4u8M5E6PPfbPD/FeC+9arNR/ZOhqEj5xjdQLE/QZR45OviQ4e72
V5JLBkOz53Ubmb1QxneObLpbdYezoLQuXhLDNibW0gXo+xbr9H70etFKspQt6o6ctGROmCLdimI3
JVCUVid70WfrpV3tJpVxPg1NjDlpL6KAVIX6CzPkplBjjLeWrYKQnUCayq+DdbUBte/16gQjiqLt
3mBu/ev9DFIbO0DuTU9tpX2xz+jUd2Wfq2DE7IGRRHX8XvkMXDdMva9NcmtMTW5yrjsktHsxTgHd
rfvl96J9j3yr/eQJuFG+gDT8uHjMg63v1J07gkuwz8Z7auLfWBrpqEmW88E3J6L4MCM3OsDO0DvT
o3tSOjQteUCFXQPIIaWwGYfIRzxgzpj2U69zUsXlBrkPuhiG2abaM+JIadWNnlBmIQfA7l6NU5ZD
OuxoY4uwpntd0NgAvIf/X4okp9XCMf2wb1PC8s5BqPtyT09a2jpatxnMkOwtNN4Jo4APyrbv2T+0
myr8x4cKdtb8MinfZT6cJsdt7NyJHKE9dOOk2acXOSNlDBjq0vuyTgyJdK8rDCQXZr2J+7K1gVB6
1RVgTZW8qoO9aaLPqq1xC3X10CqjeY5L/uhuDjXpjdLBrdhZh0rJcb22OLDgOrW7f2358HpMj/6s
Nc2E6kmJRd1aKwxDpagtbM3EzemqNkYaA2QlmzRVHyLj/Dap4hUe7fkHxJ4rV+3oqS+SF5+phQwS
vZIXr1g1fDiA+vEEoKkjimwuOS3fOwRTv1r17FRX+sttOrqcZ+K44KHcDW3FyaLDl2u5YBEX3vya
b6s/lg+cA3k0hc9ECEUAHZNtWk1VzkbM4VcUIiTezEl13+d78ldpUhsdlDnUrlxUwjU6FSNkdxIA
EhzjW+hKSYTGeDGepds3dTYLcbucUtpeRRayUKWckv3FhsnpMruiBi6Xut6oMvVF14E0GcYb/KWA
FwQF9fWPJyzvNwXbwbO5Sr3mfCt+fgzZKIMQS8ekTxYWNdOqFOAEPVMxVO3Y9ehqhQWdhJnBGn3c
Hy+3YNRYtNH2HTd1kQkbtmVA8ROby33xIGGmzpXKN4tnchccEbehciceP40ZnF48dw+4sOEJDF21
1OvPVBiY3qL3w/cnZB8fRZvx8r8nih9pg3mfieBHaIzdLwJvrs39w/unoHbariOQ0dNuqacbJGld
8hOpBfhJ/ePgDbOAjY5mHQ1dRvfKWIOM9l5F28iVRrnsYpbmXilsewj/fNZDE3AY+2BXYbmJXeup
cVEEReYVXvX0dukrIiQ8v+lNYzth6c3oftw88v2pwTom25j4jRfxR3f/OvPQO5r2bgEFwa3XF1iI
AiL6qHw7y6YkAVxwh6Bw2hOqTqCzACzFnxMR7gBT+aWxRhMyUzL93FuzY3SZL/QjXfpXAAWa+SlV
ULKsL6CbDAgavEHQDDku4sxVvg0TEkBRVDJbGTeO02sTM92hVyLIHJYwkH+Z4uMyb03FIiJwa2WI
y3iiEE6CYuuaB4lIGseY5mNnQbihypbvdZU8wqh/CA7V1tth0bwJAIK9owdawoR30Q0tyhSIQOH+
Mjqwqvu+cflXWj3KslQ4tzRNR9Ajuf6Dp8rGKGzeTD20AhpyGYZnN3rR8Xu2DJCpghYNmkB1zLM6
AKIIZQbFCfDlaq9pEY8zWJcbNiTGcbXn+Edzvh7U64v356Wvo98lHHY1HAx8L2CW3Ph/uJ9mQmp1
1zI70I/aICa2G0AjWTUTQPnv+NmY8txNn8WO0X39EY1IvHFcLpZ7mtqzI2p1VQ2OTGbzb8i7JigH
M0hRabkc7XMOawHyfzFIujbbxUIV+lOu/U7tgCOQl4q+bH8TRAaZZlDzl8lpNB/ESg+Lk/xyNV32
Ckx+xxGy8tICjqbBlza9wjPsQIiIcNlOTxKj/rboCF1TlCWxVul3nswrds7bMJ7FyztQSuQqSP9y
visae0ckxHeyMHizlG5KiZKGetC4lmykTBvDEdMkqxWn2Hvvu2VrmgktJ/Zgp4oTjkXqWyIFEAs3
VSRvq6s2l8IpX8BOXzCYB34Dv/fdNlTKHVUtx40A+eO6eGYKqKCFX+XAbQcTE0rg9WCqF3SgM3Tz
boe4hwyH6dSrcH/W9WAcPCWZZtQL7oEySa0lr3FIFKE+fpIE3ZoKgvftXh3p8NYxSLZRnSRpBQfT
/wfTGK5RtrFEUFnMrTS9fva+4Do8gzuVQzg0TG57AXr9Q/xt39Ziw9YMgxhYKW1I2vA+2Hd0O+FD
CDuBjFnwQRawJsyRfV0WP6sCuRQvwqo2aph/cXPhj0l+1WXluLrbWnRPoSZbWfmTmHfy9tn2uZ5f
U6jx/lVshjqhv5CkxvlGy9HaNtZ7ub5XLi1xApzySOcErTKksapCm0Jcfas7afICuojz8yLaa7OZ
evzYBF+7qkO+EjUS+BqSAhamAh6HH9f1nmZY7Jg8af7w4rJiM5jH8q6vt+kdYnZq7+ZPqSqs5XJo
JKHkQzPxBjt0REQn0QS5XoYaLreKu3CY8DkG4KXgFonVZwVek39YD13NPG+KlcQbM6dYk11/4Ohe
LicNUJUKQBx6AT97zRWqJ5567Wcm9ppCdWz6NZZmnz1aGZR5CQH4MO75JAf4Qw84aV1P7zA/1Q+A
gTlOfSlkXHCq8ItUhyE5Ey8Fi4z2WyBQNqQvHrZiQtIMDAC5hjsDxbOKvLeTN5nmTtO6XN7/WqGA
dLs7KZX+n9+ICVrjmQtlPZ6IJy373sPrAxn+bwnjcDY7Cdum//uGE+0IRENl36Su1loLOHiSYcmW
F1JMWU8K9AjX2LzeZrIFnDOK5a8dRjT+M2ig/E2ovSmb0YWkckr1xuZL4AmQBqUIQyuD6qJi/HBK
Yp3izidZEuMKbHQfCENtcEX96z75netM/G/V9XpeGckkKW9OV3/vLl1z2dd4neVhrNJogV8dcz5d
CT3bPbE3mZwHFR7WZEyh9QMvCLp4qzoLSMrA0i9duhsWi4mD8Mi7SICswQOTHOgPZrcUa9de7nri
lPKlB7cOUTT3BXy+7H7k/yiGoxQkSwH7H3mUBynouqbYkF9qzV0J9dW77rKohN/xY7SIaJH1oiWl
XJq8fVX3nJ19SVOFM5EjrYY53jsqRr3XH1hWeKi2WjB6s1Qp6c9fqfGpL8t2f6GWAyv/GH/JyVDC
/+INfIG5oIg42gZdDczw9WH0lKMuLB5Xxt9r9uzmc3CqQDd1iqWpVSlQCmbc2Lt7FoojiX5yFw+t
U3Z+jWZ0be6qh4+j11fgZY7Bh5idzmU5bKod2u6uA9vhEeZhMZ3kxT7YfV5TtbGKRWeCTns3f+gu
IBoy+GWqd4qJEchY6Onu10woJae9QBKDfl3MCVTLUlThdflghstU6oEwkrDGH15ySojI9UqiW8Vl
J0VhEgDGJNsIN4zEW/NofJ7OWWNwLZ/pJHpRq2SFnGf31YxH4QNJ03VFqgBAc2NXa6sNBnCklFZi
DOY0YCYlfhfcp0ZMHZY1rmDF8eClGzl7mWk8hjQ1vPusUDgzU1q3YNfl3hqB/aeWTule0aCNl68Z
ZQI/9Nuv143gq+i3KT7mmKOCl8QC6Papwfg/zwNXuyRwfUEhyr2b7tBgHkN5itP1fa00xmQmzXtw
qnEGL2A0Oxn8O3st0WgSHblNobADAbDE6pApWi5b7aCkKQeiyEOtYxuIwTs8tdELAVq3ZWz8KgXL
/fglUNb0Y/xF8kwLhQTT+FHgFQRWtThFHeg4V+EvgVDNjCh8GOHLM2oz52izMFSS7JQYa6c9PQnc
Zz9FXGIAsJg4kLP4hvnjmXz3E7AupmVj5nMxmlz+7TAEBJ7oodSb0osV84ErGDxNek2tLl+R6s74
E4vmiQlVD+is4dO8AqjRHdpmlpg4KkfmmYBJIuXirK8W+UTqkQ/c777nKYQ/dP4VdBn/9xSOyFgI
vE9alghUFHzodppSS6wf3DL6U3GFtHQ3KAgA+lA8PWxtDt9ZpJKjF68fBII4WQW0D/KReap3QGb6
BnpZ6h0zFpI2Ip/slsPSyJ+NDLWJ+HzUQqigdKMJXytWWNzSfFCFfepyPhm1ZjwTY7+Em/9PGqgA
4T9SBK+13yHtsWpbg04KLG97pUc4MWJcRYTyLa/CO4Cl6ERtUpH3pR29XbximMhCmCzwQm31ndsO
bQNAydEap3gtYDfcZxzbeN/wJOpEnWyqZsVCfodtyTlz2zhnd+uWa6S+JFudEZ8kynyX6g8bOyQ+
0PqmIMVwg56+Ou8nxXS234m76Y/t7T6Uir1gmERcQ12hrHVivihQADo0n+xm7eVvHuhU6hCnn4dT
Ssxd9ifM3C8lkpziR81wxJOULv2wtxm5+KiFyRTS7Zd3vtS/1GsX1tsfSRHNWAzr+hWbyu6R2QGz
EAdND+4+F6euLeU7Kp3zNIbKusc3cApBF4J0UrYvWYkJ+rTplQ2Jyqru6DgfCphSMlXpnziWGebu
hEhqn5OZE4wQIMwYtWk6XRuDMp6Qlnc95Ix9A0wZhCVe32gsDa6HJAN29F+3RCJ9NOxGEOYenMlM
o1W3OMSqGnBJ4ydFHNjIlJ6fwKyPcsKcyoQ3r+Kbs54Cpw8IafSlFP1UYcYXA5UDMlftuH2gKR+o
0+G6LdJ/spm6W6C54cRu28FkkJIgun8ExDr/3mkKP6iQgvYU1O/AY7VmaNWZ8JbZBiW8GPRr93gp
uzBXafK0px4xfCe/A0Qj+wgOJds/SIteswP797QoGcoxJWi2WD6z6jpiE0brnFLDl0S2Jgmlzuhc
aowrdBB5aQJiRQepTxI25s7XNWMASq4Wb4vioHeSF+LUep+I+ETV7ZB8zE9VqN07XYbMSfa11QBN
k/+Tb5b3LdqQHL5VtLqj5mQVH2Zv3fWwmOZuEBfStmgMdPkt957BmcxDCqFoLBpduezckzQziosM
eKDrKgng/7Il6Dy70MH12vc13JuJqVa+leYiO2gXPIYAMdGhun/MsgR2R2XawGPiudG3MFDGDbSd
tL/Au5SDYh0Gliyv0WJUqnvsLrniQuvChOAZbpKiv4X/yG50u9fY/VeXPz6yMqreTAad9M/99fap
Fu1TAHDc9a3xgMVfLozStzC3CdshGSC5WGteXRo9+WV1kgXbBQ3+YvPk/Y7vdMFQKujVGNH4vxyE
Vi0DMcaqPk4QO6TiS3NCfF80RbfRAXUCHDsmqYmfUWhtryVWqkdW1z1uLZJCfakkwv/pSIMePmGq
c2KG9h9bniEzyuczas70PmfE4G/n12CElbLSOwG6mGazARAQNlCUZRNUNFffKswx4+1ldF1zfoyX
Zz7RNWZ2bYKML9DwiMQ5LXAoGLdVnBPn/Ps1U9JHCLGZ1lgG6O7trbLPudUBl/S1eilzY+294W98
WfJrL3vKEHzQ6TZT0yvsJhDy5fs0R//DA+1OsMxEzYOPv5O1XwObyM1dsdFX9AyD54RrUduJNuiz
z7V3g9N/eOHSSSyr9UAVezRwssEdWUFFPXZSfeW+xGkAoGyHErIqB+GKpHHY7TFi5JneojskHDAE
Z4No/tjfpTDBgDifoK5eGUY2X2BuZvfQv/fZEgRjUlKeG6LSIIeJ+URVZFX5426v2DerAMyS3wZT
HlRu0aCzz7+SveKLjfHxj0ctTO5lgIkqoHuRYAbtBvrbbLi8hrcwJgQPM3QvWHnrTBy4pseB8u9/
0Afxtd72IwM2F6NNjR8kWaYFABJsitGqN8/B9UmO/f11k7ckT2rHcTlrwyKVJvnBDAhhztTh/zGS
zbBILipgznG4MAPOaAnvpopZt8Q96WYjp55Xkz8AT3Sx8nMNTFo3TrSHow6xZGSCpP59Btcuu3xJ
C7UXr8q8cHMZMgs2SVefP1eetkcQxJhIo+zlNftdEsped4QeTLrDPx8QlT8Igo402YqiwXDN12SZ
+DBQ5g9HltCSkgCW0wSFxATFUytiDfpjcNEOWm8FAPxttb9YFZxxtd6Q4Icz5t5Ux1Y/TKFuLMlX
b2uMklIcoxkPHR2VRTHomW8V/YWLaEX7iABXgbugKr0foqvoiZnFuXchohfbcWQxyopChPClzXRL
zKcuxjyiYJezeJ7Nm1lIZATJptftZ/JOhrg0mvhbCU/60esrvqOuZWHwlfxaU3mfMTApHLGhp/51
U2fFUY3vIjKhK/6i4MsUHCH2CoT5tInMu0IjeJm2k74uBDSXYnyXZcLIuQyzoNo1lVQml6b7sXfb
pjFp8z7yYXooTNiujBehjrcsayF7OMzwMU3zGEPzNKZgkWcT8/MjsF1irFxzkI8ItdEqOlwnxbDF
X3HixOlvDa8vFG4YMjVhM04jPGCo6LRbQxGJtIRPB/MQKHIka2VzXfmppYseJWwwgL4MCJ37ptdY
3U99k/pCLL/UOQZZt8yivxXEEllyKNIQHU15r/THbWjmntiriF3J22aEWfUGZwsv2Fg9LhaTWqlv
vDKahiu3agnSRDRIhXIFLoSBAUaLCi3UYGARzAL+KIQ5YX6/M1urHvEZyh9s/qoi0vbBXGHo3McG
qG4fE/ZhmdRdMLyufUuq0cQ9JoqVkouxG4afzrvhKA6FDQaLI3v8veDf/phUSyaSIEH/Q50X5GnG
6hOlyvvAhbCHoXqV4KIRx3tbKRcvRmMjlJeHeyTcH8TmSmk5la+F2zWOKIiixvjPyYxmbCDYVAbt
7n0hdCKPKZCqZ+1hSBRxZHGlpjfWIrcx8iiwVxo1UTCmux22+SF+CDM2B9jep9PsOXb4/zmp5OUA
wLTSbTEKEzDLR4A10pqTTLIUfiPJ/9NRfKenkdj6iLViVZXhXP/GRzlRlTTYj1D/7VMkv3v5mdXO
XlD8Ddjrv7cVqB1L4BTyI0dGK+R3XNbO/Ykzf/kBTFYWUKflpD+9fMNR3BzE0E+t3MzUf3pKDMdE
zreHewJTQ1EvEZRjWOvK7Jz3dfKRIOZdBR8AfxoQwD6B92UWn11SXtOLsQSvitR+wXwji93HjxWn
YcMk5x6PoI6nTkPC0zWl2jUS33zWkvHvpdJpVJHNemotCpx7sqt4+ZqwbPtKeRLiPssR0xXc+XUu
pwwa7efnEn74PcaR5iKr/aJ3PdhXhc07ULlBZxQbhzIDabbL5YCr6BZEZhZEIJSxt8GpDgddyKpp
H0TakqfqRfFofPySUy+BKY21fE8dD4hdndRaRh/9buzuh/T3bv+5vn+s9xNKEd5qLp7rreulIEK0
zq6lcdsu5FA+8s1zNSe9s/iIn7gJlTPI9HMOYvt7Ij14lNn9KX3MBKdTnQ6iHo4TvrQS1118yYSl
5YDMEzREB5IiIbXL0/3zsCd4ZY7Au3JBUWrtjvtjIjVQPSl+SjLZvrkWpLdWABucQT6KGG1y+Okn
R0TRgY/PtnkCC5WmFDAjZLXeidP1ovuSEC4tHnIJrxRndRWztOfLV1gh9oH++ymPHPk9kCFA8+MM
akBNPcG6WCN0r0yWngeEygwws9o4MFdcw4xVE20t0eo67Bmo1EjHA6u071vIv+C5d0i264Xm1CFr
c0PIMr1j198vr7rJPyTmA0K00+KXxUw7eixz7vSnYYUxz0j468rCtx+IcDIQ0lYlYisjxl9kl2XI
DNoeSNQEfBuwtTFfnln5v1Fk2wQWE2r4mMh2NBfYib3FjXYCOSZ9xB9ocSXFpyb6iSZR2phF9ymQ
njZ7tZSxYLJ9TowLr6mDmjc3fLPP4NihWf6bGsHMgw6jjqqW30dhWmpVefhuZSQTeaFcbY2rk5Ip
C3bDr1H7cg62X8Gj0XfQm+90u6g7DQ1msb6yflBCa8tCLvJuvlWsOruVTJegBWccvd2N6RnIpL4+
PSduMh/Qa16pVPfILfbG97mnUA6DBnB6FS1u0YjBZ/ZKG4Od4HoDVuDBNmFIdlIgCpzfDEuXRpSF
7tiInprcy8e85AcWRNU15x/eZ+AIxJjFOMOTZUJGw93D1mbdzfUHQKOWGsWEYI87+vlflaFgVKd8
ax6BEdHuoU+ydnxE2ht7V+mvBDrVXmJgS8LKIrOi/EL/D46hD1Igt6vIn/D90CSp7hwjEztZadwH
KHYe8QmpuOa8w0iLvLj31gGXCUKWyVa98Y5m7kwOqldVkYexwPdrrk3ZSeziU/hn/XDMILUeFhu4
5WOv5Kjk8AzVazjs7+6w21QnSryGTbIZ/SqBh5pP+1IETBoDMKjXKeeUD9uIEISB/pIIAhVFUxRI
lyFnxYyesgaDNApQ6UbA7Yg7uRWfbvTLa6CSscuZE5C89EOcIEL0IMZKJP8crw8t8CdVbcP/FB//
BlkbArCHciydawlKIrApLU9cfX0bLpAzEi0iNStobDoZvjcQzMuFLgs4P8qLJAfbhwy8ORXTHRKa
6hwu2IiC/bi8BEdiwW7Q8tN5885nWKEmqd08P8oJhQ2byyi5UFXoQYmxBFLqlTdpSOlHAXmqn7eB
LI1TqElePzcc5JvkaBHYGER9Fy43P/N7VGLnTg2RehfkMDWaN6v8gm11mlxI9LJbMJF/M/KFRW9b
z8uw27JKt3kQ78/paririuizX8m8mskb4nIxqsrrVDgQjZfbBJAj7XFUxjVUU3nagRR4/uy+56pH
PvypmHfExn0dqj6ivFk2/eQxdCj4cmfuZ6I3gfzWiDhkKaq/fqt35DhbpCrnZ+BZOrDj3ZyKgfBq
j4sjEtei4cexbxtvUi9TRoNr+r7VV20QHIw7JwJKLJch/uhsL/NXIL7tYBbI6hHyAdWtXrJTYVcM
t4zQAYKIkMUfUAG+vkll9w1QpzXG+vnswvKxkmtDfzTpNLO0i6jc3NenOVeZR1q2v+xgyQ8TI1/b
1aXbhiHVp8C6Toa/LdmI6RSZ+KzG6wKaKly1zhqAWjIsnVuscHzNtC7y/KbaaIRmj7Ko67zRX7iC
6SZ7bAMPd8q00lnzLCN4DwlvzMP9DcwyljkSGqsFHCryqAOsaZNie2LrGFWhcSzOx68D/T4l6yXM
5bWxawVYf9aWBHhbEFysXfX8xJ+hv+xqgcOYhbyoO48zgdhLO0UUG6pHZgS+OxbAg28Z1ZUoHYDv
OGzr4iLO2fm1X1BrIsipEeo3OjxMiiYgdwiHy+UCGtWatlgEj5L3gEmDV5QhrpGjFG0JdPyD9+Uv
2LNnn0elBh0IUd8RkQ//mQS49lvhVSkeFFpiuCl3E96NVs0MDtnCTbd8g/t2ejMYvmlidb4m15y7
iOLXGWxR9EtgoyuYT/jV0cj6GnAFCJMIxX8o8ons3Ve1dkXQNT31+L2ZaICVkL7Fl/xa4diliziz
KRpuzVGfVP2B0MjCuTeabFDgcDx4eMTPPVj3STiLuXtTMsRJzhG0t7t2Z1JDDtPz1ugeXPSdWjD/
hVGJyl6nDdSl/sw/KxGqOsDtChyJR5jG8gYQjvgbB+Wy0rnbdWZofL/p6bOrcitQuECPeM9/clUr
EsXdWMXfS6ifOBbPgFfXP6x/eqmRl2ert1empxY9noxRrogA/xZVtZ8qQkiW0xegr+Q/XmU8RrcY
d8xlcItvoYWeG13ymd+ihPBnwdUfUHDsFtHXd0oWQDN5mMMZTvrn58o9lrG9caDRRKNenCW02qC9
oKLcIPm91jr0yDbvs4U20DyAlSdzJoXdGXZll4RnJw+Z9PfNr3wwCPyp/oTbnl1mPNyjIXDoaUGV
C6C0wujS7UUjc3B8P+ZaS8jmRbZEkvpLxtmBuM6BJDjAbyZX5Vw+1dWZPbBVB+DCxpyk/s27rkUn
5NGJjSxmx8rOocCkbV82YERRK9A7PLN73UVuj41KyTpjMoxpdDWmH7f9kW0/UO8C1pTDSMi3CvZn
eKFTAXBfsfpeUJnaZ12RWJNfvm78v8wYtWhW9mvjx7nrL0578qNJCCXfB9/d/lNVPys1/vMJSCoH
/qhuSIS9VB+Rhxnsq2Twfit3FxniFJ5Vm4gzLr3pxyKhTK8Kmm63YrYNn+3tzULpvD59w6i7FW6O
cSeySmY260C/69lG46dXa9BfFZraPzSmUQatT3bM2AvlpRkCGq5fueGeYteR71hHUUv1lo2VFpiC
pNPUDt3ffv1K63Tlq1GRZQV4Yo2cjalt3G3EoFScx9bhWYlZ1rKOlcwF9M/DltUJPjzyyh0HL3gC
h2P5SCTc1LN2VHcR2wHEQQ/41COEIuxokNKOjC1LL+ch40coqvyni2k0UkH4JtjfUsQbYf2nW3Of
zKFD2eI5H7CHG/6I8j8AMk6sn64OoT39DfBC9Nq22kVgQotQNN1sByNG7pdT/RmXCQxj5pIoJYx3
HzAv0MCGjEgw9CuvZg/liapwhIB/ANXowf6tEgEshVtXzUSaOhuNr72ZEnWRBq7UCj5qp448+sDU
oW0Qpvssqjcy0D2xDXGZ6ywECvaGfMOAS/smELSQIMHCeHDrTmIlRW2urKhMDcKRmMfnQdunkruG
sfUdoO40gRsDjvm8n0BSYrzdp4nGFdmcpN4ZSSZSDCohBblbNuE/8jG0K56oY80zSs9mfBdbItsc
0gNTjnNwRoZoGIE5XCNEl9GKSkIbE0MPjFoo8WEdTdbytzI34PAR4G6JZytoEecnI/qCDrNfKTs9
WFRgZMHNm0RymQoMPINJ+/jUO5SwU05rcM0qH9BVHvljJTc9RWcx8emTrSr1nkUebfUyLMVohsyh
mCprGe4q/Wg+cKtQCehv/q2tyE7+gTqqVlGVLegvTIc4/p5THggjFxFi1oj+7JBgiJLTHT/6Rkpp
OdJgWN2yJzNcQFF5I6Pp7O7iIIIv3dA5763uKjiu5qzMp5OD3irgnFg03tqGzVM715gp2jCuww2U
3q2XCeo6nCBcEnHAZ5u+PGXzxEUY1ZimQRteVVXq4K8wC2DHmFkm3wFkLRqN8haU5OSP1laCAmq8
YKZynghmW2VJBlFa/rfrdZrxOlux6uRrB5MgTghj4d/6F2cCSNprdOj5/+wGw4l1n+sBOuMS0xkw
hy7S59sVyJz9TQOc7RGvPkc60xs9WWq4tpFoBOlXRVmBNCYWuOyZJgCEke00pWYtlVlk9WN733Cc
zYU6KRVSdvTDo50Ua6Lj7O8A2ZySTMScARAGMuEKTGXpqPKrodkzMsYdB+9V8R10ZrqXUWvvLdB6
/2kfb6yQbjgbqasSCnVMelhGXxVWfsAOGT1QyjhjW9C8kT4HS1sC1hEefqtXA2fpLwY8Rue9c1C8
A8Mz4AyrM/t7FnNR1iy+SfymLPkm0VW9RqWS89HIpCRTIGp2GmJB8LvxhE4OSAyW9Tnldp730CrL
4kt9pCl3iLzZwvK0UHJNcQTqxQDw9ibrUwzjRxYmF77cSwap+k/ZVpvsE/bu/UPj7JebfBa/h5Yg
+OEI7PcQsdWI7Irh1MwZNmfJWKLoJyg9yrs9fwUbeeSbMl+5fkWpRqvtjlCvWdeptCbjR+9PQ40n
ilIKOfdHV6wYlx++FP5qkdGx0Hnpq71eJOcsU0sqyc4R2TFe/U4s+n12g6jpqYTgoRrl8lPkfNiQ
5VzprWJGZSwrzMdyiQIj7UUQSXAfEerGR+GpPwob+eRS2yGN/ybNx27Ql8odrB9KURQyS1gigsFP
jk7KTTwUPokZmqPTywi6RFrff8Xh/c3QppQh1LZovhkuqalkzKKgAuY1CML4dBk6BDKODSX+ovqH
aGNKUorzVumIsboxb5MYyxxlVtIwGwSSQZJUspjjh164lfVjPODMcOqdyqDLcCB63/dTnXCtg9Aa
Ue95LMcTF1RMyMikIcGhwf2cldPcC62NS+kDi2YOjDdXAqBKU9zV1BTpqNA3J4VEj88zoUe4QFSE
hr90Kvkp01GG8tdUil6qDxvAZRYce1qSm7UpGzSKmFpPSiUMWp52kJEg385XDXRnY0PU6qlEfEX2
L4hAYQEuIbWF4gT7GqjMaX4oiFpQ/OVlxmvOQ7nSnb6KzcXkdsDGPKfh5vxrIN/bxc0avETFHq0I
vzqrXMHsT0rFI76P+utTGRyuVOdM7kqgIeL7+6y2YHV3QPJBDBywdb5kITCa5RMUDfTJIWUlYjxR
IKad6pwj95EGeK45LPKl08+ovPdA7g4cU43o4cSwHbGzqAec2OyR23Dqv/h1PFnuXeGqRIdWbBuz
bhhtW1xDW8Hv/UY1PmZzsdGYylFr+YQRggzWaD863vFr3A6IAe0v92BlCoUyT2BaGcOLn23Xxji0
srLxOyAnBbqJ+UOeP3yz1XqNmytdmnECWrK3l9GPNJ4DoiOdiDO9xYB9Ou7r3nDu7vKnJHpTlfEi
AU6d3K79aV0b13F0oZCMdyzoDkLQrLRkkoI1rSZpklhE245anAgNvjbC35CAcp3BkVw9YvDo4VeJ
l0tXFSrJeE1nsB2ieJsHa9ge4Ktldc98u3vXUNP8IHYJ9Rm+L4XNIUdO/xgLET6oEhSQSP3CrGSa
fmdELL+pdjNFEPRtWxnlPTqGwdYIwO/f9ETljnYrrIIqao86OF29giU8eAyl58SPiTdy7XCWVyMJ
GEQY1GFszaN6sFa+UXlZ44tXrVNBAyRX0FAM0lP/J1SLmen44uUBU7d+cgdqhpEVEXO24wWeDF+5
JmjDsZ6Sr6umfIrO0IOWX80ayCJT/8tgmKxjEW0oJFoHO0evil9gYeAqVqBzSkrKpxN5gbYQuYhn
2boQqkNS3wTpYOG1ZAEM2SE9sIMGFIsvTOyWVTcOGrp9DpfSAfSuIenec63fSsNOvXIDF+WEu77T
C0TLozxCrxniYQTXCCd9AxHgiczgUnOjxqOavZKZxEsNOopQZxQuaDEahEIY9p1xOtZAyPmm3PzS
NuQphxmGBdvLA7zPsglxG/vI+S5dPKoCiWDbtKTYhTFE2I2dfxdzVfHdoTGfNUcREWBfrDLt8rBd
ge9NnJOuBKiHOB5Kgp0rwX7xQrLYGz+ENAQjwZaK7/MwN25yCJYUonCDko+SRCDGTLaMs4iOqfW9
goxnQzntOWN0uBhHCwWSTVYBGOoBTAa6xJwBIFf7SF3Ccym84FoB1igKRNkwIs3A3h7ejNKHpRYn
0BDvQcr7/GpF1vhXdRwUf/szW8pE4xch5e6kmCuzKzL9mMJQdhH1TQ6DTww8fBe2JR1rbiuDx1jm
jUzK7qebBzpQEASvnC+kAdpGBJf/x+z2MUsIbWLM7yLCRx4o/QxT7Y+QHWtg/FKbz2yNfKFg5jVC
4pJzWFKYqt1jnodKxRINT6sJnMxydrKABpocs71fMejQ0MDI4Xx1tGVj33dIeNNBDQO+wIsnrHgO
re2mdLrm8kfsmjVuvmbsYduoELCMBSIndJWnzrzWATD9cU0ki5FePETBawRLVEQY2iXgShbkdNzZ
lyUupLN1TW2Z/zHzOVKp5/HbiWHTFmpHwo2BRTKkKXPO6wRCuY2zzPEcb8Xfny3pxT9WlIZhhEtt
MPOn4+j6Rl2V7tXHUa67qs66BbzQAjWLjxRz3BAokDaPCvR6HafLQgOva+SPX0RB1tB6DXOj/Xtp
MS7PwExI0tP38+LpLacMbnTvbpEWzyced8Id/TzUFETpMBFsXPY+vC/yD6v+SpqF5ac46beNemEq
AL/K+DxMfyoK1UBrOIKjm2tJSAYDig4UJ9EaAtaqjV7ClPBwabQ2oVCJmrlOuZD76ikNq9wwku8A
GysrMmGVfy7jXhUUHr+2b+pVTk6mGcm9FHca6m+UGLBnpSet9tl5bBrA4adnW6AZCC2pRzGh7eMc
B2AkXrtm0fYlwyIZgeayvUXQdhlYiRwBfZzXlsiKAojTTLMa1q6zaoXxhmsF33N2lWXovIOaJQZF
kqy9FnWoZKifkvdRZeJ1XAuikLyHaN+QxvZsYlNR2shDYHX1AMpEUi1nlPZkze0mco5x/OWxGocL
1luME6wnyPRDuDVQck+PoXYkmvaJ+JNnlTLQGj4r3uTX3qvQw9Jh7FHrQn15DhaGBM/aZDqCHLNw
vIVZ4jEak5fBzMzTlxMJiElreFLWojfjPydl/7fAhVpryaQOyleXDi2v5Zm6MOgEwPqhBsaqfSXQ
F2Cxgl5HxLHdpEiI8VCXfAQNQ/eHbWvovh8K+EdDS/osAoi6s+on5jPfxLDJH9KFGyVH236VCcqU
hWcdOwzCUT69IYLpLorvOVZcW1GzoC7pHnavSkuEdbhgEV+px+3nacJqMlZHfD4q7bLaTkhAg+zt
Bnv0FTkOcGdcIm0IRc+/0kCA4JM/JLFCQNAQEBO4az2At3KVPQ+wK6ClsknY4T7TjVm7ybUItnCP
0YDKerSPoZp84tQKmHRpMZaJaVu0SYbwA9UTKRPYPmftLh3AyVAOu7guc/ew79QtqmclKUFhBbdQ
E5erEV7Ll8CVmXt53qQMnuVnMwJIOmw0rzngRgTeiN8dn2muFw9PlkP4Gf+OjggjkC2biBU+3MNO
Cw375i7q+Fgcmu/9HxpYxCXBFnoUoiBXO2Z7wxt/AzCcHCn2kU8ZeQUTuL2RMxazFl+kYyErVk/R
t2gOuBcE3oIMgfDOogyD5AU+UvGZcJqaIgO/Q1T8euUicP/dpnNGZ2yRAB0BnZ+Cj9G4pN6PIue3
Uu1MCGcKTm7Ph1ZlAAhB5Ohau1YxALRcDriiKYQ9/ZBPMztPsv48WrTPB3BpYwMeT8o82Wgej6Bq
CpLJPBa32l0cuyI4x1DCuovXXCn36WEljrUtVSv5Fj4cXAKOcx1bP2VQipvAvbLLmsrbTu9baLGq
Z9JTz8P7i1oZojZVQN/Ag7L4wha1hvUyZQE1Ma8Cy4oyxur5ygL8YeFLPrQjvDqiw8UZTIj6n5Fd
31qFLkSRDXTBvJm8OJWnQ9LlXxOT/ZfsHiE/pQKQV+SgS9K0AtEOLvS3rO8z21Fyp70eaCgaljJN
mTRhhSVBpWZU7e7SipdqhkLel5mty56X98mGKT4BElJDCiyMVQKbx23zy27eorDT9YYxPJFhTtIp
ytvTmu+//3Gbgb5S4vDeqZ1utKe7tR5YDVFVlbUaSeQL4ea3CYz5B+Hy/aoMJWjeRDL9yj+Zv3L3
NcX8+6eoNPMhnqP+Mp0AVYmFz0o0fNUZJDbZIs3NtLYUR+eifIboYhj8FbinkDPevLtfNamp6Dny
DydK9OR1UUrDnaJoHoAZEPHe3092ImwuPnZXJ7TdutkxfME2QxH2n6KNBOrZF9KBgM7tVShiYIFT
f2dtHOmqf2yq9y1fXK8Ny0wGOugxw6SqTxFhmqik/8d8eKK7HJce5stVaKqeYT9jOs5OW9VZGg1h
7aeAiOOsJ/OzK44IPAD3LyIPMq5HBRiXf4pIQ5XMw3FW6+qPe7n4HE/XTM2VIh0wHmanYNx4asWY
FHkOdMOSxHtkB/YsZNep8ctGmIo0WAl3IYgB5ej3a58cH4iumKa7UtFc1TY8HO7Zn52s6cjVetN2
YDuUaMzkazQcP34lH4+BoWIoWEl0TQfXOjEs6H1uruP+NIfMHa3e7RpqSgmyE2tCzvejeQbQ88Qu
rvBR7429X/JYWm5oCox5DpZrB5XnMSmGieWtgBdWTSkcKMQeKAA3dnMQSgvqqXLojaRuv9er3ftd
YNsHDrQNPtZPBc/VXV3oWhcgsG3p23RhR3mag/8itNUdbshMUOLZIfDpIz7h6eIF8dKYat6HVhrO
9ykt0KBFjoKemPXIt03VkWWhNQnXErlquGYQLAsPIg2FiViAZ8wzS1CME+i3akwvWCzikAfc9XMI
pKsxjd0CAMLAsxlMbVubOikLTYMb0qy8WJk7uwUUoX2/QHdvwEz3ZqHV7J4AVKzD8Yr8uBg8zicG
LO4n6BF6NtLP1Vk+W2hYo6g704uBFXqcBZUPdCG2WgH9UwQ+891NGvBOoK9HYDlw20LLK2TI6BQU
2jpYPpk6jfNZwDOnv/JWCrQBW475AnZxDQffLsof9bLNQjko7SNBqnRtdAFUilD7KjZ1fOovsNY+
020bP6Z7nkwDSPZGSWVErhJbpJPKQBGjdZKtA4l0u9hCjiMSus6OLv05S+tnHTkDOvP62ngIabXn
SUANbbmnm/pO5KUyhhJL/2lCxQ+bK8EG/pn79BKcVi9R4ed17HAsdzcKRFSOzR9w3/FyoZYYzTtO
t2wbB0xso/SylaGFu/+Za6WeVSfG4tshr7HZJX/7HfT4ya9AvT2AwRvVkM1+aJKpXBZnGxYsh6YX
AWOy80VFgDHCGYp6csLDteHvpgFsuQRCInu7x5aKW3rZ4fcFmrlf0oms7rKJNyve3YNVax7QVMFi
YKnvVOGEKrtOhNS9fzoe/pNGOvlPA0bpZE40/fzu5T2pGF50HKUqZX0SLm44l5hCJnGSoJCDt/IZ
8/dyNPw4PWetb7FRYK3lKUGXtqxQ3B/OafAYyQE/CpDBE7Jt4faRPNeT+vEr2QKin1PpZTKrhTm4
4mvfbjbVxotS4Ru8bFVDqx8u1WGzhbzuDTahTxIoGahMyP7kdY9Sx9msGaTBKs+i4APEIxeKW4st
V35PMJUfsC6zacQgOjlkwpcK1lhKV1rQj8YtzbY9A5B1w1U4B9umQiNlODDlT15ds9VM3JmZzkW1
s6tsTsiZZhNlWBx4Qjz7309xMX61CRird3ybYKCFoAMaz+kX/ecMyzG7g4CO6NaZvogrP3WD2HHL
/L7C8idsnU2qspTHmc1Gr0nWhtouMYlPSjD2v82+cKlNsZSno0dskC+hrDB59f5Be7TjikfQLssA
eLUfIVMxI/BE/DAd/rmFOzZBhBKsFDIS7uK4HSLpSv0/g4jFyBV+4awy7SlkTp3pul7lfuaGIzFh
3dcJEWCc/x1X/JF9zv44WqbKZRqCAEr7ZomrjuQ9kDtas7FeqhZhV56ItFBlLfKu/1cn18n2GuTA
OHYDANHNqp7Q8kJq0Hsqo9O/15HrEce1oKlPg6cftc4e9HWmG7rPC3ZVStq1LLcQ+EquO3guPVPS
RmFw/rCFg3T7Wa+x9MyfxDVwMLp4skYQ+Wh5kZLovKla5YLD3e349mRMUczMe1uRBRZ+ipF9+wmr
OUsopibRYQgcXWXd7J9J6KeioRTK7naKLtzdq28CU8KfvxcCU0GNlGRBQzxJcgCK3yE15GyaeSw/
dLkOxSIfw53MQaMteVMaeUFCRcx7AzRi1tvj89+AHcZ/YF0tilAFlALbFh8iQX9rSODq5F6pcQ8s
6VALa4z5Ka9FKshBQdnhW2IzA6zRAcCiyALgE5y/WizSDtYDg11pWnx7KzKMO1XB3Z0HVZD/Skhf
X4LFa8kvUTF0hwYe78oJGa3WT8j1cvvA6X+FIQYQ0A+Wb0M5fl0mPNhFVjX9/iRgpj9FzW5Na2wW
PjloSzeVk6N3ntEB4BX7OHWNhJsNrRq3M2z7NM6LEWfvkvbdquYU33laAJrZMxJDGkCaGmzzXbph
BmG1G9gBLa5VHKyFxrbaNLezcacbIgp5dIJan8R3iuCMu2+QBMNX8xHFIrQPDsk7nxvUDU7KaKdm
sTBWApvQ/YgoPdCJKZlGJZvKuBOUkkA0R8un4xCG2wVS8oyBvq/IcPO/RL3ynGsg2U/j2vixzfzW
cszOndWySHNl78rRLa8LvMG6ItA7TXHk+lWb3aG/SNXe5d8aqI9tQ1L2gnUSUfaoa72n4Nior9ID
kZOKCDJzmh1FlogIHUDg8kUz/Qy8i3mdW4a7cMheuzgA3R3KjPY5KddqGfDvjWrfQV4FJ9ZAFYgv
NtvU4f6yXEIQ6k95a2srHlRpcAnP26kFMO0Ysx/YaIvCU+woQRGqLrsnQ3J4gQOgvIzuaMpU+VRd
UMecKpy5IJX9DWJHtDOuv3GG1uZYkYh4hTSzHBqAPvi330T6UDqARA0iUgWVAs5Cq8/HEMDmnlBR
1z5mpYA6GtWlMhbRGGq+SGiuJroUU1toBfrC9Oty2RRgkaM18RpYY5nPQwreScFgdsYUWQx3zJI5
n2oHzeijugCRqsMJYBsffWgCH+g39L7RSrS/1aa9jKdckqSVKNp54taN7HOA4J3xQWupmyjQz2oh
C79Mh07Q/bio5SJJ99xoXHPlIJMLrDIT0viTKLUbkh/p8+LErGxiPirWu/0cytiFgRbz7rNPtIff
6/NzU/cQSkhvU2LyDjka44Pnodk/6buT1UzuuqHOpVw8qbT8Dir7tPqZaB2psRY6/94ZW2501IVD
bS1F8q15Fjx3J+7fkOahCHIj3tqyUDAY23wfDA4LvaL//Pc5Y5w7lAsJqw4p8ZSOLoIrPr/GHvXy
34H4nSWbBl0CqMF+ir1f33RyE85+A+qZAceu6eZMVAMbreF4O7Rwc2xS9/j+hiqh3Xwr+1NI4kFm
UNwftPa3xaNUjoPwDlrfcKoP8BB+FAhcvhL8vYUWt+cqLg1uKOV7g9ArEWNO5naTXPbMDM6vsGqB
w/ErddhD7vXcSzB4nwN+VH7ixtSECR7E/sXQY8Lwh55bickKLHAp5DK8hTwXL7uGDZv0VqlCD6AX
oF1re4K4AqPGGP6lVmkC44ldBZdM/Npskbj+G64/A5XH8Oh6IA+4p/pPLcuT0TKUpvVmmLNvig8y
RIQQ3sz6NDFCHL9YfiiY4dTMhVB2E6xJcDyLDYgMGVMf0pkueU3aK8u511sghcdkgpAssCoI4ECF
gJIiKNi1SwrIekf8kjzhPhKOqVkUgHQuatKbzjj0Hwhm0pJAjNLAmDv6uTQglcnxr0kPieq5LR8W
f3ECCy1YLuRVSmYQ+JHJVSdQvYyQRD/rv9LD7KjkM0HCS7a8kOCeOJzSITQTqjQFKcpaIAkFYozz
5T/rBD+hixLM/8NcDk09DM1phJT17QUkmOhYZsFEIqvp4FyZ/ndfM26mB6CfHHWwU9/hCShblrrf
BhXhkLGfmoOIp9Yd2jgx/+4a6AjnzO2WXPBpodRgc09lJdAIL+5fKdOPM+c+E5QXuHExhdFi4uSh
cohS7Zu5H0zWitUM/vEm2PlrcAfZBV/YIxNMhpwo/Iqud8cmESd+FcPywJuZ0q5SNVWvKhyE5VwG
+g96vDaSkl4ZMB0Pz9JXPoVHLGhVgu1ZRBFVmD0KXoPUnk+RxTccmSHJPbFDMQHlNBdoGW2Ec72V
uL47qOSrlnxBaemYKz7/T/fMuJIv4XP2LRjDVwD0EVbJhfAOoZoWHJekaebMOeXCNdwhbHY7dcvG
OyKiMwpFnkaLszLiKEmOfbDHgaaTiFBoQF4NLwcWwyxfiatsQ+xMU3Ng88DObFtzvnidMBpHnLAo
14USR3wREkUTKVssAnDEoGWz3k42oECIlekWMJxRQVmSMfr350JXZoHVwfeGcu4kU2ecTptYaN19
gJcw47WeHSvcBcvf8XbWr4pp0Um/aBnPpMpziFrgH1OPQIdeobqa6DKHLWV/bNiOBdvdSJ77GddO
cHgym9QgU356V+Blj94TfnYrnLVTrYgo+J5VqTh1K1Tg26zprZY7/OjwF+lpeIqC+68uz4WB0VaH
vdCoF24bVK0xDEt1vfCFDMgYmIstArX7XBJVziXwIrtf1PPNO3Xq4euRJtzWc+gz1VzO8yK3oXpQ
VedPVkl1geimVKrxG+QgPoWdIFIU1HbZiyjO+ZTqEUc89/mtfnJurLG5orZN8OfA6IxAyLnWXyEC
tem+AUDsCc0+EQT4vroGX8LYWeLppKFUy7ufpBqUgNA4if5F8L4LPIbWG5vMBs0hhYEHmIkAlO1Z
fBqJdGn2MO/sLGGaa3YRypBTL+RVB0myJfo8jToXmz/hOD/wlH5B7EeQcrC6rfZinMjUjLcIj/hl
mMQmCGtUTTYst8pEbIoFlUWAfACD0Y3xoUHNYyzPg3cCpJyFtM1z/nvIpLrPRKWcvpju730XMCeP
toIrVBbVoe9N4iJ++Sqr/SUF/it25n9ZWMLDSU3l5s22+Px3japt3sHEtoxjS99lmxc6wwv4weQr
hAkzv7tDtfGbuhQKGK5FGNX81ByAr5OB8+T2QCL9kdn8X4UWBInUFu0lQYWH469mwEhgM7WDU8IG
Yreb790bK2jk/Eie+YiE32R2kPr/sNWDLpD43+w+ya9DNUXCJqIGxJGB85H2vnxCgRIqzFadxztr
YgTEt5wAZ9xezonkfYpcCMQOEG+v+CB9kqdEBeFAyLEtNFo1f3BbCrMNJCKVSxaz5+I0oPW12dnr
VSeY31GTEBxoCQLnnXeZ5w933jaeuJrLzv+NfOyFcamw82K5RdGM+BkZWGiVyRfNg5tN3xjf7i2V
+2jWUBfZzyfkmiPR8yQF4KmlpyxVfAnku3zn2ea22HX9NtRil7q/qoKRklW5EDJHkm0HpZg0geW8
v6tI2mEZfwvcev6pZv0A6zAE1u3p9tbmnLCHTFy0BPCVANllXD3a53jqYMbgqBN9bb6zGvH1mVOm
TJ92isl1YsEmtH/RlwQyCp0H6CY84+GscuZfxGLelAosjsTCQm+9Wf8DVUlqTUQxOXpjih9iFPAe
Rs11OgymAc8HLU15c+AXtu43+LgtxblWaUQcUbQogyHJQHZ0e4UMKxtQTNT5yZIWQV79GyKec3KA
MDeO/MRT0whOJXeKMv1zzCW/OYOEV67/mScmedApKv92e/RmTby+ztMlSpiP8WKHbsjbwTaARdwg
lPUAzJ60khvoozU1VL8Q1Vf/Za+9NwSZmJ8zQB45ejUgmcGjxuedBu+rpI65Y9ar5hIi41TcygbU
sQ5MSj6qxPn82DPC6KzfBiHHMT0yXp81Pzoe7LNQ5YXk6AQV+nVGO9rph2AJJ0AJV3+3pamQp0Wz
xolOi9zTc36mnjcqVX9sbgJ5lCPLCHXobmx/NdyMcEJJi7BJ2+6bIPJR6q7mrJBANQp/OBQpeFVI
y0ZcX/txz3OnYH+U03iGSdkMSbsfhYGbXLPqU6DAL30OoozAbDmNCxzmH0opGkpzJjVr29h/7u/Y
khHJJFoAMCnRwJ29RNJ7vfjxsTQ4PPqyCDXlYpFo27YMi7ZyZT3oRBDRcSgOC1uSsNxE9InCJTL0
5kYXpxVDASPeU9uJmqO/q0EWZYFjXRprVKHEqvp69OgDTxf+DsRFDXZYpJvDCpcSCPF7bRDa2o+U
KcRPhKC50Gn52t+XwNCvbrgkOyj7Cic/8Sl8qFEKYe32Pg9v6fjKQKF8rwxya3rxko6sf3S+5q5M
JietufeM6SRw/dvZYyeZ8bimvhR6fsTW22GF0RfEn8JpedGuusZ3ZkmRveOsBc2lkHhPb70S62gH
qzdDy6DHd08KUeqFExCma/6tsco7o0qxgLN5PAotGxMqzdn7uOtXLHM8pAsWo2FduHDU30dHXlDW
/Fu5qqR3ZlNFtgwFkuT8YKUvgS9KuKpjo5WF3pUTOqThA3xVj3lM/uuxxepCn/kcL57bVIBnb9Gb
q6qbAW3G7io66j5DgPPDojpNKscrQIhZPj7WiU30pfOo7xrF+KHilUqT7I4mpOavYuBxGqh8KNQy
23YiufbEBRrSkY373ZvrUHFz2L1arwzSBdjWRI5KF/wtF8hAjmTzd4ILzEvcJgJ4ZTEfdfdIXqcB
Hf11uep+Dd7SWzfIckCc5ruOVzsYWBQjRehf/l9mBCC4YWJd9mh1hPmPTcfG+4nNNkM4X9VH+tng
q3/87CF1UOm4yGhLdgnNB6u8mkZniLPGwbWQFNyfuFq7CW3Z2piJ6Ib32CJ32FX37sjZ/YdSVpmZ
JbxO6AWAy5mzeUyEB48/Z7Id8zIQyF1CZQ5MQrx0S8nyb//M1NuwR6vhd/T7Wt5x8JTFZGy32QSJ
FmnyWeKCpssJiMoCxUb8LAA/ApFAgwiCWM7qhrRXkV1/CaRsH7X+VEHOUScC7gAQC6E/OnvPWdhT
U00o5WmqyQ9vMpEgFwz8bW7QLslQTDH0cz10kCEpmbdLFuQkIp+BAooWBQN/kSBJO1+Bj9qaXjJ0
8lbLcwWTd1MyVm1HcR48w1V9MtSnkHYTK2woUHNvgKo7WZm2lNGeRV3y/yhjHCWYINsSAuuHpR0h
mMEemKXMMi6mZOY51RQ8KRWLTuILeesUE6tw7l0jVWldSzTgDlZLmhNVkQlcCdzEe2887Bvz1cgf
HtHTV5Jqrvx8MDZQlq9pXRuz0eSwyYYanYU5CeG4RpSdb3NOJdbJJeXTEsl/wUK69/ehwwqsv7I1
MSzgx5Q3rGJuJFcCKg8yPE106U8SnuntHvu9pv/JlvNWm77hxe7vRQBJc3HVvPIdoi8b/B6tnZpX
rGHoPMR7ztVBQ2hcTESgB7YisfCDbd69+yb3F0f2vPiE/KqIsthsmdRZzJsqJo4IC3kBNNvCf4do
xlPBQw49ctLnRLhlyz7sMdfrlEBK+K8yehaeE0DlVTDAai+gGByTMQtZR80+4IU140lXR2jT1kL4
bWXeCHSeW8D7w+LVdGUWgTFBSvcw9sX11duYhS1BAIh/yTXTsNHOjjFlKmwjvde2azvl6DWLr9rn
teqNpiO1RcL/roghrQLaJIhRBusHhPu1HohZKlcz/Bf6uNuNepED5mfma+2oDWKWLJAiRdU7l7iz
z1C/w547DIxHXhV2+ATq28xPjZUpkeSv/BAfxJLCu86JR7xQZ2Zq4MXM6WVueFkeOe8D7w4GpRKo
2JMjxNb+rQtd2nA5QpYb0VD5ejSv2AbQUU/wMEWJWPB/ReiDVu4cpQvYEn5FlmniTd4qz57PI4y1
YZXxvI/1XvjaE81KIHsu4uYAh6YfCRRIhNpoCegaxvDqnaYN6g8j89y/LnAoBNTOaOKMaFStoyOz
E+VXn4IR8xH7EPPyvxmvCZb9MUCsU3zJUNZLbrE8WgAkeaMMj8k891cptG9dDJNPuXihuWbRg/Az
85OhAxgmPnuW8YivS/xOwbRqwq2IH5hyt+Hj007uOJ03wh0QjUwgdNVf15U2eitoQ8Tnl1Q5ZVdr
DwC4mKEcsevWLR9SOr0cdCseAPpv4Nd8Q2xH+oBAsSoGIvUrvmBsx3RxzeisVYHfQHCphi0d0whP
Z5XWDFcnZykWPJn/gp+bsAOCPNB4WGE/E1OuuaPZ1pW2Oj5P1Yuuqh3Q9vsb4LiapgJeiKI1vCeA
I9McJ+IM5fbYxMhONPUyS68BXkOVvVD1EmcQ0trJ9rAckxi/Y+UvKir12Qk2LR5EfhyhQvabAi9V
hesyxCcPGL1oNA9CzuSgJpSvDAo+UUMDXHJE1ln7kJl/Ic0IdtWlDiFmZfOD1y3vR4emJyb1LxIV
RhpeOQpBl9hMbulGcHUoGebtQPQdx3WFzO3dM+J6GjLLNn5T8OnrG+wVSTJAiNgxplH1l4+hWD+Q
4kimCgvHpdj9q0YGpPGZqIapJHQBihl8UiaB6fVAswGsoCpRnp119dnyQ663EhkmEcf60X4OKraT
9RaGjk9VZSyU7XZ71J+DbyLf/8kJLD4FCTrQY1oU60tZ5l+EwJED7Sgn6pisMzhxlVac7GALuT18
FX5ijU5q0jWOq4XXPHphZwj2GI5YLRhe6NNncqiMW4tJH2ij0xTdstUh0i0AJnPr7cxx0d8+VqXe
uyVprczqUGdSto5SjWBzL2QD6qg5LM33sq3V8lxtWqLKaRyZFctn5S8VscJADbl2JtqVSFOb/93N
d0qBkrfzZlTuOV01Ele5iHt02asNx1oOBqKZAyqhQRmXCsp8+6CFYehu0h7ZHYnMbwb84VB4Rhu5
/UdP4sZBT0bPkeYR8AQ85HcMZ/B0VgFqODVrCsDn7z0tXJEHj8fPZkez/lWqKNT9ylr2ELugirbZ
vIgqZqEQepaC8W6hGREOTFNHYHPszS2wSMpR/nMeM389vhjnhDQtb4TiNwFeaJm/JXxubrHvcbc9
c2b09XU+GoTPz7bRz/0kyPyyzbJY5miqbtquL5DPEovJDSmVSX7UGJrYx5e3bjLoskmWpn7Ppatq
XpwZSymZGdajLrzoR2BrFUIaMMDN4j+nazQpAYdV/guUiZ/H1GlXoiVScpKE7quGS1fpwoqY9xy+
KUiggnVzjbq7TdRd30Krx9zORqIH3aKdu/OzdFGEgM2udDwbUJaycPG19Cfl2o0dUBD08LfkYKh5
1VA9IYBHSwBc1IPIQL5Jbp9u6OaWG/aXJ+OhBFfiSylfgVdww6I24f6dS4Gap7KW15hfNYAapf6p
qzEDnw0FFbMEm915Ut0SkU4pwsA8tTbgizvUDceayknvYPIgrdUzHGPH2f2VOE26LOxI/ky2+WS7
z1hQxCDFgWUCHt9xjBD0GCRAcfXcbAILUTJrnf1vZOKTT1+yy+soi+VmIG+B3T+QoMTfXjK4vT/o
c3g0q6ASoLk9sa3NYNp6qZO5S03JJnr0dt2tMSFAc2HwHWFZGNCS1Caq34jH+d77OB1kVRlgAsq1
BtOCrj0AmEYDZESJfNt0VLpua/guwWYoknB/0AiNM0BREa5R8ZfiTsMAIEA35zrwFJk0FOtK+IVu
IUBo7/ovIVy0jtFL47NM80DoYGPgUQ27QdGHt2UreaRCnOlN97p6RMKkkvIXo+BwZT4Ut6SMw9DW
fNnMZ6xjNl1RWGZPYbSHGNJAVXSNqk/0d4YeBt96fRGzTPHjNwqPXyuVDuMqtsG+Q+Y1P7nGdZ7V
o2GPR9uGT2DCou+hFIvZGBvfyCjmcqJOUE776A7jIHeMVtyrcFKgK/JoM8TBCZoiOxYb0sayE3Q+
t5WNxAmf9BZ8JlzSkDsB4RA3H/zGaxUvm/cX7f0T8Gs883+iGrW73VxYkcgP1XjcgJ9q7+sPRD4k
Z4mOh39jIzvMoyb4+1FCjLBvE0eGkIZSANpkWx/caNwpp/xPmBOG5WTm/G39r/jmZ5aFOTnEDL/T
rjGexHcylLJdUM0pwE2emrFHcwMnMyFMbDeC9osLfFCbUlei2R9M5hvlumHN76KiPqHohCZQSqWL
lG+Ausw7W2oOsK7NXBrRu5w65F/fSjrkIn1sZW8Lh2wykcFxTjQOtPv8ZvfzhuYnbpTI1PrJuoLi
KhfPjzyH8knqE+Z0+fPTA/oz+eMl549t5Bg4MqFO50Ml0gh6oXH5nSLlL9lq5ZQUJh6fwhx6VtWT
i9Iz5OFkakkbZ6Hs8qjbYKJ7uwG1Ur5S8JBqYVXfSFUm+e5x0ZH3mraCtrdHMb3AdkEFOXIkBsE5
L5ZQ3sK/HjAxLzuqx7NiGH4Y43A/mto+LQI3DwmXsY8O4DthqTk8b/B9ZkN/Vu9kEHhrRFXNcn4r
OaIjNifPxdSfOivtlXnYaszkfqWICkJMRdIaUWyWGoew3jT/EVOkunaip79gaSG/JfKufdo/sRSU
7DDapOJiKBbsRSz7vXmeWbw6OIPtua/gitEQc5AaCRQ4PFkpmzkUkVUIyiJoeYYvMhEJ1QGZNHTi
TRRCBx2Zoeazum54K71Rjf4Ff1NJ508A5ci+qle6B8aeVDidsPKMUlHYl8g6yoPuw3eUHVNM4pAg
HdEXFZ0Q7WcAdRuN2MR/CqksyPqhXwzHYmlslOXaNTsPYUCIlk0zvjs2i4jkdDM5HX2xsIjTKWFs
FOTFhNk/Q/fpSqyfVbxomjE/wIECkmRzbNhFahstKucVBCXxxfPdiQoZdd4JgYWyxmGs14w4AIqu
8YJRv05Ch8zH61B1b44Z+BjPeim0AIFoswMYnYMH2cRHWeClK+39Tl2giRsrCfoMXwRf+dM2FYig
Vbx/79+9Hqcqhzsc5l1d8qPrBBhLpF+4rMb0z0TGOra0rXsJfiKtUavvSWapImJIVprBL96eVTy+
pm1/c7SvkYr4unAUDI1O3EVKUyaUi3nMrxpqJFg+rg99y4oMgeAnXq0aWFex/XB91oQZUCMSsUQV
D5Jb0eFvV56AtTfUAB88WXoOA9iCx/s8yD10ug6DvMIzs+UpVf7PAwNlInjJXUf1w3J5O4wmMl10
wbaskGtwK27ic5aLS/QbsJtHWpAZo7gDqgKBeF5HwbdJ1yPQQ48YZ6UDRkx/KHS/h9T3MIHdfb+A
kG5uIgyJYrGAT1c9wusdwOB49I8vYqhGX1fS9Yv2vKYwgrwaZ8MqESrYtmmr5Ptm1dKnyx20um3x
k1B0uVRuwYOELm0Y6rN4UvLIuCKpyUIn43FhLd6c8z7Wn+2im4jIGwhr+ik7fF4+r9K0jenKwaib
OZsAT1j07yh1hG98L2szGnDJSXuIDDQyNBArQjZhkqPD/6VktiCZyAl6WI4vNR6QsQMI3GhHz04H
OvoagnjkZt7xyoZprZbfXbsvq1JOymKNPrYikbW6JsnUHcedtEIRaMcmLp5GOdcHFfWwL1c5ejkv
qzzYMn9L40cbf09MKpLfjRfBSME9BHZfoOG4yijDaYBNnufzwigzlD1FdUHHKXkwn/+LDLq6eDr9
Uj8s7D+52SkOAjSYZcBoRJIc4UIdzCU+111VrQba2iSNmT1JiToG2oPQfF6ZKvVwuxwjqKWqdoFV
pBnWEKZLECfwqEDrlYXqmpVpTSb1eUmyregoiImdG7AHoFapAYFmz01ptt5dTdp49OUh2MGjcGFs
QaBPdotvEgOa3uBRoW9gNAV6VNIjz5TCVTY/nTK/MnOlfxZvCa0CrasfkfxrvKJa2fwi5V4Hbqc9
Ga2wiuu3L1uEjwOrpETCgcI0jq5Tt+plAPhlPjkmEzNfyY9mNDUvU7SE3d98FoqGmEvVVdsXe2HW
vxfqrl1//bQL4pTSsmYqp9Yqu1LVMvnahcphSVQDfaSRGYtRMpmQhf0xUbZorZJzlz5uZQV67bP0
JoGYhhyGjfMkJPQTKdDrSce/dFqO13quBkGGe0rZC9FPPumJTqPQPPmy1CC9KjOAr7HDjOp4tNp0
m44reqecN74vJMhsqJYnpnMrHoOR7aewv9yo8ywBt7beU61CK9AP3/fUJB7J1BnP2zAuxrPoROs9
tBYFx+zmvIsHwWuuG2htVB6fGweWEkIPPCSy6bzl4bzOUfJcqftVrSdMdlqLSVJjuKDMr/Zbi9/H
N/m+46bKLwaqqI06gA9gKtJwgC8vlij/u+Wg/Qb85R4040HjZFDkHQZ9Ic0A4RS2AOsqi+sTbeRO
oV8p3WjbiTa3EHxnL2mOhAt2YEGOqEoYRzULe7R0V0aM63Bb/NgM+ndrL5XW7D+m4CDJBfByvSae
0M9/BfPywNKAz0lkAFbEJLOwS2joaCspZM/W4ooFLYfU5/J4jnBipPJRHB9RGq4Vtxk5/Cuadhm1
+7nbS/AnWLJ5pFYyxQyTPE+r+ViOMwqfGlOql66jCChd5rvOp9vPU9FQu7FsJV7EJnAOvQhTlStZ
Gyki0bTZ47Adt8AJMhtdsksIBnMJPZLFIdPCNLK6W5pbuKpt4m2Gs9bDDTQX+gu1Nl5HkKSkcmaL
vW1tVyJoTgDfRbETnuq0NtrXPWa8ByHP2vqdS9V3zzZWK6HIaW/ff2EN7aaSrKzJHZ57r8Wsc7Mq
UaB6+BbiPPkkUuBbVvHOyCC4QbORs12y+UZCYnAbgWEMRw3HCOFU9eZqLF2S1s47SRXq2GHdyx7r
1/h8zioVRU8u2O+oQowp2QXE14VcEbmtLqTOzUAY8FNC7h+7FjgBalvgrq3ESUhMTXiMhvvOguX5
JtNHKjRg4eCDh63FXrHNFae5ypfUat1/7Yv4q80DDOxDkR7cqecUoTL04eTiUc6Ucttmkef9gmIr
xii01XNc9C7YnVTxsgzQ6df+X768cSKDg8nDK2sx4nhTpGDFUF3WIDuNsDRTYrYNeFx+AK9ycU5Y
uSjGmUL1mu6kTq6EWTnCLo5MV0xh4AIEafmGL9jXX+fOxtSpvzTxUHA8Nl6vIm7MS5haSC3fubGU
FQdi3pROJN8Biae6HBLfZK46YA5PohmyjpwwZ+h5ZKQMaU2DPtm/36UqAP6jYucXhbkL7mV1o1hE
rWPKr34XCwpOgIEzdpj+AiINQqwuBcwvQCNxNSjCG7z86sbMrxVJbQ3MUzmT9/bGoVhDaduXot/d
1+SsGO4eg7wqHOicsLrMJcTTUzUTNYPeurZLRvJOVaIYoWhYP4RvENOGbqgsJjpNDtuQD8iCI6xU
JkujtD7aFM71BGqekH7gLSenBY/yS0JwhFxNWXJvdITExuEBJDPkVyw2+bZVcIW263RXBQ2/KfYA
jFb+T9wHyHSR4O01HxGCozerendChAEtqeiIYC7R5jd/O9a/FoUBqn6AxkHo4s8qn6JYBN9Bwgve
UCYPH5JSZR00CHbnrc4N+OLGlppLjhRm3l0kM4CfhAi1AezccsiF8Rwo+pGsYKGLM3wawzCg7vlY
Wyp1xu8y4RWNw6Ug1bQAnIuliuYoYe8QrdegU/ge/FQfXKo5ZiVI1YKGVHbR+IXGdBKWwMgmrh9t
PgFTb9MV3o/ktpyFlpHZJJeTql8hIVZc4lUNYOhuaj9InLfB4mO5j9eoZ1QEl6260WyLgpE5MO2T
//dgNcX8uNmndeDrXhZaaF8BGDSTKpUjPxWUMR4aainWJQ1CG3xTxCt37VPq7jCHKI/DLe14jg0m
Tzmet9wHhTvHTU69K5Git/AeSxTaHKi19+O5CHTbBrHvM6QMtQTNLNMBqR0VfzgWyC2+Fb+he0dY
68/mdiUtZhZpWoEYRg6Abjs6D6J9xQfkwiUzhOa3pK48ecBp9xhjal6uIxAnMA+ND2HDGNSDXKrZ
dmdfcLRFuQhe1JzNAhRRVvrrdGN/XYlRgsyCEuJjFbjsKZ5Vd3pUcI05I0k3x6EiBohsNZMRuoz9
0eXIS1/oMSBfUm3yDtZZOhDN1x0nRX0AerDwH78qzTmwJisSYuf52UHgCx6kaJ/HmwtlkswgGl4l
E05Nx/q6r5ZCK9Cm/JACUGp9Y7on6zXKgVdJvztDUHiaonRmWxrkSAHaoR5WJGApujbuomYqxPD4
cyrDXwotSm7bhxHm22v3K5S0LwKNoArgvH7lZNbXBhDZDVMjG1LlATOUXd8+jsJqdNZmVm3EhCuG
+BW68ScdRzan15eHoEJ6P9JoRwa4+PX/3K43x+nQeVctIE56jHGOxfW+ueBZ8vMl45+JdegLpMUe
tW7JAKA2IpnnFA3e6UXMvaBLTPWrYyRcFM9DQHa0aEa7zk+z8bDw0uQjLMPIioe/zunCM5JNKxLN
T+VdiKLj/+PfbcZ5hVgdZN+T5uAOJvSWW9Qg1r+NMORGRA+EWk+x0c/E6RomqA+NSl3qp89OGh7W
ZHOP3D9Y4tz9X9oq87vsLmxx3aHPH6int7FdDcQZ/F2+8VKIxp23BYASCGtlEa0GzBTyOvjSe7Ya
ztVkYxpfJi5U5SzVUK7wEIh8lB77ZPueNMUi+Kuvn3tl1HJuDxALXAXwHMxfeXcXJaoRYI+5KhFt
ALvxpczZ4gRTsDxeYlvuzptG4rSDeWadFm6yCNrLSdMtavFTyejx++oAlzI1S1e4d6MXCfll5nuB
Dk+eJ5X6tqODOVAUWwQvp4qGA+k354O7uPj9CcGnMIurzTNmCLy7OFngMD+dVwpt0e/Hz19GBvSk
cPYxXzfl1oQlcssHxSulNe3cfjP++DBalAZy1EHok5SPOVAkTZtsKK2+bB5UWXasS/DTsKhDeGsY
qfGPvXks8rBw3/VQeHcCYTQV4Br8meYKr3xhmS4PuLxYV58aVnt+YCHlJ7A2me6kVV7d8QUBQpqG
HxCR3a21X0wNI1CLV6ybb9rTyvtX45tmPGDAL0YSUdpqj7I6mYXAiCB26SEdv25UQmqzTTwKf3mL
1NnMCb0tWQLprwZdsRKRVggx55pisx/AKoqyoifIkB+105pTYu3G3N9KWcd+X4EDeAChyi9e85M0
IOnRadR+ZrWMcRK30fS0W+Gxb+W5+InBjGdhm/nN+mzBA2XWVgLq6kSsYt0HIltV5Bfl0PvXtnkM
A6Yso8cm6VhejVHjIvSetfb0BwdDlI9iK4RECVxLnSJNhpxPk0fccF/G3JdH9C+KvNF1pUw94fLL
+0gAzkrNUUVwHF6h9+pc3HT8gHqXXj+2FDRE9VFxOdvYAqDFdMRSgJjnTkYfhra1wWr+UD6glies
1uk/3NbB05m/0Ibr3PofqauNJjKcyI97zhX0WEvJXqv+j2k+BuLH7TD+EHvLWYYYlkmPH/pU4yGY
6eQQMhmsoBt1DCmjUlakrYTmpph2nLRrGB1PSvVn/nCaKi93o/t6d+2yFuksy084BzW0tu49IHG0
OEVb4CbdRD/wKICYbo0ZdVCBQ4yVXaXo+ylP4dB6mF5KG5gGqZsQVphHPfktwmQ9gGzrN9po985Z
/i4cQaNxB7Wyjmagv0mZVi58vNYqnYgpF3R3lga7LIhkWjB3PMz8R/TFC0IPp0B0XuqeMrE2phcn
ij4Y5llNnxYXWIeQrYHqRZJEDdBz2gcms2gAFMBj5LQrGpZXWAnn96gUZffRopxh00rRoOoGnzMY
bf8Yome4mYLzCI59jXGMGhCjBJxaeLbnklcqNptiJnkhxCXnFiprLhCNqgRc3H6+CIOUd2gsDJWW
arw1DJPqXTF+0xuNMxO2WLstK8Fl6IyxaE+JO1p9Y63GPPy/eM8Ls6mtLaZ/p+Yw64/cC77P0Z6A
2o0yeF38oA/TXOvKGxIHTEk8jXwVcyckAfybgveClFwB9aQiyi6D3EAkbMC2o9Gjpngcv/V9WGk0
2wqru/qq+PjcBqksXtss4EUowq/Ce5EZlJSa6i885t+P4/HkxEnBu2cz6lOAbj4RSOPfeSjtTvSx
dnq3anRVavCVJ+0JT0BQMZSFZc5a0lP4lwHKx3+k+wnGWixW8dbZCQyysMbinzOj945uePf+XyJ4
1HIJQa+DwgO6gfmBecs0/s5nnkQ2+W9Wf/8G8VCM72bQAY8VyF4Twer8XXwjpeQctRdjfTC76mzi
PlbiZ6caFQjqAT0aO5OQWbspQlySMseRpi7DqqQsaz4X1Hyyyrl6pS8xti3erHOefiK52+8AQwea
Lee6PZJ1esgVdRz5S0Uz/BqfxWq5fsZ/jqCHhYHNMFRd36qzjX+IhfODLy+ijf3JT1nfxArPYuW+
r8x/+PBk9uikXqy1cwqVqAckjP9nsXVP1BLPawq3UbNVbJsiQbC2acOLs6WwILoQiOeMiiWoOivA
nQa/07EOeZ3vDFfdxpMnC/5PbRsT8co05Ir5yCjxG6aGLsrYctAPxF0a7E8PUgWM6NPBz44NJWAH
4yNz19b0TYokLo+Luyh818T8B6Bs4CweOc7iKcZzjKJsesuf5QyUIWHMRMvw9ECUNUc3oM7bCn7S
EkyGdmErIFZhmjORbcchQyyU0fmKv6iBUa5D24Nkll1nlY7CsluG1nHXRAfNnXEtmuf6ED6qnCLM
Gb6KPGH3ddljAa5W4NKe3FaGgZi8ThxKCqKElKN4kMg0oGrhRd/zJeCq4zppzC06RjY8yDDleptC
MgJb/m5oadY7SspK7ZphVSDvjDv1jy1tViQnVCQLHsJMkIYQdvhPvs11s7ifL7IWHCVENcwBoPFp
TKGC/mCorAoUqlMQfrKMUCwxCDT9vY9mhPBeqyJeBaW+4M9IHnzaVThz8Dtwqlzke+G4fGDnDRre
Bx8iFc48zAB4GQairsp6cBFOLalzDyH629M7FEM70dtj+QWjHbF+2MoBJhsOkVrc/9x0Gp+87nLv
hndG4G9GPLyYZTsSjdWqq5l5ezhJHI1gpXC9+/1h2/N/i7Fst4/QF3A7TsIfU2UN8HhvGcsdbSFT
mzCJ5XIXd50LI8i6jxpHVKWdnDwctj88TTtdHlR3+mw3dLvtsty87FAwVVz2NyTi74kii4jzcMG8
bkzxKDfyPsW6KIHP/JMAIwZy3JhyO3Ss4PRN7ZNcLgD2+ThP64XJxHC37/4EgS0UW9tZOvlUKMj1
Wfz6kt98SftJW5R4VVsB3eZ1H/QmjYtPR3RjVoE83r/20koFprVElL9ZLxx6cylPSWkE8H1ysAEO
/9MIS3OVUrb+yEnIXGD5GAb4fDX6lIPRCBYbja0h19Q94MnKlTantYd/tN2W9SfKMolqiNUCJ0Ur
QMzNf+MYH95zkWh2JUo0wlTdXwKJaHoYjEl9TtwLTbYatSw1jwjjUGGu9hhNsZdb0Etvo7RqoRBt
v8fHHHv0wloj1QE+6W4KOrg/NRUOHcjh9rJtBb60Rv6gSGGpgG2tlch/Dudk+SAx8lRPbseMOBzr
79ker+WbAu7QJ7p2Xe9Lec82HFm8+76YmbuRkoxdNY4wdB2TmMu2mzDmeJNbRRiyfznIyg4rIA5T
C+gVzaIUjQOWkCUCzq6Tp9GE+gS6OXMcvE8zpNA7cD6lIIkl5vKDyf/uLYrQTrMjMwALyaXiEn8K
56PhE/g8eE8e3nY3Nkp4Jcg3jzJ9QjkQS318bhshdFV+kGvbLw5gcgVSNnVJJND/WQQzzA0XssX+
oFf3enDzjOgpkp9QsMP2nvc5yt0b8eWP6gvzTpuNj0hQC7Wu47b4iDbdcuThmahUinLwMcUOq63P
dxuXOxmh44iV5IccuEZQc2GHI4BJGV0CT/U4IKhpEVRMmlBVvGjEJOGk7ZCKzjGXzH5S1Zb2D9S/
n+3bSsBw9ZokPb5ivu6lsQyox2PbXK3EGLoKgkRzNR/LVq+FXoyCNLglx7F+C2JUuGcqmRD3NW0p
hvc2FHB4Dj3Y+J4DJbQfpChE6TYy+/MFj29pX4DAt4K/zdWO2Aps6CcO199kEAGNtXGalMhP/Wjl
ENbIMd29KfmKkf7uArTJcbwJE/+zUri6kcv11HdJGRyVowx3Mmu4LiFTC6jNaTX4qQxkO2f0ocsl
haO8uQAgp9tjJqOu/LgI5n0v8DxftzzhXsuA6cOsyHOm7mb3+8Ovl0ezO8v89o71MuWbpJUDFgeI
/QuhgDqY3fWOouEO8AoxgVEwY4Byi8uYRPmN5hG3U9uOaH1SwSYRABkQM9prHFSNSgwDIjjWGWai
/BX8UeO/K79b/9om4wxmnprd+TEVmEMlYlbvO6MAwjC0Iif+KBTYqglypQmAy4GxBgwzvqkJAb26
MmNN67jlwR8IHCa4fZrZgLWrPfI7PeMasR+OdDi5gFcpKMM4AY/IA1Ah3Q7bTehA6jiZFWJmp726
qzu+UfP3VcIrtURNgo3xF0/gqAG/Y2RwCbR7pFtXHucZBY5tO0cWtynIgtKObAl0bg3cR/hvVFlZ
ENa8mhQY3SQyT9Elj7Bkmpo3j8r7ATIK/ZIf/ZKI0hh6BpfRHlCw88umQ1Qxkmcp0dRlERUUSO9A
7GALeceQqDCtgY9mj9as2XXn2p4gPjqgJxEBy3Ed7mHE00H3WOU2HV9HIj/cA1oUcqDfaij0gaTn
hg4QsgsRAuFTZWvDyw3Pi4LKudA8eFD0gqpmTY/zbHVdj48jO5UEEYF6Y9UfLtBFSSRvR0UgGTYw
QfaRJPAz9aaL/1zICWqloBsuagPBEty4L2H81mQvXCva1FV3DTqdJOiwqNli2HI1MGyxlktlaenn
D8aNwgtkE2vEoCQpO8yUHyUvfItEA8tzxlSQUM44BhepT1i/as26dMdosq2Z2EnzRDDl9hHgBxZX
PSihnPUSOtlnKUJo5dni+vXNb2qOHfeUXIdyVC8GQ7k+TGFxvzFNEi4bFVe9+mPwtUL5r7+7Cf1O
HkLAij1u53eR3YvB/YqogPk0e6ye6/S0xP9GxKV6FLUAlY0DDRHr+4gvQ1Kr46oqamMyH4Pr/0P5
Z5K6LPwSRth88dJI1osZGIvthphZ+g3o7/XpanBMuwPwWhtt5Qtw6RvRzM0+YB0BQ+KknuEnKk5v
0DX6AnRsdqQbEHcFpLUUBfeF7tgPUObVPWJQ79SivwMTgVwZtEmuwV8yK3yoeByz7ZG8jDkl+WAq
aMcNRZOhsnvldw/ADeIkvT56DSVNIcptwPHdmawN+DObg6uT9rtkuuEZ2hjXmMjARN+ErNJ8HJ8h
i9bUIlfr306sAeWJqTuqZ/yrM/OT62VtKvRWBZIlqFBxx+LzDD5jYAJp2B961SQOQSiKJT8PbLfc
ulcU9zQJROy1SdW5rw2S3ZknzpIyiJzdPdg/aINdk9W44pBwbXvgzkAspj0GHt0k2R1/An0Ki2Xt
fcAC1jB+AFd77asuKsitnJfQtaR/eKLwVDmgSkeezlQAsHVR6fu352jJ9MxNMw78lRJAh2Y+0gKn
9L1wqlJpTn1YWHLrnVZ777Oe/xBBlMdMcAFKcWWeYfh/74iC+4PhaCCMA26blJM4bYzJcdxUpsoU
xccO0p1avIMxIAAYixNrtrWqxtS0b0QTDdu3yKFQeaUWN82Kz9NSXYwmZWkx6zYxoHUjUiSuU8PX
wiD9+kXiql+nfHbtYopzXN2Xlquk/pj267vbFyC03050i1uU37Y4CmcSTDRoQTugJTnuI6Sko8Cv
yHXSjCgHTwRPl5KJVeKvIuDtAfAk4qwb5hOoB6L3YrQgnxIbb+5ZO944ExJ2Vg2OvcnlarenNCoV
MVNDkgof7Pejfsy6RM3XUZ5Vdtgsk4t/HqmQMaQHE/30SIiBSN3soCFaiBPgg7hPscXFf+Bwq8ME
20mMbGp3uaktfdU5AjyyTUnjQEEnYEhEHBjV4Gn40MLconRgAsDPeg7KuGRy9DJjRFKi07ReXhzL
K8EWA5lwo9mH5qqKMrIQl+plK6nA6LmrHld8bopCtwNPoEbYXRwXklyn7CaW44qEf2OJbWjblXqC
uaJ2Yzs+y1D6tDI1UrnTgDezcHi96r7UdwD7wX/1mTORqEbW6XVobHXFarrrpNKCvX0JtnkYxzEa
jHH9Eha4obg2/W6MU97ipqskb/lTJxolrr/w30LS88fQT2Vw76uGmmBOPxG9j2GLo/JSJj0ZdKuc
R8BFVWGlLrhk21sti0CL0PkwUDlC5WoKNKdbhcTsd8DHplO2PA4BN/y4nHE9gfnAi6otHHVKQuk3
WIT0Hvsvdi8LkBdEuXa3XTkeyog20Az78jXprh2JU80/3XWVv96LzDIGxHVkyNei/HnT3rwjJid4
MM3hGstCZSsU7G1Z1wjvY2gDvMNLpgg1rOCQZb1C+RmcXE2S8vmRswUuOAa5nmns93iLWWVHhCtz
NrPyRrukKEjkCfMwxbsnTu88yVJbhfYNqq30rv6wX7in+I2MvRomdTk56RD/Db76o5xm+ZpOkMxA
DjIKWaGdexc0o+18uTTfmFCiJjO/7pMuIKS+S+8RE8apxoWOBwJpiTTAo3RuG0mpOibYyUPgnesz
oi3+nqA8U6MESlsHyMGxoNimdTzXhGWzFO0iJsFvsc14AhF/GGBEOn1+Wt7GrAEY71sUKUnvRjKl
DRFf5UVCOXHFx5Q9wWo0IJHCqCJprfu5bjG0ov7cyUBF2GApe2hHrguNIldMLYAsls/DNi4fMyvl
GLFdkmz3PjL44WxsSq+IrJ5mmwvIiV54vaDA/nw6b71Mv/HdwUuR7fiAkVcLy+Mb1FT5iX4LuTBh
UIUmL1bAum5BwPSdSVq27W8yE6Cz3jnExMqKWOqnxLMdbS7eFc9TDU32LMHrm5gQUO3p+eCJHjv5
N5o5eUTb/L9kEFXiXbSxSq3JeqZu5MxzP5RUVwQ/jhyfc0E0EIk7RTzIO3nA7f/VNF2Sk6zNPgzm
IyF4brUkGetWo4Sbk9ZUP/DANLpwx4qzst7HTQdBfhVJpQQahK+WnP38RHoh2smRT9X1XCXuWk5h
QZELJtXefzeefBXjrENvJSe5ce+y2/PCBU43CNU/LDZZXSO6DwZRorSj1eJ+epctp2yzP7SCoM+I
x2tVSqewRoemvn4ezanHZ+1rcWctFx0Aqg7BfwfopN/8iw8WLsrv1/9ufTdASvjJwG/6c+ROJkgL
Js6B8ltAmIW8crjlhQklT88dHtdDRtXCQ7vfjUQZQHcWOVBAy7B3hfzY2dbGGqUSzM0Fz9+x9Caf
SMtqw2LTmxx2hs9gLLVMdWkpmlEkoGFMWeQzip1KiorSJgrClVlQ5CJii48WE735HvafkZpLCYf4
5oUjJRrMgVOVrJ3ghEXM1/o4sYdoKHbaD4P3POpmoQlhYZMHNJAQt5qLEHrhr6Eji5YJSvZTvlPo
Ekol0JpNC7sYewtOfvlFrXuzaVx12L/bS7MinJw5n+oPMI4Y1Z/gf38oQzlh7Z9eTKiAxuw8CoUZ
+6gPmDaAwwRx7rb2dObYsjq09p2H6Npp/PmPIhnX2WAWwNEB6SNWm/gowi/mLmsmXTh8u7PTvhZ8
2lRWcKJu6vyf85kygU2/KE3ZKHYb1VnvdDgyhibvCR5UC2PGWZLxM+lorNlzOz6kJZJgjg+LzR+i
4XhYluKi1ftu9rDhce5/D0+ywEN9SnXbzzClORjO3FNVKARmibSdtpBQEAbeyqnLddmQCQqlN9C5
yKDQfRIpPQMKuiUjZ398meZ1aGvFcRlwAr67iwGxwMzaVc260ahNgA6wUQ98MsEXeTejiN8cn6yR
u/yBAajzpJNXg0d2CZUx3Kx8dRqb3AvZ318NKXmKxU7PrnVFABJ4TVnvmRF4fpApxGGvsswlS4JG
Dsi3QM+LQC/SuGAWMb7Xb55iKtpnBvPDAvzkNSEvX9peaCkqR8z3tNaeJWuOGs0m5PpTVg0l5GVA
UM3G3BnyAhIspNe0XfMrKWxKWoEYrhFMb3exgFi2TZoQtD0zr3nN6L8HgI9K4PULw8YD2DDAIIyn
2pee8nSpa6v8f8bu6TBHodJfD3tQym+BUlzJcnGdutzaSQ+s9rb9/1D2BNQ5iCeacTUr/1tSiNbV
9qTDluTcGsFWvW0JCYc3loyZB9M5Us3DpTfTMDFAL/vgDTeTJgGNu4O9VLC0YWbFmWNxUXR9Deis
VlSMuPDJHahKnL9aKcCOVtoHfvN6KXJ0Ey/eyl3i/phYAnn1bQFAySOk0zHcZzISR5aLk0JHUKxb
i3yqlcOPgelcP0NMFjzqWMCOqt2rod3eUtrUJHY+0EZkNcWXP4zR7CgZmybUB+faDG7/YqChwa6o
R/QprezFa10Ps39Vt1dS+CPZiAyaLDGTOsTf00k1DTF7yE598DuLtlAOUwG87BrVqLu1RbQARvJm
6kcsetW0qzo4YEuCc0M0bdfclSnBkifosCH/uBykIltXL7Fh3ZScCAfQtl8alJcS3VqqainuGyXk
gxQGWoy8z2go/q0fn2H1nlnIRx6WnMIO37XJIuu1BfAnETpUOVZ5VN7k6aCVVgdPsOoieCDHA/0M
9OA4gha5bj0q1ISjLK2JS3f9fAZX3PfxJTPm59A8Ll+n90mt7W61k4iEpuFg7lZix2p2Wmg1e8wO
CU6lql9vK11+x/2ulNHVdWhMifqaGt0vkXzj+7VdYYE1gDViSRg5Sqt7yY9/boN3x38dPZiELZim
kHXhg850MbqpogKL/hyhZtorTkN0DXJ0RD4l56WFaoENgCm5aVGKMt5e6Z8TSSLm0PlasiAnXMiZ
8Ez/w6sFRNsyt0vZHdwSljkNhCQLZqCK9mlRA2yRRxCBun4ELDc0uOntwV+yl8d6M4r6wM2plgJt
RaulwsFieZo9xo3Z47G/AKGF/t6fPLuuNouy4j/BXjyc/KdTNM5UZQexFlXWFbZJv3imSsERlquF
0YbS8YmSfSfNH9jEz42LIFC2rlrN0si/ykYJG5nux4IeXtSAob+y6P5EYQz48fZZ8Ymqicg7H3rd
w7KRWVYPWW0zHCIMNiHv3h+eu3kI6YJgn4IU8EAfZaaL+FaW+sOlS3Qod1FQaVclXNJ2XMLqArxS
qY9KpzKM/3oXkTraewLGDh2XjIb/zgG8JSHlBZ+ZKWvIWxC3cbA6gN6/ToIRmEyJQ+neiEKo9Ntp
mYi+H20EXJYk9NrM2oorL+q4ID/oi2gGgRmXYrJJVZc/JPXRwnW7HMaa/yuh2Sp0/upgP1wYnDUx
Ktmnp1WB2haTH3k/b1as+4GxSv1xZCNaFK6X1q8oK69ZuaEhXykhMpQFV6r9IXklisW0qd0qWd0e
kf5bO3CudRxmap71tosW6Ssea1yK/TZ983XGxDNAet/Lw9dMj2qo03fSVvAWX0v246n4Tfe79PCl
WCLqy7V7EoiFRIucVn1vbnJXu1+5SDvkixkvAliwJnhaCQpdSicOJ5F7QIaTLsSFd+kHRbtyNQoF
BUR7oUrMNlwKM3IA7EAAsqDtKGxe0ckdZGYqMJN5T+xtd9rs7aaO7BL2cqOkqqp5p3PhkPY4d3Bx
h0usm3gEndz/sp9umCUNkqeAKj462VP58UHnJTpc948yp2BAVIOimCO+v8mLr8pKk6zDcXpVZAG5
/eJ8CrcaDVS743og4Bi4+RNjSh9NekbQUxtClHiCe5C6lvHbByhq8nI6EB3E+vW1ISyTko0WfuKW
jcURAr7c8vh++AS5YYkHkYQD7J7sFoa3H6QzHP2Ht7ASM845Ye5H2OxKrVfZodRYGRXMKBQHfgk6
zmLncl++9v7k5kvUz3xkgM1uMN37c49ao5/FmZHhq97UGBjrSCt6qrNm3D0Nh6xlf6HJ9NY/LcVV
Bj7Ss3B5d6o4wf4XOL7rrslQtPFGlXvX4W/GNDEC3EeJIBzfYc0rPVtKoJwuN5sZ6ubvFmDfOARk
jqVyCXY2QV0QZz3wJ/Nqqwkf7XeExiothQdkiRqk0TyhKfpijXmIa1AYUELg1arRWx/YuK+WEUGR
pXQ2tRXFbIoX00agvF27e9Rw6NqVjS2Ik7Vn6BHAZFUfU/EsI+SxDdumR//mRXBn7WMDWU+MG407
WuEiBpfF8si57FfvTP1aFCQ+Xjv1m9YTuDzuEgAmXGEXDKfTNZaQJtvN/93BFmdI/NUSvLAKvM8e
txBjE1O/3muXJKzwdNe35p9uLoZCkUigzcdvLllMI+Ex2duOEL4feIe1CJikFcyjfn3hSER1rblq
5PAq3G71NSgOK5S7oIpE/pAYmhHjCGSYdKwFXdys1tihVr3GPRCKFhSY1I7HfuINK2JBJC1XPf2L
ADhQWSn4khPleq7ChH8Xy5hvqi1Fw5/W1V+Bj608rn/HZyK8gwe/0v36iI9Mdwac12EBbM/k8gCy
3LBMlAem7FOprZtZ1c6zVAO3LSnWFwNdVoUviy4Ak8gqaXkP45b0qtZbAhDbcU0h/0qa6zS8Ctie
O6MNVC87TKV8A1KHyfa5metPR8ee5lafPRRPBY8fpaXPYNWEjqwIGigetRWlygrCxa4DqDiE8LBV
wFeRrHJ9V8sbfYijvK2pxzllFjXr+nDJOxn1u2ozrkRmOyNuo2SPEc/qOr5b1CPJRW8OCH6NwoYE
MYy9B/n2gFb/ADzxxYKLRJ03OrknPFUJ2s5uJcpSOtNJbFwK6aophD6vhmTUepoLI+g/cq6kNWZp
SZY6XiVtoexFuFX5jaZt5RIOv3u1xVT0pJ1widmtsNxzHEHwQheBhiAOFH/VMoKghLS6FEkTV4nk
HXMOU6lgqFs+ooqq41YQHCEvk6ocU2OFlFYExkiJdZj4UVD71TqE7E2fO6q7sOfyhTpmnn0eVWtg
NN+KvJ00WGzAcrD1JLJA3qHn9wtB/sJ7Pf6G+84nEIwdpWaj2QGWwvQm5O5tYPJWabQocNrxsjeZ
7gL0mSH0WivYb1LhfwNeyGiJemiP67Yjgm6jZp3GLbo11Qs1krpefuS1fz2vT17U5/3r6dgpWUaJ
CV5zazH99+87Vn8FJ+VbZeJ8g/OGgVs/iaj0wUTuKRiNAKB5rM3GX5fOTtXGBgDASeaDEEd1fdp8
N0FLwsAp14w2vDTgjSWj+KXl+WJxwI37jtkUF+iD8CQpZ3K00tHhaym9IQCRanrx2GD6hQ9IRfGE
yI74i1t/tcS8YWfDjphEx7PmnCPl3916s2bQ+Lce3KAkeeVJ0xUzIXDhfPxjdC//yI5sO3sYrk+P
dlBSlcCnnwtgFngC2Asjf0HEeHELFjlE0cZErK+PkWMqZgsdy0J5AUjK3UMhftXgQIH+qLAXljWk
XAy/wz2SlQn3Vy1zCfDD7w1NXPIMMRUFgJvJGXFIvGtx+MuXPOas0o3f759eDgT9OBnud9ntiQDJ
ilVaSkXmsCzeRWs3XNL16IP6g380eZ6g7kBCV9iGjgKkvcoM8+QLzwyqSLmB3QW2JIBCeCR6KhCx
nKzDExQD3ywOwi7d1j5U+mZaoK3W7Gt0j1YvSJR6PFoubXvVqft6YFdFzEWjPjJTkrRIZTH11JJg
fxqGM3Mwi6Fpr174AXJ/VVGwmMtXRCFupDCu3U0eIuCAIPScOE89rlRBxs7HqIg8GQq+FKwBMguO
dyePApi9BuL3C4C6cCsX0vKzr1LfOx2jTbRGXTeQj68rDFkwh9XBT09qTkMtVmclWnQw3KucrY6q
L0FOX1ZUWJX9/6ePe6elej2wUDoHouzeC58ie10In4n1iQiKgrpSUeMivQ+yr1pr5nzLQuyrl5F3
slQwPtNc8+hfRxOcQf4TV8KYj7+6o1QfJxR6vinx2XI5V9CyX8EWh5k56pfYLofKr89i9zQox9CU
KjxUV6YBxoo3ZTqk1r9ZwokI4gUdvB5epPsoWlZrrm92R1SkSQTEQNO0w0NVH26oSB6be1Gzu5+B
0K0o24lFa5p90XRM0FOi+6YqSylPXbTD4AYz4GFRQ/DdFM9oaGcT3hR+8UsuCE1H77txtfsNNXBR
FzdfvliQTOQeHenncs1TZyqrjiDcG0n781MqEnRrDjIG1QKhppHO/UC8j8fvlIX4Vc5xkQGE6chP
4wnBLxzQh1d1+EMR/De1OKJ8FrK5PQWotLHvNAKjWY6XtETRkYLxgC88gKZH82C8chqB7tBLa7wn
wCceXe4Y5A7wobZzvW/cv1+F+YhvhAIPgYc5xAcBJODQ8WvI1rKPtP/nCZZ0p5RC1ZipurBl215K
nfLyAP1huaAmGb7LblGJxYMvct9vhDfXwBRh7BTZjAC7AUp/IeFsWuWAW7W2j5AGa/G1PJ4rMjSv
/b10ajLC98lVorUKZcOjL4N8yAa7r3LIgv7hXmUsBv6fv391NINQfK12Fo40IcCIFVV3yEw3wup7
KXCbh3ld4yAan6dCNoZllfdj4FWDaPeqVIzczRfcjCp8ya7lHzoGIjHqCeXpoHpVZnHqXSshlIVq
TsnqUfSEml7nlHYMb12mn0GstRHzeLiuBkUItl8idOnKpVYJ9aIEJhDnnIVQhzBisCErvCFliGM2
BuP5vsu8acAiUMwonhx9E63FzEj+LKz6EYY4YHgYgC/RVOw8lwTKLk2X94addvIFALCvcA4RH/DH
2XdxmveRyEMkyA5zTnZWQCJ+i0rodmJsf8Pl8QFRZ4yhz+u/Bj6cHv65mQpnQEbqjVdzWa6yBqPq
aqB136KhGwaSjoKUzJ5QQDBzUAmkzfUyw64CRoicdGuZzMFAAg9506/dN/jMBo80Uj3XLucgo7WP
g9QQuJljcBVuVPfW6sFr62J3lmpiBHtC9BS1Vjm2pTpAd+9+WK65fTxY1U3ZRUFbKC/mRWPgqZqN
PAOevOWeneWYfaSV7mbIP6W6KbWZP0G96RJJUp5ml4KgJupCl26Y0mlSgQqKD9tyEvvx2aObQGqt
y+OjOzXD4PtDRyvOICmfrS0HnnlNg0Spe4QxnqfnAjGlsO+YKuxbk+xtyYV30josfymFhn+4d6Tx
MLsF90srV2+Pp3Uk83TFnco/kKdpzQgETi9LqiwUP8nIqav9ghxtn6bwZP+P4CliPHrzIO2sG1vP
QNZ8q84jppm5hEdC4ULnFjtJpQYr7ErmE9ZYayYU9ZDNBTRBSAmEon3RDVmFNX2i2LyLLudOBWdi
EERKcWszH9ECuAyqonrtHnzXGG3cZm4FPur5qcR/MlaHLk4vXUF+t8kHT9deEL1EYXcqZ1ulwsBE
UMMvsnWmc/4c384E9LNaG1fvqZEmnRS3RqaLsZJfLWUm2EDKtUHyVvpNEz8BUjLqRNk4HA/biipX
6O22tq2UvT6/abUmOnvNxbWjDvi9hduGKxYaFJM+DwUjpuj5AlV9RFGmWNtGhO7vuF04TF9+/uj0
NmGcKT6ZcdmguJYAkGNw0K9aO+4Sl/LaVNIm6k0G+WVpohz9ncr5Zv42IiWofM4H81Vvm6MLW/BV
AtwGN4W9vDSPEgWhT1YcjVaeYYXYVQ4srRHXJRBAQJrj683PwtQ2P2Sw+royRiA1MlNjgXz1lmWf
GQXBn9nJcyoqI5UjQ3AHB5NwSFy3BjKqCxlh8N/kVqdMpN2FGKCuEpmtZqGgwY0icN0GaIezcG2a
ABTa20t/NJ/8sv7rACzaR4ShFr4krflpVS3aRDRyg9l9Gch/xgXBvY1MIYSzjA2aYnEb+xCYSvKf
W2pxoLfTB9MXU9qlNzMQ092MqUVHj5qVO2a+Taj/hTUCGk9WmXxalRSDeQCH6qK8wJFCzKsh5oWV
sixoeerYV1DT7wuOoPmFeNKQ67oUp54WuHcaSAEKersrRwqwelWKHuUZR9lhzaB75AHYiR2Akask
Rx9/sQDfMfJk0NYRkSAaabvR646OA5/k4OnMyrNULZoILWEiqpiEOv8QCf+3BYeG3T8U3MJdKCxi
Z0uEVStOdl1qGQNtgDt7aXh0qNCnHZiUaaVpk1uJJKKLmEPrYYx0654u1admQU5os/NI5G3jrk4D
MwnGFiHiyFW8jap2yhZRsmahxm0GudkYjNZAPXQ9JYNw9NZuo68sdbhximgyUUSIsS0ATslk+ooS
7JWQkv7WvJOx2phRBr3+PCBpB7vpxeyHeMFWVBwNoF9ah7VEQ3hUvh54smm0djQM6lmX3HDIN6cD
NUK08ZXqSwVS9qiQMM0vpOO4L9Xtkk2CSRk7pwqOyZXgWuWezqyzWVs0QTVoJX36jQ+AFwx53OrP
EuPuAGs2g1D6gqUUXrjmgcIWvvV/I6K3jLLN1c+vy+lJv72UVyDBQ/2LjyPsF7U0seR4iKrZ+LlK
oM+Zba1tY7iDAf7kqny4Nlj8J6m6kHFMiVDh0MIP2V8e+3iShZ3PERiRqZK5VFZMONZa/OnVN4KY
G2j7nqY5haC1OiYj9C1INZ/YOXr6Y2BPqkbLNXH6jJmGXL2FxdwS01Y8Ql7BupnAd8j3Ufk9XnPR
dwePgwnXs3kOPQDxAcZp2iEWWJl2Ek/aEZ3BxQvmhED0tg8aGfdpRBpMV3obpsxwGsXSqxXX/uZg
nJHb52AD4ZsIHMWt5maUmCmvDjt19PIQ5E2McmV4uzVzqKrAyfoFpPn1t7QPnvGJmkzln2FY34QW
ZYb0e1SJHtdGJM+SdndHClC/ykT+XMWXqrLiFEmLM2im0ZYLJPgLomUyysje29+6hSvo3Dl2DFWv
puVRmKjxNBM3949IJD3WFNVRT++1MGOzh+aS2cjeQSV6XRJ6oAKaSib7uG5px+Cu3PyONh7huIQa
u1ZNw3BVDJzX+9jbMCNbZvDFnwPA+NHIet47IoyHWAnk6lwhwJ0uvNsVCdpR5KnQeKTNGc3103Bi
GyMxnqjnBpgtoNGXmcvzO8aJ+IP+Cb5ZLvYDE0zLFHq3yhbs1o5sGeDPZtRxUUlXuxvWFoLeKhlN
58dP+CyxMaX8IoGx0RHSuc1W6tSLkXZXpindC4pVTzlVCb6mH+Ac8Yfwsn3SNW0lueF0cEO2s+Po
0olozur8fQJrNPI3S2DnlwAPxoinzVa8NMCkz6uNg12/aeZlluExTB5Y9HfT+Wm8eTbTggQXhLjz
VeH9FAWjWIbuF9e/LJ2Y1y+EMNT1H5YKlUlT3vC/U0VAcF6Gl5T9AxNgjPzygKonQnFRRwsaczNq
8CecmAiIMSexuysTImos3B75IujXre762Vy9oej4xUHDbo73QB/zUvq5HguTDgUdy9ie5UmeMYT9
JjX7Q0sjfLw6umy1Z+5jJTTmh9iBzJ8hgYGddMoHJHpQG6h+Obz5gVC/NgiGbiqpsmZTMmo/J/3P
CuYNAEODfzUGwAiEMwq+3uGJpqgWJnVDoxo0i7sm1J11vVh/BQeJEvKE+fOTL3a5IzfQOElXkgMb
NLozSAUaKs92nWVOms9/VnyKFR8fYNHj4xzSpsny9FLJnNVKHc5l/QdDnYeMjgtfD2b0pmIS3pPP
Ckqgqms14mSr7fVtl9Q08030vKsjTnvmzeL67mZ2gj8nBpn4FfVz6XjI99An8CwKfLtzU0qjrcAA
fQPJP8wIEyPY/99xzxaK+51JRUlEVHGMSDAAfElXfQjcSp4N2ACGAXoSQqiajIMg5GCk+lDL8DT2
GxnRBfuB/4+nFftKQCxrC5vI5lUi0KYSpGDoNA1MMVdEE1va9SIT2wEeDRgUCR7zUYCVSVNdNp9o
dfe0iOFx6as2LbwlFDcvjbQJORbSsipAWgvv5UwyhN083q51nrIgBC5sbrKVkvuMsxiEN7BmZ8wn
ZYo18Q4sbOwghytik+//ElA/ySCJ6jDF3XmgK/lskbszn5zSEs4b+3vsD+CjleHeYjmJVGnbhG4M
PNXp9bpCPP9UgafOaAZ+yAsu73axH0RklYJRVaarxC65SHOwXPMSFpGimPDDQHPDgJltJCOoKs+w
8JBMy9rH1u6qCSlBNcMyUFhghw5k735KfO9d9n8RGEvSqMBTr4kRNliJBq9uR/SiXOd2GJrnWByf
PZnM95iiC8wP75RmhF4xdl1SBZ0wlyVck+v6tFe+3zw6WNFpzXIemXzlzDsxIU/SLt3yr3/tFH/4
KHkJcNVZOcVX2RsyT5MMp7nQUPJ9AI2qP+88CYF8VYAjrP6jLSRRt8Gy8/Hqj4b3H/4ktiSH0nGP
MYT8lYMXu7AQP/k19Rh5zAON/ARhqzws4KwTZlH9qRbVMLYLcNcL6QUTa7pBai93RWiF3NvoGHj7
NQVRoQ5h/N9vm9vZ2VxzY521FBQ6otTJeO/MtK5BzefgBS7i0fQE9m9aeMmYFW0GREOBJg0d5r9S
0hkWkIiRDRknQPxNYvhotwKILt/nhdWwTaBG9cqImM9oe/TDR4kuBWWX3ma0UtejqTRH3jKRUaU7
FQhMuVMqk0BhloMXsCD5q4bxdGGCIT5Za0fabFEXLii3O5xqr7OPDAd5aFQE49XY7lyxJuW4sXeP
oheFa3ubsdMzpcA8MVJjEz+6TNRUwZAyxoscbR+dIS2ylouano6/pzBbjL4SwQS/wOPDIhxiCqqb
KyYfeFUnHqFbJnkYElM7h3HJhjjFzSiL3frbkIwqIaKGhE2LPotcLVGndFMhcSJSQihW86uaYc1R
9m4RXic720AIUgD+x0Em/EusLUHxTWQc4TVFOOFjblLcoOdf45Kvwj2syzOMv5qOIlf4QHG1vp0k
slviX8YecQiLJJa0Sr300tbGGy+dwQSrCTmlrtXY+IpcOv97rSXd9dx+dTGqotM+w7DmfSGhCkAr
H+v8v8cPWz5o58ePUje75FRnEQIB4wi8UJJiqxLzb1y9uiLxZ63E59NZTca+LUTKYFo+k/3L/ff9
v33IfrGMbcW5srXaXH1ESsVjzgVZvzJcykb8bP9n2Q5AVuFXlFe4ICpFsQPDeBpTloziWJG0UiGU
pF45jmPb5FYUI/CyuM+1wdad1oJMBEflWLAZcSWk8i9JTPkiL1OO/1O4IGyyNUZAwWww3TKq9qel
50oOPnJQzSbjIt2aRYRnWYHaEOwptiaknUIkA8fsWxSTHU1cEyCaehOiWIIJIwZWaowefd7Dhatl
SQqID7Mpj+TJEDy4Du+YMd58YmxSDYBCtL2O11maE3F3PdQVoFC8/Z4cpoBYL/1nirKYzmBDui2G
Y4494VB3Q8AziPKkz/XtRKXzZkGQrdRXkm+1yf5pqgC3RgoA7PK7dpofP93tqeOuR0UHky6ustCM
v7b00yP13WdcU8zvQPSx1qFbcWTvXdkWXIlafSU+2IUVb8Q8GvViQKhqUo/6QmNdPs/+tGTurxyX
rd3tWDlaWn+qZqrS+FNLNa9KAUIGdplzXt1eh4i7hkiZyfp6S0nfx9jszfJFkFDrt+6FvbNCQbKO
3EylQ0cVupvLXX2STCMF09y8u6RfcYf0Y2w1fG9oU5QgEpDqCS7xkjwvAz05IsiZ0DjHBtYGp3SN
TLOJGqMLDQsbGh6SnCBcLPje7wFSOLR+aFo0BZnqNXXj8dwaJYI0SsIWON6obCpvVgDQQg2MVG/S
cu7m9vDE8nJzXqfWAMGajhLOKdzQKEEinpRLIWXJN2AbJp+ChhSQ4t/R3Bfw6oWqqKGWep98S0vk
O1066w6WL7O93KBcVIDgX5U1yeoLMjfoTvqYwjqA7pV8POOaQ8mQuGrH7dC6gfoxCTFhFIp40FLC
5DBQ6Cpm1S7FzSUD4py+G8K7r8fsKfp3YP/Cka3vcSUV9CuY7ItYhguadaVZ2HvhJ3bcEW6Gz8Uj
3ocg2qGMDaN9cbZ9RUFz0LXNSBx/YEQm8DwM5kvK6aYzzpAM8foJ7j7sKxNOAJmO4eHFGrWWsDh0
ry9OzLkDvZWZ9V1PO1wAhL3VZULd2GNPK9Z9OL6biqqxKmK4ic+Q7/pAq4sqcv8Zu0c8HxvKyjq4
vF1tSnAtLsn7HwZX/AO+TvcLjFHrJiSiwI4Pu8zL4QHKU+t6gwVlqtpjEiLD6LWhG0c4csk8xef3
OgRXnSVXtnjvJQ1IfeUXVtGOoW1LXU/XKY+5+PY+8XA8rfQwDvS5vEPeiGE+xLdYXgRhEeOfHFt/
Kn8UOeyOi137f2pAkMauLQV8868KGoN0ltx1L78zeLluEDjUKnpKdpvWgVnBc9HFYLp0dg6ckNLx
wcDoGAZwk3StKBuvb+mtXaFd/1HvIW+4kMJKcI4hYXNT7jolDMDvAvnWdcPwsqGwTzuCPFamUd/x
9kXzK40mz2zqJTgR5OAMDNhGxEVlkTjfdPll/ec3rjZrwWx0rHC0OC4yUJ/1vk1G3YvBR0UF0hjj
OXx4+S2TAbtnXQRz+Af9Brx8Y3YBq8iB9SxcB7LFR7/oLgRHLeIVEtHfRv5VZ9Q/bKZRVy8TXY3n
TjJW4JNI+E6YOBd9bzRSTRLcU4Gc5/l94IxAyLtYOuZfSX66SgE1QEetLQSIqhAwuC2PmObm3ZQZ
KoS6DCqoqV2x+1QstMSUmQS3I+W9YXJylLmaO1jxuBSBR89RYoFgAt3Cd0fWQEfo71vZmQcFw4dM
2R0m6FPNZAnWAEk5d9wvB5KQQ6ptDj4gnjWbuR3EtVT7YFiiYre1gJ8aSLs7Srxp4ZqxxY3AGwmJ
kczvqmQWkhA/IR0f08NghugNHRNJIwVF1vAQOBkvtF3vQFlbDYFOTT6fITxVb7ehl+GAyFsTh/wB
6yduw+R3qA1WcLYiNTRykns8na8bgORiKnkqYtknYH5vyXiSbFinjsjcs0qKcPDrfrIRT4WsdXuD
Uhc/ep4xcJhHK+yLyNUpkrEcgYuQ7O9b+0jyILM4XnYJclK96fmyG+HsftLL0C+kIi9/st07fzo6
7wEKu8LZcO4F8/GBKRgkrGuR0dMZG0eadmNBO9VGffJ7pY89KgTpdN8tRKJLEnLKkL1ZhAl6Jnsw
SCPhVnqlgDuM0hRvKQ7oqUhfFeFUC6sQof+jtaSacWba0nHszbwU8qs9E2H1u34MXa9h6FcnvOCM
IA6H7ubJ/PVh1D1k9vA2326wgw+UxLnnL/zDXUlcBDIl/8kMs5UQVLA1mYDEmHSCFLrq/akjUKWZ
/hPECGfq7nIq9PnJONEVvaCxZfdbAB57LaLCYYAcvFfSDcZ+KWjuP3ifqEpa1l8GJta0n+MFkCO6
4SmQoMcW8J/34+IsQbeoE1HW7XhJDMroHt9BeaS2zoUVF7J+uCdwZQR5IyZXIDue0XLpOwLHGlCs
UhyKUwa568Cjr5zDDLIJ62Kj2zgc1i6zyikTCkKDCUQBqesWjB5x5ez62lPQTGs0ffxD4uCfRIpV
dYlzVIfq3aheilq68zPS7pPdqtpxCLmYSen7if2pbZGyV1zVO0gM4gXO0YLAXWJV3ZSxq0DgHPul
VUtag6CNYfRevbb7NTpvOn0mRBoZpFphjyCp61G+PqSm4Uu6xeUxRAyW8mBfVI+TXNdl3Gintgpn
ITx7bA5gPtzY8k9V6bK9NmcZypZpuk3spzKkUdIYBd17t8OtBYLviapZBFldmv5gBTxtLN2jwWR0
xhJA0aI0G7yjGdyGDaqT5SWhq9bvfLFT/BpzVjmpYi+nvecY80WpPfdYsCDg/Ybg85KGzp+/YAwR
2gYlvbq+lQt/vRt3CB+0GOMo2P+Gs2b5fm3jSIv5lhizpgJvP4Wk1W0BzrMGAY2/l4deJTIRbqWG
N3w4HdJ/fgFPFL5r+6VJxKkgBrYmRAShOI5aDu9Xp9oxzpJijjBJ1EEcmwKiHCiZzJBYweVdFdzR
WcsU8+e+REo0J1v9NEdvhjS50SJES+0ZhX95BKISodUWpIX/7PXAepGS3RrJMFMg24FGGIKpFn5r
t4CY5kKYwTxVk1tND6o+Ea7Z+R57Tm0qaKedwU319ZssRZiGkIRFk0Nv/Uj1UlC9dr43fsgFX2qd
zuLLcgmw0npzZIy2ymQmBmIYfWA1sVkTUDjvH55aF+mtHXH5IOacePZMhTHKn+hyy1SCXVvk2gNb
GkOlkSMHKu9SJGJa8C2HsylXdqTr8mbd10bYwQpl67hfmkGjOAXvm+AjhQoW0XaP+jzw1S2TwGFM
gCRh1jS4Wfz2axHYDCWQ0d1Qh/DxaDXUqeWbaOXV2P5x2wqR3w68sjEbjFZ4Zt7E9PH8dhenoFrJ
0AwmQ7Ojd2hP9veQg8j6/RE2psLwEhSw4Z3me8NzeuHVh7BumW2UmXvkY2T8E0qD2FDdD69drwVk
gewxvrjtSCPWFyBRgqOTSLgjNFLy29AoqLC4hEj0oX0HKVJZJetXVS3pnV7Xk/onw+Hnz0/GRkcH
ElnzI5H69Yk1E2iMPUWMreKrhUJZemVs3GGX2duTuVzWZPXvEcSuX0zB/p/ifP2OV4qL/K0nWqVp
sPayEg3/nNhqM/geNmh0WuKykSpkhbwCl8R7ObC+0LLg2m2ihhqkeIL+IEtmaMffhq0A/eu630MN
Xa+SEDMfVhk/onlNjwAV65KPntouiTzB38qV9m3EqU9/mac+8fv9noAU+Yv8ClYcVf6s1EBz12hT
D3/2gT68Wv+oHbbG+1pxd/W0/a8b9srLrk3pBn2OU9pdzyLsJ8rVQoTGjKvx6oMHiEyvYorYEf1L
aJKbII0jlgBCHSWRanxYD6nizMurNJ2HONbQASDuECjHah7V6SPdJbyyKWaUycz5sPVxywkirP0+
AsOeD+/F90WzCDlpgWv1fdIWYPWBaPHDGaieDTI1fgNJZnqzzxg+Ym3pSXqdLYHsnQkmU+feAcbQ
XqCqFgdtyOmoFXX7nOJEZoB6w/ZYLdxf5d9O7OYpmEMsDy1kaadbWBqWTIhcTAOGY7G7dMgf0JYU
XP6RKVD4bQkHR0JNMXXvpoBSJG4zd4VgPzQ2YmGTTRpJcJGPripRtM4AmrnQDNhbj+gkgcRicOBW
sOqno/fclRxNF+KWbRBbXnXHSjYeuxgFzqeDzRXuL54lfWAB4MrKMQ7BI/FZyIkm15ka+Vunmydq
nmXfJlP1Ifyo1ZbF8mRnBHmXAbt1UPeZistWvxMnFwbz42OjXEiLvuRtrAPxRFuIZ6KlQl0u2VWL
7+bTKNZgXDvtji8/SfGesvEbLTURwiPicNrccx3ilVVXwn1HP0dfxglooaDCtLzvTbvwm6T15MHb
QzNsrZ2zD2OsCx39FhfiJ2uco5LK4FOVN8vJxaDqPiKoz5iwN1FaETCPK49ZKYxUYkH85e0PJo/+
fvSyLTA/ag5C/GNkd3cCn0wkgX9K/PYHnJ+nNmQAVTjLX6knf4bLl41Nr9B/tTLNNjjsS9yvh9Eo
YIBYIQEVb1O8205SOPfiIHoVOIweuZQDBem+Fo2oUIc8dxin2ZkpmVzY22ud1l/yNmt3bQ4+EhkL
hMChdpJL72Ze2Sdrhaca86kMGoDerRGasbmCmKijfvNNr3OSdTBslk6a7JXrlWTkyke6q9i/MeYT
M0Lvbsv5A8UETFmH3Vg3V2W/wz7HirAk4S3JvoqiJ5ELoIgEmjdo/wqeIwOOeIi3xNvngt4sbDdv
nkSzXqIotAtnq+oG+OowT8xnA2QO5gWp07Jteq5LTFh+UBA+bh4reCC1atbd7Clgh+QOj+THx8uL
nKBSumN82BksAaT32uNSMXyYFD00CTd+/+lx4XgrracER1IL1xZqOUR9Bz/yGmBGkDZCUf2iJCRP
2H8kKMvQ3jeVu1RNF1s6IfNcmDYpN2p7TRX10y80O1tq8d8d5cgjAYnsvyLP6nZFBVqEkGV0159g
TX40VEYkeKhrHZvE12N06r4Jq/hupGkAzMhDWPGOWKGhuIL9KkH4W//8ofx7SyDsqhLNxOaw7PSt
rm+JYsSI8WKEWD5hcwhfWDUpKy2dzfwElSIsMWvXj4r2rWCKGTzviPko5LtFmJNW1zhRP9midtVC
LVlgVc1jla9dKkdsh4/mAroBjE5+uZ36J5VLu0Hq83jPYq3rFmr7URzyp7ImRqgfGeFqFHFffvn6
uB75AttKssMvVGzziw53TAfEcem/PvqPfXnklYFkhwvxIy9qOaHM2PpLKh9ZJesHWWV1sXjBrIu+
ff35FtYajvCOx+7tLvxHlbdv7mGRafiXJUXMqTg4IpSEik7wL4mxyD5vRb61fAp8XYYuFKrYvwTU
BNvjogWag9SBj/5jvkwR4FK0y449RNA033nSo/S/rEnFTa0XA3zX0Do4CgSh7zqBNaj10KG3z9IO
fz8b1a9GTvza7M9Z1zR3F2LJl7U5uWA1f/hx9DL9DIF3hluwjGMdMN4qI6mWEWn+M7lKyC+dxMn1
5nH7wifgDivdhI+YTqDDFqs74cCl4EKF+nPRWZF5JyhPyR/kGxAzEqq/ZuUERKD7Ip/R2IMuTgL8
7sc2FRSqji3PXglhgg0EE5T9eL8QcoO4y4cbke4DrxZajo8rZrZohHqkXvzB9XITwbOWP4EY117J
EH/U2rtacNHCs8tiOhRiPz/1oTc1wanCFs3iK+AV7tHfWrSmWVYvh/Oz9VjHGmk3+qxjZy8vvCCl
AOpY+yzlKfb+9QNTrB3Rn/J3cBrlN2/ctIvDUkm1uc0Wgz4xA8Z047IkpoRW/LutTGpExSMtRsKJ
HlbkX9TlxZMCxWc8bVEmVLHBdO7eHUHNdcE4Cr1E/mmBFSnpUM/wD0VaxGsybEwLcKONQU1WuM35
mRYmOf8TcDvOpCb8j/9OYxdw8WNBQJ+2saapcfdE5Mzf9K1eQJwQ/O/tRFqRPMH9c1KHe/eXL38T
1gekSBimwC/dxAF6552iHpmhUMCCMa71tNgd77uLu9eLBsfmEDZptynaS72QJKFBjumuCLGVP3VX
GY5bSo5XT9smdajVDJNU38TtofOaWUaHacZwPDERvKJJKqJGXxn6Jlr/U5c2hvLdoV+HZh62spT0
YLAwZm9KcE/mDOd3TNTIYfijL0MnGHoE9bSwfTAIO6H9DHcOCeOz2Gt/TSAT/ernqPDZ4myEKurg
EGtYDcJgkBcH/UwfsAE9dvbQcxWPuOflwSgEqt1Ev+1MfQuvNqGhuCQvoITTTt7HF9Fg7q2XSYF+
KldiWuwR6Do2Q965X2OqR+5CytmXiUFPpNQxYt8GqHAyYrSTXx4y0bTbPaWIgJ9EO2fwmsL5xTL5
AqS63pxa95GfpuKiobhS6/5S10hQXnSpJcSHz05q3qB/Ln7NgwtM8OPC6nw8qlanTl8pJaGXIGUl
/3syp8dAjmUFjKXbSnaraxCVgdAy45vdSl5vRDTwsT3ND3Oknk8Wx8jIOczpQgqMga7IDX4IkmyA
TOqGt1QOCyfEHoApOlS5s3S7EOOJWalKECv9Ua1zMeMYz3Tw/AzcoW0x8rKM9A3SsgydKkHBpiBL
huK/7jfv2IvyutdhsM3CSeAl9fm0sert0PIijfrkpoREifym0hYRD4NQIwCcR+rHS67K3pQwUnkM
OyxW5ercMpYuwfmiRlKXiv3Mg3r7KJALxMzb6NCPd/h04ZQSQx/N58f07S7rm3xpiW351DkjnkBe
A1aaNxBG2juUa35wajlrZ2zYSRX1ZgPyEpmyRb5kHuDIF7pWqdLTdtiZ1V3rAjnaUjax1Ena6P0c
DtOqZcSCy4L78ohZfVWLQ91PxIec691ZYExnQjEsab87cvcQihFdvdDdwYRliW+gmEuF6VQhHFBi
TlOHKcqP0qu92LIHtW1xU5RxRIeINFKKc3GIfe0K2rOQTJUxgsNlBaE2eT06lV5yGQABYw5tk5iH
yxaYQiqfbOQixcqIHEx1EVRvL2S8xSZPYWLrrRnqS3v3zOOc4XYqB91CNWKnMvr0DqeG6hLmWfLJ
m6hB/8+1ARHNFJ6GALZlDJOe03sUfz9KuCw7oCAGfaRc+m2PQzHC0/8Q2pSHWiOYOAReqs7UiqP/
D7VT7QW3ozpPKW72+/iD0qsXLLAdq/CjOjfrDkuci67ZsQMDFqBZ8/Bfc2TUkven9ej3DH/W8CIl
XfFVsD3KmVtPXKFF/HoRvWLkH1ja74eNkSulgE/lRSnWiXg7BMmHSxG/izNgMPTOIIeh4zAJs6c7
A8r/18aFotPYGUPVQSHqyMwIVQ1nKLJ5rceGvQxtO/P5fSxnRSIpxmeU4UOdJ/taBYSd/Pu/D7fd
bqQkh3v+NmcOLQ4PqI9ualNh12vjSuIYmb/m+LS+4MKf0IL8KLTblEWwEE3+MxCgo0eyjJOgkOBy
gGDjgvUrWaAaYWWYztsq3Vlam1eToMTLoKGeTgVTjzvavZWmjEPxE7aA/WHx+zamQlnnRNM+FMo3
lu40ebMIB7InAUTgJAlFWTYduMtTPi9aNNg4CyzUPt5bG+w4xfPav4CstLwv63RTJtijZ7jdP4KO
jGi6ViP/kBvJoqSoIBri+y+aRdYN22ehUeD++aNZJsHDUhIL9gf7oQxhgED++IQsfunY5dlxA+jd
BZib7XGg8ry96rbyDt8Fd9lYQPFFC4OeB/xtsmA4UB83tEE2mq2VUhYjr+W8dmseAWUHVsqyejOw
S4Xm8+SDMObZvYN9RZBBKUwAuMbISG+IkG8EVThapU5L8BBW5KB2GXMe3Oc+zmTGWHsELiwntlyv
+s2Rd6HPOUNTLQTHtg8yHG5W00hMQBKtH0H4vmh6gwS932s41Vh6dGi5pebSicA+jUy/JhvDEWyd
6s495nXUpaMk4dJbSUc76U+plajslsz6OBjCuMJLSfZ2fCG8Vr3gEyy7KIs3pq33jEZEfhfpaKKg
tz3K124FvITquS4Kys6xF5aQJdD9KQjFBPsQNiru3sdx39n14ku0wfyhA/WaIKnR35tiM+lYrLs+
AXVsQHQ6Gbz/fbMkn1b1S+TzZG0DDYeZBlWAK5F2IcgBqHsxm0ioGStFKJPRGSa1N/ZrETuK++U8
8x1zFPj/juuYC2Md0Q2zumG+Xo0K4a38f1jXuKUHspsxMn1p6u5nuwnZpZ06qFLUUSHU1yRhcW6h
BCJaomjUbX0U2KzUZi09qZwTzY3htguuFjWkwPPRLR/m9o9CNj3LBwrTGW1652vFRZS6fei9n86R
PBGaoanCwAzKHLjvzmka2dcarkqfL6ICPXqyCTauhuEJ4nLjIlZkExPAG+dEfXMhHXHkJ+0a4HlI
8rG4fK1a/CXuwepzW38XRw2ERn8DHWr+SwS5wcjKA1wIa3oez7E7o8z05x400tIrQVLqlUAE0Gfn
k89Dgw0NIy7ZreKddGmdBCAMk4jgtaCN7Ubf2SgXxgeF1xj+XwIk5+WcHvqL/SebAJfdQwFNT0i/
Eo30OUtE++xyxRvOtHw0IcwSHkgr/eeNDK3ewtUm4CrepJBqEewuhQ/fvHXn0sTNARPYuPTap1eM
Fo/s3veMX/XYGKWY/v4MD5Xrh/2VZ8BxF3SYAtLBIwdOmDgkj+E5AEToHUAyzI9q6kLPnkUN96JZ
eA6jq4E613B2edU5eHmwMt/svEqce3G7Q09YrP35ufwkBFmtSQfrNgBasNsJuMRT4qh8larjb46L
Xk2CrKa/xyUgW0ZrF0MwyYzk3g1ZQ1Cb/x0iww++0vYDjZCgkl3MWZdAAzt7NOPv7ZzMcPV3ZxJn
t/FrS0NQoQ9s4O17C+VAx4jZf0XRjk4heHbmbfBYlU2AvLq/BhtBxZi16Xgm295wq01Q40LriQdX
lBnJ5Xy7kBtcJ6+5P03osQOmPVRQ3UsWeIvM6FiNCCLlhTLRLWBOYWtCM15rvO0ENYbIkU+uHame
1Y0msDyFCLxwWEGTJ52nW7r7l8hXXf5fpWNgBlw11t9TDQ2e7mSdSXrLF2qRLr+NKIt6GhGt3zC+
Ce5U9COmB2lklREDiOo8TslWSV48p7o64kpG9l9IPa1tKGlHgudZCoD/kFY7JKbZyhsaCz/9WPo4
TNieSZDhh5m47LLZvT8xREk/6Fv4L7EN8FCkpJMhUrmAiMY0jZQUfiQ86PTVMWqTWXm+JBxBLQGP
ANrfW1VtxqjwDyiPLg9bGUYLRTpJC8YAGZNn6W9hJYWd+5oUZyv3enDNW10cW+aZnnUptokXIKPK
fXS1H1Oe39fGiXE4zG7/PUGecsKP/SYXch4UGCVxTE2wRMB5DQW7wQJbD6UtOceasThC280Zma3H
RfL+59qZKoWlQ/S8v+qjHldUliV2Q8rh7o7yePKPSQVVsaS5HJk4y3eKDEr9H/UEtzsksc44ex/g
BWuGr7V0nAKPrTqkd3eZWlt/deDdzTtktkZ504Z5wPkYVx0j+r9xyQJ77gREZC+JDaotSozblzUF
j7sXFPhf9zK5xRQk4FktRZj+uvlr2enc9xu5NMDzox/Wuvf2+leZdl+uG2uC2pUqct7JOBm21N0m
wOXQyjM5XSDQSGZKhsPVND7xh9XpUHLH8gjVnu9xvcfE3pPhtnz6H6muDKe0MW/ZH15RfL8n7TYl
DGBsSF2pZj4R0Th/moioIR7jtdTs0gckPvXflTtslzJ6XYb4mz6uYoGAlBB19bVmnoIVI73U6buk
mjSwFEgxxiNPTyg7x4P1nfZFjuqoTIH8Tjmz972gITieg/SHZFoDZj8z4veCXQuFhpoAc7mCYkgc
DuzrGOatqT7ERNdql9ksdweAksIKJ6ZcJdBzgUZaOQAKnBEk0qbbkVueRaWJ7U+ikdQtE+CL8zwE
RqBnhFrLEzeBHuv33yJ8RIGdyMQf2OfihgoVzuqVHKR5GN+5PD7ZTFfd0U/NraJQaWRckRHlXKCW
z3Rqq+vgiaFQ2Et06WBsfsiukvEWOZrCvn58j5sJHNo2obChei8o8r7wYYRip/XUelJcfxddtAlL
xHm7LeXkdKYYmCXxmVzcIuMkCjixCsCBLj2ZPeiI57o4o+IMU+qh6iEY4xLl34NM4EPVnAg7ofAP
vecYZNXAyDXTJc32HIMVzAXnUBduXOSfMH3q+9gwJKQRFys7obqkEv4bpkhj+Bz8i2r/qnJzuUeF
MmF0WGCGOx0rz79nbOPFj14kODd2FWi/D6bxLA5Mxzldky8nH+ZtuVAFzBeAE3Ywlzf3oekpmOHp
XYpD5v9W06HynaFFOIPT8y9dReG8VY7yHWMXlS5sKDttZHCwYDZOeATp1YYy0WwGGDmm3+FBy/qG
eJYURInxfoiq4QWpFvXDFnjbkLn/xcp9N4G2PgjmyvAldk2i8yhE4zRfVVNy1ylwY7Ck63l5eKNL
lsg0Da/0wzPZOktQJQpjE3lNJm/3PL+OO2VwHyPI4ieYLHjHwl47qSP3xB+9bVlat62rgn0zANxL
RySn+xx4K2yfAs8smLpU8FEifS3UtiV7kRaCFEVlqnzTto/Tod91131hxylUh2LvWSDxHDqIRGUA
fNeIbmjo+tB5l8bf0c9tKuaJYkkmZmr+vedNMmwZPM3Uxx6R3gy/JlaXZqe3UuUmHvTyPRF7BDH3
lHsxBHUbpUAlg6KKqgceY3o+RRYlDld0WUxjeVy3qWP0RusyC+wiGzl/cT4vT3Lxkudon4jCNUqa
LOOzLLxUCTdkczmj/D9dq2dkHC6E2BWwqw2L6cUZSEaJWyr7Slxju0my17olxz+sT6wnrz4AopOH
dYQrtm9URz2NS63tDftC8LRpD2tS99ND0sG4u0Wx7tzXnIfSehoHu6/p5wBWAcvGC+dFdIf4eBTl
RqWmmFYmcgktWEsHn0Jqwo3gEES7+d75hviCRd0beZ/cHwnhUT/8pFKz2GI7/QdvdJAvlaeXSr7T
g+qv+9e6KXMLTIp16kbqdt/odRE2cchuOoQZkVKT8nEtNIBkGI0N6xBBCxA+/jO5XEBDkMcpLCil
GDALajb+JjCMP7aPGf78pppdSv1jyV0EmBBrkF9HU+qV+ew8q4gYMrubf95cA6BfDFfcZ5MutMvG
CZsB7rSBsVUrd8Sdd05yNY89T5szfWfnhUpMVG8sf4/9rIbMcvjm7dieaCccIxx0/5IkG3Z3PDgZ
aJcH0EyssSAEfQn2iWezOIxgneqeSwiNJOEEo06/BPy7xiO7qBrxbf0CBJaIGShUOwPB7CTChyAo
+u+tI89355GUun3/KAhkJa+TWoFeGmUHyAB91v5pXv4TZ1fMUYv9j9+Chy7zSakzOKJ989CBP57e
50HENrdz5i406c5Af7s059PnzF/gUjlE44+LcwRvnWSZ6jqXiMBSkCjlwk8YYH/zJvISlyfptW26
CDaXZlDV/B4IlicnX9L1TatwXuMXCzfugpMnCXsIa7VSfVIdXYYl9zRIteyRM+CxLF6TCmWOGjWc
3KVw0bIA5Wwu7WsVuNILVKytdwZW9hYX/QQ15keh5zYW6GHelIdSAXtC6zCvmAakXHfrgNsloEZt
bPijiTQlqnGipSthx+jJ4+8OTBlpoq7MMpAK+bDOILoG+2JN51OIx+/SY1KR/iTnpRKkXyLNP9ju
7An/PF/8pPS+Xmjck4pFEoefpxmnQ9URKXI8UXeWDFVKANNSY8YHAeNy353dfCs5IhO6sDLkpvC9
Lk1K1X8HlDL1ukxdIfAjCT/rhLx0t7dJrTnlAg44vmj5XR5cgXOiepbnvJLlJ8zqR6Q28u39T14q
IhB7aoV8CH2JfrVgqnfc/UrQ84sP0IkxYqX9vEGZEYwhXCV8XT12+MeEQQGOEkjn634Z/M//EQYB
XJ700WiZ1kxJmJnpt8EXMlfHK7X/aWq4QKIJi13ZOVPlkRZ57+qrcU6r8qJ8UE3epc3VsrvMZxZc
MbUaoF1v64HyYKO3lBGPjmYL8Ha8bUqu76UYB8Qrx2Lr3hjxfCxQQVHjHBE1dd8C3sJQD4JWuSoZ
wdVpwmpB6lZAeOJ50tKT6wb0VaHQWfRDYoDCyMoyXpLSMhGwPGg80Rnnx6aD4HGdQGCNyp9pthQp
S5wCOeGCf/8ZADAQG59UnhJouxUbVq3YW98UiQ/E0UXDCq4IUfT24ufnST4f65lfechdvYyZoPy6
6f1ivLk1BdM5m40KbMDQy/8F0pUmhfE4EwsPUeZRc+6/rOxjXvRAX8Jq9B3R6JRdVcviCd0Xm93s
ZCnF6IHm9w4YMOtNSY1MhnfDezUOOePYGbHRq6B/RWVGh7soVgmxs4p4pxQbhVYjBlDUtc72Qb3I
umIT8zY+/ikuLZyiavu5bN1JPFbULI0kHkdfWFVT/dsKiNhJtrlST0pQ+1gvVk/yOFvdNZm40ZXw
+dm3wRZsq7ZGBIMyPu0iCwnQ8P/olvytChhWDTKvnTl7MibkYYJeFOYwfBQnVfVViLWbW+CO9Yny
K9xNWNTgXdnwuB38e0cemBvMU0VEmIqCofet3Cbv7z5rZ6kiJHs+VzlWB8CoZJ6eTZPokw7wtoTI
OGR0mQ4RFXW6an3VM12UZ0ph6SrXkdd4kWj65Mg/9rvRMpVAXtfLfq6EXY/7LmoI9m9DKhxUI+xC
lZNz5D9onTy7YnTPaRe/nG1CzjmtQg0nxXlvqU2u6dY2771EFdr1/V43+rptQXzZewR4gIPn02q9
Od2HqO2cUdhpAwM3bdR3EoMWuvAGzFNDTKXS08y6XpIi9aPVzPSDcG5DhEWxMiTqLVX/TFAEKhCA
sQlhxEDT2aeFNX9vHj/wNVRIhkjvpImiEmPuY8vOwwxZnQXlYQymKqrtOYsJe5rScYQ/AESm/VD2
nb2nJ64nO714udvHH+MIVOR4cMlr1JpGSbZeHFSf1j2ys7uT3DuX2OBh/5aWakcOgqS7gDXmYXxD
40vf0tdwOj9sRkIh2+HOWC15WkkPocTeGgSy4mEWH4n2yOIGmeWtCOlXe7hjmK1Hjesl0JAroAlT
ZCMWTrkXYoSvYqEFLdLFgeXzL7M9ctC6vMEGitD8i0z5m9WHQnMIyp2egmShp03KnJBf598zaqck
vDlzfE3BK/BX5aEZY2tsGAqdZU39QzBSnStjXCieOCyPW7IE4lyVc251pqg2NoGS3K5uDFTROhHh
/PG8Wwy8yhotRYZdXCdCcCiwzQs7JSuUqQV6sUG3RAPL94ydAnXe5n3jqiNKhu/jE8RYLtUAXGv9
D7cHy7yazh6DLHiGix1x4ec9QZKPZsvL5UawFBnOH6bn5BpwowBbAUPOb7dSvbF44vBGb/Z2xMnY
ZHzqH+vnCZgZaptXNk40SyLQfqaY6hxQSiw3PMSitg62IaXaeSY1XxKzkVbLd8TmezHXDJBFq2Yj
uJ0q+Ty3UI1cvBSLqpS2yQz6XbcPPAhtqm9QSJvE+ssROvuzL16DHnRqimzQx1iubgOw0BKcytxl
wLTGrcpE3uVEiMIJf9MsegbR8p4K/XVxNZYx6nbIN4L2HvpD9IXBkgXTTH2P/ywAmyv0Z+bJVMiA
tO0QuOnqS+KMppDsE4fleZif+Db6PuramFM5XKfrrzKVxfAoz5qlqXggmdJaFscP/a29W1v3+GJD
Cw3BPn3lA2Ihe00YM1ZOImiYOH6nzuOzpuhK4ISygw6r1rnmPdqxl9Uyi9VuJxZcmajyH16Q3kK+
P6OJ78lt2ZR+3UzpQzlTgEx78ooAb1tYJC1mu09lt9BAaVwqxP4hRvjZOUJyy1UJYu9WgrPkDMIt
qHLToYhnwGxSi/r+EN9kcggcN9XMzEapq6jyPXYZC/XwCSkBQQILRJUQVdhius2CdasNVtL7DjAP
Fq2mIRsjvA1OzR+lkm0FQobkSuIj6gOj0BzLKkOUvBCCMWUxkVl9Y/07PNA0myJj0U9iTqJ0vAMw
NzU0Gh0VkbjW48S2TM9SRzg0BU/+ADSWUDqUZoLn+OtY0v0ysVnkaNT+Q/QVhAoOPzDxSq2wWtXF
RCUZbL+c9totvF1YoHYBIwU5DQG/8eq3NY12n47YGuPiZ6Da4xATTwYrlnbfSwjaOuawQpKIKLTk
s+pTgvMA82Hisk/NEni6Gw/s51wl3fCozTVECjK/wIcmAGcduzsqiuoj37ZWweMAHfq1Fjgqi5N8
eMiokKoGQa+qWVUAhp87jagqNdUl/6VSVAmBuz7GlS/jNbA0pPoFEH4+rsgDiiIz/tTsidMvAVVW
YfNQcHC4YB5koNkSAbb3nL68pr9xtlHbpg8LlJ6hOFo7fZowgLHD4xxIgdye6ZXLLjCkl1dMay3y
0b3aGWsVRViKNhRm/4+UMouer+Jt4BaQX070bAfsAWchna9/ucHOD09JiTnVzfyPsVFJ9QefnrdS
qPErPftsiWDUFWEZSZyqjWGOUEAE6uQs0G3cKPHKUPT7lC5MFAM0jcC3UBnBm7W+TLSwzb5ZRRAS
w1z9CpLLfQRhjtOlPslupmXg9zZIeAchNizLkKa+aAcsPgcgGxxYC9kEs35JJhHizogx3Jg946/k
xsRMMNXRtcgSuBUtvNbewiGK8+1WqIIH3kFT7KVLBa1KYY6EnqpYUlwoYNT8U94c1Ns8VyY/45xE
O1/XAriFiNQsJofxgaDAf9QPUFARzXG8SVGjOsxVBenR7xEG4ujoYvroxugOS5gQ5l3v7WPW+JZ+
PQ+sDjMgvQxD5IQrDEYTBwURlBaqhtTMpkw2ZvYAovUBVsNnHWEjnWT/L3mFHQ2iTLKOh/k2bWwE
7dZg6MyqkmMfbUFNgSZvjMyRAm/o/gvQuGtcqLQGCSR39zqTbCX4vIeJeeCoHvqOuAiKY+0k70mf
i7Cy/3Z7bN9akINq+afRDBi3FIDk4H1W8BBQ1+90EznE+HiuToHqoLi/pgoQCcTLJ3bjxFvwqro2
E0Sh9sjEuv8QcPJ/0aMFVu/9fvr3WH9uC0NB//IP+J27+JXaTAvQvN7I5uFCo6hxL9T3DVTdk1Ys
4mz3fjd/+vNyKUfZfwiJKXWg7/3dh54xIN0oFRsMx8a8h5+iU4IB2HXaP5RQL8rT+BsSRYVOwC30
nzdi14970Q2Vq+879Shmn18lc+FrWpayHEKmzuqpJtSwL8wSGOeBYfFvIFgmV7AzVJF5CCsFtje5
yECSlRPUSd6xO9+BzoLcqu7pebAb5Z6gpCzg4vFy32ZTTdRu7s9fhtdK+uYBs1yb8LYcvmrS8P49
U5S9EtGNN2nd0aTKay7LhsOylV7WmPxyfYYlKfxbIM3VW4KaQ5d5VZiDTs+qPEIOqMiXMLIessh+
eVGWJIEEUmFaDsSdBAN2ubS4orTZ2kG/6r0JzrkRPAKhjBPElZ8D7aggMdZ2iiItKMSqkuS9InZx
YZQXXjKeULVomnCwWOoSZGMNceG4tl3IeznER2tqpKPcVC0Wue0IBmIqslQIQB3kBSuFBmaowxk5
uQAQ9a8YwEDh3K9i0jE39Ue3KBFfKUSSmnEmNTOL3EH1EA/k50y+1p1uB8+crOsJX620czw0/GuE
ZaHyHsuSmoT3uBZbulweNAotl4buts0DOnuaHoCQz/Kpd4wE9laPvI2xoOdz/p6u0VYLyDg9C38H
khiuthA6fHXnzpWm3ad6EWl031lrRa9AQ4CVJALaCyZkUo79Qanwd3aDDC585DhW41cgM9jXB2Aa
rIBl4ekVMRk33yS9RL9Y4qJ4li/yaGcP5ty2+McgShmrSNTtV6sfAmSRRZVkTVepDXPjo8SbdUco
bbKCnu7+CT6yocIVTmE5nCFiK8jGQnWH9VSt6spBGfLziH3+YTUg0ln8DsOxkybOWAfHomHqoQl0
T221NVJtZv8nSkejvwXtpuLlLv0jdoSCDtbKXmhgluA/Ka/rXIpZ7fsw41bnY0PKje1TLDBp7mtc
3Ekd3OM2g2BR3Nr18+i0efrgZL+uw3/p3JYSTvS71sPvIj4jV9OULnXhMU7oD0ZPsfWWvhrflTxF
mSl0JF7TbGw6B7MwFD4Y4SPYBiH/pnKbl4kkTkaDCN8CYzj4GioQCJhdCdvgrxqnTTKqs0ctCG/n
CL+oVBCtDXerIPbafNUIcV9gRbq2bSKrRxSat4jAQC04+9wvpl/KXHw107Gz0fzTIWcgJcUm84+/
f7HdDoZ6qG0elGEd+93OjhLtddlaDeYlMRUwgZr1Uo8HaGvPU+UEKCnJTS6QpaqUlUv356bHZTcA
nGQGPVgSerB3BnqdggAYwh1bGyL/f4h+yM0oYdhzCGCSV1dpCklzrlIH5i5nk9u0SoA/WPfxvvbr
YUkEpB3PU7AdQERTijdF58Pv0uu5428UYsaohQH/INNM0wCcyBUh+vwLQ4c7LNz+bz4DQhNkXQcZ
UHERPzxQsEpOs81xdSJT6bBQ0VNyeXSgxfW7CzMtm3ZHKDQKmRN+E2xYrmRp9u1Yubs75RTFRN8H
f9t/RFw9+B10YF4E9WEZotQBlRwMnKwX7rB438nrGU5NgwGvem/3NoNsXW/jq/F0W2fPBcOonHpU
shoghu2zXWnY42cqvciGH6wN9Ss/LwaJLGtqW365/DbGkxerhDmahWnHQGX2QUribW9psIug3Eyi
LfyIcc9KFOKdTIdWlNfMitG0dky01EcZnKuutTuM79ND4mnusLeoBJ0hpgl4EG1EB6zyLEO/wlwq
F5mFebo4fdIp/+rq4ckqTm9NTLbNPTzUN3jVxws5j4eL1SQ7LmkCifdiuH0JNY0PPN05fWJSVHSR
+lzI7FQ91EW8VSy3d/B0VIWNf9Wq3uWiWNxDvyhT9wriNrVTzHNpmAMAbFlJ+Oa7dlUjnHAuGeSW
6Nn8RD04AREVxbPO0uyBPw4TT/Pg3PY8QR1YZKropPgjC3YXk8ClH4e0nMMMGDZDDBq/Q66hqmFn
mcLr1pkuwysQEIdgpwpoFBZgEJdtinTvN1L1U6yKCcveA7m7Qy7TFE2abPPxIRaGM3OnhqeA7LX8
Vw+SRF1tf9iT/IUDC06/CX0vIyaQ0LBX4vU0QFhYAbQjKBYEM5olPCHbufpNC9OgRLNB64sHAx0K
TOhpCPUFhYqpPY5BnOGDHPDlGHjvkGipDrvSm0BF4qhNObFPpHA38hH6CLgthTEIv177sG68Pzdb
XnP0y7UwqjK8njhs5dw4R1sPNOVI6q3DTZqyot01v/G27mqS/X/l1EWsTTSiUGC2D2n0dOkWs+kZ
oa2okBR6HClkoTa9cG3CPRZDrF/BO8GGU/b4keGlvrCjG2FY1GfWTONdP3qIcY6QiGhW93joJHf7
h3tgBD2paWdR3IZUU1PIDBD2PxSMeYpqLh3r5uoG/RI+jOI8NwUgFvxT+bpzMpqhXD44Y6UFsG7u
7hsZ27ntAZhNb49jIBfj5BNqPbRGkTTFv9FwRZU9rwFv2L4Zy3c6uFLdsja66TfokcElglv12w1B
XfUbbr/ypWVYx38j5CVZyyMAJ+ZM7fxIg0ewkCsrqXxR4r4DM4lGywnUzl5f9YHWvxzX37CzokPG
A5gZ7scG8w2MoepXkpI0bmfO+5IkW80tWcypw60bLOYHyg88AD8jXrdzv+eH4C5adj9ZZUFb81hs
slpmVR6F6A/6N1/qI0vMqddqbG7ut8aE2Z+QrqbmSH5ms3pWU0SaN/KOxywBulEJtEct7L2pWc84
i5730aprhsR737jclni/0AHQ1GvYSs1n253vXbQb6pPTSrpF9hg81xgeIX2m8poGLuqcVS/K/LCh
i3xpjA3IN40qOiN/7oeHtCYlimExb7x67z/DSq+rYXqruAFMun9q8KlIAiI8Rdm4Y2u4s+EwyQtH
1cZsa9HaEnuY0tcUVe0fNha20IrQlsOSIVYeUg7jmykH4SwZaeXFJPmYpMyYUAnVXV0rEQKbqwmT
qw6V5HD+/W4sGcYEdlMY+XIGXNtHjMWHK2YBmwbgrDKAmDPxStYFCQrj6z6PZvzCkErER/tp/jwc
q4zEuV3Ztn/JFHLLoqWX+8Nc3rfn0a98AxGJCy1X0YpbGUhjkLTkWH3qmsoJBe6poBncq4boFelU
bkEa7S0ducBIGFx3wfZtOfv6DLOUwbyfk2njo1SJyIX69r4hMhcWW3fGPSdBsnDX6l2Chm5TLsEv
1FtZsyPCvIcLFDBduYVIxZm6VqoktNL8vSbKY/xVJ7WeJdX1MCFJJfvIn67mEJoJ7KeriHPkm5Cg
xTfGqOrFfDil/GPdIzN1ZqBi43uNyqD5ehGyc1K/6DeEBF5iy/9LciTxJXbDk/iUJn6aZoEzN9Rw
LJ1AFaUb8jGJrPraEoRl04X4dngY7Pxz/reIUYgQDFvpaCnm2FFJpXZjxcWNWevrwA/LKDqMHqdr
mnrhbql5IND6t+TICCPzbIRpWd8Iz8YF331WgoLwFb+8KPUCroNfPrWpXcHfrcC7biAvy0tC2hs7
t8f38pWde9HMxLJj1MyWHTEPpG/g0r0T3CgbKhy0XYgYdMFhqQJHiT9ADumBYyRyCzgXBp83waOO
Lqi9uu1gC3wo6gq/FHiQWgLgeduXaFxden4qmLKtXu0TEjfO5w6AbBY0QS8RTQIjSaVJlKLzfqpJ
6/gpxDLRV8ZMNgGmg5UileHNd619BKQDW4rnljo/nxMTTixSiJEsRSQHrZ6Au/q6zHH9GilFGOeN
qia3PnHWjsB040WtfuYDkBW08oDOwQl91IHyJSGF6MrAUvpkVSZqNMEdE3tRndE6K9v6bORqPzeM
pmTyrOIWL8Q7+3+Dm4g+2MpPfqHtAQJswpdPkRw1umtHXt+fvDNEN8FD4hFhqmQSQJGnEuPh7QIV
uJKRdH8SZB7qtwij73bjXBbF5OWAngYoIJ95i7utSlyUcCgzDDGkymdGhH0OPp+5ispoI65ZrsD3
bIih20LsyyNGN3bOHorK9FgypyBU5UFfo18oSN4WN4bzVHZqk/RCSQelNDSUZ2VnT7BdNPTJ9QFZ
s48lhUGJZ5KqP7GoBGv2Qlra/ShNd3l0ejQRrCnBHl946B6UtPf53kBc7rEFgrOv+PqjVS09yNnr
67Jd+TiVW+6o2k3y/KGvRcqXhYRW9GWrY2BtMbumIamV8n+JhHZYV9k4MmJ+P7lNu+hpDrQPt4y2
0wvMMxp7l2gDNXBtoPrhn4WxGb8NNZ9ZrYzJqB0+skjs0Q57CKULKT0UCPcV4kHV33HLw7PArzxo
CWqkeajXye2FtpHqp7aNe7hrYBB1K0AreWjpY97MPSDwLkjot/lT1QPbYpO6xkCkCPKl8KcDaVia
Ir2jVgMQKJyeFHQfpmrh0AW6HXmzp5B4pBd27hV6PKPhPb+ot+ptENR5Yk9HdHuItjvqCokIuhlD
oddyXtDW2c5GFEiuXggGidatLRXSKZg9kYvtZwRWLN77AJwOryZnf6wsKEhR4W8+UUj0ammV+b9f
hjKsWeYZI+URtpTnHOEbKSUpMqGV2ytW7jX6WXTy04MQ5JXpdw1u3+xrsrPtoOJUmy7YAYjPoDMd
d1h/6LlUYWbMEeVZw5gq3ubGw1d9S2dGCg0X5bcLtMsjp2xEQRtoebwa5+WMZl8b7Jnji2+49Tfk
leXe/9wTcqtfd6nM49VhUJoMgyhxwGbbykVGrAeEyegVSsvJ1lshaNLYadEsEBVGQTuhGQv65y0X
dKECprTihlTXXll6Fk5/Z2HAaaZrLpCEHsq0NflAeXhseAlN1n0mb1en5yLOHN3cFWWLetfn2aqK
5o9RuQ5D7NCdoe4oh0NYBsMpVjCbbr7uW78Z9OAF0TlOEkYw8AjAHC7+oiuCW3gJOMsbL0FSi3NZ
BSWeggbNsCuVIC88qbhlEWctACKjr1YPO+RL0KcyvO1HGPgfuJfEGMds4oOBv/GBmi/c0T0a6C6d
acfYGCsNPHk3T4p/oeqyngCYtLcVoGrJFz6vbUCKpD0GIlg62C6AnKWzHTXl6QVRFLb2W+PQAf2d
XzEcbjcU0bXigNkImMgEceHYOQe6CvXKdzA4LouMy2bRiFF0MxqCUtAI8a2UHxolcMM4HGGfOywN
EV5Wzn8A5cdMLRJjpWVdPq4o8cB78N4QYHVCYKHlgdRTanecrkn5COMXAvO1glzTst3Hp1H/tTKr
Wj8EZOF55PCTylWOUKhUqIvv3nFjxs4DeflobRcBqUc0AGzBbyNHnjLkJO0HQHI+O/jJoTtTSSMt
8CTZI0TFAytsvMGTfEAVlemJm6tTOj9YbtQeN+HAmhKsYG2P8tKUCQ0MwQ7OqMPkF9XoMJ998O7o
rimiHhdtvsMrcjHTj5FAA79QAwkTAbqQ5GuzUkPVQLTqg6PlROTTva2HbmR+2YYhSmefSx1hmU00
qUZcjxsDsccQE7qBAU6LYePUy51ifkQWGzy0C0cd0Doi1fLtH3RxRR5I21zVbd7UHnyHW95Un4sx
25/p9SIy6lSoL0kybFRa1hQrSm3jvnyIgCSB6xYeKThzRQ13HK7kUMitWVE5cFbIiEQGvajWgMTw
F8AlE2vQZi0tAFhuiSm6ej4yF/JuPNS2yzZfLb9v04+cuZeVrgtw0Nr57ssg9nT/NfdhZXWxoK3H
F9hRPKOjn8swHMJ4DxvcmVbv8xE+0fKsA09iX/JTxnBScYlbkk+rs67BULjLzi0T2f6GztNJuwZL
Rsq0vgv2Ih5ZTCPUbSvRDR6bHu+5LIECob/QW44vmvbudOKLbUkfIzah9GsS4vtm7oOI9kKu2XoS
5oaTMTI9mWO3srSkLxgfnSCnmI4Tt7xrJB6+FNBcaZrJPOmoqP+LFbUoNLf11741VRYCXm5U5x3V
jCObkzi0Q6tOQoNQqWuPugt775EiLGMi0KgKEO1BiWZjP17TSE3AKr3q8wUba/DsuFStI7abctx7
1aQ8Mqr9Zq8lTXaNHFGU7gCEXKbjFBq/WHVkqKWAaSRWKKYnRP9y8TwELLxSJdh4xNU/7naHe2bp
jLD3+eMapRG2NB1YfvShWVb5CjI9/LanWYkzWWM8nmNlWkh4QKKCCMuu8zHeYAv71OaJp4XgLUqn
bfxh4X07hhJPTUxue/mWYHdkk8k+z5ceaOABfMkMFPyJYG5VL0pv88WbXG6wJeuuoC2kyCWFJGxE
936A3MY4NoHIRocZLMSgd4wWO/Vj8kh5v0coDdjpomqvXmLe16qLO6wo2FqXu2k0o83qmHjbtAOQ
NMAz8ajPA2TY9/DTtSDHiFbHEu30kDHoQTHvAEAuaTSDO65whdttHw43rV6O1jByRdAKEe8lq4uT
E+BGvAHVVJy4KXnBgzIQ98dE5rzaZiSisLBUAeQ3BSn6lpoy1/BMCiIEXNwc3QHmnyIIbblhXp8u
bzNGamMASZed0Y6dM1t9W341O6HVZLtcEKW8JCDiDl9iny8HK8dHo7Jd6LL5T5NZZoKVHNUpohLU
NvEYO8kg+9xEq9RRkYGdkVQhtdgOUoT+2ksBVoon2HZG/Iln9A6TFAbCqLe6OeJybksGdjMFwfvf
WRryKFh7OPmHBs7GoNnH3QWnnBoaHigTDnQ6tbQ1Xyzmi7SLBrkHZ5PCC2pjccDyzq2J/BM7sR9p
yYKHniWxT+fOZNxXNxWGYtRZ1s1X2CAmYuT5X9FqbLOv7q/GYuMw3fmJFC/ZXiKuIrPbWq19KVt2
ehah3o5SHBid6XE2yJfynpKXFEQ/kJFBezKNUdkM1p2jJfqITNjLR2uml/+C80swQ9QNJXeazzLP
nrhACauOTMNU2dztJNAVEdWu+dQLhGn/oM6DPPrKSrz30JMxSvJqifC8zYKFA87g5hHQ7c8XPuSf
VkbKQEUcIwrGtDxuwbcP0rUoPqT5Ks/kEDScizFGK4D4Mz2ii0wq9W1ee0s/p5nwq4FryL+oNjW6
rLSesJEJfjHpeHpsNhvjK58scuUnmNLIwLZIMNz6fyNpG2xJlWLcNFTt84apYwKyO/un0NFA1zbE
UdgwTxPXbhelAeBGaBHKKllm5h813qUYw2SNigXBFfzc8U8FEYFwlydwd4kynSfFe0qJUeU/8He+
mOpCwXlXj5eXam67l6724TRDFqXpnIaq5f2NMjGu7s3rM0UDINBtdiOU+O1FUbgdBU7DvKDE8k0y
i91uXr+eHGhb78bLnGNZo/3WvztxZ0zI6Xu0yZp/2HF74kPW8HE/0yydelplcQC2ClBslW+MQnNa
NdCNFOjuCdBA0AhO7TEgsLaOOcXNx73S2R9Za7SKp7YEBWQE22BULx2VJi3Gy08ANo/XG+H8js7c
RBuczlHuMkwU2BlhkGbt0G2U+I5dEOjhoq/NGfik8ygF1saI25CYgvUPImEAgIATrv8hzR8bo7dS
MczYHV4phEUSu5erRzZR/3dfGTClNdg+dwBdkds5BDcTEHXNszzergKKjAvkUh+ESKY7UKtIQoF8
utUQnNWn2fSwYcYBTFWrBbnurFLcRnXg4CDMjEjTpX4WGCz9KxIPx8llL3vWIvQ/uXEEAZPjbUPM
OlbtQRpXPyf6+FB2T+WR5mPTBv2ke3TcVXIMf8mRiazsftjf4qF2BJooeBAGDgiz+kOHvb+KmhD0
tsyXdxMd5HLQiC/uWiNjjI9eUB0tOw7DeQz7EfdZ0b+X5yfxMFnCSqJ8uYKB9iO4LlzCSg18CcEj
osXrqFBvKILPLtDDuXXhAGbxQGpMaVAaml34OCMI4g73lzsOoiArT3VPDM4seuuhkUg7eCi4V34z
ysZn0mkkNiVvqpnc5urtNaGWlzD3gb6QT/0Vk9RBF6FGmWILQYQJYxf4vWsiE3t+8F0X96E3zg0E
HFS1jaxSoscY+iOnAFF8I6Vwyfzp/yuPeB4FxpGY613b/Pk8uWBGmMeCxqDq0+gdXLgsNB6ixLlR
wItI0pvx1YE7DMTwP/SL4gysnLnloiaBFpPCaakD9ABRcqxwk6DYujDiUoE4S65OrkTP2FGrn4Kp
zM56Y4ct3bQPdLvgaQ2ApeUp3s0HZ/x1YwKV2O4yIe2OMOuLDOmbVIPv5X70pfSMNO8DPOb5qWbI
tuoRr3V6QDN/fbzCqzv0TKuSIZXNAXFO4gCr+GOKT25eEhZaS0xCyWn2thqzav5lsAmHPhQBzz6N
ZbLxen6M5bWzf9lC2HJ6P5zs8E0Pwc7wBZmEfFmU21ZMsGdLSp05uGegTY/iXZT4ptY/TK2LRlal
7YIGeqdctW37q5eKkgMSd6yN7CMjv63SZPMjXER+d/2oQoeyozj9YTLOLghnnRjCQnOB11fHr4m8
E4IvZ9q+jR6QQ8RT5x6LCYsJvzQB8lGW/et2ORVZoR3AAGKfNr96AOFVDVdSgTvh3z23F7I6K3v9
cNczQMJ/fw2Oi7HZd5Jyoo4pynLCU88A+c+mdZrVFRUfk5S3tCCNjnbj//TXY3JISWQn9RiPhYCK
+24YTGNbf4H2I2Hj94ZA2yBYdjFNcUAMj4tMz2MzPTepo6G+3kIiqAS5Eancj6F1KgdBZIJRyq8c
JpSZINZvzL0+jI4OY/VYxHcnreAQfEqQQPpjlLKsc2psRljYL61610XmtUQPkB+wvKXLz3qDqgYM
u/3uAbCJfjFEIsj3A0shTJG93TYGslw/3qIdAx+9kzlwbHyK8EmKsxOlrFl1Een7Yuwt2PUYBTgd
eCVc4NBNP5EKGlda0Ds+ye8y+zfdqe64kmT0iSvBpv1GvycoEjxP2POLQNPuIcva23bqFQ45F0tV
HNFctXNMLJjhAzFYtlc47bqFafH9CZHBjjy2urtLvcTVPB38r2MmXYqmbMYzM8UbBD+MXlIxbn0u
tWTTBkhhqefrLSkDQNGAymPq3CSPZu+xwxwitxI/RwRzuVOP9sxqmhLGxwalK8pI9/uuYwwEEskE
J28hmzkIzq8VG3GheMAYYglEb3tdVGaWLfp+G7qfCbot3OW+zEDoR1Sch1FwHZN7q8BcVm6DAbjR
oerIO4+KemZ5Zh+cnkmis41p16C0SruTN5WsV/t1RtUXRjCOMdN31nboGROJLbL6QU54b0cHMrTR
wW8vrWZqz2nF3VSAh66SdgopB2+3cl4SaSFqJ50J1kIcdLfD4aADbS0EHkofznSTy2ElyA0zJcY5
9vQKkd+sRs6kF9sgWShuPsQhArL6mWlJyNwsQvenTqG7F/gYIEF0DYmPKafG2gqRUUuaM3IlUPxI
L8/cj47CQXwDts7DZMNulMMv3DM0FWs3VOQxBmFEPT/ZhFfRyctJB+fxOJBMuB51Pao09zZVsymN
0aFoheQ3MjLpClB2ria4LjsMUjbLGsU+w/JEhTj5d6CfZcmR59UjS8womdIvCCnbYCkLhbBmgP0K
jJBi2jnd5FqGzGKJJDpZoLFpFkCCEB+xdUyAM3x3ZpaSnaKxx/T2clJjJsmYSMiLTltuCWqrK8Cx
DMrxVIxjsSRojyhtLX36kZfzDzd6sQMArGCSkDOlKFAr+2SSq7wpQm/Rg2hbm1sa6ogLk0I6VPcF
WooHDojx2HRWfZeAF6dCO9l1uAGBFHJVzMVEjSOsMKKtWH2uvQJN52V0pUD+XRmILd0EFl3d0Ors
9Q3zN5f8ae9wXnW3/yLphMt1n5Os6JwpZMFzqD9D0aFDxwOPKjHutseqX3Fd1ZFONSFEUs+DQLte
0OR5deWIzgXRjVNhdrNfpx68Fk0J3d77ge1ZDdKbbzHMyBBSVuDoyd53dr96L2YknFfeFMwGFI0t
bcsZG/fSEPuVTbtFzYCIeIkpD2lIZJ/lbg4/jSLRcE1VpsAh4sU3sAAIpFeoxejjg4I23DRcVBuU
OR1Iu7R3ML59k4m0dCWi6OaPpmJiOT0ABq9cscwbWyUB54bKNTp48H0486OIL1ur/JgBTt3AvWop
iajgtz4zJpaHZn9nzPE30OLA8xXUIHjFvSstNxlYoHUUHAFEOU5DM3t+Q3CMkQ7M8+PB2hyVSvd1
JFro1Q+8be6HyyVtfT/OYbllhYILb3jd2w/jzKKdXHyGjkh/HPTwd2EzpfwhknFyUZDdpwVbbL1d
eLJ+Ip0Cw6KswP6iXYKe6l9moYHwMwrP6KhLRlZsFFFZq9GfkWOIBSm+7axj4lerRS+NUoT1+fxS
rJKsYvi+nPgp+ozGJNrsV3iiGLGYoAPuMRfGTHoJFodi1ekn98Ph8wYo1TEAdWPKkbGhtwv9LUMa
rrbOx2YWA1Mu2KS+CdB3irtvRu/zvhdowJwJVXdQZIzJO5YGjjPgFQIyc3KatwJJYxO6TvYqGbHI
ybTA8WIT5HxGYggGIsHuzotG3kALyKuXToRl8YiLJHGQ9srLh5I7MKpiyTXTuVjjV5fRj7uUREeG
mqDCEKg2C3PexJBpNqyQu6LTRWrtZR4FZ/lZCAWrwtZsU+8uRFAEV2Y/cnscj7mr3G/9LHHUz1WZ
+8CKpPRAM9QHJYdjWQhVboaYSD/2fqj6VEsFaNvSo++VhhYED/zFszv5syKdcAGYb1xDy1ZfqgRP
u+KliXqZRNtAejwIJC9L0YenXDKVPUMIUnO4hotS+Pg1s51s7JO9lI/DyUSqA2rEIZTOOYBaNrRk
WOOxljdTpVT/6Z95DhnbOQQBvDWoEXtOf0+Kj3qhr4CVqw5loj+juZkzj8Uhyf3q01rx9scmMk85
pi57KJUigc5tqoWI2RMrnItgg9d/9qwZBFL2vaPQVGGtbHZO4BztPXu13aLUcuw8l93tliOSU12A
SR6rCpCzQgDRPye8mclzNMCqcloXym9dHvcZAgjs9TnjkSdsd3ySmISZtb0AMg5jCUthnmE2geK+
px5OOheBFEIwCrkFTuIDOSirXLpqHW7Suu/NALOXqe8aM9Spqf4UlJ9NdiGI577H/qpCOC2f7VZP
v2b5K8XdoQqW23OgFrr7V+vrdiHI7TQTftBcCZrGgubIZvgmhO+KJ9uz3+pK+xXE4r/uOPI8LK5i
diDxECkujKJIYPD+Ll7NpBJgVTzJGWzxzsZYGDzJtBFTW6r41SgzlFRYQ3NGLL6cZgUxu8Qdfy41
6jaKAG8BBWgZexnGOFcn4HJOE4fnFcLsCvfbxEXBUCLwUvhHbIm0OkObhak9WHGh0tLmmX/OjduP
2t5se4//i3au7Z5j6z12ypT7rY7zBTgbTMYfwdRyyZF0B6jelAhggYmXHjm+LvIknWBUqz1C+Svb
5zcyf87cdw9PQZubbC1KsEfMWi6vjcfXNQ4jpsNi7YrZUSPpGtGlb6FuP1roU8nEBlPDhiY3tyAN
6EdbBBTKzm0GpBFbY1mSKV1yUqHM7Obon1yjldRUVTTeXHjIX5kf7qCLgXOxXfB3slwVoEd0Ho9f
lufHnAU+dIKqKzAmcWOz9RjzUoauN/ty75/LQC+X7uFoRUrQAxZe01/WNgegLk6jvy3RRFbyh+Fj
aDc9ttiio5UF2j8QKZFH+qw3k0D9eMrG/P1vbz+NFLHsmUj8/OAEeuU5msSfXxUjN2RSLC/1pCKh
HEd2pJFKw4N/gdo+awuIuS4F+VRpP+35A1cR+7uaJ/0RXCXFshBPav2LYK+gvOkIgj8nIPX0KNnF
jkgAKm/5oEO8xZkAqZYAfX0oVcxk3YPLxSoI7k4XrNh26/C1LgkuOIwsEseduW+dWSb6zBXzfSKN
xa0IQacWLGismZLLdcOYusYDTxGRt4AOGmxstn6PWdRtv5+BnonhS/0oHHITpExegIQmCVUH8z7X
VDtrQTy0NSsixbt69YF86iQ+ftucMNfHtP/OmAN7zhEc8htgQa4gTEMNW8rqRZYb2R4AQ1oTAiHQ
hmdJf4qpRO+JmkzsY/GPsaL/B/PcR24DlYFDwkK4xxD7MEi6gJNgZVDHAd6lte+TPdM881afzKMP
1F5xOa7dIi6cIvKqbCIZZCjhDBQgDUEtcvogwSveD/+ThnUFo74i+3ijzCCh7AIgqSiUu8QMSHrw
MirjZ1Oh5GYnFEuXl6vJKzK225zoTrYy01zqdSBmqXlkZPA1Jv/T0FHSzMMD5q13A75B7CCvzZA4
ELJbmfBHtuNEDSqY2RIFJiwQGloX83DH8vG4i8bNWXVIrOM+WTZfsCGTgrmCXVKKT2+tfZSBgk5H
1LWq3AK+3HWHqz8E1FM8EBi5JBW3BbahJwKHjdFkEr7lnmiXCHZnqVeMQ6CTMjK/r+4ockjUL48r
9Xjn1bnBWGFsf+q3F6h8r9s2PK7Q2Ksf7LQ91G88aSEbhS1e6aBvuR81K7gdPhVBohfbA3r+tfgy
xDwVUzob3RWv9AKCN3QWl6nRAgKoKVvQkTMQmd+OuGaCuEzAAjXbdDPXOC8hxiHHPHLHpCt5Qnsd
5pb2WSbeOEfpV20b/xqDOC/sx7Jbrxpigzv53NewYdV5Iic1subu6qEmtpBo08Tv6ljX6w/k0Msz
KDo1C3+ZZMnIvbjYZEkz5rh4aafq3zB3jrwCrrmcGv+YpRG6/hoOTUpHD65sWVuhQe7ieb3AGWFr
0C9jD7lMa+RbugKht2hSIguRi9csAUR8tgyogsGR0jFQgk+C2hx2fk+CcOOWJ1zjDdc2Pg5GS3HZ
25U23FtV1fTP9V4GW/HrZ30nk68eROpNxChpxoso+Dd1sIysPSeXoJHbOStdK+H+kuUJJQsl0cfJ
G5NUeDDGMkYObcOCaMm5RH16eXVWdA2sY/s9TPaJZQPHMV3mNwcjIxTRAb3CGfbiHXxVTSZak3BN
YQcOJZ5X0FOXiZ++v6xxtZFYnEQgUhlh2vkELtAKmg6Jp2Q3GgDxwOonbwZHuvWWLIGEETAQlLxo
1yQ6j9q+pcSvt5b0plTrzGAeRPRBBB4VZy07CaGwV6dcXz2AjfEW1U2CIN9JVNr4P127n90tchaz
U1/q+wLZRcL7eq7852kRoCcbEPuSPM6Ql8ZnLb//VPegAnVqURJC+kGS+uGS6shSRGAXwRZL5mlY
JhAhBYam/ZGPbOtF3SsDeZ1qAV5XwH8KN19bVGCgWiG7te2dc3fpB92/FSHDxZSSDG0SeHG0U3wP
lKW7UVVLY3B6rR+AkRCMAI5Img3F1fkZxXwymD8iurMF4DAD1ViM1PA5b6RT4J+GLD7741GJJRCX
atayL+xQYdLw7vGb/0mvzATpbKiFCL97xKsOYOiMpPcNtRT5dSAJDbRYkWYAHLQcH63fUWhK7ewk
aXdrOzVWOpTG1e5UqsF9qjBzNgoVROA0oJBYPUgxjYPsrEux81eHseGb1+5UabPs9dtZkHSrHxAK
ILAt/faNFBMF/Ul1sv9AAuwNyA7Ox46fXtl6YuV13rEQucAV86GZOvoSTaU7FBG8jltJEwOVI+mE
r0wTg+lu+8V/S8LRCx7s+t7k0b59CNHXbRj0w8+XF/1KoIDz15ofrnQFrMWf5c4bFE8fMPklEWNX
i1c6rK49O19xpRDYZVEVAbdrkYqDDutBJebZP5ynSEoYJgQRhjPD32vxCD48PORrCVqQpL6/2Zl1
LsETDgBiLklbbLuLGX39NJozfoiPPyWOB2kVQRtlDxcme4Hsa0WjUieXqSHZqY9g/NDNPu2LfAZS
q6Yzzak3rAXAwGdls6mxcVzFLDtWa92WRuDo+tzJPvjdhdDAC7NCQW3sjkO4p6z6U0EdcBQju2Ok
rYoibl7zzf/KB3R5TGGep36M9snuEozOepfuEg5Wby5VdeshI5QO14oz5gURKEJ3BGakJ2rtSua6
Q5jDEbmKDD6uKlOIjfXHbtljeNzUbv7LUsgDwDvCSkE+Ts95aq8kzoPTuaIuUySzpeDBYB1jwfD3
RYSsgATFTFawwVHCwOLlKm8eyo7BPxgMcNMm3BBfeveIPwgqrC24lrqdxccKwx9q4MmhORh7Rx/Z
p+8SwIFH2SOQtOLycBoDyU0v8NodDeDsxAr6lN6vWNp/vdrl+SagpcoqN4OBuAD/7+9xHMmmUIe7
pWxs6n5JdBYxhMOH69q8lz9L6AkG+aLZSFb4kB2bU39KAp35glnGZEDZWaSs0IWl7Dbuq5dqzSce
/P/KgT/fnABjQLlFy3cf3cVFW2/H2TmEp99fIBiy672EkNZJ3zkqaXtTKJMh1Lrz//eaNDYajEWF
FYzO69gGyfjn6dQuQME87mJf30WUYHoBmcs4vju6gD485ESY6zqKr0KdJBmPbUEBxutW/2aXsXxp
1C5EFGDfrxCmvhkd1Cu0tgvWT3GFsxfnnX60j4k9C9o24f3n2+F0QLYgPh6RPj3KhbH/Ze7ln9/y
gNoEpGtpTxKNWzXSf6phT80S10LLS6CzXwmWRdyTyr41i2ipty4b0boPYby7vPRhh/tdJRJASlhX
nvztQE5I7mcEMqmGikdw/SlArMrEwwXa/5DQLcRlu8wpC1LOW7x+84MK1QHcVjts1N8tDdLMKSD9
W23EwfPz7Io0wzYKFnRSVBD0cNe3o1Z8RwXq7Row9Fpx1wBzrekMYSXLQf2n8hVscR5NcFU8RV95
pc/89OTesR427plL+27t8qM954JSlxLL/LvGqdssYk+QsxNDUKwy0HwWASSVqITvy1pkDtLCeB7Q
GZQRTpdMcnV4UCFnkrcfLpStsWmbCd6ZS39sNFI6D2eJtffNRxQ4B11esg/XMHXgo2NVb7S/owW0
+vYNVe6CH5TigSOw/EwF/bwS9z/TucrWAK2cZMigZJaiNIp0ZPWdPZmdAvkRCpLhaBYMK59boKOq
qjhsmoiR/GbGliV9o+nB7JaPLejDVndZpKZErKat2QuljxB3twefdl2649qkhQHZdatheH/+VkLJ
trOhMCcmH837ESQ/NpRXmziqbVXml4SBYnudocfWE0y3xI+ECWTInUW7LHAuEZYcqZQbUJyuR/JD
xGdEzCeG9bl+Io90jxf67WPPBIQ3djfZgxzL1unhVEdSNEOGLCvSi1DcTMEHX06sJrmJxygunfRm
etpIdSifk4BkUq6DR8BRAtY+UuoPLv2E2me9pPNUAVdoH3LdnZpKHmWVWyfN0zGP13AjInqc9I68
u1Ciw3SER+k/UoJEOQhm4i4MKW/lt7atr2NbGzoJq4P9ieBaY5BSWmuZ3WKzomTDZiFTS7GECKbc
iel+P8i35Iy9wFYgQSj0UfNk05UOyWRfPlMC8Ww1c/zZGklG1QRTjbb9HmlxyfbJPMePPdOC0y6D
98JM+HWIJsCz4zo7JHATy0ho70FIO+zPFJRpBWOvOX1I+QKwOuek/OFYbU5uXd3oQc6SUXtqECnM
y8Ajj2PytaphVkYRcW1GZQiDsHbfVLdsohWIr+0v8tEXifTGVMD4aotBCMSO2KES/XIKGPzl72xy
gbFYum6KPZmfhN3JTlYbvxfOulhvRb81s0EM5U0xH8zfy6MaEHan3MjHbDnNoBu770vjn+ncZipN
8rkg6WKNPnJ2cs979HjDltvifIyC27+uDn6m9v1lJylRucuB/FN8pfkJ9dRxhVHjARDcuNCODtWv
7E2iXiw4oWXt3EuKsDL9xWvHLQIoqXX4v0s+S35cl1oT+tA+XkdiHgLhJL96EFIfUb0yR35c1WW8
4/Gmzjohq2+Y6Ioj0ih01YoIytc69vJbj5YQuPBzZ5OuSUuR1ItoY02Ai5mHJLwDfHRdMPZXXFup
mR0l5PpVSpeOfXYxxT/hQN0CR6IPOMVFgQTvKaI50WgBdMh1xRcWEXJWaBb08IhkG4RfSLX1oe4I
An0WaOFas0HLemZr/Maj1i4m0LWM5YJ8P6NwbtKwmkfl+OmvcqFGLepRwXAWJSVxeVAgNj2Q81xL
ekn/bnkrxyRvNQwgXIFMq46uTz8KEDnyP4TRXE/UWrVIDrM/4nge6XjSDT0Zin4T0QPECYvf5nfj
e+cEEog5TBsZuXKFhMgelJB3RN2icHwNfAVBrbpDdT60VybMvIhlFjJIAGCKzVr7fg/JIZ3Q0h5q
+/14nBLVK74vXWl8tY3+scrtlNr3Hct7duGdmxM3vpXFieDad6rNnsdtWfULDNp5eFkUvamlsKsn
93PlWkco4yGKepW7+7nUMymTjEPkMdArTjyagedU0ZBQe0aWpP7M1gIwREv8y+pFqeA51cuQHlJ3
UIvC+tSmp1fh4EhyINXvCju3VkGN1/vEdpRjzdM7y5TMxAL4xWqeKYUQ42E+MmSmN+RqB+hErIYn
ysqyMdpjcY1oHE+8Zd5+LDy9l7xu/CQI6xZVGbP8VgwF2J0st1jXvYIH13ohdzd2ITVjn+4AWLbG
NwL7IfERf/Zk4Tt6iDJFFiG+HZXswnejAp6pn87Awh17GC46+Z6G0lIH8gywBeBTjj6VOSYK/qnJ
mP6z9xhyZfuxuTh5OFP/MXXpK8BwI9PPDocf6kAV+CK2sj1Rb1+sltaSMBi8dBB+cfdiSXGHHVUi
Jw66YA0Tutobap5SdIjWZ654ttpOjIeRes3bfNoz1H80HB7Z5MdhNknWdhXe3eryKVk3cRCHc3zU
P8ZYSa9z5MKMxhvOVfUdq02QxgsZiFLjBM4Z7LzMyXkpFuEHx+zwiGdb0DOgFQIfVpBsV19sR+S3
d7rU4bL5eZIRDcZopE7zzOSi6LdLDlh3LiYx/gRWwroYlYL8qF8My06WilV+FWzr8JifuhYVBy3D
vedbbuuXyY2UpL+cnIVdE6XSRDrNvDIy4xUclvlqc3Ji8+kOdGrk8NftCqPntQJT+IAfRtJsg1e/
aGW6UYj7JquAe53A2ntyTYfii95eb77T8RPtpCqtvDv7WUv7lkxyDLjD3RiRhZgdAmyDhaeRHQqi
kU/rC8zhLULr9fGaZcGuZg/djFsd/XJdF+gc7rQ2n33W6CduP6D70l2i9Cmz39xKVCwfo+U4kVFF
HMKliK2cCuPDC6BDvTmI0KmiOyCSqRZMKTAvsCAPgGVr70f/bEaCryBdQALSq5wwoH3FICB4IlfX
/FgJW5D+i0OfGAxb0v5WMLNOjgEb4oSWYboJX1n11ieTMN5QR/9ZR3NozaQjzWV1ZjCNyoHDbkG4
ZCRAZAFXsPyqHETaKUAOozLbyG4+w8KMAi844RFB4JGaGiuHdmkcyKVw3vpsvU015x50E9sp82MJ
KTXfewByLFimJQKDfnv8GjOCTflLa7AD+GTMfww/prwK2dQOwvnE9VYu2uSyZUAwNJADHKfIOQLX
QzgoCUlll1XM/UqsmLyBEu82Q0q8qrBYOjVJAerTtGkWBxVIyjr9stZTO2mWGwD/4WzVmpNBiDoG
pBJX3mDGp5MIZjADnnddlR6JDM5DY/myJsNtEnnrYkleG8L+Vd1GhbJDaAJCYcpkCjQMfTju6Kqs
ag8v/kOpzvQokpMtpml8B5WnaLNbP2jbVZ6vDGjmnVc5iSe3x4MX+9WvfXUUhjuIJKW/Zv9LvOFf
dVx8+XdnV1bR72p1zQfN7tPv83g8nB9UimXNRnipwE/NtuVfTFiOyhhdTOucIIJ5AyxyloNm5iKv
W1Wt7/Pe7HnV0xky1fn56AMjWnYYBPBa36a1mrWGSDLVHz3NCH/oguMdKkzw4Q5x91r7Qe1jEa+m
EpA9WpkML/RJ82a3pC14x/w/CjBKZqg/IYXAaXTkJtoq7HW6Wqv8X+zT32FFfqXXifUM4JYXGiRm
4VXhqi/Jg3Qi2KVtufdWqUw1mFITKoT1QsDxqimLBMjlAQyENzJYOPMW8t1lwCIuOKujjn0IGwtw
4JuGCJXI9KaDcVB0QGc8G78LPfdDBnGJge0gtz2oOv+pftgNJE200Y9KcCjOMp00T7oPjGIU5XKM
wLynlUK1S/oUt3bFDqUc/WO38y7XV/uSec6qluLh53tXYuvM09fnQYFpFzo/RvdvH2svN2FJsULA
JzrznA8iqGQn9uL0W7r1MioLJPO7albCsuH+s+d8LYPj8GLKVCfHY4gzLQ9SJwla3sMeIvj2aG0l
kwTjsVLhsGli1gciEo25Lvo3MNDJ5u6DtXMvTURFPHn69bq//U0MyfpNVR4woFWvNHh8vr2jxTCr
drY6iaXvFpTrKKjBzbRGN+v5T4rWPazxinxmK6DWM4rjCFZ0wahWiUoornhxkvwPDi8yOwN1/y2t
fWbdDS1TlhQNiNcSgdpY/neG+xz2j3Y+/P7rsQCs2mdq4WPWtLlIlrDwyNWzUpPVNdTbeV62hdj8
BK7ZvnGcHcymP3XmLcvC1yGNuY7RmFrpXcaKOVQyGEdPPt6KOPrGcdoRnUQruVgBD7xr994msgsi
4mzNVx25cExAR8Pw56DD8keV5qsBavYRRUC+Fi3PYNrECHiFRMpzzlBipctysu9Jzs7D/sL6HwKH
tFFjbE5Z7YO21sAss+c6gdP+j76CCoPSkAMoVGUd9Y8ZhWh63s1YIbrZg5vh6kDh8yBmDpFnagG4
tZGGffS1esyNU4z9wtwNZo7wL0xZITUDtN3ukRMSl4MvC2LhP1PBzSGPjqLM6PaeyFvSGexe5SGP
3JxiO7fPDiV1wHL/uaftZrwmytCjcV9kANEDoRPRWq0blyElNe7JUdELjUecCyn75Vfe4JzYdrs0
Mw8CNNlYYKrIG8Eded8k6gpSQ6OY/UjG+t+i3x6Sf1YffAD44+G2giU9i9MpFLsaREAhRBrhONW5
oB3mtZmVuY3+2iASy+DptJY8u8VVeeXMsCY92zXJllo3muJNRcF9LJsZeY/Sl29yho9D5VTgVkWi
e/6FA/G+RRe3qlEeJP38BG6qSY94eqjMjZ9AiLhaZO0bVPKk+9rf04i+q08RupUUxzvARTPxEB7r
P9iCxW/pM8hRvycAyFhMR+ZJvKDbGzLXQv9iVS/cYIiMQNTUdjZI1ksbh487XieC6EPxm9AVy6qj
1homqjHVODoLrqnXmlUCHEab2KHBBwkJOtE+rulaZOkqGCSihCUipKXKwgy5ak20MOABseb5W9PX
XLQjxCiMdOGk9lyIRPN2alBMi9q2tVPXd2WwD5SIuhuAozavYU3d4dB1PMtyO4L8wWGzhorMaffg
RyZDHw3D3bTPWFlONTxo0lRsFhq0kl3QQJq9pebqZJc8EMlkPXJ3sw5DeIBG6aftGIZOdtL79Db2
7AHUQEMEOyduO5g7qn9VI31Ra+AjHkQmYynaTpotFcU6KpdFivzfR4jO5ED4vSjgpWj1/T9IMo4T
I6NYmDiyBcWdmWT5Vyh+QK9Rj3urDCp+5QjnYQ8/TC5VspqnD3zRh/DeqwJwBJgeDh4dP8xsGvK/
W7ZJewpHbqEN+rVY1qo3P/kwuVTMaWrAM5TpkUHO+j4/PTa1nnkf5KzHD2p7aGrBQv+0BHBmjw3b
3D11yIQwEvA9eEn01ZTHahloKyIiCyTw1ZWzb4qsQsSQ3pByIoqZgBG5cPCOjrAJKRr77ruFhHyG
+dipgDwcYOl4Wv1Mn6U9FfpMQQ/mgc50EAv+76UZRmrYs7mjMtJlcZ1oCRtBuB5O1hdqkJHaEO52
WD7gzTCn97TTpweVLXqUOzwdSY8dz22LuoWc/DuKsn0p5CvnbgbRF6K9UUB2Fi4W4IzQSmV5F4pQ
kaafthKDRXFQNVGX2JJlBqjFqeyRmiWLK2Vl9YXRxUW025CE3X1Ee2diqcUmxr1TH+M1dZMedKlX
0OLTchz8XqZSk4Mt1rq+GodKziuHRB7JL+/nvODm7fS3nlbikjAuGVeoOP9FUOVthM0DUNwjVD2p
yFHDSEziTh9+LVqD1UFbVtT/U0TV7zFNZCjj0bxZAiXKtqAJ4Q3Z4pjGMieOQ0m9HXW7MjgqLTlm
N9AM8nOHoW+sOiqeT1jjIuDoxSqZyHaRmZFuJciPk3z3jQrmhDMUkYinZziwvVDYCZ7aMXe6eHkW
hjQqJMz6JsbnrNWPOU9mTKiYnx3jdqZt4CGj9zdVG/LnpcSKWRUctmeRJKmYba0N8g7QmFIcMOkY
7hJBAGIoQg4E7EO5SghIJERMl1szRZrwMozkF4oXz6k3EvBkKTGuSJjyZ3eBghg6HlTHRS9pz6gg
EPxoaJvLTNiLUPjOKkVxfF9ciFCJykMEL6byrv/ki00DWBk1qah1qr/pVlw+wHuj5UYaRIVb193R
cqXPhfuKzWHkZTsK88SDt9fTFLJGOXAjpOgnlTOWQkO+uzxxMeUCcArcs9VkVi2/nEc1NVmGvvHJ
Tyl2h+rIyggkzAVBfpxtWQISQDRaTOqbFtwSpamk2Y+4dYGSk8ca3XyvcYyif4Cs30u81Y/b/bZx
iGwqoD4eBCUAkr1iWL/fF2QFif9+d0aXkq+B5iS3LWRA52gFtLJ7h1Eimr06NUCB4QTkAvlQBHZr
maVNMQ8NnHeF0sXy38Tg/v2zuSlE2+E5p5YAzs8xSMA23CEgcNk7TDvamojTa+5APug6HFtdHCRX
T7YMcGlLbY8dFHQO0Rg9LZLNYkT6ukogE6bUjRjlsToHJM/pdDXOo/3fsvUCL/UoWRLAj0Vt3KPB
ICB+idf6+xORFtqvAsN9AjzS6wzfF7/oi77r9oLhQ4Gf1UPZF4kkS1iG8+EvF0DIm6/nECSvKDfZ
bf4Y8uis86aFoTRmUa2IOHq0Rb9AOLp8iGBsScGyqTAK1aZW17z1qPD3faWdPfIrtq8vuoWLb2wI
3D38BC+1VNnXUk+u7JmEc+ifnCDsXJ+pItyhbMI3Mjk0S2d9h1c1XFdc3zi8iYDFw1+W/e8wrCIv
3ujT7re8x/eiGSWERKq2YdvRJAhhqPZ90hS7NhEnoueZb31RidHwEgJgP/2nEsZxoa0wwVCf7pGS
ptH8MuOcGSGqYLj3GLrGBFMwCODnYyfoRgxyRi12zI6Dfm/gwWI1XRlULY8m50n6p7LcMfEpREFT
HuTKPFKwN+zPEmr0ApYebEZiNUp0fkxKDJRU28MHxc+3IX3OZqIkZcWIDFS8iX75MoXGEEVetL2j
KQhJ5NxmWK+rm1ZMYt/YTstInKTHZSR6lmnVbDe2TEZGq6kSvnrLn1fuvG5gJbXvutG2MAVA5FzX
8gnXD+unj7rpcAcrfHOd4mMCusiIoZ2Nm44oYtaCsfZN1ouX5MYEWXO4V+nkku9OWaMw7+XqNDFD
KuFkZCMg2ee5eEH+1lutUCkO+OY745o3bEw/pIHtLjlDNdjIAB4a73tWsdcB/+ibVU1IQmP1qUem
cfwvI9MQjC0ijMfHR5TqvrQwJfdvI8vdnR9mpKCHMcss7OqAWh5hDlZbcq2+SDeNTx3Lplt7iiuA
wMoibH4qOsbUVM2EnzPFxUp833z3+K0+GbO586pm2QLlMjRoU/Tw8f/rQMG8Mmk2/1x4wFPFepNi
sJJaPNvuSp5Rw4du+V++T5J/f2JsvaX3+kD3ERNH/J75wOcerVFQTiSqKtTKK4rBD5mJqQv2Zli9
lbJJTFuXAKYo8cI3Ss9pZQB+omo4R7BQJYhIewIbZZ1INTqkQV5Ns50ztGj1XhNXEWUPrnJjK20d
P8m4Fy6d9IbTQgz0v9oJXDbxZWREjn/Pue5NWx1I4vYzZbHbb0zIyyVBk+huM2/Tg9uAuMOtuwAg
QCsWBK9WY38I9Fmz4BIMmetl3wAzg1j9wuiq/8UjSRsU0Ij3iUHItSqwTOhn/cJnBGkkCyvssFBg
bBBbf+eiwn5F6Ea3TaiUObILxRTMbb2LAKldhHnSAb3LDaCw8EYESKri821xk+QYPAgVB/Bmqpvg
znzgGNCC1mqR+qhxfhpQ2R4GuF9EThvN2n8PPtTKutH3rXKpXAgmGkW3NUxb02WOYBRyxh1+insN
bY3yzzk21H3bNkHFQMKpm/k9hlp1XydmTYqkwBO+a8g7Q229ncvdpueG8J0NxOU8miJbXDnpLzP/
GcD2xH7cGsvd+mpl/MPxpSyLcQQehXqp1rVc1WyRYSPrB6M0ievWimAt5mG5tVOS/sS2RhePbXHR
n1CAP0pJuKUL4WvzKqJN+WxG93sgKfunEc2Kb1UMRm1j+KbW4BS0HEqn3ywbrJV069lzKxQFV7bZ
LGHdPZmO7FtczKjeQi20ohoWjPUPKRxza2qpyxT/HOn8lHrTvbeYzY24pA32MdKmaCzxGYCZh7YQ
rLobW6b4zIoNg9HVw0IP/9rxTUpIbOX27a/4DQ9T5GG9ezHu6vHE6H+rXt5qnDDcgDKnGketSd4V
kE3YPeEtbvW0mhApiKoVAt12NEchxgb5Bsu2+Q9W+emmPL3jbW5zi3wd+CchVFmeNocY31w9wIu8
d5oZcdfnsRfhCFaqO6CUoHgbTVkQjCOXJWqRUbN0RbBdeWSUj5ER+84ug2qh/JnNeKUDQdS47pM2
Fmk0HlOWYf0lA7yMLEGYKYKJrmBIEPgDXHzHwArJswHnJWx7DEunlnHLZjmiEmK3DcTthWuVewDC
p0Pmqrpg45zAx0VYRwdNMB/U9l0M4Kc93sS/UKJpnDt0sLJ8ckykmtmSeCzY+J32ZipxnQmxT+il
9MIQWlC63CbFmB1f5uWn9Miuhcmyvk4Fevan5rIchV7r7+xDcFZu7KZPP3TXAcBjt8rhqIqr62Uo
qYzz3OAf4RY6eCJGj/e1/ncZEI1NK7fW1jQAvMHu7rfuY5PMQ29zUL9rJtLukbKSk/dxS8kSbY6D
5n3Nj1RgcQEz+egxX0att05CMaz20nC7MvG53HzjFSPeQmdyBy1My1MkjXdL4rK3LQVj2ODSm3cZ
QAwEtCw+x9yN59oPbVr6Ul+wFiTjGVbXAUvbd2Ovf6kKYgm5LQ8PyrG1uJ9aR/5ymgTZ/yxZPFyV
RXKd+4VkpoIoFZWrTwXIAdAA/hlWnQkdeygRHh9oCbCYjoQz3UUnVGdkFjOcALXfK9+v5HOQvFr5
Kt50YgTiHjFxF4JO59/IfYp170xz8PK0gOvN1a4zhju5mB4Vy5N1+3C8771TPmh2M6TkBVGoSvT9
QnNGsW6VEfK7p2aAoLJ0Uhz3666nguwpEQI4YmzAaOkd71nTOa2UgwhEAtxdzh/Fc8cHvyFWOg7n
IIecEvhRYeHAbjS2crxsgRI1Nb1G7ILLJl8O7xy+BNPJ6Dlm6exDwP9fs9dKTHYcWD97arXaroqR
ueBUTS5hOe85+HE2qmt6ExQOCxXd5zTq46gtrYlYh79M7n7gtxiQ38JtYZ06WX6/ArIbpKyNhH3B
RT6HMy3DvbEcxng1aYmR0dSdvY4urJVtoPwip432K87GxGuRjyY9cQQk4JVnWdDLMc7J4F+IOXp7
ZfsmOLgX7LEKLOMTE8Mto0WKOcv0UGI2vBx4tK2rt5X9EkKDA54//sPyYs2WbCF/mvy19twm93So
dlUwTcqpjG8kSvEDx9n7E9cB2Gr4ZVhBtaHXq81BjteG13n0sKVK3IUGaUVA9qGXUarmCEN5W9wh
5dw5QP8L7cEGqUZ1ZvNVxtzVpTbNnCFdcXOsvkblnJbRtkVquYArncTz9Vh3VOIHnoIEBDcrEyVF
RcniRT352YgRzHXUEpTKljB/DLWUogZd6Yj0Cxp36JdNOgAzaxRK/NvecB+H2WqI5pvZkBb0v0aB
dwl2L7N4+zH/yWYCIoYEb2NXaFs7zvNjpAKnLcNuD8JVSy/FM/+zsl2f2/DzW90vSKW2bOSmF21q
TRpXOJs8dLKGueQeMR7y2nouv8UXcPes75zVfh/hyMgKYlJa5LbbPMuVXF00xzNyXcu3gND90+4i
1+w2MtMjW4RChwFvRFST9UpJScWc7K8CO5eY10kdABgrRfXWnVdwZRVPAeikLHUdSXxuQ12enVV7
0B6tXi0CchoNTxrgq1r6YL13Fw/CInQTUKA5VCqlN1fqtXt15G/RZa5ql+b/5SubXum4V/IvxVLO
qnu3EVghJb3k+Eu6iD9fk9v1ovu6BQBhKWiyslS2plLdiut10g8UDHZKJQ0E9tyoCpJ5arSCA423
tkMkmJeLUWv2xTYoJDXsTykzKouFg9FTXWQn0jNEDoHdsgxXANB4zfQsuBxD/NcecnfrHx/NXT3t
6SGQwG7/fMdzVvEPo29BPwbCIhPTAnZJ1Z4HdMOc/8dpTQ0zQNbx1lNhOxjdYkI+Oila9e0A73RV
OC5jfQ1a/o/3BzDOtGl24+udS0RHAgHntytCq93FmzSj+xx/n9RgoKTI1Zhw7duOef8A80XTND85
Jb5/w3a3QDP0pXd47NnwAl5iW56rtemikw+qWCdYU6l3Yq1FrpuH/RIEqH6uqV26NA895jrw/4Kc
tRePIZAG4EEZjN36TZpNBE3hSRh9xRKZtH3KPwwkvtzWFJjCgijhvs27opwQ+mNkJiWnTBmTuPQi
YhpVcBa5jrckY8VHNh7cWUNNqBko2O2FZXNTzzGFt45Hj/rt0K46HPl0x1faxYktFlDJRnr7Aj5i
YsqCSKegKSvycogQ9MOPrv+Nu5/Lrkf5XnWSgkgK93t1skO6wt9celOeAZRyB6GF3yhYyDvlBkx7
ve2HIHB13xwPJfPsa+Wb0VBY9GG7IwneC1JCzgNbKy6AMosunY4SZjZZLfmKpcr8xPF2Plz60KkV
VrHnhKDmBZ7rMcsb2xuuNq2db8yLg66fzU8kgJHOwQz+ixJtsykAT/+jPbOrStksrzROWsMs+CKZ
xtyZz77JU8Q7I07ITjgcJ2rIyGzizCHWmwbrSQNobHN8+dGBPslfZMFlRyKnpXurPMjqQYs+zj/q
/x2a/xF4eAjahLH6P8B0tC6zgomf5+2wspBQbF2UB4l9lCAmlDEZtJOMa16qXoDWbCgEqfZtS6bT
vWWOQJzbEE4k93R0htNVBBuEv++FSc9G45rYBgkUD/vy07oXUnyzKdZan2SmYYZwIWSewwa5+Ose
3dLmLwaCrLmn7uZLgXdoVWyTtuzITtd0xwXTRfQ8M8AwZT2z2T3JoSIgBFCsOnsSR2YUVeicqG0k
iR4+wgMCJqYc4l2EDK1WolFuSmC+2ffeUTbfKkpnAfzZnRllEaxG0kACXpPDQ5HIvuusF7X+x/S6
LPj0JpMa9+VT/HddWKE52VQFmqn/L4GWRWuZNsnfU/QVzpcGt8ZCQigjcukNTu8hYcUu0Q7Q4ZtP
+Da8uMMT3+TDgi7j393DHfBAQTnK+h1PBRM3uCKu3RAf3yaTJXicYAFeldrZmzfDakXsFMO0xyGM
lWdDSwZuTpSkvKzeKI0GFV0Q9b7XupCUDVfgFQwDlLcaoWlimkKBBq7AULiyOZPedtPWdo1ukkL1
d1e63/HB7P/BONqn/Y2pIDiKUvC2ZAq1auj/RUYNp9Iws7GOW5Sdvjae5I8Pe9Tew3lUbHtBte0L
g2RzgBPriyuEGXA7qXfirH0rmcCZ3YAp5JFsxFsyKOjT7XCw0P4rnMMJSB+HNqUmmc5UJuYUi7t6
cmk0LrDXoUYyZbWCZqxDu2bVDPj8iHSE8CPkF/TNUMPLhn8KkxbkwBC7+0k3Xpn2MkexX5djhTgr
4FMb8C93ma/Al2jqiy7hb2+aBzAjARfpBU8LGeWJA+BqV1vXTfhtTVLNsW4UbZ71seSvvjj75DwB
6rJPp41RfPs3udogBaPi6cnKLBI2Ny1VwNsVp+AjkGucfsOgC+sVqSWMw1n1FZ/+evrUI/5oUNDk
29HxPKomk04aLWyPIGrh4fBhEXbuuNlnnHHiAKpDvWjTF4bsYmZ1cK4RYKt35KOCpfpHbikWqku1
X6Kpj+TuhBNsrGNia9rc8OBROOr1AtXyB97SlQfRNDEuDVyQQww7PJykC4TWWybdNlDKUHZi5Jht
pg06SjVW+hyus7ZHAKGS1B8x6N2d9q5KdzDZrSLGu3JJTmIJRdhzlckaZ3xKCwR453CSpO+xZuii
+QKLqxjPxo/CO3fqaQlwOSy9XMukjN9X5LgBX6X6L6DN9KeahVGhDqJJ/80UuMtj5YHfe1I6FwB5
EM/lpweBlHLJTrWhPvi/Qxjrcz98qGAq7YuYo3W+oSnTBrjxNVOUYbnqveKnkRTm0rgPZ0+X76Ho
P7NTVEERUo4FGC3Gl7pT+ms1nK22xUNfqVl41SAl+EFlyqHlSfZY+sxFMjqiGwkzoX4tWBLrprdw
2gFzgyTrcv4oiZP6xR55iJAWHGOjzbGB0eY8n1yrzsgER4bXHnsLxSSoPvyaBsKD/vW/S3IZA0nl
PPUCjVdJ5ihRxatNOXQd3D4b4UVhgKlSUGWztb0A4gFKsycbDbi/FhkVfW4IsFLjUjlAaOZ4/eGD
iml/uozas8+iKSIGALyHWFJ+TlwzhAvIwAk1S4ac8vT0CcggjVJZPeAm/OsnJ5sMkiX2NtV8dB0D
8VYgPQIYqY/iJFq5+vCsceZjb6vtSfF6fj7Moy0D/5+BrXhnfaUmxO1Z/HI34h/lcBWzxCWcBDUz
Jp6xbA29iFAAtUM7rcGvgPiGi+eCjIkvN4Gxj5ObCQFiD9bm7bb6YjUq/C5v++zfi5ppI1aUOKtS
sVpuyyUDNACBvjwOx4H/J8Y+Ajh20VY9fbIHlhB0la2Gpsdna0xW78bvrLLAPhMXEYWqxiVMPrNY
ZY99mFARdNTjSqAz0RFEB0UqS3D1WEB+p73C/oF7nepauCSM1pS6MdRimO6v4pfJlfems99Q+l7B
O0B9ErXo/Zf53ScXuTu4E85pUNeqacpWC16PBUzd9fBHQBHIgZ6/2Fqft2StjXWAj7rz3CWcRxNO
78ODuxtqEIJ4DBjD/WFU8FVNBoiIo8Hfmrko7MmBMpdx0/53k3B413oFNXB3whFiuV1dvfexFQft
Te39acs1VYIC2uAMSTTgpcFw0I+1tM2bJYXO7L1zmaVt5Tk4PGG5qx3MQ1BwWojnwjs8PIoaeYDI
XhHRvCaKjL9yB3htY0auXLlOKoYoLEackZnecnkHycCDmYX26zGgiWGf8fIVezW9ndTW57u2IfuL
X7o1SrQoks/bqyGQ44GHWQ6UcLy2u6XLs9KUJ5QMtefqWmnh5jAE5y2gGMk60BhGcBIxuQVtanNX
dEw3HsCeqsyNJ6rVSya4OJXVuYQX2lHmSIBxgRi4kD648AGKb/LXRvd2xgWHzF3AasIj7zm81Fhf
QHy5x1k88VZl0OvDK+wRgZPF/IvaGJCLtsoXbEnnAJ5pUayVU6GDazB1QEHhHjtjj0aCxxy66q+2
MPtxm6Vp4glZzHiwO5miwzqvpbFEvXHwHheDpQEOgEHt3B7AeXyJy3qZQG3bp2yCf354T5cgQ/s/
spZ3NJ+FKVrIY7y0TKsNFY9lTFfdBVRzF6LhIEFVt9W8gsmNdzctcsKTshPr62+L6IA2GlL6v+wh
vRqVzrva2N93D3ygDqEB4688I3R4N3tJakP5uptuU0WVcakpcYwwHQIdxBgVUPrillnv+DA+29Ru
FDiX2FFM0RTdFOff7h5ZJrPJYzGAF1wfprHBOO4aVKeThojRjoirvWsmMVEykBMVj672ZploWb/c
i3lXC7zeaq8k3slMy5xmr0878G8rnQFIeRe1aaSg3Rlo539g9xzJ+ELpfoqv1KfMTzwovAlRk7DN
5A+6HqhOvFFDRS5lJhveGOpvBR+1XpMH+GqW4d5DvuTfMmfBpy87SJcr8D8Ih2fGTqRsxGryMqNK
Rp+WG2ZoPMJ6pMFhIJGbZtiMFSRmQdmceppuGEybSWyWZKZ9op85Ly8DmnmMl7GBr7Cy1fmYd/Sp
hxO72WGHNukgD74iUdLxySjei895/1UkYgAut73oDzaZ0YswQqvxaKFIbavhe0wUUKOHKcgeQ2/N
j9PEBRn1QmduFyTMXw+UroDs3qpuzyHXXWvSUO2r99Qxd+WqBN673IGi+cqcBydFsNdbALsPu0Nb
OBXpt0U1HjlvZAuZO0il5sLT6/iqAQAI84Kf9nxo4KgiqAhGr8M0iGmA6qal4I21uTZ/4DXvmqNj
qAmnWvsJJzD1gb08+wQzwRBEdpyWxd4QXnoDR2nVvzY6Kqk88st99zlnm7ghHYUpxIALvAYi+paz
i5cSyP5m2O2d2UTlPwKxOTC1eZpaAiSg6rtj1m0jgPSVOE0JpMMKCc3wgRJaDXQS3LiIGWvVZ4TW
XKmqceejDze71/A/7jzJ3H0UfXVxDt5LQu+MAPj4BWrYtlNUeYb+HTDAfosMBY80Kz97gWCXTtdu
spvQuM3mqwvquyRpDSmI1rbn2m4h5MVRr+S7IIwnP/gZxy4I212nuaD2JNPewVt4cDDv7T8IHHyi
97bDL7Jp1FhQ/13/Xq9G33Ul0AMffY7pg7HHnn3yrshh6lE4N1O0LyKF0JbWIZ/MjBoq5zrXxSdU
p6GWCzWUMC8lhbWqzdpBW33P7eRvS92g7AM2W/x9BwEHm0ioLdIw0ZJIKjM8f5LgdNxUhGcjeWdb
2njdrqX994lHX9T/9NNWp2yL6Vyq3H5zm10QpLfFZSiqM07QhXwTif8pIWfur/DB0HZrOZFDXNAf
On6Z/7Q58SQhvsdiiKxAXdsUWs0kpPEbXQh5ZC3WPUdkActF2yFfWfPhXW8XVM7oVSZaW6rn5boh
R0kEZ5OdKPLvjq2bJQhg+xtGKLncpiozyB3iHSgZh8QQ/UQ+YycKO29Ah32nRoyjoLRz/SqdWzWZ
gtX1fv6r+xgtk/UeIzqIKc+VGitU09WAhGeH5WLHlI5fDrOFv6U5DEduc2oKvubc7wP3HV9u/+vr
pLP5z7UG/JZ1nVXeHaAfpC2KUubdqVs8Dkr1pDqMNX6WGWW2aN6mO8b2z82FN0kWJSBo9ESkYG6V
k7XY29Uijfd1hycGCuY6XC12HHGR60IExt9Evl+9MN8Xjb1S0OjAAcWApossv8i9RFEsZPh9OjOe
LYTHWKXiyy3SNjn6WeUhicgSgx1LOQdalgAD7HPrmHk+Snxee7p+U8YyAETOZqRXuZ8jbzqROVbA
hXUlzQTAuVlW9cWpHjc3s9akAw+Gdn3iRHC//EQc/GppWsdlSDOkhhIhYTZeJzORJnm4YOgSbuhX
0NnIVCxirUzvmTDyIdg/lgA+mq0w2pCKiNMImL8quTm1Y3/Hak7FEe0cvzjECNyJQmWw2ZFGN0WY
ULFbXdyAnRB84sVGAJHoFpnOMRNznQF2vQ3riEsd+8pemUVXjh0F2JJm8W+pVFEgvmFY1LrY8zDP
okNIUEUKWRIXjZe6Ck1CIvo/v+alXM52CEEMtpNCDKdOs9D+Ghkv8dba+tkiD7YQeco0vRJYElQG
WCT5tMENhzBmYweVnLbzluv2E+jTukLh65D3+JG2JJQbvTtZPsiFGU1E5limoR73L41nuER0e3QX
TwSK6KMp3xoNIyBSxjPGmt57IOlHlnmbfdmUheXM3HONof9Syv9uY2WTr6McXHaHFChhWhijQSaf
gJJnVqSsPCYS9IIrTJAWuqpGIMZbjQo3TdtiqHsAMX1uU/3kq+MtK0uMAtBoybnoSMRBhz1hSKM/
UrUTPrZ3ZEBp5lZNcHY9wq4VJnYL7BeiAPAVX19xp37QVgD5qdbWQaFK0vKb5ZP1dLUsQpJ0Ljnp
38YUqC+myzFjXtO7P1MJ5X63+Je1ZL4usHt9Wpyx4Kjolh1tdeFaH69wq0DnpPQAJuAm7lksKIrR
W51d3fp97EuxBCJHl+ViCaJachY4lgD0Z5tC+YmlztQhPZ1SFuxV/7RX7QAdK50LwxWqU3fheFZo
4xXc1YF+z1m8MynAYMy6I9cZu+awDbSDVhvF+TxVdsXwglux7/RN2ZbkkA5gMg5zwsIaLndUXfCH
E6GOaQenL9MrXNNXElqokFMePX8Bz/zHYLSw8oWj15L4+mXcQTGqVJKeaYIsLkNqjRcXs/tN0tgq
/s49yuUHoWER2jGP2bgUUZcQqDcskkCGxdRKJrxTzWtfC74HrtwGhYuaD/jV5D4spSF/y0Cr+48y
+B3GtCAyoKVFsXM+DZCsIvjD4cBBeUOWIPUbNh+lXb8Sv2ZWtqTDhfe/P7IG43e1Y+MbqN7iScDn
ur4nd6ACJypbC8QoS6FaIaVRR0caZwFYqInQE1KeLk5Fyh76hV9nSfUQriV1/4EIJWxGZcvukbvq
mewdFTuoUZrKP+eOSbZdWjz2cOyhumykf2gW6Fmt3TTUEht+IvuMlQ+WpZs9R9qbEpxDnUuVdh9v
gcMgX71gkt24aHpBDjQUrPMZPXYvJt5odob3pFyM8eeZH7jWTXrWNXhMCSkrozniU77mA93sarpf
neqrmHFC7V6sw3aOoywoOJid0FXQkrEcxQoPHAxCcpactC3Plhjo0LXx1Tf7KqKDE/C2hJp46q5P
ZR4P4H2AmVGsiPpIvTizd6F3iV9NIubhZ222m1krkYCV0PtKarTEVOEH12qKsT5cD5UOIve/0z85
yZXbZSHZSQTVPMQss6k1LBmzTGkvOnipyPEMisKCXMgipR2Ou8XAidnfK0Am/IbCpZB/OiPH2VjO
+rmlHPv3Qzn7uJ4GQNHmV1f2goElwn95IgIuHBGrrc2GAuF2Y2hJTsLuYDwEq8wtQS4rEeoc83ee
0hRaMkTTcMFcQNdS28YlSNwPZSX87/XRxUP1FxG+AP87YdYv/scP1ftiLP+JLqCaJ+Wh1e8mpawl
OCr9s271XxqyyyWmeGO5Qpuwhnn2/FOaX7bjfLX4Xlt0Q/BWjrv6OCphHDNA1Zb+MG9l/dGBddFA
fzLDSpnHvYWfCLwRK3B2rydX3VzqtFyGUYSvVUcjk0DGekB/yhF51H6C774MP4dbu7phFuBBR5pd
P5EKRDg40CKqukuCRwNyz2lc5DlHPkkkKfHLJrkmevxtT309zZA7amgIv+nCe90MNB6MDhvXfuHs
REjXHCZDUSpHwrGJ1yIqTxY0kYqiwL5CZsniV18AJF62gqn2Aj46kWBbqbULxKOnsG2tm8p0mQto
MioxpmZEqD/nm8JYKnZyh80LnFi1vJ5++QQd2E5+8egEQEZRL6sFo3EDcfztyqGWatwkZN/u979+
+hNnaFHowY1gdqMhqXIygMSYdcjOx4maqjOTbH0aPo34FFZQq05Fgr8tH3AkodDZqH94DhuYVayT
73jjLjZNj1bsqeey++P/B8hKWMlXt5AVYdrEcx23GPI68zChK3UYjrLP+A2ReMRBWVuQDGql5/AW
8tvNXW0PVNF197K2WUgB3FL1wwd+uhrv7k5BZsoNeAPbyhOh6rmSd7As3kfciJxNeBjLI37a5DjQ
AxJizyL1frSoRVdWc0mpLWmDcMsTwG1flGvcHaa5TeeVRXByVBZihMDKpSoKagJ59CHVcmUHmvfh
3qXkuMr7XV4HdE07tYxZjBpOwsKKIdL/TN9aUl0d1HM5J2eio5aua++sSRhhKuBAS7w2vcRvbM6E
lFXWK+aOPzymCA3EvdrFlZ/nJ2xHLOBOwhU/HVhKmz/INPGECfXaQA2Vp4U0leW2kCK9ECGFhu6O
hvgjRMvbZFcyiPox+nMMQa8e/Tmp53vU3Fx1UdmVbyJPvLIhBGvX/fCwZUIV+KW6oavIWDan2g/4
8R0z5MBPKMO18+QvPuvIzQeLm8JZayGFg5HZRFalTUbPNBRuctCs3eIK+Y3LoiyIkcqhMZLCE160
acVu4TNv1334tKib5khv2r1M8ErKyAweLuBrRA1eu4/RBxQSXr8n8IcNfXe9ijMHdii6HdVlvKkn
A9CNvWVF3xMXHvLP/E+JTwxoZYTGBnSQj0buXti5jcmie7dr4Xhv7bl76n//A60yuIOHZv+KEWSN
OcayxD5F098tkML7RbOmlXlu1aCQG2BMgbCr/eh2/VU0JFRA/r+rUx8BFZT+P3EurxqqwUfqXx8S
+HI/hh9wA0avR2Q1PMHz+Cc+wVJW7ejB6taES6RClSeuEPlNUj/iSEWbWW+VqD9BARPbxmd5znud
jSSUUjKZ/glPvfQ2yT1yr6AvTV4jPAMBVJJ+5Hwo9y6ZVEZzWzD46+mqNG4IPYVNE/kiPcbULUoy
BqFW+hl2woq+NeTrAcViT75oUF989xR4Hjca8bkLmeQurdKR5IYKRgRm81crpGDwFmsaZYpWZunT
YYYyRjm6BI3iDoSLsOQet3MKkk5REjWW4Mo1lntudu1IQR2vfY/8ZvLTs9WCTJ+2oK3jd1wRlqIf
jK2D2P6G3drQuTaq9Hc8/Aa4YiTnqh+qtLjbsM8fIQR2BXXHgGctzoGSp5BazVzgH00u8fHR79he
pSzmHAyKxNajcQa1e8tTzpQLecctMvSw932TKklK1xuCWHlegc/xktS1MVhES8BoVcc0WUHCBhzu
ozWlxgNwWcEYdMg4G0ZMKchJV82/eYsMZhTNeEUyQzdtIYbsIVWaREQVrNahwnuHoon4NRzZ/5ss
/AMVvAfph+49fSVOeKqS7Ol+eUBhGvOyZazaRs+dQyFzqv5XCgiWmG8mbgh+v1ZKTAZzcAYuI2yX
GXmsjOGgicv4M5Qc92RYfk26vegxdkA+QLdq7+dCOPfWMAuM8GeAGpFHPvVMmMkpR6BJzqXgFwNo
Lrbg/BJIfo8uJt4uea5G18TAgdtfxUII/66h6dalDA/wGPbtbJ7cMhXAnMgGan9TKFUQLpXoGEOt
T5NGsQHyM1XMBt094RjzIUNpnj0rkuvYcnfGrbLTVZs3xtzTjWqyvQ2u+lq23C0clR8xMXbOPvkx
q/ie+1GCrALf1uhxgfPyyBE/g5IJIgK5MogVkOaeXUN6l8WEJI/iR6TzhatOU7ls57ABGdk7iLJz
UJDNB54ECK+SN+DmPY3CjLIwV/8NtEbDIZeXfYxQQQlZsmUEtowd1NMmjLhwo+Y9GAASDOY1szVK
z5WeMcbvx96CBwr1YIZXrkAUs5ANnfZG7Lna21ngS5DiXN0oCzs++t7OIs+PjmUI6BzSP6jDN/uv
Y+G27Zh7qu+Nj5e4TcYOHWTvsDEnetZQmH8yGnNs7cVuUOaftSpFmetBpeqOsLeYYfCKE7kmh4lS
ePZsrfm/7otzhu8xyRfBp0zPOHQh5+mX20h752PbnIJffreOFpL0gVxwYsxJQjxC1tHBPlKNiZQB
SBpnJacs5yVt4jgo5maQ/Rze7LS1gjMlK+BSWT3mVwraYaHNWlpTRl4dk/7nybQiMJRmC5WBJSRY
apPYDIAws01mcCWra4Tk3iZqKVbE8Cv+3hF5PVd2+beU3xIiazQ4HBZsgRaCij8zryxsLQa57FH9
IzFtS5kmwyMKRVZ4avf6fBLiztxPzSw/5hyv+EwTEmhHi+Knde1YlEEIfMTYS/9xx+MYrVtBLdMf
VoOoOcUpBF/wvIIb9rEPpuDghoKj22nO7SJdkQZl+jr+NjxN7szvs/qpGUCAOGMwasYqBHvgiaby
L4NdUPVSVIynwiKhAP7J8gzgNdmsIJmK/+HXW/D9g4pSmIUhFjMdWp1QYRk/vrWs2DMXnfwB1PxG
u8giDgQjHVT56FTCrnmjqhg5OZPk3GsgTjT8oa27Blc2/AM+gShzQveGBOU3vr+E24EyGetBcofD
ylwfENimIF9Diov7L4Jwwt6a7UaCJwcyBqzs05thsUeeXS5qaYQ5l2gmCaabTKTsf0FGz21Nbkqy
WjPX9j4wIyfYyigGAfog8iJGzp/fWxjWnxTFIGQA7dDAs6ckaccu3aPsQlyJ7ilv/UgQFXhC8jkg
Di3kt2seWmbqx9Y6ccBQnyH4mBmep/U/nMSsiHBQFm/cEFMsd/TM/8iD6RE2uL+GdIniEmHWL/vy
64/bDxTIBCVfXnKNDahAjBtxO0VKXf+F/f3+UfZpACgcBxsZS7sCci8yRA6PdejYAhWFKm6KAkVY
+jYHLK13wMEhnMlpJfWoNlXGa+9tpyfgNRAgeHl9AH38wwUBJc7zJZ3lKPk5FqnB4bNHU9N9pH4Y
aydcCFHkFd7qfjFAJ8m8w605hLsQhgVm3fQivosmnAqklJZifP+GrxytJbJ0gesVwwhl3THohEJt
PXOK7PiJtM8foEauHeIDfgsIQXkFfCU7v4j20IVL085HWJgSFQt+X0bajLHI90sPhVL903BClTZk
MiQRQ1BZ9FBMRAvcBL6cDhAL5GZJrSQblPefTU9HCu46OXZs7oyjtxm1kuVmRaGIQU1+uV1ZOZuU
0JZCbuBQufUDIm9fFX2CWZNOoV8KO1jIECYCsxqsko9lcmAf41gunopNP8EVRZvllhJuUjYCVKP2
8W7EK6OQn7ok9AsXoAglf72NXVQH8zUUj/bCnSl+dVYuP9OKerjaUZfeyNUTOWlDmmJ8330XpsxW
Jdf7Qob1OOFRhY6gq0NlAJKTQrp4Y3UA1i7kWflnrGDR66EYlg3zm6qmBcUsCBo8tkEzfPUJcwiR
H4itsxz7FgomjrhKSTkKwMYUdEMBKDffqrnId82DnZ46e383VXiArmYXaugVuA7sV8JCm0CUmM7d
kkXH8p40yPbe50Ai4+YauIGkblbrbBYuJeyLnDo99h9qskg8pPoDH5tigxXwmtIH5LEuYsjLTU/b
xbEOCOqD+LgJowLeRxpbfV6Fev0aY9y2v9Jic4EaS2McAfETwPEPATt2Giubapild+n2f5SX7vi0
Ezmu6GQw2IAtfH7iwZSp8NY3TVGX5Dt6+nwGp67cLeXmX3aS8PNhjkSaDjFO4iw98uQbrYhZ5lIS
gL+iyK8+KWLhlDRV3XNgyybU3NmFB1mnFZoFrXEYgMVTuNOo+wF8R3gMy7bOU75p1CCK0Sh/f/Pd
mvW83WPOcG1zhldEHJ61OpBjpOsx/HdRVoslOG+SOlV5JAli4xjZL3GCAzHQ4bBgKwRG/MwdHeDg
IPj7ficJMxIe1cMwxpoBk12qk9BMmgzIn7FKuU+JHz1TtTgUA0HmeFV0oMxZa2vgbHX/RyM8axD9
84LE/AzFjjV8jvAjLmjUWLmPWZPgLSQwMDfBpi2t89A5UIZMSEGXc6NW1+xo08OI6EEBu0WV5N80
c+Eq8AjAN95CYyVDJpEJBPfcK/B+qVA0lxbau72IToPFlTy7ow5upxv2lacFGp52QZUUG8fc91gS
IQ8WoaO5J5nzsNZOC0gjqqJHk1rfeWojrZK6xWoNTDkYyalPMohDu0WBzsRj9lbn593BVG6b1KMn
GR3SBxrpKbmksznhq60s6EPTIBZ88Y6pOx3IDunUWbsd2URoTiwQJAspHpdwgXmSv6oi74qFVYvw
X99TaCqAmDk73smYeOhHcmRS5X4LYdIeum0yvol1ZRmRs5igRGG1LML2nfBPiQYAyF/Uo8RXny8t
BQFT0RyiOJ6ss8EuJ/V3JVtOtgA4Gs9uqcRT8mQCps+wYjuQJCaAmmpC9wibFhf+KlXWYuoHSPFP
uP/+5J3isCNd24C999WIlYWmrmfTZ192/e7AFxWNhrgf2yYggILuMR90uKLSd8+Rz4/lY9szVXL/
s3UiJWHD9HGHkM5ahjr41OMp/LLPh0JYavdkveKo8XTL3CWGIzjq18jhW113MQRB+Zj9lT1BIyHN
BzDXWjBjNRB831vLLbOzQRwDRhlIwQRlNt03wezaG4YZJP963u5iT0c8VopyTKOh2shabvBQezoS
wtdOKkT2Oy0ozye77v1Lr2FmKkRIMVAgWV1jpmHC3gE8SH2xBEJb7l5Mzh3FgMHPQGgW9AXizAyQ
TXyk+SekQ8tX/02mxOdedynDx97eFwWPwcehb5QsDyGT4IxKzlhdY/98asjt5qejN0EVMdORZpLf
dSIQa2Hv+zxlfYDneelO5eZKSneOJTQBCmwOkDp5/ejBZw0JStvtZjOdW9iAjMbmYP7rNqV0bSC2
mJL7vBi2schlYCw2SEiopTo1F+3pTc8a8Yu4sZzKfpMrJ3Il2vqBexWfyeOzQlK7f2JA6UYaMYkw
zDX4SszldLxHgu43xyc4c46HNnWCJOlRz1C15wjg4AqIIyn0hW3f3mP5uuBbBiBJjOXiGOSCq2mL
MDUnPwK5hBLVVT5lKD9g04inljRwZbMKYKy07vM/xwoEepo4+MiU3ogMKCEfH/CzZMiuVylczO4W
RS6qk9mtWofcp2IwiPOgsf9Iegp/VbgAeY4hSoyXMpeHlOXyGNDrZU7+J6iHT0ktsSuiO9X7u42n
Ck2djBPMfU3INMJb+hNCfzAkGzrjJUpUNeUdy4P/Zw5oNrs6v603Gzm5diMUwBsqJzmswzm/qItA
eJq9fucQaxPyVk2s4njlpFQFK6BiQdPsAiiFQ84KS3lF5g9EAOyLzdglLS09y39JKwaZroVAFX3V
FP5oAPpaC23BtGH6P+V5eE9hWjR0/8A4K1FcZfn80rswe3Us+VD5MHI7jq0pnDIp3I7ADR4lUet6
ZcjZ4oS+Dtva1iPuEJvuL4qawWVCCnnqs6uL1nXKQD0cUkK0TGd8iFOYo6a3o41rkPtLEMCqlXEu
TV1z2fC4ZtOGPrPDVfABOsbtmRFjU8x6W7zwUsm837m/VxNvKiqw8NxsJkGcy0qL/ubNM6mY3gVb
JMmY8vJxMDcj9tPQGfrDZlIRz5THpFdi+shEbtWH5JY+6wNxsAAVglio0gmVYhlglPQswqbkENx2
2+nIXbeDMeEZo0chwoDBN3vsnfMY3d1cNfH+4nwc+jOIwX5etDR+qq8BIiHJOhgQLNgiTRdO0hsX
80PTydIRm332TauYuk+bLoJuct5kknNHnR+rPPsrn3EXhHWnNxfCiPgtquvmG/4xlnlkie5SIpB1
jwba1zX9mPXu+W+MhLStOQhkWEglOCGyHzMtV4TPclKWwC6WCw5K57yEzTHnC/Oj3+V4vljbsMHe
c4zDgDoEH16OhAJh39FJ5K0GaPrlzvI0mBVKqC9/rUSy6XNpXk1WP2QPcbHgz3f8yv8xIm+dqRrM
DfbSNS6Qb73KBW7TAZNL/99Xonm2fNxdN0HBxbP/vVThXSIz8tiGs6QbgbDey/NGv4HyJ9JqivQz
zHwoD824rXrekLHsECWo8ML0payJY8K6y2r+ylhHpKr4ZIw+bIxOUHr9n5Vjmw6YW4nH2xu89db7
a5fmah445pU6382urmCTOalWOkphfPs6zeZYTLH/T1hlKUH34LBzleTkZDQamUyy49Pb8DiSeYTg
0aFxvy6fJRXMXS4ivjplXvAgvNNN+jgQQACRRrBStcnq0bCtXQBBMpS/iRGmSFDjz9EUxQ96j0+Z
5CX+YYkFpiL72JjuliDJGv26sPbnxlmbXrJ/XEJBh+XZZ7T/FjRmenRawL+AtEvMjgKtfgp+JJSU
dKRSd1asevcDXnJkgSxhi6XEgaDeuDKsUB7qcCrOQYHi1loH9cTPoPCZHDyrHuzyoJxzfM0U9WEG
9ps4kk0nnFSx1eQ4Zc2se9NUu62/ngdSbwilsLG4QkPAqomxxHE27/Qu+iGjoWU/9Jn7BpSPVplk
bSdhM/6TZtedC/24R/3U7w+UtoJDsaIN914OxY2F1Fe9oo4yILCW/1dU08yq8MIbpHBzb1YTzKRu
N91n3QezeqsqrmiPkPa9sH0JyaLa8n9tGYa5ipKam1Kh3aXv8xQMvbkU01TuMb+ugcM6WHAPSobJ
J/mDZ3AbJMYF+5e3v7VGGZCSrwP9R4FJ8yszZ1prWnFcC2iZrPFLXKST/eRIiS0ZDTpyS7184rss
NFQk5bY1yh2f/ypwnDvsvv3C6QPh391Ej5asBOYq0bDdnqStRVdQR39Itjs6FWBBA1y+TBM+1m8T
/25UK3C/dehWnAl/5mGU/CjKG3a5j4b7si2Dlz0HdEd8VG2SYhJmOLL7gGkWtBBLRRkAkw4oZYqm
xsenwiRwzGtPQwCJKK0HP6ogUrxvZepI5EOY2UzjmR8x6IVkDcqnhPryAymTVTHt95rm89qlogER
MsYM82g6FPXYVRIdoaRgoBi2bLkPS7XIE+pU0pUhw0aB5q9y3XD6lEUVTwGg5Hkpv73zUHzdrtVw
uklDXGjuUXfJO5QaLDPHRQCS93URLNLRKqEkNhCastlcZD5J8mzWlpfT0hnKw27QOdiGM7437w6T
2vWMDCvNHrpNdLlZQqJJ7a/YnFCEfX7FJh24GKE+T6lifMBeKdI9DIK3fA168G578sq8Q3rkvtH4
MvpZWnj1yIje8ykhnHQlpGugOreCjKoNjY6noDK0X8vCHrcPH/FyxmRc9jjyxeD7VaTxZ5BnYBW+
HTzrZz60iKU5rlDXO8XZ5nKB+x8eWw38cKMDj0bPoHI7ImEu6RWiiiwvTdMMJHBiS7ZuyNxGGavi
y/5y3Hd/JR4l567LglJCnZbizKQcRBRy6PZ9+R+YlNYRe8RBz+hPt0/P0/H5c6nJ2ItmKP+50hYV
4rHKXef/uXz7+K6nKwVwkIg3o55JGr0FsGHMRo5sMdRWb6M3sOAeGwFI5+IdmA4UlyhvPQHosHjJ
DgUT8DjZIJL7+/FN+IPMO6RtQnjViOfZ0c3LYPQSbhU0Yu+ViQFbGvjHKc2fhOMp2i4S77cvQSAn
5ZsvAFaqzhwx8aTsZJoS2invfM12ZVlbOAqgUkrh6BUa8ukQRblJlhi73eLRiXAfmltJSrqmyH6C
Mdyna0l+SVl520YI+sfRHzfE3qVmSldlCTG4qkczWhlXVfDqXTHPVwCAS02zzfVDBTRnfAwh0Kp2
thSIFKtY53vz0r+xTIxbieA9N63JZ6l2QokxNj5aP/xFHKCGkjZbM/DgD5w82D7nwCjyllseUgce
r+12UCkVo5Spvs5Tu/DE9OUHYwjvr58CQrCKhgKBKsuJBA1dvo3DMbvvEJEED/vHnazfdzXwHUkI
EIriFDDMbY+Gf80lirtqfUXNvM6EsVbBSiypBvy+p42iW8Wci3CtmZ3tQe8aL9K4Qpisgx0bJ0Vj
mRivLHKVMoXv53QgBczUTj5U2Bwx8eNjfzm5jlmf5DwAjTU8XZqN9TVDsEeXj6ZlCnGMDPwpZTNz
iePPNHB6BboUO73lYmaBALGWi5Gb783VnOnqD0w/jH2SJvK0yXQpVrkvxF1Ls72jew0pdVZsn2rW
Wtcc6AEC0MSM9oIPX6n0JW7jSdtBV6AeaqtleqOEFjxl++vE8DX+4nHmqpKp/S2lYyFERZ7pDTO8
IYKr+/u2wr4zBJ1gFfrE45zpVJ1irzocF33mC/mTaQ0vnVMfXgvtoxed9YHsB39ElHN5ndNPl8wr
tZsCVYrLGXO7PWNsO7RwIFC4KdZ8cFE9xDVaZpoAuN+rc1+zMFsWaIwui2u77iCkcFiCkeSHe0Sv
2V+NLYAHMpymbjZC2taZhbDhDIMg5OP9xOWmi7WGZYMOBsLf8UjrjlxA+Tr9SUTniVnozl7HJrgx
xDGA7kF7tRTgnMFveQMbAqgeA1PbevlWuRqC3pNGEZLG+7pWxyGW7ksCLJYsNwICL3gCaZ+Pd88t
R7olq30vPLK4kHxtFzsKvwoXi/QAcqAgBW8eLCBVcm0hg6tuFOdKCGQ8E4It8DSEAFOq+/GCbgJc
6FFBUjygQ6BbH9RVtmO+PSmOsbvy+UJiqwwp1RZVp8DqodzFHKXddQC0sfR4YVt+1wng//CiyF20
64DzwY9WSLI11R/S+4SaEV2lM5/vs3o+8Vze9uGy6eylmZ4+hctwv8Yz6IBGty1ASWXkPF2Go2tn
nCU8e1EoqB/tIgRIxEbxlX9Fyj16YKn9mFvpNU9bFyN31zxE1qkVw3uO7vKs0ySWChF8ngp1VMkk
W6RoZT/z4LSmdpY5wyRLeu0B1b7lbjW4rCkKohTwEGYO9cp+vleKHMFLoXA1G4UELl3nxRRV3znK
2/7lhNYmS+ODHpKKXEnUbARDuabymYZwhIEaqXFrocN7zesgEIuyvNprzSGOHf0RU9y1UEwKvn9o
eDaailfC0CAy335M5kl5lQwZ2U9+Own+GnVFIM3lp3FYJ8ELuquKm1fT0EgUQIS2EbuNzg5HUMgD
3Al+BjrtIHYNZE/fxjyyYa5OWuSgmn4o9HlDmuWfprqbS3blDseh7sMfdwur5NvgdQvv1koCBegb
C8IBSZS2snXwzy6ru9+NKZjtSRf5+AvAXZiPAVENBRPNMflntu4e/nUIY3OdmKGTalyPwixWIiva
C2X+9jeFKkhhN3ssgy5c4MQuKNsqMp2HVEmueqTObkbJlRlakuTtcwNi3ip+3clAjZpr+gz7tkNK
7UdNggi+QaTExKVGtnNJNGf3mQAToTekuEgM6byRNwVfCrA42egTGyW/e7UXET0qp0nIG/aDqnnE
IVmeyRoB9Q/5Tv07ZHelJ71eKV+uwHzF2LnHIaaVgEuj0oJkqoriF22o6qP5QCDUpIWl9NhfnV4F
I5p+63YVJu45FmYUy5e+FjJpD23FZ0HmkNwO9IE+KmytB26GYEZkuVB9ASzGOZlYxpoWCYV0bRTa
+xQu+RAgBBt9e4dSb2Jlh2MaBwdsDCFJGL1cu+NSZ9t6bP1S3p/lnvVFLIjAdArbGWCjo/BaXVQn
btASkClt8PKF3uLhEQ/3T0nitK0v+AZYCOrecUdcdmRjxZ3Bwze7O8WqxEGpA6mumBg3xlXVmFfH
9Q6vdfTpHf1uzVoIiJJXY2u4YffZQ/BJFjfNMUHj8mus1F2beSc1+9fKxwlLpsr4yE56R5X82V2Y
G98KXpC81U3fIIDU26vwAxrWmsq3lYLFL1MLwWn3gKG08DbVk3OGr4P+hIAUkG5pvdQ3fgHC6T5T
nSdvrKpEhPRXukNvRuu4FBGb7kl7CWifQ68AHEMnxi8vK+W1vzGhqWHowLjV27iU+htvSv8ZNZNd
ZoEkoYdFwKky9IZIjVCTjr+ztrIPsOmTFgThrbtWcYS8S9LaLyDUutcczKxAuwh29TRMfHqdd8ID
W9Ia6SkPWHfbsKno8vAUcuBM6aHhxPEOMUwcYuBsE0YH9COJlTSnTJ+Ub+tJH/9De0xxuk2GJX4E
l9X4indMVZtxHnAq6CskACYh/47kv0/eUDxYZ5PCDp7+iTsAZ4bgbxNyOwqdpI0KCe12CfvnLITR
b3v/90l0TJ8oaCmfIjrjhxg7jj0L6wl06KajMwUkEnB+31TLeB4sm30w4bmYeadWQ7yqPq4Njfk/
zeX3Hl3RZ4mCZNUY5fk7UHnN3PVQUA59V5yPnhAiYJ0xhy1kQaJdqklY2h+z0mhQV4KHkfgshFLX
5i6qlwcTnPy001BNPtqaPjrXgbzYCgtxwD80RLaFznEhpo0Q80KIHc3aj1xS/lB6G5S+zVkWdo0h
3xjr64AukT3YZDcO5WM7X6O5X/s2zYqg+/bobJLiB6n3o3NkXQSYef64mD3KlbHFT3RnmDtz2IsG
6vKpfANlrt9cgt32UDuwjlFKi1wcAZYv7B1ufNdssKEuYnWrawZvAYEcVto5Xeorq74ogv4Ms4zw
codCxcNm5LyPJ24m5fPTU7byPrxe6kdqclBmRg2J+LRw70xF1XtzHATyYkXtzahi2BXs/kj6Kup6
yUCyIMZVph6sw6pF4Esj25LLiODk4X8ppzYCHpFpNBFBKmDIPH8SGG2hGWRQD1YKv7se42YqHgij
FAxAwXMrrVqvNz6X7j3jPMMHoO+4t6If8H46whjLDp/zZBElGxx4kWWWBoRg+R9o5p8KuDuZK8bj
ssaDBP2H6WoKV+mtr/EIUJyRYDY/cfmv2xti1qC7UXD0d0rtN9At5VGL7J3Ko/0Ae/QN4n+vX+iZ
aPGznMsVqjItMaIP6xPuOC8ffDIwJiGZC9nJgpK2mUxdiYNzxedLsooBHlvBPINbqYiUjfG9HVdD
93+GJ8ooIkNPntN0dZiLTN8KSomHtONRKABzvjfIU5nM/X0uOs2KYJZQwxPF90+Jsgzqc/bs2gMq
oCAcctY7/e6r2SaBPToJ8X4dhx/iKGv/a2x/iVZdsyPd38ZUUGhLvztvZ9fbDYkyegNW9Cu25Ba3
yn5bKsujGXokYCJkN+oNS0MRKVu+0DmuFp0o0Shn0HxtHYDImO9sW5anPLuJ+UdPAnFLdB7ArKfh
TREqTvxJw+ixrZUkE/tt5FcmUERwaY6vJcmy7RmCzHimnl2OwO9GcK+5AiETjCpDacfVuOZnrSWY
Xt9+9bnqgil68kwnbVllQFbgHkqeG7X8SteM9b+yoOKKwwJnwCYuP0injXH02Co34CiwpOm7Ehfd
HlxgDbvFwsCVcd1dfaG5w818tpItzTR9UN5Nx6kDaxMICMRTcq19HDij52gg7kgcysETs/FZEXwF
i9eDZYAZ1adM0/8bZ2LcGGwO9GotmReeREwo+i02GF6niC4BFAeLo9vrOMJBW9cdLBD/8fGliIT3
bYdJwri8X8SrxaUbJTj0Frv96GQ+NoIMAjM5HORa6cBnl7irIp1/gaIMUCTgKItA50D8sJYCyZlQ
vWfp+KTtp79dDuhvp8ZpZ2Kio8WYkpPD39FDwgo66975ea9n2ggUtPn9LwKa7BONtvOPFOq27Eb4
ae0OXk6r3nwOsf47WC0T4KVzJILVrrronb9oup1fZiLwiyN2NZL+AtqNEtq2zaUZoeSaN785k9lW
wjHLCc82ne7O6/e+sF851z5E+ich//dLUeq/eJVHs+hRUQ76Gevij8PzMK3PgwkkwE+ExcXDix6b
YvqRJwER4lqxeQA8CncDzWtsu6H+zU3//Ng4FXlfE3r0R3+/2+9DLZGA2u7vvHa/UGg+Dl3u4kK8
nud7cHS1IWBj057Fhjkd2LRs1JQi9C49fkTrfFnsD6KTQdIp2NPWXainr7fk2RzOggTv8SWcHvgI
20GvqIW1vYhisO0aeCHb5ALLCqRIaldQ7owlR/3Msxb1n83UW3kN9zDVMDLXEU/gvsc/0ILZoYOI
5M6lNv9IBbzzhbNeDcdXQ29yyEDdb1q2IPaIbz+in7A2sXXDhsD62MXz17o3mObMrzboHz0+egsE
ps0vRxehiugh9pYTQ0NmKEGM7MZVbhni0whcvLBUlUfle5XXCIMMMgo2960UNg6UZbpVqUYuxYLt
1bpKgQLsC/JNF5aUIyy/16R7f2SmXew47l9Piwfcx0PZUzwcTnt8jQHjbIxXuMDMyr8XI0HZj7hp
HUesocaQplkGSuvQ5QvrqUhHn2UcviSjUEMYku62ZtnGQst12wGgSG/n8LnJrF5a0jBaTVggO3ja
OyIV/NIUOXArQznvhdXmMyvn4WkFg+CLXUTq7Yuoz3P0o6iuX6Y90iVlkDbVCdBnipTRqx0UREeH
tnS9t1qcXUUS/Tzw+QQ2Dzqi9OkWASET3MlP0VK7JuHEWd86nKLb9OMLsvH6081VbYF+O11UUVjM
s/mCNGhDeKNkAF8VMJxhRXojPKjX8htKJ4/MO6+My2LQMQXzHvPrtc5iUAtuPO5rNK6Z/xeI0BLw
LKABoDLQZ+8N83yc7jgwvdWb4DvforL2bq4DtypJugVNU9FQ3myWayzspd+cRlVsevG6MyWxgiCT
+0njpv1/zuE9wvDh5qNL3IKkgzPCacAnbx0rBJ1L3SO0IdLS3p05jT/nGqr4khqlE9TAdAfS19MM
uf5YyNVuzcCcmHGQMyvX3Sqg5DT7pkWFqyHyThpOunGFw5mHqZaEDCGY5/qlAbQDGUZe7TXsIR83
y6HV7oG/b5Xc6P/uKsYg6eqsX3HQgz8uZvTkxOSpbgBeAn1jqcHBUSuyXUW6sfIS+vP9b/I7IrQQ
P/TrGSmxbe7g9727ibiAaVLCG6KqWHfCYELL0ep4iY/VyZrlo8ykaas/2c2/1khxUHKcqw1Trf7j
G3CJ/hvhz+dPJKMR9n+q4E24ANVp8u+++o6sDiYtfg+L7BCC8uA1rdlWwbjnhDCBn6qk48Z9PDue
EOQibsMYbIu8vEp9dtAyGFbQwunM+OCI49hd0g9RojWvQu+jW5Ve8LoYnAjTTy7lxZOzw7Rj+6Gk
QaBQe1dM7cruFoKB1MN3SfMCSuEaRIdTtS1Urxz53v2bjDhn9KMp1uIIlTM4O56rkvnRQqqKGNCB
w63p0LTZcRP7H3RK8VpEvfnUPvjJu/B3t21MvjRJzZhj02TnuzUWBdsQgBy6FO1T1uOJ6uQ/lD6f
9SHOt8xVmJxd/FeL7u9XUB2NPN+L00EzV3M7laN4TZ+eYVRW9pg/ab2LYA5T5ELlmvP8lPy14eik
1wG/qy5N6B4DFU6MhXsLfAhaL7Xxm4hcuqVxjsFQdj0UQ1wegqbwgSWJ8YuE070ApqKLK7liOJli
6D7fBZMgnmvDb4bBX8K6VMqA1xW0zwAw3FP7E+eiy+uvS1OyiFzweRascoRNCXWI+pnfGXnenmeN
TJWjkce7HrprEfpYH7nhM5SYvF3Qz/872XbyHT1ZKUwV4ih0iPRPVx1trhWMlRbYb2jZgjCu6Unv
SLfYuBHUhUAdRwKRThHTHIvfpejmaWCL4ogM1MsG5OkKTXY4edvi0RCTxe/pcZOQRTsLs6evqGgS
fICotRNq8azlw1zO8oFqmC2B7mJwp/mJiBos6jJgsFXCGYsfRvdZdAOP84mhCa4qf1xLv7vXOQ0Z
4Cm4fhkUjtoL+KvXjzpEXQkFAjmy0xnv0IgW/cKum+x+ZCd+f9qvnlHvmkQwHCCB5aG6LOu0EW65
iG897EgAcAvPJEprbnA9YUoEbjJh8eXN3oJhfwkPLmgJd5Ue6WG1+sGHoMM+itbYzzO/Qof0A779
qbyuZ4gernqigjdicSN2fBbd8wRbtdXm84QaJzXZBd7ZG8DibgyDPKq2GOj11/w+axi5XiXmcAVO
k5Pm6Zlkmlai3AM5GXDo5Y+nsQLMR4sNq6P91DgXClieJL/DZj+lQ31W6akTNIgUEXsRR9IEpRqF
D0Y2TdjBkNyNjtA5vw3eb5utyDUby8wCUuLzjwl/liqRuok5usXrZ2u7Z5qH6F20knl2NZz1e0Zq
xK6Q5HMahGrEXYGC3ef5kQFBgNFll3jY7DdnKSnB11cpbuWr0sUY+7vsIgIqFoAdkXE64e1ApDdf
sZNujR8+mKC7shm4L/BvT/Ai4KRbQ+76RYAeEbJdAbEvVutokWXfTah4LIwI53FVBHKnv0x6wV1G
YJdkW6b53G3g6BhmjKxbJ0kaMec5o37lO9S8eu0rxewNK5YMtjTZ3rOU0e08gmAG1asMxVEal8ka
WtDfDmWCuRjcAuIAG+7AKDLTJYcalsKlEtmCB7Ho1mo8JDiJfEzKyM5gvMILfxfg5tE8Ku3inBcw
P9UNtUGy81GD3Br9Rj9eev8kwLfm9/16ZUW3Ulq+QRfjMY1dmuqA0dQY4F/D1uE4LehsAURBnZl4
cloQZLWuoxC2uW8d0BoNx2ynILk9CWlVpauPaJui83CS5R/UV4PaQZ42+eWpITwgIkrmpaKoZ03l
SLuzFxwZzj0+dmI02IxV0khNNb65BItE7RXxLTJ2VmbzkCUtV/5586xuQVm+ytnaXPW8KifmrKyn
aaawQ4uVQT2wax8iKFveLLv+VGVEjjXrIX8rfBgOS1cG+xyUovvCgPa17VGK+hk47XJGhfj5mll+
NGDEGLf/Cukhr8tl51lndsB96tOSwkqfst2nR5QntUzjjbc5FdUkMkc9JVrY+IvLHfHBI5xl+eut
B9wtahR2mo8sUGXbi5zMRLPaCHZpCJ0Ved/elREfN3C/4ofYjgmDsjxV3a+ZjTNowb+BhD+nIuv5
ntlIThBREbEIQdmRYPFLV9WLq9x1Uv99oGfVKux4xP3M2ndXw/AA5kXNe2I0FGsa5+ZYxgA5qOWL
BWeU62qwOh7FsmbhaSg+qaLCoCefbstXCRi0QzMCoshCA2O4iIWEQAhna52Ty7EFaPA800eXpMe/
rrYwhOave7uavho9BrT3qt+7PzTbmCI94w0uje6+KgNxzMRqONgUQlpBK0Jpmc0uDf8UUEvI1Nw4
xJcH58PL8+BMe3RtRk3ERG5NY/TrwdtIH+XfcihixoizxYgIqmjaAHDAAclAG5k+0NFULBMKZXc8
VAinsRFuRPmG9p5HJUuyCwcAp+tKLwfOHypGPtWB3L7JbW4sOH9OBeusOfmjZaEgJDu/3vdPUITn
1PQB6XBeYNPOVbfAHvx+WIwJvLKA2jRQ5x8o/3ZXlPjgLaBcXgQ/wXM2UkdC2jrImlqtuRZ3igyB
PU0ebrFm8IXz0qMpnf06EORTTs2yU6T6Uvmluy4r6wTmRlMvd/Csv2L4J0zvF9F00GRMREIBPN7T
9R2u4YoNNDHA+lLbORlNjdPnB5eJcvTz/jkcyYRdkYXLzeg1tnaMBZuQ9R5Bqv5OCFuUw3Yge8St
T6XqHugw+ZNzVl39GEGadQOmhGxHVBvcegnNzgKyfB5ArVVXqxurvJCa8ULNjn/KeTvelOBS/GQU
tNJClyfVtxiw6Uw+gSPGVEyysjuT20mRUNSveKkfZWivB5tfLeD/FPJcqtixiCYTrm74PhEbR2zY
gPKo4AWqQGvlDPmS4DaGy93HLk6v0/grBbIKyG085K3xYXNWFzJYoXCaoaIcNakayVrW57eAEgQ6
fpybXuKnf8tMt4cGStL7XMkx0MNU2tQVXs+kenSpt7wS9SbDriZqOYSxkV3/6cJDEVU9vaZMfMbW
KgPPCr4Ucd2lmobwxrH+2leC/YYBVHEkP4UVUuq8zD63gl5ErAyo4aK88LLUJ8QTF/uTWJcmGEDe
c9SLNRTzJGO8P2XuI9TSvS0R4pl0CjhjJrS4IztvY9zH8HyTnowEK/pBg6EfX1JTkgnfWbpZGsAe
JjyN16wX2OtLsp9nzpOaKdOYDQZILby7n5IDUtBQkKbADdl4OmUAypMZTIpwScoh0vb9SABS45eR
zMlkJ2Ct2t5X/yKB72Y9BN2zQD3DQOtEzlhbu6Us3oejrev+zfv2v/tNyJbIaQfeFfOEso857tyn
Y5Htw4fZUZ5Tu93GvWBj1gvoI4DtJOfnakwWdOA2aUogWcd9og1NQ4UssO8JnHS46zt3Z5sUtM4Z
lWrfXOcn+9/o0mjBP/7dgCMA+gkB2Q/ioxpZyUp2jv4NV0yXJPmSwVPEkoWhYeoWYUiHgHPzyOJu
4AIpuTLljjQwHLJUyIeoviiWVPIuJYjzQEOD2OA2nJpB37CQItupAg1i8C15qzgS46b5VP1LqcUJ
/54Co7HkWHxrCcS/0YRPRBhBK6hXVbIx0tb7qBaHnoxGUpQsPm66/Kd7/GFdyvKdXXOCipBzo8nn
MlCcp00n3b3pbvz/DvjM1zoRVGo26pU10rNGvHEazAwRS2Ynz6n+RVIrXtjTDwGGmO9HkegR9Znd
Jb6Qt7bKeTZ6PC/IdTPuSGBaCwPuzLoaXF6fbCSnpVfUDflyleXRjFwGLguDRM7XsP0tKO4vcV1T
Z2iX/HH6Qph3KczolNkdp7P6vxQ0phJUUelhakb8fsUr+sre6VR1ldcDlcmwteBfZr2jLag0Kcqi
koNYUgjBKp1diQG+H3VQp1g9EGIE2XBGyQUBn8qnT+GjPD8MCfV+nxFJZpK7VGcWVW2YgEGV96TD
SblX54RV8Sg7PuXV0ZcOso0/OKoMNv70QNXCAAA6+46oiOVIY9f8/ziftY3ishM+9zsxO9lsjM8N
PnvJTOIWD976M0pMdFGDLWdowjhENxdhB08vln7MNHa2XBulAe406LxEPB0w15pGAxBt5n1KiFMR
wcg9UG+ylYilgnjpNCUrRiqtu7x1dz424khiVhgMIzPsl/4T0t9GMVMvRqT1aJqrBAPeHfhs8f6T
YtK8/Alw2aeSnUTesIpTjJVQWlNaCBb+0p2sA+FE7WdeofP6Hxp6OO8NlOGPcvk+DVQcXIolFeli
rJII+47rrrN42MG+u3DPMz/JKSneONH0DVtfntaHTbYLBEqqy4Und2ITAOm+p2ClVLRtgy0xLcAd
syeB71bIiFRps3g48e/voxwGJjP1EqXXcMnoxyldWF0Idhzm15S/UWm/MZ8L36v/vmHj7d46K9VM
HPUxsm2QLocaPhKzaIkIPZMea20zeYgEz0WsEeABqgnq1afa59Oksxqyl/FhBwQJbA4Jf1C9/h0q
yXf0jKLDr5UqdgrA21O3aXO3F5JTOtCEnI/8u3xYpXba3vHizKyWtsXSqMOxE9Qr+qea+3EOXOA2
euJfj3H3Z1cQlAulKAvuJnBfKWyryt8EkVmmnj2CqmU/UkWhWfkiiS+1CeudmM1oADeDsWkQ2yr1
qCmFTOsQaApvNbnI8BvnBK0uBYkgLX/zzT6eU6LpsgG4hCJOyvrbSNn+SnMZsvhy+ZUKvyvibznH
NpISuTGH3FQ8pIJHtA/RZajwZmH2M+iHeFtIgGb7me9UzqorTmCFzFZSxAFz3nMIelj9VXf7txJ6
V8PR/UAyHUNplkpEMOVBp5ZJ5tSS8q4aJJy53HTRvTH01uLOAAheFEvpMqckqG7m6Z93+GVYsINP
qKu4cELO0YOc3A13IIM6QBCIa+jLBisbW6oBy2dl59uSNBtphcsqUZubSKcPyVt/qjPoNkBV6gn9
faWi1BO6Yu2Y7zR6YL1thOrQGevaDUnjjOFs0kDwpNwYAB3dKhfVYXdGCCkvxqhOxsCnnn45TbGM
OpMbCjSDFBDCaTHLy3WDWd28JfDkqTcdXBWkAXaxQbdVKz7VWvt0DMxcPw40broOKQ2hwNC7DnF1
42zLN08QytpN5iqX9W9P3l1GPxqW29DS9VWFQD/lW7P2flh8GzPebfl2vPRcPuV4fdy6KJLwNW9d
LpOifns9rLqeaaJ2Ld8pNLZu0RhTnxSMvxcf8ZDKQZQfgw+kmhgM4SirNhTBN8yUOS0LmGHbOJ7T
aYMoDkvuknklTnSytlGlz3p/eIcr+QKKUGYxcFBX3aVFFUtZHS9xHd0YaLIYL8bnRvbPlvEI/VEs
3pDnu6+T8BTivnbNpaj/yymV0Wm00sBuDJt7M29kuSz1vSHGFyrzOrkHxQR4BQgZeLvvqPRPX52j
K46sF0odmHcI0GOwZAPlYVAfuzzWqmb0zE7JHcJlTDponNyEoyTck+tUnrQrpiVKO0djnm1gRx+r
Z0cuoClYC4f0K/km3IO1QjghUAh06fGGJg629wKFMKxp3/G/SUf2b3wa1seCqGcU2Zp04YlH1E08
txFGVfdPPfv38qJrET7eCiph58YqUlvAnvrpeA82kcSBkFtPrM1EmkG+vegKth0E0jG2gjDZHvoZ
FsYBNZvRQ+a39N6omTf5xnRezay5YdQD3Qm7ty58uW9WoMMzqR6AmSvlU00hVl6a2ubdMB7LWOl3
gu/PRY9VLbGJj8wfFY/F4e4SMgBAFbAC8rp2LLdGADUfBevZWM7RcHDwPj0f18P64T2Xuq8myfRa
CGsoFhrw7+gQ/bCplAUljK5pc07kyXYS6lj8OebaSyZ3YHiSjxH2jjFA2CuNdy3j6TJGSe8o9p38
7sJWkepV+EeSlzaNtOe9d4INkG5+V3WmMtTl6E8ObXeJaZzk3vmTn2VKbLYP7tCeJi7f7aYfkfor
kgQjm4Q+rASqmjGM8qztMnOtujC20rh4JU78MEPumSvm3/wS8sO3UFUN3wlYnZA/x7Ran03BuXeH
tlzGtJDW1c52wP0B80/XSbxJcNZSwM2Fgq7ALGoBUnHhh4w4eINYqhiuQ2ZJRHeTzTCXg6Nmyv9C
ivHI8rSnSrPT8iqBYSYOpWpXWJ5FGKdalf8sa1dCjEa9OelYcL0KgqqqZGNY1F/vU8bbP7xmWFRC
v3k4twrzjJrk40edOc9az5kwIHYzb1DIVheKuySvBsIMMOen9zyX5rey6zd1i57ZCN0t/IVJiVzJ
63Y2U4TLXmjzevfuj6P8MDSWqFge41kg24/y6p5fBdQDrONVpIojwvwsdKwwOXTYgA1AR180F2hY
LzQ9WbIGei8fETCz2zjHeSCdUEhVJcRqSPStf/4Uc/PN8qqGI+TspuDC540IW1FErGjZiFshJLEN
i4dapW08FAqvxI+ZIkbPHDuemTNY93ZrOeqJ6A6Cq/+2BsC28ltfXc1SMNFCKatbg0RunQnAd4uv
9fvzLXzzAuSCWMhhTE9htmGYgHFwOWvdym1TrBqfnmMNag5YU1zbjNjw8kCh+Ct+ysgLqYzUl8bN
auMu1BkKjOaXNb/c0u58gNVuzXgFNrXrRGpZgvBmwI1hsUzYLU95zmwib0qjMF7XpyDgC8WrklcJ
qCcjD7ZRS1gA2OKMbiQICrXlSOKYxbT3Ti+xHOz4eCUomLxuaSofad7fez7ycG2mKBc4bC7CyHP3
zq39EjIfdCO7+4VfBefPkUwTY1MitPjpQNiSpZ9bCb+k0QKrcoGc2MrTdTq8/ANKhaRSx+R4kkLw
EjRW6SGPjeGj6rTxW7CCeu5zqhdf23kOXPjkqhkUlWXr5aeOV0PdDeH1q09Krm+eIOM2CfAslvrj
k458Vb5AUqCNfdfk8DafnYUNaRNeoxcUZWLF/9oKaRLTbIcW7Nask0Ar7UF6ISkYsxulyY4q8d0P
jMhmPFpvwyeo7N3OTDCwOK+tDvX2db8xIKE1AQi1BUOIP8N6U4LK2vZuHm+YRm8xP4y55+E+nPGj
zlZ8QLJsV85k4zCEU1NI548gmfIyzp2l7onb6ZpDp+pchfUnte0dnKtg9eO6JhWMUw7KoCY0mcMr
jtIbzNgmPS+YVwO1/ZwoQmtltkCUZHwWHxY2BFbEnHxhlgifxezR2bRc1djVCSH6lhrufVEEZCKv
epTOSPb5NVeVlg+zXZ1YPxDy/otijt5Ml1nTJnNNgHSHr8oSu/gj/B6H4NcnybPqKpQpJ/SzlMM6
3VU7XaAgIIUWfUnZRfFhC3EdYVBRotdDlmgluiePlJe7zpbkUyTT15+EWYVyPWFGZR0DY0wLcrFd
iq7+hPlZZxdL5+hxVZ62J/fNmGclk/vQMDf3feAJx7njnxWnh+++KmWi4RsQ7Mlul4ViVp56k026
kjqfTtIuyfCPrYp0iXqWMzuTMV0wfqX2dAt+h481cgrN0B+SQHBT5Qkdn3BIWfRV1dBX6qnQ+CcR
wXo8zaURovSVy08QuJcbSV2A4UI4IsqQM5qMP0DPuChyByiQL95XKdcopxPQnInP81E1TvApyZ98
DkgUw4VCeeVFp/ZYsDtIK3JMCCnweavFF+aHr5WT9SNRVVN7K9DlpOi6yx5aTl01+FJ1KwIJGP3s
FCGLICxgxhrgLLVlEf3BBm8Gw9ZD/KbMmJQ5aFSDW9RArEJW4w8bCg5ZdWXSIA2qsVETUoEfREpK
pCrykJONEPunmGgbtKgAONZvi14hl//j47IZQxpbS8LdbrL1N9+fIYh5mGOudBdngnthDpoLYyeo
RnxXhdi2yK09qWTScKnnN2sM26zUMnNqrPAeb0LqnQwc0ob5A9INTjIhVZk/pHtH2hQHJixKxde+
PcjaszgWnrOZ2isiWunu2PMB1WffFBIO4XcNMu+HRw7+KYwq89udT9tzlgWeeB/UKPiM66DCqOun
5JThJKBq20+P/JKahq5BF8RX0Es0TLDQ9nmaty/mUuECnPswSbFeb4fINPhzMVaggchGllgHb7e3
ILmOcwStdCDcVvQsGIvNJksuZLsYe7i8qlwzMEBDHW8l6AFESWIAfkk9Bg/u1jcC9Mhmu9sk4eku
8Lgko6HHaCBxGLG2j8y6SzbdqnQAgA0fJeGxO7lgirDWn8DX7H2abq3swD9LCDruypROWntQrvhJ
vVUDRO8pte1nDiFtKlWOAUcU4btlo//+N1l1uTCjW2PQ2OkP71yStOO4kpefs/42TM8qfO6mfbsT
eHd/rxl/Pw9Wue1u4V8bxS/kMmK2cduAZo8oH1zyLZrXzL6Z4mX9NQzH4Y9qOUD7eOxJQPtqlp4J
Y85GkpYeWSXBDef1BKL4Z7DCiNdJ7zBIMl5y0BnZ2gIVd+n4T6NzXMMHcrr51i4vnfQxa7p89Wxh
P1BP5XQMSOVPD+IaNZkCkFw275B7b5TaUEuoav940CajftvHE/WyQiayjKInfFb3T72o2m6kHme2
OIuT/cZOvxNkPYBUXTVJRoBo3+eb0Y9HUw5HiRXA94Lz9Mg6VNNV3z9jpURKZqP7G5WY93qLqyG2
XCYPcJN8qYOQB4aeVN4RE1yqb3VZObT+zTr8ekKLiKEuBhgF7bLZJYP5XJ+1xWQs5MmRJlEklGs6
32b6yt2wBpg9GKnzx0joBYB5ft37afHsgYjU3YfjGmJ5TKW4l1uMggvMLQrvTgjK9mEUZi9kxHiT
XXFMDBwuUq/XxV5rhQCXiViZuhdmkZMwJJGQsRLg3CA0HwxepeDaU3puQKO6ShTVNhTjEDjxMkY+
gXafN4bVzF5fLZRsHwVzvNRu8ejZcNUcS3Y8wRwpalzwAJjJS6W7aDPQC7MvKLqBH+AiHXFw7Wvo
hriS+92QC1ss9vutW8fJnrYgR2c/u+DRjrBHrpweeE5KaipHXc/HZFHKDWNIcAVEacMTWX5kcCeZ
YcsDEmIlL1xB1rymhLemdEtteTktGDfcv76e3+qH9tqBzv4s9s5U55YmTZV1NCkMP7vhewSZMZCW
0/SgowAudO50v7KUWGh+tILyOg7h9/WwsSMW9BuNbi8+Xhnh+3D5uixlZrD0qeXtTCk9axBxTOCf
1ZRVCy0G27PdPOyZ8e8HNd+Z2ukz9cCLxC07QrXIz/VIkzJ/avoKQ1+QK2XWQIgpBaRBGuPYHLl0
dO2nrdypLX8ihsMnTlUMbaggluNVA6lnYqNWdVrWu+0/FlJLMJxvQIbGFfEfmI6PpNpORAB+oQlt
xUlcS3uD4RQ7QEDRNRQXVSVvfMLpo8VQ58H7ZvuUubdmcDTg41/lw5k4/bI/oVgZZFn64+AA1wFl
jhwLwACsPU/Ayg0my/khbnBjibftZ5YL64NRZmI0Sg1Xqijl/4/teeAFSIa4xyZVqj5gkwxW6puS
IDweda2LuUNbW3435IbCa0cDWYlWJI438xMpIdWUZ5WXaLfhSMGmFiyuWu7nyRu0Aad42RKapP6r
FGTBDeH62GwklgOsB3TsAFrVkWsp9U7SqAYZPXLFKrtJR18zTRG9Tm24jUagGXYShfPR4wO4pp2V
9BY2fLRYcLqBVVboCr5ul0sFturnKF0p8sBpQFScMph6MnhpEt0Y/N4zFD4zNUROkK3m3FRMe5z9
hfQY8aynMYOaaEcK+CY4QLDiOapTvGK7DNZjqS9MlYG9bsVMs9ZeXEouNybfLo30UW3NgiqIFA7T
h808EH5zJq557cfeQLHFYmxgAZgwC3K9E9rWkVaTGZUEAi9cc8qiBbLO5ErO7Ys2gnZzoIrgkNVy
P0Lln6J5/uUur5lWNLNdm5Vz+DKiB/sKQNIpYxsSqfO4uvtiUQ9KdpCxPe/9DWhDf87RgBK6rObF
xTusEHmgUa0Vk9x2/o3Y9QiwZBgz1fHRUIftzEYg+DI0gZD2xQwEhVI5c/Uz/RZglMmSkr3Dy0FD
mO7YLyWm+91P9kBVUnqo75S7hlGqeK2kwGkEr1sazHYnZ6gBgHi3G2JOZthZa2mSK4fC0/HhQ0+E
NmHUnI04FUrhLHK8SPV72XKn5mcdkf495LU/2vWg6ylQaJTtvXocNkFdJeLQICzaRCvxdRLEYAVQ
H3WCmrFyAtXhKcyXdTYuaBb8EA9xl/7TJVP1Da7qvXkoIkvq85kLUrKjdimWWuA3Rpdn1mSq2AJZ
iLL3ZdF2LrvSIrTwiYe8xoCv/hVKrPFpslQxo12zNghhA4E3RdYupyFNRsMpr9mOPNExx6YdWBDu
IoE39EHHjtaiVaZXQmZ5R6X9umfNe6ZVv166j43tYiSfhelx1AYlzkgSxM+AKDlyA+qR9vSeZ2v5
76Z/vSHKIdJqN/E1SyRRbWZb2eZ5wMjunaX/hdgkjamE5zIQ9qTOnvGWk7FtubuSw8KoAY+F26ZL
LrQB8CO7sLp9ldwLPwnx+8iMxtKgXoDNBCi0QD3cJcaSFs5gX/sr/loOXvWo/ot4epZgXPZXzssj
Q03p91+5eFQT6gk1g9gJtnlUDIkTM6WWd0w8sEibizlBnBZeFXSvBL1vZtqBYlkKpVV6H8R9BekG
oEM8ftfpkPobISh8srhmlARIVc6/Jq1Owx5gvnJW96IiuCQ79Jt5Gyjd/KmlVUs5bK8qSNfZH0k9
XXQWsSkFhAMhXzeP7I+ab2uj+/Uqh71lQmEkiW+XdDFhCPg4aICNSJtmq89X8K/rVceV5u019AGU
juMrlF3V2qNDyCGBQf1QVvYVd3Ip+IXtH9Wc8dg+MA4hYMeaJQFmCsX458xW3xId8zjsYiI+dBoN
ECKCQKptN+OeakrX+z+OIJWVl7D462cDlfU8gDJRFvtNDTOUvobZab4i2WhSs/17dC30UX/AA5Kv
D54LW7EI1E9UJZYEMwdb3pu8JL3Q/hkELA8jZGQDp1xUDrfLHJjfxfOX2rjg9PW3dWGYn3Sd+bPc
LSDL5OMX/YJDaExc0PgCBkjUcqoI9/fqp1dOvxWO/A3OuTXUs/vxCGV6UliOsLwFQDZwTJCpuMxC
e9Qt9od4J//VSmbewkf+E6MhPSlRN/dzQBlEjBZirJgUSH7j8AAfxc1XeZt/EOge04SYQ0C4D0VR
RBEv+rZNL/hzwk1Ri9+MhUHKe78YsV9D6ZQ7OEWaX/GcRdrKgZ9TkbAkLW2x0ASPBqWJgSFkIuST
kkyCWkxq+maVPvyUPCZW0go4qYoodjtJUGNAXoh6go6U/yokp0Q6ZrBiOXWUMswF+F53C2viIOX/
VndGp0ux66volGHVAE4kGN2FLZ/ld9Vl/4ZOg48j4MQEXemtZZ5Z29UoiBlgYQpG6c5aic8IY9Sy
L83ZHFZYUnUUzkbHj0DONBKmKIolWIViO1vZ2HXXuM4c5q79pfQRfok7Nlh8R4QnydTGDnUwZcKn
YM6kQe08qnwdQ5VWNwcUQkQNb7yt9KbwzWXg0EuBggcVW9MZCzN1dGsrxHqfc/heDAzUpY+uuY3y
67OAEtsFFiYY00NHFlGb+784XR+hHAD9j9iIc22g661X+LpdtE2ub47sgvX/+WOzRKi4+of/lwRX
toQyzIi4jnjE9QDx69cAhw4h65CTEmuzNvAnDODHkQurkHeCgm6FXxC3JNPC1xeGceAhlo7+zWjg
E1vfTlg7Yn56G+/ir4bx7+STo5JAy37FbTO+A1dmYEmsu6HJUadN695uzZYJuWxJbFQ0wDu2mnmL
8Snlteim2KY7SRte9YeAcQQVyYyCC18dhdUt3gmM1l/Jw0n6oj582SAO1u6BC3Kl90c71UabV2Rv
qbVm7gd3j+qrSZBul9oIhme4SxapqEFsWKZ+AaCub3DJQ6jO9oeFFX4pDd5PT76vNEHG8mwSjQpT
l71SQgTC6k7Ka13MDCzda670SH7bhOB/OseD87UlDVtDQrtDByKPbb2/1f+r2/OyQQ+HVo/4YIVj
bK5/yRXkwZVpGwNZlst0LmBlY9nOz7JpiROMhQwYZ2zALQmTfh/ErtqABBXurek2kby8nbOSYWNI
XfPlX39Qj41qD4bf394A/txxZpuHapvKKPpYptM/vbwHgUCVokf06U/P762vxNa7BHC98IYqDAdt
QbMxJdhty3mZMkqcmuSfRa/icJmkGHsKRSK95yMDVH2dSSgkOEpphTjYaXFfZzw8HEecKbTrQI9L
ezZbVDlta1nVpNMv1slt+F0zbqIvQY+K48c69LpVpu+INSvjUMzB3BKsjXO9HFXPkwZg7cYKzfds
2auPMFKGZ7J+JxrTG0jSmeZizTn1Rss75o5Suie0dkf5DdtyKEHlJIb2BimwSyPIfhz4uEY/FIAG
06Pid50AkMK7yNYs0qttFnVBG9tn+Isur4++Zit4P/z8PBOh4xbANfO/r33xT8lU3hlRY79bbkUa
iWDhu+XBVxfxmA0JYvnDCTVQa2pMAmj+UJUdSNvDr5RIYIznBv66CfOI8w0Ufk0pXhUCivro7WxF
wJugwP51BgEJr3JtAxXbpVP+tJ/4Di8zR6jidKM98RiunNg0mEpj3EDik7nkB03TUjWSqBYwXdVX
caPxXQXxrMWHVWcsoM440YMf+apHx8LvRzT6NHBXFRfhLNYYkqal10I/Js4E0KKGPMWgrSd3owLC
SVIXDOjFfy89YrRl0RBmK2XlrfAhWlyLqktrAl7a15eZlYd+pPj2Aw2RmklSbJEsa8NfvuHMpZQr
DpMzMm+CAcGE8WVt/ymy3RSSFvR5pETLgFJgPH94GOKjY3MucKHWmgqKSguT+/FTLcHX8zZ1O4DK
j9TxEjaEQaX1pFJ2b7KZ6xFPOa0VYRxR0gZdOm8mlrWEq+Q12I0i692eVtbra3857xu4mXRhQ3UU
DK+K9h10wkQdGsOfBDOgKf5HAV7O7rlVrNk7ge2G+NS3rJUrw7fUe/LeUtUVbcziXPt/VSSzigFx
d/GGM3SVwwb/OJcFnFdW1NkWUVdn/LsKCmtD+rrhDaUDh9gb4V+HJ7Qx1OAGxiJvDR5oJvjpqjJ4
fj030y9U77hHKM9FscCCdTCVWL8R7ibBzrzrIZzqHrcFRuhAPxke/E0umM2xNipWGfMinujXjIGl
igCk7JNd+SXW+638szsh4dn3opkBOpF2cmSUyuiHZi8waJULWkCbE4o6DDzRhfWHmufICKjxcGeR
u/5XaBHYKse8VjaLIbEbgQWEXGmUWqGvkTS8ZJ/ZIyudyMl85FlJUaFU8ysB3KRl8NoR3A0J8uFL
ULd/y02Wh6TtRGyKcioJmSPk1MLQ/OX8FkzfVOSPNmrvkxpQnMT+AhCBSlshEPLizu2GR+SX3BrV
zYt5q5jwxUS1O3FlGKXgL7eX6KYfzHzMi4b5YlZnuA7Me0oQXb2OlLqzn68c2pARGe+peY53ue1c
rxO+45ZOAnDc80OkPXho/9pJWLMASuhzk2PyzjdOMwSM8Y5Or2d+fjYBI7qVmHtup9lQeQbKl+V/
sy3Zcvc0awlETmDypDqYA85Ljs/Quw/lP5JKOLq73YgXVrRc3UBR7HvBXCHGb9WKG48kl8aGXflW
b52/cMA6KMHH7qrjgSbo9nnta7gYtNmsKu8RqaE2mKFk6VPt0tO9gaum4mVvXcuE5zGVJzqjNjH8
aTedXH1Vb1jcHXgbNQje666as7m+WQZDxKE96NrEG1nD7Yesex2lTEXS81jDuIkr2dglbBi+znnH
+XCBtD/BtqI7jXjPBN8lasNuY1kw3NbRZaS45s76Dt9+xqfUd4SgT53+8/LjyKBsho9qcR0p8kDu
trIpS7HouQ1V5D5nSZcVFMB+6/0nY7to2fkuYbE/HudTNaLHozChekF9LIBFn2Mrs1c4GZBZY8Fh
HT4tNtD4SXq7a2596us7es4IfhRiiXIHMhM1cNi16/9Oj4k0Hyrc7UKmzsz/FHzMXCe9lKSYdGm8
vkfxm661lz9Dl5Zz0xHHd5xyK9N4T+xu14Ov9J059YyeqQBvjTANA3UuHCR9nfWAbAq8cc72meLA
q+UwxzZB3ckniXL5g5WpAYhNwQtyuupZPL/Hv1JyvjNBVN6zG8f2X8u2rYLVd3p1J5/NjoQ8TQgB
KnCCISjAWnjWEy3RSNl5C4vZyWAYMx76EZxsJCJ1Yel0YXz3a1HZptXkner9/G+jXSmxfF3P37nz
NxLazl+I4iKiAAohzDuyCOVscY5tkVPeXWTgNWzAfGas/61Jw8ZuNMJI7r7TPJtjaIRVU6KESUtI
1ImmVT9tIXyv9DPq876SWlCEegy4fQWamQwURDgFjtCbib/CQpzQScfRPYF+FV6pQ3/Mg2dzU16B
knjerbdh2razsvwjai1AHB8Rpbjq8eIsNc43mtYgO3Zkc0SlGWTB51ZoZ0h6z0g1QB+ziMIFRTKr
Yy/Ctq8iwIxUTPlzDgUq4oTRBkfOV40odssFLtDu3PNfJpun6z0pN16d1AIsJALEHUFGdkOU2zCr
aug/hKMHf7HFaTuWwAjym093RTM3jMSMomH0VxavXi9EKsaswCg75UvlgN7iyLNJXyNJRUaDJr80
PLdV5d1emOItrcwjzQBht2jKdIGEYSnT0GvGcXyE9xZvzD9rXwbEG3AOSJ0ihbLSfpHXFRK/GPOI
XJoZUMVrdJq4UGfYCDZLQ+U1By++rqqsULPY/7ko8AFiKPc1vm4rvZOPqtrpZNns5lKnsJDYFeIg
m3wmkCDY3IQWjPR+l9mkX7RIuBU8WA3yzX8AH3VcpyqnkYP1Dm/pIjNFnCwUz8a7X+59PODvWAx0
etK2OPzpGSgkJ8LyurBssGjx3VVNB/9gfK3o4YEbGN5nX7JWowTDOfzKxpcPIhrWXeFnY3VF2QWK
24w41hq4UNaKRj+vK4SU/I2YvfuEwK7ysr8pb/BNTcSm7uuVa8D4CdivfS4Y3oLEDmqA+2PZGp36
3RtFflZcCpqV8Yf5v/3DJ1K5FBdUkjESg5clyuo+VN51KU+a8TVTvz0GmaDorSEDEiEvSphnn2r2
Di6ByyTC1NMoZRjEr2YqMv4WatjAEHDpOGj0xqV/yREGDKag5ah1f9myKuFQiN1GFaRqzVChFDCy
f+9lWYUq0htWSsjlnusX+LMBKT1DqAXwoOoQv7BoHhRD3qFopfpUDY3g8DBwdke3N3GUjftcLEs9
kyxiZAeIXrocMe8vpIWXgXgnxBsTxpLkZSsZVtejgx6QOlOdT+noXU4KLNZd8N2CeYxk4GrY3Vu4
YWSM4KfMvjL0isfS0rj/LXgZB1Fm1YD+Sl4WXYhcjs3fCiQBffdqmqifHs/RMV6JQHlKM+JuTJ3c
K9pHJuyFWWCBtcR/sdjBvvvb2bH7yqYbdUn3J7rVLnX22Izw4UKCJhOF6hTF/YzzllD9cfVuB66m
4cHmBzLIdxqBSQzwww0+IKAE8LX/KxsL0wZSIKzws+D8ZRBG/BtzzBMU84G69X3ObINprCfPFKrp
5/YGK0y/j22gy1oRTsOCXeazqRWMjlKKUMUDZefgJrJ6i5PESzBsw65FjfB7uunzuJI6ujPkBUx9
UKyLmM4avVzqUnYUZPrSv8s2K59y5ECFt0xxXOkZjf0CUfUjknnKfngwQst4XwbjC2y+/SxDuGde
jm4MPzMdclTlVNSt82FUTDq/ZCm3OGuz5N9eNC70RQuoF9E9Mk6TYQAucLBc5m5IWPWVIEog6JsO
gGx7jEOeRHorlC5K27S/VPCILHuENdtVEDr0mQDMXH4x6eimKbClGQy0dpFNfn7/jattWj6BI44S
NYITx/l3PiL3dJNEANOAfMHTX+Xj/ii8lKXCYdlUGsOBYGgn2DTPqnpqnvP8QuI9HrDlJKKsbi+X
Y60v7/I8uKjg1LdHX8CC94w0tN39luO4sHSjaClkdgEGSppDRtj8MeM84uEkN4tKCaJBMwOzWpvl
Ij8EhUESaF0imw2PADUfYgxFEY1yUvSvMDS7Qpt2B6Kq8WPQ9qyiquLvmO5GYx80Meo4IMgIUhZv
IbQnt6JhUb1MGinEhGQXPkfnHJqHAtG/beoMrZbpjvOXf7T4Fgd+b3HNPGAtO/hffeVnFvTi0ckX
pieNukjns41dEt0Eo4Nhv0ANVlg5lQiZ1OlPNiZmEJOIHSs6WxxQOxS9wWQvCMtrOcIMweTyNBtj
8E51/Bb/T6EP0NdTOlsq5a6Dl94SSXVnn03WN0ZHWYnv6nADN1wcrDfKlrV7EKlI8KSuJdBfKtV5
4Gy4vrzLenr4MkgwmNq81Wavof8GrQWDC6hOIOEnuBakU9Ic44IZ9qRwR6WX1QFxNNCU3Rejo4TC
hWKxikCqXJg/WwNiBHkB1cWGMol4/sAn7YM70+4vMV3J+oCfCnNwqmRrqsdHqjCPUgDND/DOQRLP
/Vxq2cGZYtzqMNevQAsjouo6DWRWXPxfD66jv7qshWXbKILD0lGUsJyzNB8EO3KHSDstS2WFVS0c
TkpEWyDCW9aqpyCUnTe0uN3+MSpfUVUl4JWHLS9P5Cytcd7pZOR4dXCYeaoH/wV9mSOYUwoJIyrr
t45i2I+MrrlE/J07AnVceytpPYDkIOTCTIps3OJRGdYG8xmDQsOal0F+Iw2uMEuOCQLPvPFyIW0B
kjChBVcxXz/nMGZ7eD0Lc2vjUxbaOUFB7MdFwHk6ARk3flhfAlVvjoJ/uQr8ogiW8/OF4f1RwkXe
TKp+tfK90k+S0jNn9djJ+ukZ6cfJVe5VnddKkrnIksXDPdiSfceKB8SU2imiWGES21y9d2klFBWE
S+tfey/0LT6wEaPjm/tAokJPc7MxcIgWKk34L0cA0qYiFtdmTaAHb87nFC7Zt92+WCBWc4aoSiat
Gv3Co/sPhNV0/WroP+8HTNn25B0Ywy/qZ8RToht+bs1+CF+VQm4iYkRti6QesEOpxK+xcXPaxh0f
bCI2r+5l106CZK3KISP2dQFLTyI3iV2UPxKnMDcAWzt8NfCtyvToF9sf+O0zEL0gHRHq/70dXk7S
ZaMheryaX8Pg+Xbb68cSo5U3WqNlgJCMwYhPodWnQG7BE5V7VwBhq3sJqGRmxK7Bm82RvgSiwXLO
O7BlCyQubjTP6oLHrYVZVgc4JjH1DTDzQmAyF1A/1hu+jV0rH5nERYuf2JgS0oIe3b6H3OtX5oaA
OGCNDCwTJOr6W8YhML0aMDSf6m6j/00NhQ8bNpnBWv2G+XC6LXFUGIlJh5glKQp86gMWhCzNDzMe
Yh93QZU0JmQu2l3p4KXABGmTC/OtYz/hf1v04QzbG0ZOUdMcLvQZAZckiLl9GrhbzG6NXVbcLhOY
9X1fkc6fzYdiw0W81Z/6vtlfZlo8Bquz8q1pIWOjF90OVRrtK1hdTFDef3Fe7iqoDdx+eu1eV0pA
XEa+nu7/7V4m87raUZha5u5YZi4CFKD9Xow6q6p1GiyndMwaOB6UyU1FpiWMtskXtPUSnXs4uhlE
1Qv7l+w7AWLkaFrHaoIp2i+5HewuW9TVuLq8jPiI9//3kOwCnVXb4mxc1K0TIDfaqP8a600d+gEE
+2dyUGA08+G/SWN0JebOdp6NnhCVR7eh/3e6kuRRDBvcTw7Igq8ZRnP462BjoU7VAc4BGGn7gOEH
zzc8oPDae089ayc3hyOPBFM9JCntcEtaWqJsQe66x6i/GSdgFZOnan/pc3X70hcBbjnPn9dHSHbu
LvUr9L07ja09JNPif8jO8XedqjH953LoV/7HVaTddgRPQ2Z6pfLOT1hydHFJ5vLlxXCFw5fI7LlQ
m3kW3FvMHZ07CIUjv3ye71+QYPcJEEKh1BUowMVYEGLig3z3Q3J7Ud19MDK65QBl1yledpCf0yo/
HLcpcgUyR2YaQ89y+EVUVH04vyySHQDy2rxUAo4CRR+sWIsBACu1+/famTJseRbjUdWKSl/W/H0A
moRsdk9Y1v8cdaw4Ze+JnBymVTb2gPZORC6QmY/70M/8LTE1+QcYKfafa4wdBuhjduHKqbA5oAo+
qyB3KjR+mG/5D77zsCqszSevZQSSeqIeHzIoKBXEa1jCTTbh1EIvSt16O/XjmSvJRObZi/9c3yiR
+tTo+FXLa5SwamspPk4F6wBiX3M0TihA//eVDX4HRF9YjLj9ZQ2lqADT6hJicQGRiCtuZQXYsoP2
19j4DvRj7QYKvNgVk5IH0sfM28SQ6YiIy61zMd+o6NAisKpk3d1aIaGasiPO7v8tRZN9sufy/1+q
6Ag3N63l9kU+h6eZ4Ztb4sYb6M6jpSPF5Vr6OVatZuRHE7Z/hHicWZVrz7skwfW5QKuiconqpr3Y
u3qsUO2BKsHgN68I/BcpTdgX+kocZx3jzvHR16NRV7MhPWYq0hiLlJsQFg1mqXCmfnfA9abdh1za
1d3BlZiQ9l5a5zTwK9gMYAXs+kdVEi3MlzdsXRLpI10PAnRex+em2FcoM/mSeyxxk3It4Bg34RIe
Z595rL+L+VAgRrGNQkAkcUsK7+FRlK7PNwFEn8imPqkiEl6dvm5/dD46TuFuWM3VkwFNHo6S7QpP
wuKZN3scHkf9WvIimOqoqSTLgdJYZzdIKvD2NQMGXkgJV/nknvP2GGBxQ+HPWeTmemp1UkFXAGUU
jKz8hlEfgGCgZW7fkzjzFvMlXn18xA4prsa5lBy6dQRioirTFdA86idT4cZrHxhjvJZSQJDCe/zn
xRRMwAIbM6412Cdt0i5kipBFT39oOzvZcPVnKBSx7ix9KJ2A7zw+kFGEXGy9eUbvqk4x5sQWOOzZ
uFSKKcy5Tl3mq+WUaDrLTZkbKT5o7kSgBNBie8bidui8C8igQSryapvswomgVP0Qgjz3DJa93pgR
JLkq1RcB5+xVm0sXkgsgWsXYs9qjSrGpPYeXEm43xN9KSYnLiClYvYw/pMDKxDCRjvweO0+VnYGJ
Wa09DziEVvdYIQAgIqnjE+/wN5wNsmCbSYe9XvLKDJiW+ewxTo2c5nne8DzIs+bWXKoyjTOo3MJ7
boAJOnBCeo6n3PQNpKMithrh2HC4vs42GL5Z1n7g7KFGSrEATbwMtZ2D1sPR8siwHJ+oxenTiPKw
LKZ+SOcJZafitbPpW0yIfoVWlFLyGsdT/y6AXol+Fxh5dhglig8VYA/nKqLE7L+ZwGcPXb62erMS
GfJ6J95ClG83ZPHhDX+PYwr/gMji99AlkIehGevhpXMCoPZ+rulh4KWp3rQveCkPtrnRISPADove
ZxeiTu0iNakLeCeyIzPR/uBbBdYv/fTbtbp5Azp8LJ8Expcu5gIApPuucoo+l8wUjmZRE6V1DhM0
44U3cLEldiomPbVbBELWAswIPDJ5VGAjpIpmPhx0ybplMo+fzroWk5o5LrBlMMGijSkK80A6VvVc
6hjqBM1M6Du4eTuxyApytyIAS3W/lHBfMzSAnD5LjOyFGQTvdra5Ts4bX5bi7W5se7SynLB+itzF
0rwMIZVEcDL+ppmwtmG1bocsI5CNTxJGmrOyvVk/Bn71zGRh/Vd52T8j5gRlQlQAqbh28HItaaLt
4noCxp8D6aaB6+H5cEpt9N/Rzh8E22vgqcjpvQkQp/IhFcrQ3HrI6hCNqaSdQ38l/adqt6jy6QCD
/gkW6UybqEnWTQxJXOAqaz0ZlBxv2DwnwkyPgHN4XdhJbTOMo0ejqVcGYRNcEKl9Pgtgnug7HTCb
9hNuBYPq53NQx31W6lzXBRapssTZgIE7ZDmTCwc1FztnGNpwVzwCvIlsBx/+K5RgHdVNSlZGoMVH
wl5rWWDyoOijsAIk+3OjvL4S5umvyI2Faonj1okY6m8/98c/2xoWLS2/LAmeQdJ3Yk4OwWjNBnJO
x/y9ZPYKvqtH/E3znMOFYDI0X+i/iE+3rEi0mXaBqNWLPswo9vvBRlbUTmziCEZEvDPa2s/HNFPt
CG4suxlq0X9KEB5PbMquDrGi+MEln74orMaIfwEDjX81CCxtV3mckCL/zkCkvIKoEEE3YC5fQD9P
oMLOQBOFdHYJapcYyGwpPj2WgriY5YR6dqm78he5UxzHB0hwO849RRN5cPbSdhjF8XzW1hT54mI6
ePwclIaBpx24Fl9b6KsUyu9sfeXLDxVdiaUCYswUn5kilrLo66Om5iJi4U1BwcSsymqcHY7T2jVU
bkOfqoYErRi+sKi0j6idM/L6/S1MmxciEFZD5ia4ooyVt1ziT8h/IF+bFssw7+LnMu55H9JdUnPd
YPPyjAw2ZKJHbG03zJfUMDKhhyk8jSDONo/wNyzvgyMQ4hwD8H5adASWA9NDgKM7hoBjpRVQG6Gs
/DPG+Twze6Tm32QR+NGtg19eEGzmmquXbvnNNvleGVCeEJpiSVDo40ZWZso12Tg8PpeHaDBrUg3W
gIrXFeDnqcQQwSFVZmEp4+OSBOr4SqWFwjO5iRyTVkpaSW2/4hpSdf5vDxtnbtT7nCNvNofomRcd
oZgTxbVI32HfOZXebh+TsLloACU8nXhjo8AtdueWNHpgMV5DkmP4HH25h29B7H1f/s+RN0WZ3XsD
LyCrjEcdpJKfot0o2Yf+RuxVKvu+3XPbSltGGpZWKEVehB2mN8wafX0r7Shtv4kAVFDxogoZT4jC
EwfC7+JzRJ+ErwVhng2WHWk1pjNuYOMMaED2vCO5eeACOix0uUn9uZDQMFN8jPpY+YM1YwCt7Srw
uvqRlMZkRuZqHqSiTuv+bTFbhE9NEHWWmTXS+4PR27pRA4B61gKfyDdRJvjMC1Y4keeBrnSbrs0T
4Co4ofFut5fC3XZ9JcoEaLYWzlj7XClvUPCEoq89zDGxZyDK9JRFhqzVxEeW+tqY3yVc9tEXI5jE
cOy2CsBQoI13kRWymxeISRCu2mSgqhcWKACmzGA2aKHlTaLbqB4FKO364T0H4qdMit2K2Goc9r0t
k18nR2CFdzS2cJcYrKWFX/nN+uGaS76S15iI6PfHC6R4yHAXcgKcwygkZGXvSul43rcpQgOZ3FDf
N4kuPBqcjjM+x3LES7JWiagC5skeRZU91oJnNRRZWuJg47y6T3Ew5QEbS4MQKKLUwl50KPzYM0vU
PcwQFMGRCURfTo+S+XMpscKlaENAkPq4kGKhGaQht7qtvifJttux+jf4bqVYiPNb5V/UY/N1h5LT
srHHe5EhuhVEjA0J6M1g0F363zy0h+s0aTKEaMbVToKmJ939lfmQHJ4+6Bw7BqW4+apOFET+9Pgy
0lIrxi7YVciIdMyJEkaLZ1LD7P9MLJxtWDgzYIRsWm7D0XKlwRZW9RyK3i9JvT738/dR9rWfGu/f
DCYaEHCZZg9bRlkmRBTKN4yTP85LBp4mha2TevlFVRNlZ/uUkMOZjzAzf05j+Q2/s/LISZvweZZz
Cwq0NRdlpKEiuntSWhcthNCfphP2VCrByL2DozLIp2pDCF9mAlSw7zYy7bH683NJp6nNIQMn39xX
/noXTVu9JxV1zIHNncZjUBmshQo6aBJG6kw9P95kI42nNUFOm/JxU2S4rzREssfCUm/gNjie5rzT
DFN63OL7VE7q80AavCheqPSpidI95MRk+O/MD/IIMZxD52fEd0xbiqICLK55ilZ33O+EZTUIbukY
BnGRDIDYOA/qsDOe7USGnxIY20XlpBMyCmckfw2PljXsfv+MkEKIzXMP4MFVhkNHbra6PYMGRdNg
5xALX0nmCWVYz6Tq7aIkjoxtoUloqcZ5MBYuGQaqkrsma9vYWXMT1ICT5jeUwuRwQvKhAVb1LvVV
2ZSs9KzLXxA3XDSjh3qnzoWYG0fqqGXwIVNZdAU0rPbIPb4LHVJK2ciVnXMljdvigGaPNP9OUFrq
HjGCj/xhYKzupKNMBycgHxEZEao5Hosq2Cgyj6jAZZG1t7Dn7mzz8d5m7OLzG4w+uNqfjIWAmcoi
JFJfJqYms3D7hM2ffIqrUCdokUkCyBKIFbgSJZM7cYkGIztbhg7FkHMLERJqXr3NVXOP4xHI679J
OE24wJInXyfusFH4zbMw9jpxfO3nY7OZvBFLV+Sn0eR3IV5619XWnqhwckJ2z9XOw3LEF71Uv2M9
+X9hVjbogVgL/cIGKbGVIK+Z45CBnPeKoFeNv/xF6zTm+gpm3eI+P0x7NvUicNavn72nURqkmKc6
j4QfjABGD1hdpNp0mHWj+DmKSvrlc+Tn78BKejsVbDW+DtLn9JKOwkrZSkAELVoc8vA01OrH9p61
R9iwEpFkzOgtVSi3miP9+xBu55QZ21OWNuus8fBOrRPW8KOg5EmNevxXLz+Sk0Hz6vf3iSghvrG9
xmcpfTZjfBvsefrXYHa7q8jokMx4xS8xDLXYQatwqt0+mELnm8x8rp1DCLcssR7TC2HB8cRn+rbo
YG/d5EUf/lD+uyOdb657fSuTiy8mxctglhe1SO4UewyaWoDR8lGUxNAIG3R9iKsnJ1BaZVOnozjw
Tjwy7p8KuvdDaOYTAfGY9e9vLpht3qQQG9N0p+xyOQVvPjZFFp0lUEC6TlmYFan9EWCPll/fzrsd
fjiRQUi18prM6sB0+BKIPFWTF85lHieyaA/pPicTQ1RD222MBC58ltRMCeOoS4/K8CawyP9Ey9Cq
LqAoz44dh5I5fowjYmBbvX2O91a6IzhJ38EiDOi+e9ncZMlARaUV0KBDk78zw8QRo6u5DXwn9j15
8o5zeI2+O+ias/M6uRktLiJFmhhSZcfkotuBRLzT3fdIiGKl3O2DdohD23l+te2O4B13x0W+0FP1
0bCmmUdktglyfYIwabMbWSAEHF+fI18Lh1DXJ5RYmoDlY9wvL+NvgJGE+H0cDUKuNeVYNde2pWSS
6l8c7gAtlU/uc857fUfmbnFw2vmR1aUcqCvJlcpCafqyQOWQDcZgb0iEff3hkn7N7z5k/r85rLj1
M8lbe1AF8+EIDlj+0tlCKUXPdQMoifTvINka3hPGyK6uXv3RhDcVnemsbPctx0mL7uN2nwJ5MPnm
JLqOO6aHWbg7KmVK65n4usXkYqUKRr8dCAWdVz1uezWfzqDwXiBQSw5yNHb3YufYjkp3RmroB/EW
Am5Idbnz3/PelAT7Q34bpKlyTFmm8QeJlA484sP+rv9z3omDLknUgpJArOFIiBxGb2BQLitJdU0C
OfzhgUEP0z9mZQieNPKoftVdDSshZpqkW+TMASKjP6Ew9jOwokpTXchdIuSZHH7ibOwqiDHfHN0E
d9ggbvlFjuGP/i0EYpcjAICRd3aB9E5mVpmv4VDTTE2GLqSOC4jUJHY84TJ0ekh1iyEMvu26nOyc
D2OiZ4DtFFJ2qAo0Y7pOAb7temfBlFiR1letxXMAzfggMCsc+9ZDErNMlV+QyMPCiRXwgARecnlz
LEr6sAApk+Bq5sjj+WgLL4vlfFTWznfDcP3O0OAceSeHmzSsqpWYIEyA9oQ7kaEsAtUUSITMkk5O
swUcBlkEwEfykY0Fw701nTgnHPbmY9POVc7/mda4Np825k4hYCMiVW553BT+EzxYugfyRuQjhU9z
J/j1u08LrLBuwS5KJP3pHHrPwgO70gHSoUljjrFwBVwaSP/nojNZS/UYGXFO+1UpLb0sC7+4OQ7+
+bGqb8WXvasq1ePIXO5UNi8WM47oapT4es0EZoV2vp2jnXnw+XansgzaBpy39ISV1HPEoKPxMxsg
eN3qSmdtF6uexG3UjNNDdd2cRKyrER19x2gwOLkweJ+TwrMSrC33w4ZytVBv+c1rqFG5XGQn9Clt
IMUOZ+XP462MZJqo1etsDIYDJUSRglTqxVGuwBAl3wImbJSkHiMSB/VBoR2VdiXt9aQs9tPHdYlJ
Qg1Q80qBDKat7cuhpn4FiMTih+LaRLHRqZ+i1TztKDv8Hjk8IhvP6xjRQbesCwE2Trkc3r5e4NNp
AQLSJB8zLYpkqze+zYNoZoW9NuaXTQgx93VtjOSZo3b6SctBo0zaooR+ldpZi32JdquctHpoYubL
J97Gm0n6y7tqHnmtUzRJ+yResfZoR0EpiCbZ0a1tdOpgA8aBQsO+Y4K36ezdSgn5GyAQ5LMd2Usw
vCUct3TlQEN8m0isi7K+5t9FO3SV+xDTHWecXs8jlsQJ9vjuyMvtNcPndKIQI1ZJcsdJPK8LRqC6
NEOVrHAguKLHIz11bKmIrZdBkKyiQ3WlCv1Hi51tc4xClOmn7mQcRo1/DCVKeUGkd36FbZcFRlVL
T1m3HJIO/ph/Ns1IIle3pEw7teASNBhRn7x3b2S2PUf1GGdsmfWNHUFFzOkqqutDj7fCJ5dkhfty
JJtDkf4Jn1HpRnKBcdC8wn6JviFEwSB+idCWiTbGFs81H1hqFFegH6k7wispLIiOx0wsFGSaZPCZ
JrAhhM9l+5ctNiEDmgTauVxv3KD8R8Omjr6ykUYAk/nwygHpJIyt+4aw2N7goTbKKn9RzTdecNZ1
mfIg2wcweThOUT+2gK8fqN/YdUp3TLztmH3/UVzmoUc+X28vLca/HbHf999LxzlcDeWVRDwBS7l7
j4Dp0IIP3qwDaHsVZv5IQLZa/MLpzQ6j8c6/YyFlOgpz359b+mB9uVXq1SPk/fDqq4dFueEwqgyX
JxzWcgZ/v5N156QcXY3ozDOxapG/jTnfQadXBxcikrAt+Nq8u9tJORTdVFrrndaSgPe1Yr5eG4zI
wbgJs3biAamowh0Pl7YzS9wELo6JAqIPe1v1oORKMr8LLJPyJxM//6i1BQyPxSkrKIpkv4QNIFjz
SA/z9VeuCMb8ZlVGhK/+/00Fa2DxlI8NTCxVzhlvmAt7pXWGz2NMF/rG4/hIQTd5yC/0VhB4FQcR
R23ylua4151dowmLWeMVGTRfCupnlt0WyK++CHmOPwFRRtD+IseYtLMnIqF0p0CROsTMJEiby+Ax
E+DebXinyE0JRWOK+5iQV4yeWiFgrbvZEsw2/B/2YRVa5rualO+vkNlzJEfi2U1jOU2d415DRsSY
VUeRS7SbIe9B8Xv4gDfmHM9mfGyo66L/tpp+K4eL4HKC+WERo/sr48oiTLgPnBsg0gOa3+g0oNu7
VhTTGlpGSBzne5HcvwoEzR4H/haJxsp46nw6TVSS9SAhpCRiNsMvMfn2GShc+WyUVvO1rVhjsxZk
nbH1ezJmlS1rgj5VXCIjLe/lwEurZkAoC8YY+3urCnJPafB/a4eVf/c7gqlHetVaEwgKr0ZywKz8
4X4zRLzsl1E+fws4IW1QKAv4AxVFZMm36GBIKc5iQ4927BVsEH499CzeiVnY5u2LMXqv0An7rqwk
YkkWhDjiMva+3ixmJqhnvuDRkbHzbOMNU1Z+lP9O4JU2blgFpkYlqEBe8hadHgQ9K7jFsmdfQ1sL
DBBanEalTZIIT6NCZvFeEIi8Rn+uxl6j+vb4ST5XSOHbpQrZdajM69ALnu0ruvmnOTT3z3QkkAyl
pxlzK1Lj+VAuUC7gsVeAR4KQZhc3MI3algmrJi1Y2PGSalhsYhaRsoPb13M/lF6iO6X4gDTc4GfS
e8DX+3BIc4jErpPSIxTyuDK8tjTb4eZyF3GXSMVeD6/cWNFIif1xYk3QQxGcVh03EmiVqBn8Wckc
QfNVuPlRU334VFFjdF+suaBhvVsYm2IHzg/tfa4IPK+4irErMUjXbCEK2HBVFzI0i6GLjXrXyH92
XHJczbNiLecqBOQWSHHi4GEvCaXHrfWvDe4AZXlW+CXzwbjdaz1fVB7/fqZhEIErD16lWc/cmV0y
ZtUTF+NUtX0f3SECQBnGwemtc0iuQMKn2vPvrCJtcMAXTgF67iT6K6NJC8DrGvF1HBBBF9mTtefr
I4eAiEqU9WwAjtkZ6f3xKD8rkcRJX5XKkGAVn114/+yYZozjAUrWhVzfaVvaNL0Y4LAHbmffDNcg
3pnzR/S8d6e6DUo3nl99MfAveZc+myrS/Qocu+Tg4iX2QeYB7gkNgNLEXL3vELX+pva0gsAxk9ZT
aWtOUHVVkW+LsQlky1suMjzb8rTGNZd8K5vWgHq2ae4Kv+GZUCnQGow7uiWXmp4wqT/xUUqxk77J
X9piUDymxzBc8uq3EOslShmDsuxvcZiJut07xBZ2/jXQ4rx/zfyU/3t1pdgXgXCLVx+yU2/c1jf6
zSdFzErosqQCUMEej30vJVEszQXa9oR/tEse3nIdU/fIscjOoGPd4xlrBox9f4ZJu23qiBZRHXye
jeOJTFTAAx4NnNBVD8ZRPQcl3bT2U3rRwr8UgeiqhAqkSa/55JcZwXaGeG02rX9FkUtDSxcgCB8t
s9vd7mgRJcpLV/A27HtVmyVH7eFAVQP0dkoacSGZrQdt/1eFHVyk5WE3rezapmE4bnlKl+gPFF3Q
bXc/QQXVHh5sIJXNLIPjBkHqpJ6Am9McuTzGd9Gugpvy7EJlpiN0bCaM05yyGNgIdi/hdrnb4Wat
j8eEjtmWFTqQtkhyilal6BSVRJy6b3Ah+OxsVXg598WL5f1mAoCPn6NeZbKknIoNosLYTv8a95aq
MZAem3zZqAV9LCzkqt19Yn7G9X8q6D75GVrtHi+5iMhbgoHR7BNe5MWm6ySO2NkqtEz9g4ZB6riD
Bq+qAVnny7Gdewxk93wqZNHgfC1rdz2XF1MdRVxiADX76i94fbMgCE5wZ09lzNvniXV+FXKP87A0
sLMs42WzwoccE81JLtzZdd1z/DfsDxQLWO+oJUqas1j/bueuBAT/WRgsL3S53GOC6jM+I3NT/P0C
8MJF792bUAAsWgji0UgY+zy2DSfq1Zf/aeMn68SAtICUgnoYZP/WwqIBAEugnZFwRdmJQNBp9ueh
+Hb3P6enHNMbeEhMQVluarP0MA8HNau6D0fc10yHhuLfLH7dKP1xC2kCk0uMpLk7/351OWzV0f3T
0n/MlYMRZl2q7fpbZppThKScX2JrwwbMyyD28KHCa+BX0MRpC2/rv8/X1g1ae42jjzt3Hng1noDK
FDEFMpn6tWL7gjQ6kOsLhzfHD0x7eE9pHhab4UuZykIPvllHqLHsnGTdGm9S4sBe1cMqi0tk0RZb
kmlWgBxP4PaJRdTQDP9A1N78rMiVnTJbITzeeoxrtaAr6ckPAdW/uT72RBaTE+D9drqLQ/QlJ18r
tE/RprFzYpyIq6+4dxChkGKrzuQDU6+kBjt7E7X1c0+H5S/mczwn7kQHji4LiVbJ+Wz+bezC53oT
zTx7G8UEhXEg8hElF/mwTOzB0zpTpFCkf3IpIixfEPjlenQB16CB+t8VP8rWvguql0+7QZ4N38sn
JkxKw6UmuRXj9/1HPrQZMFV9RnX3PREmUhv8Rk4mh65j9/XA8jAqjHj7vwJ8KFH4klmkRsm8GR1J
gK7bulJ74Z1UXkS2WF6NbsC64du0I94lPK5YtJt5ldcpoE+lQcozkmpEi/yhyEcr2AfIRIrP+BhA
zYvWjUVYgy58TKJ2iTE8krRHBLiDu4DIMdc9Qf9UhuIhDzFpq6AZOF3DF4ERcQFXbikyQ1JbNmQk
0yYg73vd8NkvGJVTRl38xrj34TIMODLvhEdhsJZ/4ovrNyv3x344Om/mZl1h0o+oAimoQano6cgN
Le9i9Kw+kfaOKNKKyUYytfEKqpVaitXzM2PsMYOpRRqqT4NKF4PGnZvbqzK34dzUYAvTwDTTA0Nf
CZhbsDcu+g6hSQ1X+TI7GyfdoNMLUi5UbRZowbX2LGI5W2hZz1UpMck1WcYzL6iLpH+hNUrtqcWS
9i8Bj+7ZUp44GxKhn6/pH65C5wHm2jkuqueNBoYHoQNUOj/xOFe5XkXjfFBLtU7O2frQ5Sr/Pecz
EobmjwfqpHD3WwLL3qVAnyg3e9Ictji8ZtQopab0A0rzs5yAAKY8HztJ+71I4thQHz/KadZdM03z
HZWmIPGQ/6u9OKnXHzRARa8e/KLJ0hA2sG87Xr2cKRt9i1OE0PLqJi6QErhM2n6UXdDG1pTdLbdx
iwx6qwjZI4sGvvFPaRHZirCcK1sk4ih8jfyFQ+/r/C7SUqAMFGZgS9Iulrb6NLx5/SYRDCZ7OZ4l
S+4MNI0Tq7K8oaak/p/VEExvd6Xs1q5eRYvFelPJ3/Rqw+IinUNJhJbrn9uqhh4bsB0C1vFcdE6+
TCI2Qqj9sVy797fmdrTsv/0kdQvy1GuMzOcj0V3Vx0vPnI6F1jD2kT1Fr00a5b+T5eemhL90B3Cl
Hsp3n0YANzIXXKYk9GlLUW0vusMDj9bVE6HTYmuatAYYpHfuop9m7M3IxggbWbPK38+k5/mqi8yG
XjPxPXvGB/WAeKYWp6AKaSSZnEbiLyY4Pe+k0Sp9DhLEPpy7Evx1Behdum7orzZVSmcKfSKcKmuQ
U8N3b94s1WZAJG36ybvqIk0yuYZpbICZi7oJrgUbJYAIYUPrFx5UlGnIeMHRD1q1JQuTI4nSRxHo
s3Tda1LPEp8OZ0MYAT8PQ2FNQwCwIIYJ7mGyUnQVVyM/ZQEzEsg8qkTiie0rwJehGsH83R1oy2fY
kKaaiYmyMFBuFJ5/Yq8WxBhj5kPSfECWkIy//XiP19lYZqxBa8GLNLgCFEev7O0SdsYe/erC0DEZ
Adlm5kawUq2Din4eiWLlm3ezu2a5lDw72Hiacp4NnydnIJ4ltFw9uYxVGkqi0OSjEIL8llLxMZfa
WdxOtUNbA5h715E5xctAvOFHCVdjkr5c0rEkRtLf9M9TYCXZL9dclWEVUuHaTGeFkaF+Z75NtoHu
vcxgi270QQ639+6ChhqNV1N98GnxV/jy3UQK9F7mN/C7FDpBkg2l6TUJqVh9Nh515I6rBKmKhVBT
HoEJu3x77OypjJ2KedN0z2CH2RJ/gre+GltLxguPMSorgiaLpxkbBkdamb0y/NqxgYfuUPq17Bxi
FSrDfmJZ4V/XnTESwElglJZQo9FdVMgYSAhcHme8Xl0hQZw8cHG3gXAiYUrNMp/q8ptN+597Wa0k
Drbq37ViT9dGDhz8J2qGcmC19BdXpSiqVARsGArR6ehAbku72qbPIBReOi53zguePcpQPeZeb8Kp
zshDwKj1N/TV/GWWEPZqse2405aeKo6FZ4UJvKITFYJZoDDVC5gEzuAgkJYS55SkMwFMJIlQm/l3
zgG1MvQI8WCIst1zEG0Z8FXC0C7RCN+lIgJBwtbaY9amLn1EhWMetmojmNNubGUsRwdx6NgX5Vba
mzV44z3dDID8cAz9zrxR6+9gG3AgSWBp/wvcX2Shxl7MixG2zGUDQkDfmaR1BruBN3/OC79Ps5/9
J/dF+AcUsYqy4RY5SKoVAwNhQmymRLWhRKywrcyjMA1lHU5KfWpO2FUXQtvrG1wVgYo/7T+1g9vu
u5sX3AbmQzNimBb/NA6UW/CBRnet0ThB0WKB1SdMVCI3ZQ1E5zDiISMxwfZbjsjDywD+UN/aiMan
u2X3vGGxmv4lqOHBTYaCD0/Z2ezBGU5NM29mkaOdXbAMfrh8fNqTSmvTL9IDNKUfzMFImKRwZkHR
jGBdN/d2KsAj9cG6mI/5qvJeWJu8m7rLk02UWvEvNGb1gFM/gDYFt27wnz5zKQegeyvke/NPYj7A
OhCGUu/ldAhn6+7itzNRW1k4rWVzOvPvq+wo9Jz/rcO2QohNLYsaBLetazrbv4VQ4Rk687Tb1blD
dYGJJOZhwsZd2e8BgCRZbxHvJNdEC5QHVBSJTcQ9oBFjrl6uaUHVCld37dT43jLGIHByVY/MTIQu
N8SrMx/I83cKCSlZtLx7kqoQDlhl0F8E7aPQqNGZniJA0EO0VbJj/wJ3cHp74IbzfE+hpR4Rfawd
4HPs19DJjpO39q5RC7FgHffqwoeotBn/FUFKs3SMDXThdAj2L+VdKfpokBXDIi0eDfY26RZfiQu+
pwqkofd/Eze1+x4l9F/MV34wuadXzu/2GEn8dUdNW6TyjpLIg5sIAYfSpoaoUwCMbNj1JbAgaNT1
AEuZ7KQTZOuIel3L/9AovoKKCK97y1lxSvj+iKgmQW1F/AlVvmaprzRi8f+frUMZAjZ/aIxF5SI/
U7E3Pa4HNCvFY6FaleidnMrawg4lt9p6P6KektVip8qSy2ehYxopJyjfeC1kgbSE05jknb3jj07x
SBCiFxPV8J1InzKrkpJbp85wFMLk4C/Lr4pHpLGh8yoiCvY/z/ruy5y/9po0P1iJqotV4WNUoCZp
B+3e4Op2ciMk2l26zA/nLCUFrwYdD4XOt7vXQFKDrsAGdhlyJd86MLLusmbidNHyDv0GI2nSc+gK
xyfWQ/76s2Xhcm5Nzo18+aGw5eVXiP+Hb6jbAXyrOVEVTweopdpFucMpSG3lxbI5T/l0XzjTnKJx
CQ2H8pHeTheoR1d/ZSjuz3tiVz74BpRuBf9yypOYAbYAp7y6Z0d2WcAbzYj5bvGguu0Zt3Yc9lsU
YqcIw8OKvFExqHGCUKnrZG2I9tfq93PjhvOQs1/H/+tCnkeDKyp4KmHpI4cM+7OtxhSUuS6jPc94
UfIeLRc/EI/rfXunRlWIu0xUV8mXcs6cl3sUJzyGwPy/anr1JlN/JwNpr60kfO1Nf8YFJGe2hmRg
vKa6Ve92B8FPN3yiaDaMvZhUdFOSjJvhWzgmgm+D+HA4cEHCtHXZn+vIKH//iKgHZcJ+JZM3c7zS
L3Y4vTrTH91uLDYms2cTMazi/+qKIAx3dFMNbDtpUq9heUb1puAe9IDMjCjxVnTcfc+Ky9cdKFko
PVRaTpifGFRAt821+D7TvkWjzXjtCYWUgI/a+pHPXGGjWCGaAqWw480cP7opuU0BwYZ0GbGMzsua
rcJzA5UH0mtuzYPb806Q0DdSC8wZI9jDWl7BvrfhFZqoQvyoN0ZahyxC9ihHrPN+By459Qk/q+in
OIFcjVuoMT4E7yo9TpUhL1uEz37DFLwE75aWG/5DHZFO5JTd9pc8BDg1vFDm1AZwiXwrH94AlmdU
+iaWvloOpTE6Z8EIMjUx+pGSIN9sAXpWQzYX/goFCI8YjRxFIIlGCLu7R67B5ig9Pr5UMwIiZRO8
6QiqD2Kd4MZ55q3ZW81h/HTtD+88GmV/sv7b21oNO2T1LYnFupbuWCgY7jkQ6QnfMJ7gHe/pWwyo
rURGj1XrOIk8gWMdlnIaZphhpnT071V+aoeHioriQZ92CAsuEg74Di5g8GYGC0rtSpt5JstfDLgA
vLFabMbRbfeXuG5v3VI/1XMLG5FTgpnwsMqDRNpNlzk/5NWLCyBQSzu0YPtkxKWnKT/EcWnNMFix
QmU33qkMyBzJqD/iD5oHC87gLZltkzAYdlK+PjdJX1TyJI2xEYvYCDDSHnonrcNuJqUsXYNDZKud
aVg9K9+5lqUqHStlxbQRIqZXA2eb7aKTc04ouflPGCxWzhxVaCfRKv8Twg2lgIH3XG8p9ciZcsWE
xVejfp0ZwJW9qqMLYoHQL33X6gycJPmZDb+qwcnuqhX881toXHg9X+wCKq9WYPpWN975OjQWXJ2g
J9qS7zDT22FmaMYjG9MheBt3/voozawhVPZdV0xKxiX/7lCAoHOhO+I/fyX9VOtx3lEMIwzitAKJ
tBe5X0lhgLLYf9X/vRg9FD280HchvOr7AFUbpf8cNg+B42H9U6WISj4aD0mcxCxFn2qJmHpqRab4
lMC/p/VRuRM/pPQ9YSW4GFM20IhuEUZH4Z2uj+RYojeLKklP15o8saR8fQxiVh54OponpdsKcNjZ
5ZoWm8ioFC3jL9+h9lmvTpHAXd7QOSy0FpX+4VzKWDJ2Jb5b8oHA2LRJz4Qgq/tZQDKEH3C4hbTT
aJVkpqwtZMVJevHPLMjA1n+t/hegm+r9qoCzRpGdWms8vSUZAv6LISEZdm4f0oNi7g/HNY6Z5Wth
5JJAv8LlCMHF7thmpGHWvMj6OkNnYCpl+n82FtgQPh03dEruFurzVXLaKu+627g6Fe/AhoAr01TJ
KWOD3qOMzg2lWpj5pkvNOIZhLHzFQIofcp+5+FiXHY6PYo/wwe5fta2OLKe8od4VMKYA3YFcZ+7k
OHLHjBnczEjPym38CRYfP7C3hafzEBTMZq7qzD4nejjqpsQ5B2T8QgOYHLVgj75Baay/Mtj7bB7p
tO/lJY2mElLMyIKPH/FNXnfvqZzjFJ92H2Dfhym0Ew7an42A21gc5tQeNg+FqSJkbC5Ez/QLD4eZ
TMLKIIsN7gIzNCivb8MEANgXKMuue+r7bKP/CoyD0/eIAWNspoLgyDTmIcExhbtJb2s7kVIURPGh
nujXXhx0r4rp5foRConRzr2FNEfiThYC0J/f/zGNeGTAF6XW0/RdQI56tsBY8j5cKExwzwsuN0yv
wM2w2fnTQGk6rcifVawT1LABqZY9obtsj8465CkrhohqShFbl5vysReyyBTr+5Q+LxsSHAAnB6oq
OpYCseR/oQncx6xuwPzMGRN3WV7q8OpeWGe6d6Z9Yj9id2NQJ6TiNRfjfwh6FnMVDyTCWooWHaIB
QRGFSbQWvZKL3BuxqVKgTpLd64LtUu0c/mU+e3ZqeLTbimkaKL+Ru0+hfiLj4Pg1yN4S62SPnrYm
dwgTUOFGBjnZrQUFpE1otBnh3r+V6sLTBh/n1CSCdtO0NBojtdsftRt4XJks8HLOr4nWTb02WL/e
7QSTYdawnDpnNJRc5TDZVmg2jl77HX0GVSHNuKYBdLc6kHGI5IZ6znEKeRSHhvQSRjSpndODTXp/
GINLs0TgUiaChu6T5OVjk9MeE6MnAFYpmty96OHTlZAMl8Owqq9BIyrDe4+5TwaFnPMJr9WKF2nQ
EhW5VzeUafH+B1YWAs1KiPNvETYV4dnfz/t7WU+AZeYgnyhVICEPBop50ZSLJEWUS3CAxl6NTQSB
L9D8zqcoizBhPeVFNklAqmeqYXsp4bEURC7SPx43/AKUFU9kKHBSuMaqhC+HSGlD761TF0vc/cQ1
fBy96HStz8WGwsShg6EgLPVjQOFrNbapmE3deiwfwV8ZNRvtOYMaDJZjGYyMU0gHM1UacilqSrNT
VvRy1cBlwstVKXFp64hK0pYjN0C+1uUix0I535Vcl35BtI3EluI7iRShAZ+FT8Mpl/4s3bquV5GF
ez3txvqxns2hcMKIYbHPFDNsxFXs7DUkNBYUPHTjNwKS1ftqA4tgoihCXKA9er67SPhKp+rwbv2i
Jxz5baL1K9DhxovNCgLln1k04Qk3ls+5b88gpAK8OS75nv8BNVqb8Jo7CK7lvdvBZgOMk75E14QC
cbJ+OP2LjfP9gFcYyIwDP6zs548Efnum6uve2npmODI0afA2ObC5zpRBiUu44w0dJYw1ZcRimaIe
55lFAVRb8rn5uSx8y9EjRpevEpN+gEQg6yTQzweNvQOvZ5pIt45c0+tlJa+mUK+Oe4Z95khAykbZ
UqGkGWPmlfHl7imdLjJ29k2ak2TSpr0d6bBWN7UzYBeah1VEpgqyfNyBpmoP8g6vV0v+kSb66b7N
Va1o7V8S5B533MWtSWhmsw5ADRZtvon/Wj8qwT8QXUYNZcJGXcG+hNyNEJQaCES5918bzW7cG2Se
+/2Da3QCRpkYYMDpdBmFBFAwcyAvoqFFVcYb0fsrVmyvNxnlIoVsHERJy/o3Y6W1/mbGJdotrHTx
aXfgalpvsjGa6IgRojl697zaClOHdAy+/9D/a4WtHXI3dttOPmYDP/6Uc1KF1ABS0+23E4DjQKBn
6giis0itsl1lTCK9ZozEhjWQ/iBRnGXdOVm0T/QVqqIre/BSE0CEWfpaCrPcrYaD3ph5IapHYjHN
5+CTqTPPkkOBATrCg+Ctay6D8KdT5iaZWcIiHlJzocSl1f4wjAyrY7tFqNSiTlaSTAIimGMY2NHG
M9DJEP90BjsXOyGuDlY5Y28hLbNcZsXbt+yQywp/RfgszBRhFuBO0Td/dacjABFOXFyh/+vGcRPY
ixvj0+YEjZkEqgr3Mxd6YDOdxiRHLMSKeokaZLWU8EB0OQjqTrkg+ImGspBtY472X604DwtLL47a
oatfx3rjciG3UXfCU6igWgoRnexJo0D4Bw6DMOkC7aYRUlwpVuK7/BXjWpjFhgCQK9hp1GK+Hphw
IMKgAR4855Rh9GPxldEW+0mGI/Po2BcBNtEnzVF0DpkOLh2UjLuZ9Dsqgxzn777L3U2ZQRO57739
rJCeGJDkjJGbCGGt6dUZuvrxUbGoaaQGOJgLuV2A2Ku7NG+ir5g017eIgE40cTeECI0f8W8uYaVp
w5wPgq9e+hsrZIXpF1pbGJtIXIALwi+/EcGTM0hVsErGYdVx6SVavKMBDILRdKm3641MRIzTqv+g
5f7nNiMOYN95pjfSHl2tNPWH7ykX6aDWzUTVCYNg9tK6mrm37QFjEM+mey0e3R3ivRI/tfwcSxkH
9Z9DgpiI1bwur82p23ew6+qCSaZ/ELxCqRWR4KqHAzeWaBtovHWgvJvN7mG/FePapb4XQGCMp2z1
qY6AfsOduR5YAaRL48pcQd5xAd2SlzyixBojjVgGNAiY7Cinka32fnbw23XEg0hNxZfEGSLV7/3s
n7o3CZe3QnHRia5+lIblJ6u+TNLk1ef51B227Izx31RmrfBAAP0CfbVCbEQyfJHhL5aqUG/WWdiM
0aymO21kx2oe7A3hquBcBLmhflx6h7RfIp5ztoYyl8xuTiG/CmMVtxCDoYsmePFbyKxmHv12/slq
rzXiqaE/mTaS1U5F8ChqVYpf9Ie0r4qLlII5uhYJ6Kur5jvgjWYxtuKrwDisAYv38SrN+tR8gmra
NsJ/SZKaAXPjN+2mE2djayxarQzUri1auCBuoOdS7TugNlcXc692wFVZxhxTdFYPbhbPFbj7BsGA
p1hWuGGCpfyuoz4V5aaKPESNgaNcsV5SiRR/Bm5Zgn5yfolqirNSyvWmwxGJNQ/P6MsCJPM5Gpog
qZxsJUDz6rcaGV7MUJa7gQp/IAzdEZbU/5FfYoQeTn9UQxy+GR8fb30t2Oat6Hd3nA0+MOZYWnjO
hniws0Ydv8LgNuTnZuUFH2VtvHtA+M+l+GjJZYd8UWRyRQW90koBrTiwbsXWNTKxM36NjpJVraZt
MTQaw5lawR4wxtYdZtedBW/JCvd6TspRbUeHK3Gm3f3fstWMajWKFAKOKfXAoWa+UTa9dzzViINp
UEJ6HLwJ3TjTvm8T+T+ebepBSBM1qtDJZgCgb5z7t2KduJks4xgbxIFdCyMKC7L68wr9rsF60voz
yL9L1p1CQnyN3TGfJ60pAmf5rcEyajhSGXS46wAQgmXVvsEWXYKcfFoV/Q94JXIXbN3e/C99KMFr
PumhOZvHxsNyaGqiJFZCuHU9lFsALC+7TRQ1x/hbrRKZukiQYbrJ3B6FJTIn+aFKTJuQt1hEmPo3
bdEz9yeemgQPajseoOGeWc9z3eShQjD/aQApnkI/9/1HcuUJ3nrVJnHprwqVz+z3LswJXVw9D3Oe
AC2fkROXTw+0PCgmfQvKMSTWWs4hQWIb4xrEQo+DAATi7G82Cd0BjN/cvOHxanGg0SAthrGyYSLt
QAWHIDnqlp338IDBSsInk8GQKXW7ZVve0VOyUNNAoPY/v3LiFdBS8N3UkDu/G6oMq4w2D+DbPo7m
1Sa6FKvTVoJh7XmbMbEZMmmkF9v3nJnwtsWxa1DBDuroJMAq4lyActLLN8Y1jSvqwKZOtnc7EfDo
dzdj2OGSfH4kUKpHtBvlrDwVLyZKljfrPbPtRZlxTItzXSKRqulEw4dqzQLKFzeDnKAlgZ9ajEna
ttBMg7qaM2ril3DsovqiTznPjK+gMb1LptCHPW05XMaTEYBiYXnHzl+9Qs5WWZ+/AbuxaEnQsPOk
ma+GcgSYiA90khs4JZ1Jse88k0ne5NyIz+YzIX2LmMheKtGvqh7XwItEeSXf1X2b3A6o0zbjRRUI
ReEF1/5jCpKJFVJsoK937Vg9x21nVP6z2W2eVaphwoQm8opHrdX9fqDhQzZ0SOUemjbbKjmOATgz
6pm41z49IUgiQKus7z0deS0xmEPcOYbBxVb2OkfKmNDRhAYxetYFQ8ceb1HiCe0WSVuARGiLfTvc
Als1mvRT3A1wTgMdGsJmk1j8hOSDS18zJqy527mGxPILBWGy+kptFhARKcslKAOM8okdD0yGKSIQ
I9nCv7iZU7yXNbVkRbJgaClqp7pAFGlpqGTOSVK+yn9tRoPqoG26THSxsSIDlICqLYX916eGWxwJ
36fJD9wxi5hKwekf4eCj/sB/q9W9FvORK56wC+5+UMg0Oz5+7aZAtw5cODgtqRL5QJ2rTkUekMmm
rEuhxk8FGSDmMnx3aZZ67uBiJNCa17RJnkK9q3KaN7KxizfB7TWWFljZGkxAdIdXak4HP9MBjz3M
qY9q2B/pHp2kciMUZMr7ME74iJcYO+snsdFXd1+fMXI37NmbUY48i1YLOTCsC/uyT7+biB1rNs19
sj5+y3LVB5lVB4GumNI3zuMDun9hRNsWkOszeEVaBMilkE0AnQSQbM35XJwtwkr0FriRga3fnvXP
aZmv42d7cIy47kKwY/3L42j5HphdRWb/WMY28OtGZN3o8QGPN6KhDrcFDGGsZX7eAdf/Xbp0DWsP
G8URDRnW3VH56fWAgcdvB2IsvFD1SwT1MNDrA5cvXKWFrH6wZHPGwh0ptSY8Ewuh3f+wD/9OE0g3
uLEeBbJEY0CxkiqaI6V3R0cDACbDZQ4WdZYViv2ApN1+GhWGAfmakoVat0RLJmx12Ltm3MQWgE0z
Zxe0GAJRyA1g9cTRXX4XeLpFNdt19PIr/U9NCZCFZcvBi0j+ga/YIUjBonvB5P/GncKc2B86Pq2q
tQHFefcQced5On76H/5LFY4o67UlHC9iP+zIerbPt9KZPiw7ZvRI62wfu1S39T5JKjaVoYf7dIxe
yHTSwpj0vpU9JvjfthqkVyNN3icv1881ifbb+R7TRvx2KhM1KpeGvDc8kdbKHHCN3YCc7Bd2Jhis
W0WmxzMea0KFK6PyRYZM6TKALDwzHxZSFP7nRm3MPucITX+DMgSDFqHG3pUhjMaJ/MYzFN/ZSgfZ
hd72N/TEtn+BVYoEJGCcmfe9M/xxoujJFv8kt7S3EbhpB76QaqssdadaiVSWfL/8tYIY0q5UopMq
8AW59FrBIAio9xeOjkZ6jEMrK5HEXtJgZFgzO45zxyEn6s2VLfRw+gRNtAtyrQmZa3BZQVmiiktn
KBD7pHsf3lYe+K9ky3MU3e/pts3V7nyp+M68N13U3RMqXZDMZqP4JLHgzGbJTySUcFDKySSStqWh
iJr3amOYfqBR7Byi57y3W0Um/SSTMA9VbHgLsM31MCrc9gjaLH2yfDBtTawdbt192rjbpJUz5+Co
Wdi40rMx0UO/Bz6j4PFdMNPeGwRXti9uQfBlfKW22wPMMdTZ+cP6Kz+4Lk0NgA14yQ9wsFnw9bho
kErTbnIEEaDtQ1WIJbZQ9hdLT4YWCO84q/6J6eow55oOQej5JdGmWYmz/xlxV8i5+camRkR1jTY3
CsqzD7J529opM4Hx3OXG1PakhBXxpfvvHITOnIPOOTiw+ZgiwhAG0G3W3RbiGFESFp9LJXNjmtPa
bCHO5olc7/tSE3YJj7QJgElZWeQElTpyG5Edoqe7HaqTEL+bnDXl4lK1AnYbtS5IYB4bq41g1hvm
K979mYxQ+hlwKKYE+ew8BwcR1OqG9hitmJ7+leLXRzklOlhtl7iC4GjkvxkzwRb3FWef38y4Yo+r
Ptho66ZU0aGpUzfxGN7uq0jN73HK3Qc+GRR8reCcLdA4sdNYzUTMLXuh9uxi/VqisFo/c63uAsn/
5blAV2llenmnHA+ZoImCq1G91tEm/NZXfBc/ji9BxPjHTVEwiQ1M/yxGXyThS+pMFSnvB1I4Jjda
PRi3o9IY5Bq0uhlPRxZCzlpMctjcfFNAas3FbwCrsw4MgcoqMkMudDhIVSpbed73kUjkk4UXajJZ
gR3YrhYbqnNqEFGSh/sjuu3RKtcTGlanIMUXrP3TucuJ7c/F9HY6NOa6hEYvVuh4hkrX1IFrr3Jc
Efs66VqsZ34eazpgqckWJyqM1M+vEw9tw2wJmgxJalhMYUCony8rsHVA7ZB7DYrOY/ec/DYumJz4
bHUnorBby7jTAlbLiwfcX0gun8r2Ei0oqvkgSJxq+NLWXM8Xu+CKLYA+Iqr6hXg1tIIIZqQQaP3R
uQ1BKsprb0454AdlxrF3sfrXpTbBud/yyTYxzLstI9RhNH4NCfGyKCaZay4zRbbFiHYL6AYGdSos
Q0yj7d3TfjdEE+3dlZhY+O8E/zP/stv0eRYTQsE37tw7kLELXm7RNXay6udycIzIcybLTSu3gpAt
ybL22ZMqjJAj2fAeAs+HSfseKZycHZSqvemKBV9jKfbVjv9Y9fa6stS/cHQq4MK2cRa8iZ//EkKH
vw8Co+t1MT7gXohH5Y5WooU4KTK7w78DDbXOreX6FYQkVW4/beQy5XcPcNd/tv5FyWFlcfe2s5mM
lOLlENAOidRoGj+qH9aDNN2ssx15bzCVVfHf5vjKemJRBbV5DL7V4cAf6bGyMyeOxBxp6coIq/8C
iN0XD68ejZY1F75DzupkrkWtDszgY/5aP42kK61GhCPgWbmL0gI7VDbUqxcDf89SvDbLzW0yZHnU
tTI7vt2OPF69Fstn1dmpSvfb7AsCCmTnCr162yS2ux0VVbBpP1RFlAKF11P/ygpwc+Sf+x6nzc4Q
9lJR/3MBGbRABtlAK+RsR3ApVnamalfNSVaMSYMY0nIbc0rvphNyhgHyna9tiC3TuubqakcyE/RD
FR56vFlGOyPSEwhL50xKo4OmvfTaJvyVbRqFwrDH5CVZ9uANs1CPVujYum9kNejHH/sM0c+3cJdN
Q+VHF5nqDHY003nUhSfkX/4WlQcR2aLMLeTs1gbkrfRgV/QRNFBVixLF3MWMGTCg5tTRwn9FVTkr
B2C61pcUSU69Myq9Cx9EAo6eBIRNZ4LA1xPXV5g2erxDfYLUoC6mWGDPuRIN+wBj5d/rLaNZTVs9
ubDDcnhfybJvkaKwcGtZbXkohmjuLBv7V7GKf2dWViLPMc637nLOyYxVH87FQeAuGZb0D6Gaupf+
dBPHu/E8S6GpC1544aACqCURRoku8PqUl+uwKIEs5GVyxlR+Jhx2pT9pqP69I4ZRLtxFirzzyVuY
3RA7bQjCrSXddzcjhRypOafgphed/r2jzBZVm7VFGD3w7vBwug4GmdFZF71paAKfbUWCKnHk1f37
Cv0znMDY/EYGPYJPFxBmQV9nxfpGSnCJ4imcjovWI1dmZxvwbv0JndM1apXl3ORpDbQ5GHP1fO1s
QQ2voxeS2vmEoh7i+c9/nOWNaZuQYl4y+O2ClqHkysTZPQrj3Iyf8u+pQSUKapFcbvi+T6VtLPP9
4lYAmAP6384RWjxyNYFbrpjlfdEq9ow9SlTm1DYIzDtnygbVGt22Z4KncA9gR8Qv9mF5EYP9YVvs
OA52HZXXoZlD9HH6XnzRSDtYpeMUFpCNLyubRhtYVWmUPelylxON1tqlF2d9yhQnkpi+teT4gywY
+IwKXY2w/WYv85UfMu20cr6p36hcavSmbviS9P0YY5gw4vk40f+Wq0ClxWCFXzu6X/F9kFR1AQYt
Uu/6v4+KAlfdeWeknBhtvpjIu8CGb2ABHqRsns5TdQfGNdDsMENdy63AqeCUjCIORWaY+ds5XNjC
DPpKGRTvcf8QF5z26PtqMfNhQDLO4uQ1d9xKE+ElzgcEFZXxhr/LAXzV85olW3sxFJorT5mgJ4Ah
7wYSv+fo4hObTswo3jPOgg0R3IuffkScMKpefGbde6CDsORGOzSek2WgCtITbZKQIiW0jmtBjFWQ
IqKSIK0XNlUREhDeZu2EfWJNchpYuBd8GKKMRYTNqYQcgVYa5E2q9+Ssl/9f7sC0hFqtWN8Y3wfq
2sdzAhsMcJTz2OFTIIMp3scqcFgkVjvzerN1u1nQIfsoPX52iFJw2MBAGQoF10p28wK1WoHvLaCM
+FlJe6CrRuNZvrQQPefL9xUR1KuEqdPJZCl2FivEF+/YfML/3515t7nwCcnKWFGrDAVhGBW0IN9n
k4dZ1453cHLhqgAWxP+S3bbObFwiioGPcpeLU1Q2XmSkbaeVy84i/whz66v6xTqTSrHm1XuX4NoL
M9Xk8rX8V/zJHAQQkGw8CdfKOHPYd0vOabI/Wh97PsaNXSCq7Blg5sE0dpRdsliA5GiwnCwqUmnr
MqJhLrt0kZLo4wi/pII9yeJ4HWMwl+LjE5E1BqDWAGbHZqW+R6sA9mth+yGd+ji6ADY+Xd/Ui7rD
51kpomgzP5S+ua4H6QTliYHabqxxE3oMNgq1KWOPlEcZeWe/uNM/uIeSRUPh4oCrX8yCypfnjygL
pQVcQLOikWDk57H1Iwae0MBtvkF7cHzA2+v9XcjgL3PwDOjCtX7syFsEbEtPuczjo7sigSkcBkAe
EYnCRXtCBHVhIjKTUmSSfSpRE9Ywab2DKym6Dv0aWQoGShRoikoMBZpbVzuRgbjvReUgD40ikPZ7
glERVIVqCivOix1AWbqhXVk00Ujklg/xC6RozuPw/LQNUN8Un83cVtzPGCpwmvaDc0BxFQ+UD0en
XEWdZQthsTr/45Knx8l0g/iiNCVlHBoBI78rIqcUWsAR7dfTjEyXDSSAFeNNS0e+v3pL4JSy0HO7
TcZUrAdDa+4gktG3bwA1LDpcZytYCB7sJXKTA7s0wcVWmQxVg06BPxSiOpt0IURZv3igTooN0AGM
53zSw0WxAJoXpm7S+WyUB1LpnOf0h3gkasln5K8oU/Q8e+LLy/M8lKp3KvNoEQEvYEIAe715R5Q2
r0tmF3j+dAjhXPe2tLsDVelrgAJ6isHMuPCZ1HCSoljGvtfCu7YVmIoY1GgW1Q/08yUUBp+hRTir
GdufTGHQ8D/c69b/ADh71q0DESAWZ8IvkWLOZZF2sdiPkN36VAZD02dpGLPrsnuAAuGQCY8VI+f1
br4OBE8EO8j7vVToVRyVeNKO4kKusYrOooGR0fUdIyhN6Ta8T+5tz0uDqb6vVhelkeHezWtm8O4W
P/Iv8eaaDd9HFEOoAmLGdvb/ywDPCWAJO03Dts68z3CpCAKAn26Z/pEpSaIIndE7aYmyGGCoHjIC
VZ4EnV5vz/+aL7Q+ZUVjtdpGRYGSCAMQ3uZjRHBEopzx2Zk7GWdDW7HqUl0v5b111OP9/aGN5oHu
vsGZKP6aMBdrqHkpXn7zFtAGmbXLyBX5aaLGeTKeBEVa6SilpJ0rXh6j6UOpXbyQ9Tmnpc9Suec0
Ky1Y1b9zW9zX5RYrnIdEnKTE+yYkDTef3C1rJBkAy3yg5fRwTe3roa+Up8/ufbVzK5XEXTOTz6GL
zqTCTAmx473pDR0P3Y3e5F2iFDEiHFSemsdl4ZkrSzy3tgHvnTbSom2zxMbFnYwyyVNXfXevVnYs
nXyFuikT5X+PO96OLL9ynP51hG3p97wmhvXcfNmkkWNiCJPJ6AbDNUmSOBFkPCY7aQaD2+Bd7MLL
yfutJaWMkd7geEXXC/u/a8LxR7kHakxaL07b1CjY5MVJInZMeJkB+3Wd3vh6IjaTfOqAQWJSqaMa
A4PvkMlXGt2rPanERZ93lMQlV6MytMCN7/16iViHsy5LnWT6dgKHMA3c9Nj0uC0W5cZo/g343usC
AOXaTgMwr/mb5xW1DXEL96nI5WaArLhFAl4sBt5oGQWBYFYrz0/Y8I1smXmnQalGeI58vN4yD1q/
5ql9n2wjf2NLqSHu3bLItJfmYcH3TEpkevKHgovjjKekuwoPxkRNMx/4qI0wSM/UqBlUYbKgjfG8
MtklWRaHPyVfaHW8XgHrUVDcob6aM+kYFZU/wDqmar1PKCCwghsSLp9WfDFhllddJGLs9oxALmSD
cWXVIlni9NCHD4GkI+Hz7nUlnlecruRlicXNKLn9rV6QrDpm5HL9PJKQHxRZx4McMddmpR6JwwDl
T1kcWsTe//6r3H+qE5krtDssWk8ZwzvNzqSJrW0rwSBDQ2bnVXHtlQ++yzxMcNEsjNEYy376B8Ao
D9sTv7GctHp0zpA3BQEwYDIcWXBzJ2ySugPsFBv4T1iS1bL7TUi5mnStDPEaj+nrG8k+ZjaYDwsL
ZvbAQpcz/H4M2p8Csq61u+00gmhV70p+EDi2v4uK23pD1QiFsyKxmHGXvdC7/wc0ZivVwl+5vOlU
rncFi+ChudLp+qEc5CtrwXBCMI7be93FNE2u9YHDQjZIbmRR6oWDLm9WHHOKY75EWgB2OpwN37uP
QwyfIoHR+ehoUHhyOBwlUo5NHWgWtwL9B7FkT+sP8vD3X5beM1QK809y0SGXsjmsIEXrxt7UUBEK
1FIjNO6jnqh24u46D1tT0OCXuc4UkaQdkhEo3sqFMkSQjXwSe61OZWAOtiz4s8MpnIqo/Deu9Oqp
09iVF7Ga3/eIax7odF3CLfs072wt5SwdwVickVJWdHHhUK6MQQzIYufloT+YRFDE9ySBjbhlHuWa
Wv190flN56WGY3Y6Mmvxp8xsV2s/QKz5IXZBb051d96SUPzvzcitE0IO6BTS5xN1LxLn49ZfZKUc
nSIdmywcnuwYtjo8NRLqn0guglQpAKnqA8e82lEePVkr28M5CrqXIEp+WVoTALNCL/1xPqM5ea4M
Nxz8w7fGclZkCAHTHWFKCr0z45c8wcTTQLFflsBC6dTifAVkz7LOYqp9IRuwd3q4Yl+yFdno1sBu
y6mNIGOLLdAsEXfUpcpYu9A16smV583KTGmDTDO1gC7LghBue5cfZTJov1D+dLnpcupCfJv7Da+o
Deoq8ikdm1jVPYkQ2WJ42ScN7V7vxwYqEmuXvL8xwm0aUvQKEJDLs3muFVbxdNGssIRrG2BVQC8d
/EinC/BExZ6N4M7FlQ4Qj5uSXKCr33rDzalOW4MUykKYF8bC/NbTFbiasRUXcbTkWcXOEmQUqCWq
KSt2cUtb/8JKH32hMC0UHXMmutO0dhT9Da5FeNPvCyRXU5skPX2jbnzt+2K4Q8+i5NS5Gf/tvyDC
Lf7//7sEDCtll9qJs2WU3zlbYislNqJmHx4HDL1REvvghrkGHaGGPZMABgBP1A9XfYKBD11wJi6D
YgowxosZwzgCZpR+CIEsVUhSr8msS+zQBdLxULnnErqH1cBIlz+TQR/lWgVJujtj1hgv0h70HWyB
cthduYPk3o1eS5pq8vE6SOse+wGD5wMyfhCnbB0TLynqkYVFtz1EoRi5PHA6ArYyaT3LJFlBcaY9
oMugyOubAo+7jtvXkpSZODGc+JSTi+W4Tu633dpEPwbamDfQVTxvmXcq7LJg/rnqLRfJknZl4s1h
iRaHI6Fj679WzsiC6naWbOEMbj5L20JdDrz/RPQ09kcNB45mZj3MzmEK5hmX+wYfFRj8JPplkS0e
5r0pfhmYgT9ICC7JkncumDlfS5Dlbuzc9uTpvExJzrIFCGxvkmO2uGz0VHgRfHt/ZYAdR9zHdHKb
ZA1Usw31dlceyLMXsSSK/fH+LXJJrg3WYECD8Ko7p7kxAk7EBBuc7ZxQ8JFbwcQMwyLcrK3ZpEj6
BQUBMFpHpwUltKgdlRWlU8aFHbdXZgGwS651saDOQSCGgx5UGsRoTB3RvBRFxiDYnnwhmqF3oVeh
9fBAvLz2vQIKvwlj49yYwIhMn3gRWvMqUTS9+jIYaEm3IqxnO3/kkuatmQwIJhFu8gBl3wm3itON
dOU5r9BGxnu6cAMc32Wrzgc7ZU/amJvsXFgE2hWOBZYR49gi0aH5eFs5AhwKg7qcLnLJrKRzL3HL
fVmXSz5AsGsWdOeCbelUSp3i4ctUuLCKB9al7wU/mmfNPrtMo06yYoF3w8hsQ+rKGraEM+4RONof
07KkcvTVrJ8dgAXBzzZp+E+UAg4AwEVcGbiwYn5otG8pwaR9uRm7lZRWb23M0EE7U/r5rG8dD9c8
kNsO9zctMFACe3ktZtSQsgxvBksU0tOJjn72Yi11Q6SKgydQXfRORw9V2ZFwRCLMGLr7JXu7AzP8
V8lmoiMeeD16yGs6X8giIL7hn22sV6JVeFodz4VSR10kT4DXa1A4+PfK2m9RILCD/UsNeYmU6kbF
vAyjIXTB8BKa/3tBXYYhJMBIWy8M+Grz5feYYlW5tQLwQ3uwjEQvqEub92+8VbfUPkrK169YLUqy
whY873s2ygEMv26UnxoFGFgedwznjiMAcurWvAHfD/xkS8xw5+MucAR3LtIzCAbr9YesrfCW2IIp
H8T4t2lKsiKvOnazEcmkRtFKwLLlCxZeF6maPj3rp46E+C4J5m3YTqxvSX83fQ51F4lot8kZliLN
2rTw7PnHd8gNmHWkk9IV8UHfFNpTAV0sQ5YkQOvtOSq8gWayw25UX36WNj3QKWzuFGguBmqeaJwo
Xi7sLtEzzBXz9Uab5w0Xi1X441IJbk6nOVXSEeO6Thx+y6mbOXI2hOn+9jicnGbzuX3bHMNQ/a54
EJnjj4M+SGR9zEl4NYJRUCziEABg+/RSzDv8IJ+CW9RDqLm6OYIpsJdj7IyQYF0QPyeSI13+zrJs
dB19WqbKFeCR9fiRs8FLQjUELxOmMsiWRewcwUBw7mXOLEVjpTNACEaths86PCMR6h6yPBq9E51v
Oypx/4V5NgTmVeBwIYgRCgrUp9wFT0rMPii6xp7IeINPJ3S41LuD+BjVTXjmsr6lID3FQDLrfTyD
HFh+rCI/Ag8cmsBKJnBTGpGQQgKoVAnRd/EgTVObw9wXCC4KHf0NHLiphCI0OmOR2PQwG3+ec2eA
OU/u6sc/fWWe18QAHzpEwywSCu14YV9/cQmMzrWiQpgAxIKdfklWpYoN/XIJH9wErp/e4uLmfESM
7wM1gD59HcroeIh8yGZrGp+4C994U90LrFiFOJmShKFJsqNxzjElYRZtY+/I4b1WJU/p0vP9KI3I
rHtqKRZu+A+tbk3sleUsDHvWIB9iY+MiTpMemcvZKz8xRfu2Tfz+Wct5BwY3OEOjnQLDXznYPB9q
0AHINfn+TsdOiaHjekKX5OGPj2LlFVgD8fi6PQGcI83cgeiYUn2+lDmZCOHXUSod2draQBcQrQe8
ycS0HHoEVvoM8RNL0Y04YcoDWJhUK+G7RGnIW910NdSakbv2ojIlYu77JRm0vB4e+nvglPqFtmN1
CUO+mwjDEkyLz/4BO7I1DKyJgflXjqznvHt0PnYmlZLNJozVCEJuURA0UFiPrS8orjU1pJTOTgtO
xuB7l0FkLePMoEURNzBoboq/4JxHPfRcSnTwMY1nlBEiSvjOLhj6aococ/ntDz3jeVNvnbM4wpvv
2zXsq7FSP0QZX7EH+spECBrmV606Bolq1quJ5fk7bqqkmEStsm6MHRtczPMQ20A72EnIrxEzVm0a
pY7At+IbkKFr7gQzDuDnemxCwwXm9Ozz6qznP5fnsTr4GY7rHJO2SfmC1SinZqPtpq86MlCrVQj9
/dxLm3SWjnhu3MDzK/b+lvlwWY1MBAEo6NioEpLBH0OgQi4gyqvKnyJmerxSspx7aYR1/ajEVlpV
/RuakHPQCQNfuHAKn9msHsgAOHy2w5kleYRT+81KIHjJ++g4hdu/0aA+JfEvNnMWKCVFlWptpUDp
Xghmwh54n8A1Jid43058BKUc59r8nFdRTRerfGetoiq7jl5Gm/941v+yQtZMY+NpxQZYQJ+zmf9e
Xjjt2B064mRJ6vbttieSXVS5f3Umm7B630CeMW5P+L8g1jrNNUpolfdk9x32zGU/ZDXCC9YDwgfP
VO4CdI0xS90b9TW+4eQbjpVjcLvnvtTZTxHXTQBBHI6+XuM+nTjFzVLJlSBoUjDAEjsq2VjGbhYi
daOYlE8nhS25nxMh9vwZilZmHuwV4aJ0tFQxBqpGdD+3yzbhV6FihK7kOSsSKLsqjyW5ypx7J7cp
Dn+XOc2B8ICiISEGZrWaEjb0hop55aVTRhDNFvZUMboskFftXq49dk+mG9ErmRpaBdzhGntsfN5l
RKmCQPou6sBfUrOSYdHEZJ7IkbvzAU5mcAVl50fWhqP/ZvCfp3989tYYwfXZyH28mwWZobeYcFIk
TBWm6ZpM29qYqmepvPzV5BInpURdcrXfYfYuwwULHCuZYTsydkR8lpBa6P76vUd2whmzyoaY9hjZ
6DWjkOms3eVxFllMhtX3mrROl8P+0RxZDTE0g1fHVOAbCdxy+73qpR+aEGRMzyNe5eq0A9XCocvl
esj8aZdBRxNDqNuN/kdPjGuRpXsqAzlQnZd/PkHlQmSrwZUaBdKLmCddGsdAwJaFMtYUm1XRSBXB
i52IvirO1ca97FYoseASh/CocOhGu9m9UPyyrX+FYKIfkb5M+fBqDLsHGXqH1m3c88Q+1qkreDRr
1aF3c/zCZQN8LElxdInOTDiYVPaVdtYo3LjAHslBd4rlvjgsoJ7igFZF/ZUY/v0DkB8d3HVqZB5t
0JyyXKg67VT2v5MdERuI6Beg9ewPNyferUB7PDXAoRu+FsTCcyiY/Qass7mbeROoMiPPhKI2cA3d
qPbMxuiR4cbgFSyJs+heVOqR6IJ7Gf3b/01Jo4kRoDSG6Mw/4/xkE83mlhHb4KxsjkYWIBEfEBEr
7Kd9BBYusdBMm3lGzOYWAzpt3wYab61SHKL9DX4/gI2ERa9TqqRghQEBwKJws0Zhr/2jPSgFxDd7
pv1+qX+9NeFSJR+9m+6xsLQk9xEIlz/omhgEGt2dt2EyG7xwdYFVqKze5B0deIwTTZybqSv3KLep
zmD2tpUNrLOEihBhl7ie8TOqYaW+08VsXY2KRtbbAfag3CQjhrqKsshJDVrHJsnbasQt/zsZDLHx
pgPR+doezsGwjFuUpSc/od6rmH9dibU1uJqssUmY9LcpZpPdgj+Zp/khcKXQGpy9wiYRLkaAh+ig
J/zTOLYZraIa1CaolCkTZg84jw3kYM1G6N2/We/LZA/GRzUwVU2y+b4RMh0zz5tdlqnLnaevUVhZ
zFQfCCva1YpWhX2VaImheb0sTy4ll8e5RUdXY1J4bZmpglvVk19bgGBR4dRa9jE43W9G8raMxG/O
sUHuSYvVtvju6qnv9LGHpGdRBkFd4vAO/f11W428dqaqFI5Xe0wfPBu7Yzf1CB73ZcwIxLud0k7V
chpu6/7ePXCYLHXlOYrZ50M3f2GGcWr7FfAsONQGE6PQ10W8shE9dMOpbxLth+9uyvFhgO4tVRor
oocfZezEm3zdauYFt++ryBf6fUlB0SIAkoqjiArqCVHdW6xNNKKmiMVIRGDqCjt1CZjS28ErIJs+
OoIbHesRuCnb2XmkBxnqvwLOTkg69av1K0GVv9vxWprWZwHOB7E8UyjleqTseKk9prHRxYKpOFLb
uOc+iaX8CN0n9iqJYqOWrnQZfDT4NxUUP0Db4pH81gl6QeKoY9KK2KWaNtmr6qM0bInUlnX3I+PP
eDNMJSr5j4uc0pFeLfLL9EGYPRBie8NKSLe3PAuHWbGTgBYgtJDBXDZbYWRKSwryM4xSVohEtBYH
51UG/1NnClrIJPhELl6tM/7otYrOEIbV0ILkiEkNcuj7cxedwP5jE4xrXIiCTQE20mBwrmTK2FUd
N9XjDgCZ1rFHjJI2t9KzLjsX0Q3IqLOULWaCUGqEPb8U3QYOTMEy1lFs3Wpjhpzf19r2+vWf7fDp
ptO7iBJeZZ8ngLOJo415eCOgPZ/X4PTOayK+mnQ1TxwIrO0pMd4InmH9IJ21X23w119rj2g5MUhq
+uPc3ZOG+uHXMkYRANiY+vcTswJQ6bLVO5njtSgw5CQmg1gucqFbrcMgFtNHTtVeigB2qnDfxJx8
h7mTjhe2ZPsVsrQ0ZknZdWj4OVwCscPwCebbCioPNDtgn1C5BYgHVdjCI1xfcYZYP4bS8PY4yGSz
NG6IDzMlhCUV+BVo1njNksENKPCjhTCbg04glbU3WAlA76Znoi5USyvN3vIwEAMdZg6IHObzIfok
JDyl3BkW6tAsIdcNaC6zp7fpcO25OyuA78V3fyZipfikoonQRAsTnBpLxkM9H3g4ra+2o6pLzcGi
LynURECNvnHHS+U6HDVGhSx7X3+4t/hkL1xmYaYWYm3yvnVeeE4P8oyAbyNedSIcDmEws8a6ZG5G
UCn4uz7rNhSyvvGeE0aFK2lTtQWdzOmkhBAksQdXnmdjOvhahB6RQ50ykY/jvvGmCQZ+xAKTXOdS
bSrHQnS7liN8s8QXGpDppyxqq826Vp3alEF6bJ8aRkwjlwXkFv94UCg7MVftz6WKvzQbIBjC/biy
8ow/g+jq/gLI71OXKQtnOiDilFsZTRe8A6pu7trr27HCkJzEL9M6q3UwksFSjPDriB5KfsU9ZsmL
+hZaMLGlvpSVT5cczbHNxsC16zaDclzFsWjVCFE+ohOjHaRlI+xAaHVMbAJBzQZDM54gs7rj2IOH
0JfzXER6esFKytCfeT3A347shdb+hN9VHQFZu4HwUmRbfMKIMzmBJPyjmooiBh94mAgfCRiJ2Iti
66zpgSmDg8upm6pCwJDqx8O/R8JIY8N87vVWDvEAPlyzUv+8IMvPyqd3qxhfXiOC/PJgyfsPgDyA
++zsVqdgjFscvfJH/FUTw/v/NtIDeQozqR2jG+jIpObaKr5sid/IGYXxlUFPdaNRPO/YW2aW9qmm
QpT8zn+Aw18ZRaGDTTQopn5WuXqWI5eoPVt7fzSMUpVCdTl1XD2YCZyGLLXt/leRLbZvHSvQm2mU
63m7Z1SLoFD4ZuyoEnfOwhWlXA+OtA+OuXpT5RWKIbCIcNyj4MUvkAP5qMpeM3ssS4IYrqab65dW
5YFVwS0OzyZbPd/UzS3ym8cYueP//9q+E4DBFzPDpkHFcXQm9+4pUkCUf23YaeHRb+Zib+yrPprl
KLt7d5tQGhpepOvJNi6pxqssl2CBVsuML4sKcuFqL87qm3ImB//EPk93v87AzQYDFdocUpEij+iG
xLPm07HGrfOzZE5OpF8/SOpDVmpTTAAlXomF0p9K9Dmk8bTFWEfv4xbljTqt1+y9Z1UFyrRgvYeZ
BVcTo/n6DPyEdfjk0dyhLjkWZRK41D0yq6NKWSXktdNuZaKviz4gjDls1udSi3gski3OECfX+6Bm
0eP9NfyiFn74EVrAbaastch8swx/fa6uhotmM1q36Qcf0XHrfD8V3BX2V6d0KqH54jB+8Cwz5uI8
Ve5OpyPTd97ZH18xGf2knmE/6E7Y6fphSAOBEgLScP7lk7rwMa7VYIvkLlPnk3W8l5ybWCLQv3lC
mlPxIXPWO7EhNDYWuM+ViDwu1Pe8Ny7UBHJwN9gNES+5ENqekdn4cV4BA84rfgxsVt4ouOc5pKc8
QS4UyrwY/sIAPL4/fWiIRhebXh4yIDTz8Y8MhLAHNGQkCz2UBPWx/tMcZigfiwYho7bpPvWoieiZ
bsdKjg6AEw2ISqJFp7bWMHmZRh6sirTDCt85fLC+IX7RAKW2sEwKcx0M3E8E6Ism2w7V9sUNJsD3
9KZ7fk/NMa2cjNJkLroSUNfGvYfo1CAg7ixN016O4LRHcwmrHFVN7MpCZdRWC6ycNic61g2nrP7v
gAuqvW61FbFyocVAF/qUeIjZOI0DpEc5aVj/WENsw36yyanRjzwwBOlTh1cpa0Iebw19KeCzaujt
BIGXlQG+YxDzb4tmlwMeOrJji/ny8yRrtGSXEBWnwg3IhaBAVvR/rG7UGffaAF8UGqORuQ9LcSw7
eRTUD/fX/OsQrTXAjvILeJCLslRzumzvrZH4P9lnjEUZTmnjdeZknw0CXeyFIOjZ/xK/ydD+3jaZ
Lih/hAIb8NkvgJT+xM+omLnMb+S3178KmbQFzRGOMtADf3oiLNphbWmFfaQ5m0be/dP/BB14RlzY
0jTATBtgsHKLT9P1xXHTPcgB4j9o+Qb7pv8xTqLVmBFunyq7gDC01ZSO5lro7ImMz81uuY7kFTiQ
gC+SIYEDNuIX0l8yMRGMG3QALNfRVyL3bkIGDb9HXVTLMoue8aOXO9sYo8aAltIuWq9JVfjRLvZ+
W1AZkjWOL+Ap/TvW1KW2wWaQZHp+js1rng6yHiaW76P5/RmdAV8DyLJCt3pLWNzDNI64exBmuvHy
AE9GzK9hj3KbcoeNoKdMn8+pArl8tzM8AYC+HjPXwaKZRmktuuFkrQerH05Sh7HrwgzCeigpuhkq
IUrvdh+r64eWnARWJ/I3y0Cd8b1OTDFGF8/spjRF5X1P0X8gC/w6zF42K0EQ2XnlftbYPiaYHugW
yODlJ8Be3sS/l07HqJcuJgymryGQ6N/uaK2Ub/yNTpmXS6c+A33woFmAlPBSyqJSLcnNe8zZukWS
rLn/NYpblFLHcJgKgUYHDBRnnb6o9rizpKkaRIwBZuUjvvFqI9xZNuXHdOiX98Eba02tiRdaQp6i
62IYfVt56lh9BO9rhRQJWmg+y9Q03GlMtAs6xQMG5MVa+NDI2YhIKMfKEPMFmh1+8g30IwYxBw97
QyJgDDthFeMw72ORcbDIBLMKyO8gqBWrzpY4jppTD2S1G38wyL+cf8Vw9z0U7jxenRoEWF0dt0t/
aBAnRjw5CG9C8ywElD/4+jkoY39NbxVFthpGHdrmTzLlEwfaiQYvK4Sbve0PeaRHIZhJlUc1Bh2D
uIg8d+z4XuaU2F/R+Wg/PZYPFENShLRAODWe8MrImtLZ4IgjLjpUmKtM+E0uhq2IxVhV6lFHCZvX
h8wRdP5ernu+yJyC84a3t/lVXPVk2v/HZP0G8txq7/Qi5MZtJXBYX8ijJl31BdiTRFTDPanocPua
lBG8wU+RSZ+xI5D12NIYBniH8MpajYxxS5RHu6baxZ0h9QePH6W7VIoHb0tKjtJ2rPrIaeEqAlqq
pTNnt0YdLAOassGXQHR8DqQnjLIDxH5Ew9R/xvChu4Vwctk5YfWJMXCXQyfXNMuqcUOaE9Ws3WBz
h1x5q0vIIgXtl+w6VDH2ShYj21L/kWD95/vDDYF//eOzH1To5/JWTZkSx4CtMMyyWMFa2nusgPY0
WgqS16foLRw3xHhkSN5i5VstoQBZTt+1oFdpCdy3cTRiXLJgKG1nJXMKiRi6kNlptyHLH2lG/lp4
TS+thwPl1n2UxwQgSJBEdZjvX21F+RILP44EWHudR+CB9wSOhflDw53vohBwdXsc06haJEWyEUyg
6FjUk/aihyi+Vdk6JThaQr5vRyD6RvPN1YIbh2gMn5bltRoUyLaz4t3inA2EHCe1z//IljpSqkTj
jKN3WdlpAe12GhBnoZqrB32a1KcKdGV55QVxAarTneuRE/HBaw76XG+g5hJwHZR6/pTmJBfoDX+R
qcNUM8Hxdm16lkELbE/Ppnr0e04PcAh1KOm6o5M45DSokfxanhRQZdHsvxRw1dPmSfJT/F+pTjBy
uQ/DLlJxJIFMPBeYlbyphrMYpCE7Mp/9seDYjrT6sDpAS6z4wYYco/w/Oe9qDyRjv5KKVbiy+aTv
4CCCmja7hy2KJ2Y8G2ZaqVm7M5eu33uFOODZAhGfs8JzW+mY6Hq+uKMU69eN5tIav67Pq36EPmSY
qpyGpphOtb3sAXDoYvKkUXWRZaXwpgsyjAkYb8w6T/HfWFrBPecub6YbUhD/MTRnQiY2Pfci8+/w
Lr2bZLbVpqBcvsppQuXsuW1VeLGiBp0Hy3//0jnFsWYhAuslvt1B10om4bx2HRSzgO2I5qx3UYW5
qpc0N5hfHcp+xl+Rn9ZDXhG+97E5zkL50Sfgo1ShPS05u5NkOuQgNIBZFnmlmnw/NGyMGYAX09Ae
/uxQEn1RSptZo0cK6Ze7yifRz99yGCG4k7whQaz2/TmuaL1niCZN/ORXa57Lk/2EN6Uawavg4ls+
CVR9Ri0uXxTfxgnGo5gLhgvuI60P1XH0a2khpyeIhgcamViY10OVZJL1mKzyE/jBS4INbDsNyLyS
cwg/1Mr1GvFdDsKxooe2WSrGLOXdQoOu9AhiNKeGziZ5LsLCWhJrkmUUKbKuLA8RFo0Re1OfW/2c
xI7jk6gYKaQHWfOViGVXGh4u0yiEFFoMkxK3AyzfgtK57MwFckLZM5gxcUqGuS2UTZUtnNdL+1xL
t0LaH6xuPGAIiFr1ZqxVNa57eyavJ9wi3w1i0d375TFzUvP/YJ3Po7jzXtHFZ5hTgsJDhvy+jC8w
wmGHKgyA9I5V53rj16147V/CVEAQohdIW/uNOiif8M5EQe/m+E79vikKBwHiY+0cXt3efikwxip0
RZvq5z+ThFMRe+PABtDc+lZhvTIHXRTFxSc4EOks2hEczoWthH9R+b+GM4MPai/2fQwDrjWQNyRX
hOjuINqavOk03/vcpN9sib5xGVm5d4Y8vy9DXb4i3MP5fQScWNJOBOVKsaUCf1GVRJ7kI9F1t2kr
2zYrNeVbcwH+QeCOM1Mh8/GYs60m9e0VBj2TDeFN5mLzzgQQ6ARF2VXp1uIT5inST5CQh9elpeo9
g85nEh6dfJgyQFvqnFISgnZ8CrH7rBS+Z/01t5eAtIM9dZMyU3SpOApH2dSlrVZSiRi/05ZlY8KL
fN0LitSXMXtGhZ8YH/l9NPczWnSpUL+aBOWYPUuIFsvNCDOm/2HYXdmFm6DaVaFb7bRmiA/0yl30
SDe4mPSr2RC8TUiG1Q9hMmT427oBAFfkwV3q9oNIX+MMxHrybQWomZe/dftuUOTqJFToS6vIP9rl
fymd8ypS9Z7sAQt36VsLFiYVwgF2oYdDfmbn3DuO2wLP96uBf6lonbQXS0SauNXvAnz8gY4E/QKf
WTrJDgePQ+qCD6H+69APd1nUi/6tf/AeUskoWQEu+N2MfCqltfDyg02XjvMZ/qS8eFpBlrrQaAq/
zftrJ6d3J6tS3zzCT1zRsmTSlz6WTt51Y4rWyvXtmu9Njds3WfcPM9qYm/u9x/wJdeY76Eb1HBnr
mNukMsn/kQhbfm6TXfYYkbqyd2AVZ70FInTIDx5GPIS/TvvE9N7XpN5TY58r5t8neCp3g1vMU9uM
yN+wSusDaLF86oje+8FMw78NakN7mOcWvxKjQUbrP7qYfoVIOp8tdW94ISmTeTLUYFl/KctNEgdQ
vm6iVOQ5rM9icXkwHu7hWra71iyQKMhCIbnALVKtW3CLd5NeF/6wF7KjlR1c2fPG2aw1ORLNDZ9f
ctLH2NXGXPG/AZBrfF6SdndekAggnqgYttbwJK2YcevIMzSnOPJFgxsgq4hGDvoMissxIsFeudId
CufWGEQMEUJwaL3M6738SfQ3kPezji1HKOsDHtWR47MrTEg/f6WRT3ZqltWyD9LyqNZs8nUnqtum
NB+bUHDPlLeBOE+sOuKI0Kq5lvtuzqTunB0LORlI7PCH2ZEkBZnF/BbchVIjFzax/GVnz2dudOTj
OxXq/yIqXwBwrup6t3zN3nngkTfFXI8BOa+P73CA/C4aM3DfCLR0EKOMGnHxPGMTL4XXPibgKvjj
jCOoMWV/XPbit5UKRGa43V3ekbFJP7xONAr9/fAzn3RczHwOaJZEybfrWaByHKZx67umjV//zj4H
/0eyYcXmlK1EBYWM8WjhQP5EcGZEjRSkWwybc2XcBJ1poPooC+a6vnbtHKpjo7KK+WX+V5wni+ei
zlLwxp929E4E5EscugYvyv7XILR5fcx87UR76tZpDwExLhQURL6oSyxAM7qAayDCDke2yd/hGHRX
EEwAicDQ4eJ+HpHpSRnwWCXkvurT3oRJQlHBp+gFsq0xIgU4SbOtbLIeVmmTnpEZGIcBOjw8V1dz
28nn1vWYPXnCPK1uRupHDqkwQ74xhRx8h39xsJC+ky/6swl0CTxl6lhIgnnyzxzEwVhNiI/NREoU
2e0M8uuqChnD0wx44z6mWWddBvEeJsF/XDGp5RJV2tWTbTaZgcH+5AaaVD8LT0nnO7rm3yRKaEBe
jlShlDWR+MXl+4qe5T00wZDc3ZyeCQ6v+v/+542hD3dRC68FG9BLV5K2wiGbb4DURi/8yCdW4sQe
KPKIVFKliPRurRXQNg+3abzR0vyLYaD5x+cfYd6Y9t+IMWfERH2XDIxC8upNp8hIZJE96YilG3Pv
1CQvfywyxDVvTl6COo/GAatgooEkD1wG/tIvtd/Ps+1dt3SL/t/9XzNUVcxP/1OpDbSfzbe9tWEo
atme4QOcHHq/y+LfPbQniB9mm+biuzSZUVmC7HOMRt+p8+/XsqiuOG/4RgieRtdUvAjtCIOBwP2w
YwoAVfTr1QjMNTChGdihrk/xYy4215DIQagnwXn0FWTwosBe69L3KzkpXpoNZKcYmnueZ7tNJwj6
eAJgzs0FqPXJGvTuqHt/6z3FBEU/DLv/o29ggGFFh23NEwvGd2N+bUNjag8FPfqabGRIA+M/rx87
ySyb27hNh7jm6jsj1VcMGEOysg5L/lDrF2UZTwYpW4g0xk2iIH0mPyg8exaYW02XX6k4XsRZqVks
B1IidLaOoJWBp7bytTLd3yszs17N9cZVQ1lnEeBo+1MdY8mWMcKS9jOAK9PwWxZhAlbAR8lw9oTd
FarfzhAUVUwx0fSkgG4AgLt/GF/Evh7pIShI+JQUxYp6ddLPkXPnPPrULNScvZJm0JUBbOfU7eSv
BW2iVDIG2Bt6zd0EVTXjC6BqnWOLtOg1AEQWInIubIseAxXRpCF1xRrGN+Rc4QenvjuTKEXc8We+
5/fWSiCTtP95f/r5FyUKNCE9IOdd4MhaEQe2zx6VIr8H8Z12Z60DQOZMAX3rglC97fQwT1OIhd5W
AU3+sq8B5P6o6Lj7rbMkxnyDHSzF8wNgBVmgPwdhXauxd9TMHZTyQOJhOWnPBFx70UI+xspQ3fCv
QDJqIHQARks3O4eC2EVXO/Wm8nnzspfjKP6q1i8pcwzMTJl+NXaLpf9+gfNMuIGf695wN8oZcQXT
bcDlAPUusYcJHjBPfyNOtMAJxzWjCf10JFOqwcDVg434BFc7O2PeBvcM4X929UblRoCZ2JGfPH5Z
aaLyFtrNUrvpsTgZ/GHXbkyhWHGgJVbmJO9IkGwL66TkgIboWGgrQNJsMHTxmsTMpsjMI9QvzsMg
tgnR7ksOwj7wXUk/IdTXW/knwTTuX2IOgVSsYFBwYgCKY9zBKiHG+7m6oYk2ebtwRNyt9eaJtM9i
KJJOam2JW2h1B/Tom/8Lx8mPssurkFapAOzA9WHDVsKLVaJK+26UMqVRHUScnC9OvjVoH1Ec2nDj
QS6mliPmdXMnWYesQ4Me+2QQ7UL37PF+jYFfETVcJBw+EBhpSzjgOEi7R947K4DQjGyloFn6C48E
0BUTZp7QetNsqlAgvijF0NIOGF+EjKpHVGq9TsjjR7fIn5M8bV+zDJUG+dKul7V1Ij7AHFEWcOYv
VdaVukPZAKFriAU7ANQNtgddLogz1rp5QB/IWV8avflp43JJkQywJAB8A8mB960HrXk2gJ5Vppt9
YJlBHag38CKpYuVv1k0ODtUBpB77tR6Qt0dLqnBvFnI7yx6P45bUy13/8zLVeBZLR8IA1PRQ25+K
lKbYsbwAGHemZegz/36hTYI0Dp1EVkb2TWfX/o6YF9xlblMZwIjnVlhnL1rP7BJatUTdjZ0/C823
3puDmNtUY1A8ck+oSIUhDyGeP8/gQiTKr08u0ppZAZYBpkqgCs8Oq8yNjXGhZvKDIfGQ9yWSaTdi
k+6fgLF80qB0uLalkzCRi5LnIeZw7KrdyCG+/p/wYcQgn0CCCHcsTrjQ1RwH1xEYtt5F7RgfsqLt
BKf1GxluYuhE2wxo83t/MochDJ8EU0g91hfESswfGq48KLnCByLwSU6JuJObLuJTNFijgDocM3CR
zS2pAoKX/tixpqF9bjs4IfLTXH2apjUTSRleiiVsUp5q8yrtPujE37uiB5oxiWqPL4UmclIMCotD
BWXxxWsE8ZMPitSB2BNlQnTUVlQsqg9jrfkrDzD6ZVsYyVm/pLHmaZRYkspPZEfAgUFPGO93OHAS
ngQspY9fhiSFIt9CgXFWBtdB2+nbfGvHjFTCALVzFfJ16KL7DvfZve9P84ZhFsIqCLDqGNoQd2QH
CFHn/ehj7vGCKSmH8sw6Jr2zlYPtqpK8LH5Y6iH4MQefiragUCBmF3rnJ0afhURHmtv4+ddSMR32
aLjEljY4Kser/daaGw+jTimhSaXOBrUQM7phemrko5MPm7ZcNhXOLeQjG5FQFiyclJsqC5L/jili
T8UH/yPLMMybf6TH6Hk32vim1DXb+UvjyRUQJQc58aC2NrRhKqkk6F12IPWL6FTRkQvCJB1q6FfH
Tp2s/l/lelv7Gw45L6tecVOuC4bafD4/2EbV3JeKGUxclR7QneCXfcIi0sjSbY/VCv9dIHLL8vdH
dgypxpviFbRCDieLzCTT05uqZ4R99S3kNJGPmsiVXqRyo0Cb7t+mD6UCMvAJ6C1fzhOmr4j3DiIK
XeHzpy97mrrwf5RgpbePa6Kte1P48q0BuCODk1/74pHlWYzQRFtN2daFn4n2v6H/95bWXlrvNIRv
ilqS3AQPWPmg02ey6WfJSsNaeVG69TVh2ioPpcul7VnOFp+qbRy7IFLByvdVa0oNivT/kYXZnjUk
e7DkDqkFSNsG8IfzMo6H4mRB6eVlOFnnpi3P4oGNTNprQX3YBrcU6+1IjYwmIZ4dI+ei+qr66P7E
6w4/ehbebkDdB3p4t/2gZVGY/TaXv/ohm2xgdci9YXDlQofJWS2L83Oo0aR+zey7Lelgf12jZUrZ
9dbYUwxPEPJ0t+LurIwogx+JAVDJfRB98s262fjRHYXyzYdyFhA6HuVD/gt9Q4x8/oZN7pIFCMfU
JuGm8a6vFsiYVOwd4UKeHw6arO1aCwVHsjyxSQo2shvnMpl43+iUQghxJwi4o51mck459hi2wXWK
jFtfVNdFMnkX2lQMTnQwlHbQZUHSzX6iGSd+DjL4pP62zbAFFKPGd38NXLaS1Q6PhUCH89gVAUAU
0R5BxZ3d5Gaqb9lf3XuyXuSRwYsOuFyZnrFDLoe0dMJR4Wwj2EWPmzdAM7LrFGkL1hS8D4Adg6Cr
i6wgEMdpR0v+kj3E7w+2lwoVgiG84fu8ZxhRXF4itNY1GRJ57m1U1iMv71nEdyn+WhDGEO0Thvlh
yvCDhwCYd7oIErszHc7D8VE6ly2eTnQ+n+rDsg0B3kEwYM4r7iW2/jjZ3kp30HDUpNysqDuY1xDd
F2+kcuojhU8b2saadDfmKrMfbvcaOVOnUU3zIkoGKxIrdrFc3rFG4iK1X+S44ZzpNqRrrDTrZtxs
cQr9r0rK5T8vhrHKjWDNGaocidh/9gwhUUEaLwkv6pdyWd/1onLMg4qP/J24RJ9bLQ8bM7PRX2SJ
NSytUADt4U+vRnJiBea8al5nSbo/g3q6cmU3+NZrCPGK6O8H92uFMKsgQcVPFtnJHZH9OwtR23W4
R0T9BcszH7G6QzLX1mpd/cDz5B5+ZGD6f7hINkySy/LgdgXXqnP4XSEE/sh72VUZHTdCLauvQLJK
kjGX+qa79ihDiXhm6foWrde7Yq/mkminU4bTZwzNy2ajYkFvxGsjc/R53IxLrExpfcl/czFeFXhb
rS9JFAW8oQnRcicqByydFA8fXoXvjJdHVifxUkLSjcIwufnfh9w3lUszxseBtDm+KQ1aNQ2dZRbB
zqK0SECQmZHrDTdebYP4lcZwEjRRJcR5DGp92kTgDwKhmAbgV+I+qoIC/ApB+Hox8uKHLwVDpXOq
MEImsEdCRBwQV1V9x0eNSYsp1g8NpsqCQ0lg/Jw85QDelO2C7XbuZqOtChl0JoIfQBkBXG5oroHF
HAh8Hwre/4T7xUfGcraANF6Qik91VTbV2QAgINOt29zoXJCvnYu/UvrPbUAiJX2cEae4B7GKF0Pv
B/p0b8f/JR11s4fYP26wI6xloPu+8YLus73jC5A3wkOkP5k3woLu7i4f0AqN7tE2drgFuZIvGBHN
cHD+YNxUiG3IaQMqU6OOQsVrSNG+GKj7Mlk1l70WZxFVUwz+F7c9/P3poWUXoKe4PlWcJgU0+Wsj
8iuDPapUkNvEu3YYJXynxFPTnLmnu9M4YWTT16hVD2uTaNVbGdd+/MBF9whEUr3KtpZuaZizX3Bd
wQpRms/V+WdiV9VIem/zFgggDh1rz4CaFSq1Wn7isYgr77Sy+Z7mIhAdJ1EXhnMfpbOnh+VJeIxM
a9Tgk+DG1nE8hZubZHs62IUOZhsf29vEgZqDuFswiKWeQ8tU3eQrVAO1dvKA8x+q6lg9xyDxD9qq
QEq6c00LEQhAZ6JwwRwPClaGmNxSluZ+jU0esCjdKo37uick4yvuJ8X4QbiSv4ycY7JKuud53Avr
Q8v5wNhflAovnkfw4iuT2aMAoZ/u2EWkKG5C1opI5O5EKioDWfBmJM0UqTqWkhsYjC5wgXFj6A1t
pPzMYEPYsFXOUJFz9Ei30gd+sUv0C/GGqwoaKtZTUSO03QaCkEbwUNl+yex20mI5bDI1ifZ0KoaL
EamG5iK3T1Qv6Wg3hWFawvB2bSjM1zC4H5Gdz2xcMUKBHJHDz+UPXuAr28kEm4+e24i/wX1Y+Kyy
8xY89VvFP5vuH/skvo1AXumAnD7nPDoIZ7RgGqsK+DGDoyQThN0uRcAZLSkd7iiaqMMM/IAsK1RJ
QpJ1ScV3II29uUupjIO7uuzPqRSRCDIi8MKsrT/7E3o9q6cmxURuQdbdBSYcsxM0cQ4rrc324V22
1pwT2CCVysOiMwv7AuxdAVhSuaCjLjzHG9zgS3SQzSIPB8YOYIDv5gzaPGya0mzq0za3CkwinRNe
+i/gM0W4VuFWHRDN+Z5vNhpN9qPmhxIBciShv82kmiSx7dI7E6R7uHrxBFslgFwN5fE5PZJ5CoNV
E7+j0lrdYsvR+QlGoU85qoTSGLX/lXGoWnqxYq8ItsVUo9gUnZkhwXpV0DOmh+stxfSgasXgA8u/
PqubqCZNYrmD3I0peza/RZIopU7ki007HJGURKtEHIHE4GxVfZNxKF5y/kcAhx+8tsDd5xHWCkqh
wSFPjFwJd0M2+aUefKZ3lSRy9EB54p1K2RLAFfSYKbsrX/A77DI3sx6sIlTTinlHEPIgUR50UeDP
s8Q7wPj6zsQ6XC8fUpDbhvo0xFzWl3S5z0aULR2cTyMiGJle0/23tj5p1xXMc64cSS4DoPLmDjBA
IYpar0mkMypJj8+eErKvEGKT/m/43NR3tMhxE82H9GsHkQ8dL28x6WLCySRqrur0OhFm+4btcmqF
I0/qYCVLs/ySBW6h4Dn7WR+dHZPmFXsQTpphdNlETPPll1tq/unTksolaGP5mK5Uih/zEU4DgXQY
/umriJ3MySISCJJrEJnfZ6I1lEPtgfLapEWJB2qLE9r21jCy2pxlgeM3mrtNlz6YIqeQzurGXwKf
rZQ3CQOgZSn9AuxPxxJnhir44yucR4kK5AxAtFXTQzpDCghx30Z0Vq9J1V/RFW4hxux4NtJ3BLi2
98Ph6+E+53Wzi+WXjr7M/zHSzKzvCwVakumXBFhWYSa7caw1YorXf7pZkjYzN/TPU2PwOFGuZOrh
0W8XEIOJQQ2eZd/7D2i++6xFuNJIWXdk7un7fBapgJh5hDgtwNqE5FiRj9DbOo8W/0kqUYDY9Kf2
EWcT8Re/C6Yh15d34K/buTgKvGCQW6ajXxEY8MyfTwQpot4P87Kwv1bjr5s/nNapTHTFyR7maosw
O3JGbxt/0caAIOjHYkbWIXg1zVlhJcCGgfgutBF3m0nHZvn7yH0TREsxpxoml0XKM568xTmhGKj/
TKaR8eszxwLE/FzSwe0kftKYJe3k0XP17stNmJ3SLoTAqEhfGgZQk0hmepoPXIPPR4zDH2h85GGb
cS/+fr/ylIVa3EteEv0seDRC2tiwK52TevbD8WiCC4MlxHltj5dnY3iZIo/xFvcbzcVlQhpYWHWw
eseuAmxT4xSwIFP/FsWUphYGFeDGvupsdsRnhwA9TNkjnpWAY3WpwQ1qkROYjngs6IuaBj5W+2cp
2TGE9jKXKum0PMCo+bqqJcE+sh71DsKhQErytNNqTllXmRrCRl3xT1DtWVkzBfKnXDZt1iNSwSm9
1RUIQzlcBN9JgAIootDqir571SBrgtZelUpaNfmlFqBcKioRQQqixe+nLUCXTZXL235bxlc5yar/
zW+4IECFwfDVydOmLXnSXzSgycWr3Y/3f/o1slvnlCKaGRdrfVxPlpYG0dqUnBs5uST7szMgHNyC
QHuTXgjdmcVef89xG2TtcnzW1fkMOC1sXZXiOKQVIW33DzwxGUnMONSGZep+4K+t8N7I7JXmwBe+
AWb4nUvIcY1y8WapXxSKjitGoa5pvSH7NWvKOteuRDz7a1v4aPS3Yn+KH8RRLZ1tQRpbPmr0Wr5I
9LmRLmJm8g1AbOnDeuLsyUXm9XuW3cI5VglvTb/1LlZZa3PQjkvg4F+AvsweyXVjEx7FCmTQ0AOf
cIWpXzPk77+X6x6R/8rgjkq9bXQ2mFERmk9cabm7i8CunuiIu/NMpjq2vfEkUdIFK04z3qChh8iv
TKnmNtlQGnX7VwZWZbmA8m+cg4h42BjASM68QLNR/SEdoURuxxr/Uvk03yuCeOf/QGITA1mhfGoD
Hoi85FtxWrqGOMxsxLL1chd15jDeHVjxEDmDSRE9EBubY25pso4R7mFCyV0jVf1aas/cm7pr5YLe
21K4dqeLXKffRUWD6kEoAak3dMy//Z/0ptSpzjBj6t4XIEpvXh+k/u9R+i56QddSn9qR+cKRyr18
NKyNqg63xJzZ4XPGG8ttpKUV6RY3Hi1g0QnF60qruk2BZ0r7WPZ7L6inwJggu12raWM59ZDed2Mn
C5Zju+dotkhcNKSmdgQX+ZVH0Kwwo9GmaAKRJuh3HFYN50npx5vieA10c8o0tDHVFcDRFyFSJw2w
SODKux/Q6BAXacllvrQk9EL7JBtYn5PCfaGkZK8iDwTstBR0seqAv6Iw3xlOjE+LZQwzgjVkrVaP
zCGtV/4YhsTjAoUm/yGT8z84qr7FoJwPdpqSvGz3S+/XnjkdnfDn29BJJlVrpkPJe7tlzwB2UJum
QYMuI9vKWgAIoXXEH9gbEoI9F9S0bfhmqgvpMCAHAVtwA6RM1UNiEPKe316FSOQBmJcoljteCIVS
Z1CcesH8nyZDMx6qZ9ZDKyskUhJn+cyNV6v9/tTLMVezTUuRdGmsDxjbQT7t1KNLUKUYVWJ29WM7
MkDxIDubLJu5jKDJrCOrxY6s2Ws/fMA6lqjcaWyfTo533v90SAboW9FFWvKd9kGuAqx3RRWJD9ze
OHIWQizKlSNyq317V/j6E/8MHVcWlvH7jQ4ZFcZVAab4BUAV/vfTn49pNDO1sN2w9gC61vVDMdIC
PMKLyzmrV5sAHskvS29+uSTPwxPZxi4zUJC5aPv8mvbE3H+MyNbxUFPuUgsqCcH1R96DNiz5RjZD
e+XYsKLy/6pFraNc/D0h91+LkZ+ALuPlR3uaYgruafv/6ZEraerdTxDxsP1FW+vEC2hMZbe6HYZG
G1/DVyjWdfXGrbMXqKChT/fbxFs1jfxxNZtpiX0veeeahwlJ8y7gDpEwmJsBdcrxaIvxjb7WR0AQ
2eE42s4qMvlyJRepCzAgtIrPt05aZKMumVBWTHHLhyH8qKr1uOwHRnuGBvo6uHT1JdYNTbLodKu0
CPen14RAOHNsBWbO70FpUh39e45HWDIw1GoywClXFQ9WpqbrfD2up0Fd4XcpH9qTlXN7tfkCZw9m
j2PBNSLfir/C5Z8SqSuxmMpbQahzk7ujTN5Az3AWnzMMjKZXglQcAlh6P2nfiy8m4pncbCYvEF5P
tV0+NXbyNNS5MecifCF5Rc2BS/RxknxBeN/3BEXD2qzWvvdlE1EoQUv/qyxIu6QQg4clZqaUwDz4
OCqrzSQBUHG1wLa1tIO4KsZ8XKOPSUPhaKZL9nOAX0xP3mhRm0dCn8um9tZMaXx1sSwJ6e/ETgEM
jYZonp/+Cc1aJuqyKVedMc3FFA//SDe8OunqJisuWLEjIsB51c3Z0OR1fWcLz0kRGY4J9liRTK2K
Sx6ial4qNbhVPQZoSE0kExYHMWvcJirLEiqAJZfAaMI9LbjD69/i5WLPVEJRsEyQRsdUqA2AoVp9
UnHA79hvj7BtSEgTlUByCAvUMtZC4gBFChz3GElKq7KrDagi53G9f0rSuBC9WweQKcBswYB0mOK4
4dtHj1LjBG5a5KfEJnpb9nt+noDFy46kwYXe+iNY3f5PlmoY4QDiEZiYKbR4pgl5iXPe9wZnk8rj
Q9/2QOegeROhOiriuQCLWdyRUQ4vpOYIDH80POzqnytHj52OEaQ35Urnj94jiVRgCvT26Z+Ym9PO
YKEOQ1z0IwvjKre/J3MQ1Tzk2kjeZVKRhmVs+HS9N0i8JD+YW0EfKHzUYPcsnXXWV78Z3ojViy6m
SVtW++pBL9XvIozfhaDSwEI090oOGqU46NskBjV5FH8VzB+3tKvNGzp3cJfDjYdsCHwF30NxNG7d
RFx3FWOAliTOvB9SUddYZErfw5FWUWI8l468Yrgj0g1x0Qmc1xXbIEktorNlCaRCiX7tULpy/S5G
rhubVOJ/nwcGNNDs310j3dPlp3/GYh6jPwQIYmSMfdQjNgbCdfL1UdJ98ppYDGabeMRHMbTFLxXI
EbpgvTRhs6ILKnRZqk+IdBbFJLrA8bNTaAjqq1C8aIFuIvFwepZtic4nZD9ipavdCd3jzxHsyBE7
07WhiG7U39/LaLYTVR9onTQjb9hWF80zdrCEwB/MwCsmDwMDhM77JkY+zILM7g/C2ka+avpSVyCJ
2u2gBH/4l/TVDqyEzI/hC5+HBACG6ZCjOpTxlsQfSKHvM2ZwjjemxrtcCa/Xg5SVb5+LcxFDUsyw
aiPsowEOw3dBrsDvmgDxq2JowlaCBBhpbLh3pw3gJjRQQ0QCKFZjFdl6KLl18vBPsDqygFwYOOgN
jIfeAqLGsv0OfkNxbhafjPNhetCDDNkLwHM2uv6SGfYFHCh/DCNW3r1ZW0I6YI0lSP3NdQZewTpA
YyeXYMaRwhEZdF7zvr/jwXhWbS0fpLnyhaL3wTVcDmdG47XRz5Iv/MIPR0zhHtAr+9vcX5dOyVk1
qfYoyQQ8oq8e9lqQlWpV9DEH7X8yYEkqcqymM4S4TUvDea51LUrJaLMEwurqbdAjm5j2imFMkO1q
nDoo5fbBwLwlrr5P7rxw2p3xAVPKWPvhcGB5MgbJmt4nY7XD9/eTWt/xjH1jozKpgsA9Tb586yuO
e7BxKmxrkFfigL8uwJy4Qn0tCkysHUV9R4PFHegy0WWAQA0NYsyj1stXtdRlSMwZjEaEGPuWbaIY
EMw7xqQJun9c2PZoB/x6IBRhlDshdppJbiTr9ICvD5XbS0XGpbtcJKXTp5wXIZ1tpYX9QQ8S5ceS
jQn3hieioBzqihhoo+p2g36/Up4ZF0HrVg+gRW67U3sUmocSWbhy8tAovBlysDuMBDDipJN5tXw7
3dNbxQ25xsxU2pUFLL71SOxi2PKRS8AfhB0Qei7bolan9Q0TTZniy3dqlcPVWjSC7TVfffo7EuDJ
aDPA0ThjCX3hu/1wAAx4Lq0l4LLWwHALgEv/MMwx48UsxGUKge6VnrysMJPmwhXZ+qccxDmvVG6F
84beYIIWWpRgh0rEzg0vxsKXxom/bUrGGdqb9GMUyhM+ovVgtLWeWA4cn1X+fr27rfUX4s0WZTYH
5qm4CHFV2uub52py6jHXDlIUCO/0KSRB6Si3t0P9LyW67SF96wiQ9DoaV/wfhEZ3V2NqNTyDYFkR
1cGcMLGUTAlLlKbg3e8YRjNNl5/73lZkA5q+IRG7mcVLO11KiF/zCwr3RyhD7yzHOxBIfBwoypZD
bYEWADC2VbuvuXXy4FoV1sSRgxbt49xFW2wtakqZ0j3MtSvZ+BQI7YKc0aHbCVZr5Fgr4ZwxqkNz
ihnZKh/mnJY1AWYCKz6eOA+OTomZdudBBJUrf4S9rOKUIPoX0mjchvOMzpCIuAhGr+BYJGrssGvr
GZhIeI7uFltibyz30zeMqjxV0I1ABGgJmDhSjCd9zOxUzeMT8L8KAXQbgXXZ9+5D7RMXFXDr1lsT
fFV/AQZBUHxSr6fgCz1uVmFAzQg4jID4XIZPPMTvvH/dVi6kM42R5A9fojGzjJOE5uU1PsTXmR3N
FRqHF7TJt6h7IHUx/HxfbTwc+XZ2kbJq6nGFhZTqER88s07z6m8fYtMCI8Q9B/7sFIweK9n199G9
dA/qu2IcivnIy4KjeFSyF/4E89ldFhDg08NIOCSJsvgUriQap0tOT7YMvt85zAQrAHhFgZHm7oja
6kafzCqEqood7ft0dGjQ9E85tk6hIEC/J1B1asYI4Qlj9pb4RHgY3+pOJQPBzuT9CwpHwUMWQRPv
6M/OvF69w9Di/ESSTHJblVxMCne/sqCvt/zJMgI+5Rq8YtfMsRQ+1Chd4YvwRuD2+GTYQ4rNMhU0
lj7nYefx+Vxt6M2Bcb6BMSN1X43DLIR6Edclr7K63nV9QkEFerKeWpYUCK+XqMe/5lFAFZRY9Mgs
GmWJBwUedQIlUOu1C2ePEf9tHqZmNkmorvzTwzSVIiHKiDkB3YiQeflbHc/sAfLGsApo4HJfNf6j
9U7uzXaH0QlDLR9IstDpyO39wAK+saCnnLK4llq+ZsFjp3R29i+2AAmHretfWnz2188rTIfrjg6F
ehPUUG4Sfe2VjDuHYuod+hp8+Ld1ljnQWwuKn+Cai4Fx4lJyP1OINEyD8YgDUAhFa2iYXnFYKDRk
R6JpHDtP+hgpJxk3D//aI63qVf+xzBAOMxBCTa7B2IpOW8/lUL95mnDiTjFWhpX6sqx8KJ2cmxiy
x1XhT0hRfVAvlv+jt14W163RazzNDklLsTgNsJZ5lQcWj97ZulpaMVTY3BNT9nBVUrzONi3Xnfzz
RE5ofJtQa8JpqkCV7Ail7rwfO7Nu617VIYmH/WTqQe0K+K70LYDXVOjpVbKezWDEBpcFioM3SGcd
d6SyDyocipc9r4zkyfHEcK14rQlqpBUbSgChdAa61EgwP3FPS43/eNpXEyweeVrmStVavgxDEKRL
t/mjzm1XlnofRjSJbKBn4a+WTLBebGTH0O/LMC66niw6mkFvq54LZij876UG4G5Y44pB6czooiX9
clFqntN7KZrV6fvQi5UYNcLW69X45/G+SkqextvtUgJKhZpdkmZO4vX2i+bk0QW/LXfaujOKb6v5
+rF2ss99sZcTvHb/s8k51q2hPp2J/VCDwC+A8HpT2r+xe89uspkLzCeRxnRxKXR+S/9TqPdIKo72
+DgZXBtcCw35hgizZPXNuY7B9A6FZDohazSVTtFOgmd4oUIoksECk2KE7hSyrI22kNVJOW1Cx5uu
WwhyCXfHvS8RJy1r13UMPohBlGLvAEyo4h9alLMEQpwWuqEMnyN888GLnYo0LH843IqfMP0+n2DJ
5Ohvxi4sixNQCcHH+RdAGgI9vDU6aJ25gOmyvoT0SflpTHm8p7wZin7GrGBpTzDS8zwsYFviND0l
MpNnG+lJbYsqHk4yyEsdtiGQuKxCiJzqwwsr5ks1SgnjBViRycTw+B95F59UF+xGDgAV2I3CFoq4
v9Ty22z9tpS6H6ge+OR3oKV4it7KeNQZepa84ZhNtQw2PbE/DsMdRfqJQZ4sp5VF3g+RWswPBJmP
+u/VFiGwmMRS+E4QcVc2pDFf9vLppoxkS578qLRuN1WjW0Ft5MSLK2wHt/0pJLvsSZHh/FBuU4D/
DEMzCy+GFvBvGos1n7EKsqw6ZwP8390K2aKIlJOW1pBC0/5JZdp1EqNk6kBoBwVubfssuzDxbgqx
f5hVBfA17RQtwWYkjnlGwUVRRFls/Omgxv6txcvRtlxqXUUW8KISG/tMDNu0f6K+ftqF7XquyTGM
ne9cNKQgcT8dmgEKVgFDGfQJTTJ05z5WMObwQE7jEyd+kxsXJyLU0iM4aQgULkRAFhdXWNHR80+p
efxdiomvBw81jxMgqF7hZBoibt+LESmcSK7m2Bj/m2FUipwQcIiPCvg0G92zLJsfGAwYxfYOUhLK
4nyMl9TdjovhfXL2iqhaTx26/8iGWk7U6MNhl9050bF+xmwAI6KDDP/RFYDR6Lpl6yzgaqZFADey
T9LleI/HVU5uCh9F+H/dbZIY/OFkklPOuGOwB5o0frJeJ0NFjHvSxjeoOyqVYIKvhRhKGwaOv/cC
Q7IBCRXk9iK6tPdhoyVErsdO5eyYgNMU3NvSr2NuQHdoB0ALdAmRyn2CX9PziRHrsYBNZ6Icg4JG
GHOMhOD+sPtaCFaYMFW9MehIswv0vHMere8atyb/V+ulyd2d6z4h2SZnt1KRYOndUVAzgdr+2oE6
6ikrnJ/inL9kiG+XkMrMxim5Bnwk7UcUf7Qeqlng+731dLtRp4krceNRq1e1xlj0hO1Rr1dvwsf1
ZEvBN/qq+l5eBZH6QwTlKJ4ZjRyfV6uQFA8cMOeW52klUiBRbL1rDW3knp6qqQ9WZ34+SYmmu+yh
H0w98vveW5pLELD99pqzlHYaiaTHhnoGaMdZkRPZfNaT3C4luCPpxNRk2a4IP2hIkQI2HB0CCBk9
yrQCOcsA05vcHDxlBV159DHtYRbpQvTOd1l0cIuzH5szdYJjb3eE86nVrLDQbrrhjtk3LkZOsksP
etJ8if0N+MPGSU8TdrKzUY+kel57OQc29MzVxisRxS5uEWSRkk2U/idNtWfMpW+OO2zHVCRKtVcN
qMOMVMvZTpBZ9Uq30nMVE6/tqBAMyh5QI6iYQMggj0Lga4eR+5pwy5WuYEFpcbnXfO0f0CJiIBcw
yKNSO1AYtyZvvg6+YFmRuVqgpdUklT4eNbifS2akqO8644gjTfAFZm/28Y60porjs093ig/7wcd/
hKsRO4I4GJ8NdvcqYau4S9l3TrJaoiLyuFmbU7GiFmZlFr/MvOFGQf4oaNb/qpp47OPlSK5PIf8W
/PCIrO37bRK0n7dQvOG/qV7n+OTx/PyN6aSwAWF6El8ziftW6GVTam1nosTT4q569bwGzlabkGdB
/XS90aIZO3XTFS+w4uhCocA/BqjogZ9EoLpSs1x4Xa7pHWxFiPvYcH9xtPwRIjpUSTOc4QAUf3yP
e2L2KfpjjBibz5o1kPDz63VO2e2qtYbosxKhsYdizBriSNVAIoxkJzMZyplLKTJxxa5FC6kyQzaI
0vlKAK0o/fJ+BhzNDu51+5vQKOsWb3IwbbqIYtnzIzJlLXUg0CesEe5eXe4j+t7hMFJpBKPsPpUP
NZgwd1QWQJYvmebl19YvVlu0+/oGitQwk2/tWBuHZsEigYEFKXC+mcf+RF2V8GHA8VIKR5KajEUc
OqPM2UD+u9LrdaP2HiKH2gP8v7soTOO/im+vwZXvy5U8hLu9RIa7R1EkQdLK7OouR75dAV7BYSBw
OUK0oJJw+c29k3E7s+/UnTJcmwhWyWqIjGLgGtNsvVkaIcnS2tyw/3jkRBi7mxGOuGF9gY4Desi0
SuwU7ZC7hWZne3dmygUwuhoeQs1LnvgVAhY+mfBnwf9ledlk4OS22nknSJuWEQNvYkRMFvLHPIxD
p5f5U/PLvcu4wU4c/0jhILa7ZjeWImCNoBYBiLHOEAbrsZrfLTbAfFXl37Xn4zblVxIuH1vnMIdd
ZQqUFHMOlZwRMZIN1lWItjT8g06RnDU2cgWa9mJ9wFU+fmjBjjnVzGfwH/FJBgco16SgZEILJUxt
1+TcVQVBSY+tWoZrmdAxA+xLWQeiAoZHwJzzss/KkoMO0AwQ3Ml969oyyJ13PtJvjEIAHnJnd+Ir
3xUXnUArmfWX8AFCsmmOlvM9bbnc8antG1TwTQK7OFFxcCXrVG2EiXN6GghngmrO+YR6xUAltm7w
4DuccaH3Yng9HkDVIhinn2L5mxNot0th9U5HzH1EgSRhOjZwLo1ZOR6sOwcv4pwU4r9FihpWHRZ6
8d7n4eDIzB0p3Dm2Mkuu6vrI2iGgUcO3J1pHobslgbS9faQ7VNhPlZ7QyYIQLLl8w58EtkHx0imN
lSEd4iJSUPbTAy6jHZtfeIR5UndPE20i6yGruTu5sBYdP5YLEZUve1oXporOR1DPimbsJwynpqab
+ZzpzeD8gbhM+NsFEuOWC931fCHkgtnKnft8/c6IEIxj536CThJ4s19M09n/EJ/Zg68zZSkP5qSi
vskywUQ69wFTOYsBcFXrzuRfKPBlmEHJ1ZafSsTCQ7QByERkO9HX+vg/KmSeQuVU100EmObRBsN7
CICCkJr0OLfhPVdNXWHtx6V/oEVfyfVozg5ESQgZDWObxJEQ5kxgV++Z0dHJjU4xR5FqFXPO9jav
UVyWvls9ZJ8+bTPgtI8iDfVf/TmKp/vprzgcaZ6n89xiUNl6NhBZiFEFxu+8nQVEjTGuzn6Vvs1Y
ekN2cls7tf6zTKKPqNy+pEEPixxsZshxSTh3GCzodkNuDEJlb/tY/Kxt+MT3+nvuyTIhuL8IM/x9
fUcD7G6lw5UfDWeCWAvSBh1mharWovdMIC/Sb5/ACWJ3Io+jH/MS05IgPCXhkxg0XMOR2+xmG9w0
75khMEGahskE4P/4tKXIVub6i1eBUpVvKkhsKg8P1eVbHiVxcGOeKv9H3Gx7QE/BR6rSOrQXalpn
aOo7kwTmTnHobEt9FoDRfrIJszGOBq8MMaVmxMiFfHh4az1uDvQC27hhyx6p6TMiNwqMd+nkfSoS
+KgyPANLLbgzRnmPeE2BIBCTZvWC1GWFL+UdhEW07F+RDsU+8oyQS1lYHWYWseslKWEeFzVXRac/
KbslMWlwcm3z0pY/1VxGUAlSz9sXLUKVk8++WI4d7Ne3pif5xsTqOy6YkY7ZzENC3aiRisAt4vxA
nr4WTpL4ZbVdHrrg9Z8nrb54AE85eIyJlf7KXl5Td7zS4oVzySmxwQgUBfgDlvjPeUcPa7mVaksh
GLmEdwumBeOSfRffm/ElAjbW6x7MEJvzqsMdJGSZuJ0GfnBM8oBN7YZBbKFZJD6ndInM9CEZsvRU
6cuXoLX0FNyoETlnvDk56PR/K468JLSZc7uyaLSrH4U7/fj/xFp0nOxHqYTdP7cGUnWWDzOcifiY
PYr1+3uzaAnFm2Gb3BHIpoI7Ko4WH7I/NFyIDWmF/4rzXPGTF50j/IEfoCFlKBBwqDR4e1tSzJ4F
fWaooVLbctaV8vQKsqwSVDLOdwFemyr68Vu12VmMJPTWfQRnEWaJ575Rte3wRM2uKlkW/y2HS5uF
pwM7Swd0MWB6OFXZb6IF5TyWtn9eWAsLsFp+n/TScWlgpm4857LrSY1G0uRKSc0ZgTeOUGeji7De
v/c3xQLB6kwzS6fTkxxKdRXMWNNfY4W00yU0E+NfSP9EeO0b0DaEvnLcXWQLPNFFgjeSjsT1ZaCk
yp5bzQ3F94YY32R2a5bLBB0K0+68h1GloPuCn+1esTnTJ8FOF57DF6wn7SGUU+nBnUvc+Cr78bWl
VGR+rEpuvcDZAiDFu/rxwxqpJ+9Tb0BosM3wW6mZKW3oDqGdxWDwx4Tf+zlIIEnFSMFUV0a0QcoC
3Cw37yM0AGhkwfIbsF8K6DQH3oxHoYK5Roeb9KFFVbyXYwsBvCv8j8wgKCwOfz6WWpatm5/0s9Bf
ld+3q1TH6yt5eDlSFsLCX1FfA/tbzKv39/ifBBW96GQL3ej5a5L67aF6BOVwN+aEV5T1xA8kfGhk
5D8BiM6U5OLICS8rn5Khi4vh2Snu9ox0YPth1t7n5pA3PxBcsUa9gfSKVhiLzizPrS8Ok6JzNava
bjnx3dhv1nYe5OoL1Ml7tTklnS1L0tX0qMHW/pydKb3+rfdsVWn84zfFIfkkinY7Y5+ra91XXN2s
A4yVru3JR/D4O3oAKUD1FgUVS24b+UBx+Bf/smlfhdnWBu9uPWc8FyhVOWriTnhd+qaQ3J9epObk
vVvnvztBUIKp7CBfQJ7LXtZai2VlY7epIA0II9sZwoqgR15nAEoWG47w1MOYOtBRhWWcXhtSK6p7
tZKfLFCVLcE/XJG8rE97j1HIZTQY09MnvdKxuYR1JCIsqlx7SXGA1IfNZWmffflMeGhg3U0e1CVZ
to4VrMUP7YUxOXmwcKA1MtevpU9sFIp56fArA7KmIbfbi4KXfjMQyRRCLBBBt3BKvNpsp8dQESPl
hRlzJr36PQM8dT/i9xstEtQPCU9YHPtxeUzTF3jz+Hxm42OGPagX6okrtvFvJLnQm693hDaGcuGH
wqQzZh0oHojd0yunqLPs8a5yp0vbeq6Oql2pfnLzJq9DIB5pytMGIf7pLaei8jOgLeXRtly2ejWy
vtwq/SXUokN8k4guNj/5ijzzaPaXbnDT5LqYT5Tg/ygdFsAViOpQD0SI3U14YWI34Lah8ZmG6ayR
BG3DPmVGPOYXHcbCER1zpnVxM1C4xK07IEHt17ZvQGMqzEFpYCNDWAmCkmIb9Jo0cktF0Fmw7Wdu
RSm8e26phedA4BGFAA2yWGB3fmlWyBcbn73sKnm1Mk/09E8wrVssUbcDeh/aM9twFuHYele7OFov
xg/iTkAEIUeyAXfMSp8b+0j1b7Lv3htMiLACOEM63RhV+3VFdY4T0IIQ+MXWL78p10Ml1kLUyJHG
yjgk2FvLIcEe1/eCIEiehcWfhx1Sevz0zr7HtdBrvJnscURJSElwgcJ+xLPbvkTIyrl0fcHgr19M
EfaD2tUisXRSg0CMXnAlx3w8uloTPvBrzyKIAk/5fc9ruhQGn3Wmzn2y0hd69/AjmNbuxLDi42OO
niaVwq2WQio4f4KVNpXroPYpQAWMIT71KzYp4XwtPXcfUnz+ErOwbw4EoPYv3ej6SGbWkV3n+mdX
vH6N8IdXoFXJ7OK0M3+KznnLfncE5vJAsg9N/hrZLqYHeIz4fGnxmP+vjrCCTZZ1yUa8NgB5+tZ1
gbS1Bb13ysFvbt/u1zG8Y32x9woztOegoLZ2U7Y9TxQRHHdrypASnp4EZLdqhiN0ZoCkPmg8y+xp
pxFsFHVCPnoVpDZr8BBbtvLq5vMPFfu3Bl/ASC/+aensqxKUSfgoWNjKyDClYhTOdxETm6MRav4t
a6U9PQ3n+No/GM3rFINLkBgO+7MSTSlpQYfDkm7uVVBjKy0hVIw99uS1/3DChM2f4Cphfuw3VOIm
ca5i4B87w9P4aEBrrf7mLsyeC4yb5hG14nWotF8cbE1n4ip449Nv9vxSSYGNCtvWNg9qHIVqUqFk
tL4q/DUMRwHCWOFT7ckfLkWvV8YgqY5F4VMhFJC+k2kRQbqy/TN4kxzf9BhEd9DtSnAD3nDdWLhf
4fkLjFIvWqXUaz6OfvCEGqBOanpN4s58O7ToLqL2clkXkWqQtm70qDMWmq7i2vfgqXtXNIByOM9K
wIMwlxeKQM0a9zOHHCtr8y0/r1EtcHHKZZ3NlBtjpAe1kYj9zCL90v5bICEBB0p9G2Yz196g+wQr
K/V/KIEKYWiFeuAzbUtrQ0xJXkz9/8dmm9cQ6PbW08Xk4jCLzvpwxtiCkE3hujlcOTCWm1zb15Qy
g3zq2nItGOTeM4wYi0HtATbV6SNYeiGoafLvEDS7t0VHq1kfwXFYk+fqT1JkxbM92+ldmpOjw6Li
vXn8Ix75QJis6EBEgKHPkUM/jJSBYx/g4adP3Hx27j0fenTC4EeLjmAuO+u3pbJcGMEoQYpPg34E
comYNjEQr+p/2Q20q8vXlRmOLQjJ/XxCaZXVtMxgWttkyXg6k8o5NKBk4L94BGw7/9dRY9kDzeLp
b5wLVh6OPiwF0vLzUFMfci0MzDstK4+00jxwH3OWwigaTQ8NfyQXp8ZQCbdeflyz6R8hMIU0ZOND
QnjInxJt/v7k7RkC2teBSWEyJZvlz0v+dS625NbpdCQTQz9flCmEPBUizJx68iNjvtrme9Pm0cUM
WBvRaNf72JkijgnqpYOMp/NadZLFBsMaSWJ6xaRq3rlbJyIFBVQsw0U8RC8pea43m+XpZfUzZ8Tp
YBUMib5UOC87DjbSQXqEUz0/l7xhdlEp9OQCNSHjGv5TvDqDp5zf4X+5T4lOiKQIHePHXoQJyOgj
/dopRoMDzNe1FKPFaMGlgZlPwQnePzARHE7vr0QEMTZ0/0KXrYT78kbMELO4IDJLMVb14dU5hyXH
auDjFEZLQ7vCCjZIpzyMEDDL+7GDb5VMqBeECNEItz1OHG+/S6K7XtLnMYVBqnarfK1pBqPNkuVd
UO6lgdMe3nYuumuoYQ8nFzrRefDYlTN9DRKNLug5t5tNzScIVwdbBzwS2mTD2dHfUZy+GJ6Wx2mz
H7IB0RuCtgDeD4RwLbwZwHDoq/WJ70llbV3SL4Gom5DGa3LelrGBaYX6GOb0DUzHwSU37hR9G36A
DcDBTUARZ1XxwrryQL+Bxi0TsA5uxbD8tIHo/Xqkv8XasBYM47THeiXFUXBuX7F5tFLtZW4wUpuC
BSmTLAtF7XsuZ2m9YPlQN0urPAxkZlLxNFEb7aC/x9jAnPIF0vEm44pqbmIFdpjUWOG2Osn1jhfk
CLAo3n6s2xvWah1FZmAT3U4ByVYzHHdMcAf7J9t6yNBTSo2+K3n5oGxieLmDZwlgFfVqgjiZ5vq2
tWSTHUaQyDzSPj978D7G1DxtGblruaf/PruMHP5WvhBRAKMTM/NSBnMcbwyIqbvc2sNjNFu/Xj7Y
PJMUwM7JmNIRxW/+kBwS75gnjqP/mfXO0EYlFG6EK/MWXRp/orAaMszyqyvP1rOkn7ihZWrhQuJP
BHNINFzRIbTvjpYR68Hv2Llj/epkw9YcxigP6i16TPPVshW+YCqZuAz2sPZC5JQkaat478EKzxOk
UCKtcNtO+Dm9fr6qIABjVRSlaU+9tHDFv4KLwndA7Cj7KfkDB4Hmj8XENgt6GtQpG2QJHAKHDWkH
tCyCraDJmaAfw02+IxIDuz9kRxC5vG+6wWugG8Y16lP/Qanhjp0WwY8fBVk4r+mLLsCFPhu81keP
lU5V/DOGuXKBey3p4TpBpMuZ3Pkv6niArVx/RA7ST6z8k9fKI9/rAeynzTdmSL3n2FCugKwDuPra
B+nKuQt1IIPoU9vfGCYWx54jU0H9ypVkV/s2wNP3W9JLVom29e7RlxEOln8EqoZpUYeHvjj11W5g
I8mJlHLloEq4Rv4+AhKSQxpaViMSgJjc4+4NjoHiy3KH/aTsSUHCHtvTHZU+vOEaT9bk3yoF4mze
5s3v/LAuLBK0ReZf2UULDA71OUFfcAh1L3rI+6Hwj2nNxs+8Io8ydFOt9r5zEKF7EsK6KCje7GLW
vOhUecWDiz1wrFSAGNS2AZaw4cUpW7+6WQMq+R5gfzHeeyI3KzgDUCmeFQeqgfZ3pcjL34LZf/Xu
yxoMjHQxkMAyXMVsQAURSlck550uPixDzTuQQoC4RNBdIuWiUPr3fsMiO0+hkD5Nskif9dHo/jJy
Q7txWqwiphg7lQBuvSnYJVYYWK2rMtSIdgfBmvKUzxIe6ETdoyyl3pZEWF19yHV5jorXGEUJprq7
6eGhBH4a1KxBFyuf4WZdIUgMfZTJd37MDLDm9Zk3y17Xd1RI7NGgjLmJ8kgi61F+SrJiXGEzx8r3
MzDx9A/i8ROF3pqdNQonSAmNje9nAzNFeYtkdMuw6u9gezIGBZHdrU6CBx0FJ8hBZBQrkSRz8kr6
KoaNbXcSf9fwgPg2CEy7+bFp6FhF3cZBH2/9auJy/sSuR1aP2NB6jstR7pVnuzaG7OnSeVFolP1A
HsZOzkQlo/BPvNIJpytTf6JZPfkkqPbZKLAVWJy8Rf9VZYZkSbyGVgGfd/EAMHkzoya/UQQyquvp
vjtri6uMR/qucT+32mMw9MYcTZ/EgnMGcrsWq3xEAEKWDVYsK3fOVL88OiwPLUpa8AHGVxv9Torf
6x6p77McJxn4p9o74Xsf5JCI9AD1Qzlxd8JpYkyaG2kXzt6IFv0U6kWAVuRiBJ42G1vWfBzT6+1Y
cA6b3HLWYFm9mzPScVt1EJkirwKn5nsZVJ5AiZtFcljZZ19Mn8w13bUyqrF2WxRxoz7qMLVyWLo/
xP21O/ID2tJ+GIgN9UIZfYFCP6h6yPGmVlKKZt7N3rFmLxLaW56qzhJV6CTbvLCvW3jby78+4YhC
QjW8o+D7DN3WhZfdjPNRYB+PMIJ4EBZXE86YqEgWRnEMxvYT/yIrLu9ztdzAmP9ZeXabyoJJ9oty
ITsE2XvjJ1kfz/CwPvGYIkKqpdbThnD7TWxQHNzAt2rqmg3LwqtN8YiFJvRlXmkhTY+dUtOlnSaO
q2k8XVUB0CkMd2SVerA8Z2dPh1wsgOzyYMZDgnYL84AtTdBMjIv8Yz6VBZASjTMquFs8i9d+SVTu
ZbAYzskklLmenEEsT9FT2EaHpiZgLAuo8731H8pfUDemXViHyacSFiz03ilpnBbsgkKA/Rg3M8ys
WQtId1XDBPBB7kn7afWGryvYAblsrutSvqYUnJAqTDDqrT3K62eZ2U4NTq004cQUdiwMu3W8jbT8
iuA3uqMDfNXzIHxaqbbNsZikb1f4r3ysKYOtJN5Ob6Fvm1XDKUmDXA9X7hyiZDUW52gjpSlsu2dK
SspNL6NWXDOUjqsk9G/3LgYYpi3U7+z3eMCZ1BikfZmRxuJqXsLkUm2Nntij62+yWMKt0CaDWhwI
/SrzTA15Q02ze8ZI7QJE/aceocqe3zNgA1MBygWwLZ7wpZc9QDT2HrX7JxSpFeiLPt4wc3o6uZQ1
lcrqRp30mup7vXaAY29zIIpKml6obtc1Mf6BkFy4PNz8CZ4AM2dCc6FwcK9fz7FOugUfI9wlkj6v
LtLrHQuVuAcU6wBenOOsge3eW8HPKZeyg3Bju8CcISDPj/dNSGgXOIS7y43cfBccYpeg7ZOsyhDf
EWm6Z9WcS15RrYojmpN2paa9ylkB/50hpS/FisB2stqybMlNtqbv++PyhzPLOQHQubsgT0wCJXks
bML0y5ioDtW2WFtA0AtAMgEdywrUDSe0PwwH/64XMsZNNuqQK1/dEZlb9bw4pTmlnFqFsO8rM/RG
Z0zty+DXpxMLgFK7WtSYmuUpBKIOlH8fPFbI9EIuSyZXDV/W7TfPO6lY79Ej8z4x2LnpjfcUsOJN
mK9XR4un29E+YMd5RKY2KgBboO9cDdoqU7MHoji1o9o7NlienHYIFP2ji4WMt/LnQ9HGMDCgfMdv
lLtYskPYsRDuWi9kXaWv56aweftakEIdHWCh5kfYfGVq93SIjSalxVEXowkfEKT/MUgqUCc19kfA
IzDii604AFdJtGOCUS77rKq+8FopW9E3cFoyCkqDtaAULYbUiv1ldEOp5Imjwfd7SKzgiGjJgvs1
x+P98XfcvpFlzsM8zbSWC7Vca5k3UwlchFnJ0fDXPunXUW0FYrYgN4k12kHMGdTAhoiFGcoSOOLl
I1+Rd4UCBaefCaqzRubwJTE6rK0zLVBa9m4M+k0OGzmeuFk2IDWT9orrYerpK4KE9M/yAG5zY3ZU
94/Szx+/kye2hoiVyybwmXKiQ6laCqdkQP+52A3gmyJzOHeuMzaW8MGCQdFeU40R84U9teUiJgP/
tjJ8nKwnscCgkTz98xrB5o03DU4t5Ia2G9k8eVN+mPf5NgUuNIRsSjKRa6DW/Bq8L/XRZwE16OjM
ZbliSbukqGsRoXD5IVV9qlgtOC2Fk30trZsDCA9Qrsod7IV9lLIS5YwpqPGMSwbeFUryt8IXwb1j
+7pvexoijGNTNePChjEH1Acm3623NH7hYP4RuyopqJOc7cqJAqFs6ghdnOrG0IZ7H5G5BYgfaOGB
9ciHjMNi4SSzXuugBF591zI71fR5qZQyvlaeIsXITkOilpP/DMWWwSWmtQKWAG0pgHN1U2mikdDf
Am1YVLtCwgFRNuQ6X3UjNK2aw90e3v06xy4cYsq8912k8TfEE17rnIl+Z3qgufSZjxyqcBNtI2jr
+n2tG3d6r3sMhYE9YKmy7bN5D7c37pyWUPa+kkj+v2BGHJo0mzzXOJKPT5xKaE86KMElQTDCYR4k
oTTGmFdm5I7MPRKTw6xhXJNiWINx0bHBUIT8ErcJ0zx7Vg/oXiMu29lpPVDoW8swA5SN+oNoS1rp
3sMB3wMQrR0xWDcoAtBj0BMVPk1eOG/PSnm5Wjav8EIpz29iVOqrxKhBvydE6siNRWzn34y59Sus
PwNmSx3wWRQfyx2pYEj5AuW/5Ro0BCpcF+lb/pNds1739pkJv1qIuNdRWi4JmFpoAKUlfVumIv6K
p3A+ra/ezj6abJ48lSHcDVPvojLvzri4CEmckAU+BBXxrcSnbSkHyUFIkECswQISW55dYUCPd27y
wx5GA2fkFtQ0vUgWu2+lLOz/YLPThn7LvioGq4vbsIe4CD/h1L05wXJiAUpi1V9UoVNkeDOK4UuT
ULJBJC6X5QRP5cufhK0QFANzYQSmXpj/XSB+hmFuV4Ushw5Muxl0tzb7w6SHF1MJ6nolCmsqJUwX
/kAVs9Z7wUkZtYvAgtjgj2njqCJeBzwvwHGLIOHVervTtb1lnP16l0U03oemALWH/2tPczJJD7qC
2ASQM2dhKWdK9U9fx2dBQu4hFiIcLd4WG+fsTQ0/fecJe/oQmnbA94n7bcLeNQaPR/ZU5iqwDOX7
J54UvTYvuZbjA5uHXEv3v5PjiY0v/hfwnfBG0QEYyrROlD3+t729jQQioyayVkAQZjcEHCcJghQt
6+gGHBbV7I1NG2VcqpVey/SXHDOQOsFXmO3hwyvNglVHu/AerCVCSeLmHDY7vDRivM3/gBW5Sc4m
ucJhM/G3ZINiakA3GBWJJysCs+EUvms6enFtWHc6zKsGBup8jqnBQ1XptJOGucplln5jMoq2gesX
tPGT6bgmU+Z5aEiu7kLLIlz5NUfUFoKZGLz3p5lVDHTHJfdiUq14ZbskQnQbwlHxRJT2YcddwkCM
31OdtrOsHNipEsasXX2VJQhWmt2rSuQH74Agsr74/MUi926/Ii+fo3M9IzrMPgFlGxwT/4AKvc9I
v3VKOhiAJJ9hBIVGElnrkatAhZ8uNgsHYLQKy+wev8hS93v9zGJUCeARiRIzvLtcv+/lF8nLmb6x
J4lDSMnDWVF0xUB4XuOB6ramoFWxMNO/87QLsqpoH8rNXa2zLJLP3BQIbDNIsclpaJ3j5QLUb34O
wVhx2Prtc2e4S+6fQ8l+uBG7SvpW9aeMkL4jA+9yQjPSXbMwYG6tDmZHQLW65P0S01mwqeenM8DU
fDUfjzTvbhNTuGFI4gsfoHKuOPtLMODACUCNv36Ho7ha4LxB6R/Mh4KnL2ZnZAMs6k9YEBmmpMKK
UEZkaI0sa5WPDlBGbSK2YC1rAaUAgiUNGOHCzk9Ou/tRge3s2vILsstPveBmO23zU7MoWIG88j+q
fD0MqcbpTmOm+EknRe++VCpo9XKcR6m5MA80C+JSSkgb6MHDRTbYczKfO9Av6aA6repbner4XIGl
6kfN5M8tJBJku8SPlKmSafVTyEjVxOCTwhiZHIiFXjfXQ3AfoGnAyFG6gxZBDxhI7QY5Op+ZPqBI
pYLDmwAOEnFxZ4/ND8I3s08w9KhKAYmayFHXvcuIoyW9Bv3WUw71VVeJvqgpAX9tzunYd9FwWTaI
Fm4bDzujrHW0JQVXRSjmpCZWkNvNJzbUxBI6FHY25v/JcmXJtlSwugNfOUdPDxMcgoMnMXm3QPnp
VvBEjPygBdBrDqJQmfZ02dpw+Ncla06IFpwFO6rcJPEN46Z7Ed4nczh0ZxXwNTWjjwbtNVkxCT8q
D4XqWwrVJhUkoxqH1RH9LbkgnablURuWuLlukK8JT2X4wwB/d1OonQrbPoopDqmCqKop+36Md1bG
pDw2mnWaecJcYh7OqbbTZn7PwFlIkRp4Tf19WRmSExy/7Urr7bm/7fcXzG/FiGds8fVDSoxt8NIR
nDac4zH2beex8MpS9L/VjZIYLM/MWawnpqLLJxWkMKP47JleosolwYiCWwLrtl725HRSWfpUeVo8
Jc1I7gh4XW3gicviDVW2/MlEuDnbiLHpgvisT9xfm767QolylDDlyg+YZcatG7Y2lBUB/fJR2E1Z
J38vxCM39F93M82yfEgivqR4rmlkNeiczjSgt7H+G4skYcyVak5epV/1H3dNoBW0Np64B0Gm8ngk
LgiyV1liDnHGB8CTsgLxPU4DoR6XrZEbKaQ5IRYH1KpYPQWBmmNmRLe4Fh/vvJU1qF6aetnRhqA3
dvHaX13R4xTzyANgD5LFJBx/nDE+txrruE6aL7K7hl1voF1Tu3/z2rddUKN69CZjVh6eMxYfTEsG
dDvzbzj57UL8jjH3XnwEaWwsNH+o4M9c1y7DnUtfo9fCEfdixEJYJUf0dE5zVPjdJYYAG8OhjYpM
oiUAAnsiO2Okh9mixtC3aMswajERJeoLcntc3STunuCJjEUgrt2HSkEE1bIEyzHKixoRbEBjVoFk
IltmLmDAh8c1mE1jMYrE3lsMSOYkyUsEGzTsipqEXK29aiEMdRd5obb/SxNQcXDI9ICD9aHTlTS6
Y7JI3IutSK9KDMDr6+RBUMCKkCXvSXMxJc2aHcl2aNDnZbwWcK1B3T+EI34RPkSGKqzzPZZo8bgM
Cxu5V7qxMSuDhUu9jwUpLjHst8Lc5nsQ/4jYJqB8DeK/N5YJRzWIRFtkHTsjzgRXr9ZBhp91Bchr
h7gkUeQ9QqAMRCnGUleswlx9wfC7ZwELLZDLWRwJMX2CXCZFLLKLA97Ii957g4rE4C7ar3MRalKV
r1Rc3htpVku5KNiZgcRwOTvoUb3R5xfTSPuy0WxjQjrC0x14mICgKkyfl9RpIltTziMr0v78MFPm
Unt09ESTXq7DLgVf3v7QmAwzOVoS48t4GLMtN+iPZ31lDAxQhvJDFfZ9xraXqJlcu3TD/A+Q+vEG
SX+9aGyqvuDi6L1cDSXQMMvtKNq7P+nkoIOqJE5vOHtHxobHsW75SGRaQnPh8Fj46jwhqlVZA86K
dlQgzVLnT0a7mcM8jbJB4E2xDAeKqmajhv5OIkmBd6fl1ctUhIlSjIX9iumDojzMmdLAirMYk3Qr
aqTl/ao+y2qDkMA/sY2r+8mqTHp/XgLbEfRQUHD9XriprpS5SUfyfKfGIjers1DNR9PXZ/NKWd/s
f5cEaANVjPZ1krUdM1NnAlIUmA2HquMtMuMBswauhunZGFld/dyAxgynIvmJ8ocm62TPzxa/vcKn
bkRS5qDqMWLgz1T1zTvOwa1Z9PXu9jYI4viCgcLF0f/d7ByAR9WHalevyZXucx0WEJwPCxVgB7DS
GDxRGa+Cpjf+UfkStP72DfYRJqkZvhue9uyCxJ263uDTAJIzEnhniIz6QrR0BnpeWBN11VrkuB/2
TxtgEPK6texMkXiTv7H0l9MMIBLqER87hruu3DADuyxbwsmviOQ55yQR9hXctiEjGDcNM2jjor0r
LMn4flLxNUMw0eTDfots1lpW506adSDEoToHqSBCKUW1PWNl1FpPIm0ptCKplzn1c6q8918iMty5
6v4gaHRBnREDUrWdt6AJQMle/qhJXGB2pjTNCrm0SxvQ8lTfuaUciOq2HY2PysxrNWStENlIma58
zRu0r1byRpzwaSejsfRr+NVhV7f6wS8q17cLV7MXA0gFHfynbrOd82pxWMjqebGmPJo3TCARFnLQ
0iVX+wSHHlJ3+TB/m/wGMDfuU+97papsTCa1LQbPxGaXhYAXcqqtWYrM9ITHAL71TuzRygYcZX5T
BVDJryuQrjcbkOx/I9ThlYROMwd4JzFuvc3HBe6nJrAXugHlzEH3COK1nBJ86Rfzv0Iqi8LY2ea/
k90D3fLBcAXgpC1IWxlEOPM49PpwE6x6gzH7SSddP8TD8mUrAoTXlssfDXZTX93fHfKcPswB8Vn8
mRd6r1VaRJ7CpMNifuBxuD3qVajntoA7IR9ZphMW0nNbQ/fuqPDI3FAuXYTd7es8bxpuyttxGLn7
3Zcrz/Bz/6z/G9GL2bo223d3TP4BihoN6MkhUQRZiQ4Sf3ehn6TnaqzV8Ii/KJdniBvCxWgYrQgq
smtsP2/CzQMuPQkHDzktdPCcmQ8VxFd3+43txXXWH62lTvrHYkQXxIalBC9+Tf56j+aXOhYdPl1R
U0BFi5NizIUWGtrYkVmy3jlfHMcOAzTMDJZg3zxoLFGspgTFgH5Ysha4nOPQeoNj5XhNeiXYn/uM
9u9SRutaVKY8Jq7ZXcYb1vIImYnw50TsL/cn3TQB9nlygnPV9uf+QpK0pmZW9Agyg8JdjNsqSEyM
r0krs8I7+B5h4qh5th8MlUQRE6T/tsy9jWX7QMafg23g10UmkCGoWJm9FW4EYkiCXBPyKJRjTD8C
rceIgSzSfFNVuaBBhGzMPgVrATmHRPkpCx1wVjM1FoxC7UXSUGrGy6w53Uifr/xdxi/kK8wpn/Ib
qZBsnYtQqKOVjwUYvVvsinTKxYgqhO1BM8obKJcnxDlNUtJ2V/P0pHHxJj3tGZ2rOX7SQhI9bjgO
7wdwQORGq11NhauweWLriZVKwcovlQYX/3hxVcTzbe0L4hfKG3Nbdin+aXIQ/5aEWJUMMhb0rDxe
bHOVhlBLhDPrPHwAt57M25Nsv2gh7dsFR89x2pqjRuv1Yv/Zq80r0gJ6KP8W2wilIoXnLKBARyOu
UZnCmPD6jXPaou987rtktHaFhNtI+zW4OlgohQbsrmIzs0KrGonSLu6JYPjRyyJPa4/Hw2W0Bej/
tDE142sGO8cXiAQCrebFVnUzyfNLlx8LmNmUMjxci1h0HDtcQUJng6DAIkZo7CutplUTfPQz6lPp
IN9zKriP0eMQXdvD0KlRR/fXdfrELp8p2mXr9JZJ8soKw0QSHG7P3hi13NWxFL6UjznVA+BNKNif
AxYqPSsID0BXqEr+EjfDfQIjATklvauKkPOnO9gWj8nr2SUTTu76IT3+RWhCZ+EN2op9hM2bljab
h+bNj2T6iU/b57YJuPmjSyHWmv0e8H63z+S+usVyuXEpBY8T3/jxJReDcxoNXQDlJxfXDkcH6tYP
2WpvQ9U4S5AoO+R0Eg8Ei4cEcCZ+gfIvXbCtd379SMyHPpupNgy3yS0YJTvUfVdVartCQhEvVtHZ
FiI0BqXAPXlQ7C8mc35b9EptzMiHqbAzqA4neYjNMMEE9Y/Hlnx+RTuOHXIJO81E+6oXS7ysYHj+
qZJldm1E3Ovco5PGO/liZtuGPyAVOMANAQnYmC4NouB6jOLlyuFtikUNcvKn20XTq8tUozZN9ayK
+nHb45NjUoVH8joJNpsTx+6L1nhI9tlyL2doq2d1aA/tfpuffLPdp8xjobY5eWcFQfzBcdBaLQa1
IN9Yjm1WxRM/kaVaEDd4wLsyDAOAkjjss6ruSvA38y5lQzmJri8vToJAymkuac5FJtE1kQgY0O3Z
4JaZJVJWM2yVe8TGBsnhUJeQ8XdYRjCF+QjZfCnPNLGS+z33x1O1t1g0aXPZuRzcPyRMaUfgEMmL
PfXFip6PKujWN0mqo/0UoKoewnk6cCC0KEdlLdhmcgoARGY2h0vBrqdl+iGDqBdTF/xr4uekI5ju
ixVb6Qm2EGuGAGim+B0Y70cjfknNXyMUns5tyLXT7U27rdE9nj7VD/WYFLqtwnlm+4l7LwBLmkNX
Yf/NhqnS+OySwq+8zOqpovxOo+svHMh0qVcCcZKVrUo6D35ULI81dpaCFZyzvRnxiR8q6f2zuX+c
L7xa/LTP3vc679ZmJgURwfbTynQcw0fT9pK1qTwGDWgNhMrVla6yY4g9Lx347YwkLx0/Z4XOk7lP
HfWPPYvcnNLDFBt255TQpiUjY81CAJ7JXhzjM+HucYmXs+8q6me0Bunfcu0WPNfsAOSVpsK8megL
vaKqUMkZpo6nWBhgmo9F2MeFXw9xc3OUyFqf0DhWcp9105rEEMUSYfTsGh25GIhBkmezl8QbIkR7
X7OjPRAEbbQ4VAl9qL4czOU6xuzZbDfMj7WkhnQX09nC63e8sAxI1ucw/TCAfW9J/Yx/H8aB0Lns
wPEyRcGV7XIRfkNQc/rp2Wkpxv0RYZ8/PDxu/hEnoXhJFfM8DpbOOZ7sNZwOHvhOsIAeEwcJ1BeY
XRrtIpj5J6EHt5UpdDcaNUFX5viC9Zax+BbK/Iwt1kXaEFbPmToKvpoCEJQ0cuUWrDr+Kf5OKb9R
kwpqunrDu6cAmqCj2pJhwOXKVfAyVmYOvadr5AX6qkr+7epdptLD0L1lhkEWeB5tOTutc+Dzroqi
Wqg+ra5HvmeKqDvLE4nTPVpOmYLk9Or/feHDcQjYcwZ+6Op96kQ3SsEiGbVAUbOEEFUceoyfKc2r
rUlmWhqW3p5ggCZL4jsWSUwuPwNzBn6rozCG0/9Dzqg5XAnjdfZ3Ahez0WkFbD+6/a7/AkhY/Ec4
lY+9PYm5m0y+ESKkqSvR7cXv6sy37dkXBKc6NoFr/Cut7VprBYQQk0YlmfwB6ahQtRs4wuE80UPn
Iyxx0wDSHOHCIygfDoFCICrDkMnFb5sUbJWUgzin1L5uqWR4/NqmPJRIcRfg4JaztRBFfqlB+3Mp
Pwci1pC5JCu2OMMxiN2MMvBhdYp5qCELldANkNZZEYYE6f+OrbTQoV5UKCAfDi7vRCHLW459eLxq
yY/aawVkfKe/VDv1ghroU3DdpU1xcLENi16CUGmxUHvYgqQxmNvhjHCCWVnt7l7qMzy52zQOFk0c
31fBture2TkvLuUu3A4jV/kVV8WA4t2n86dTaXc0zvDP93ikAFMZ78OUFJyppIpxkm+Ud6VTvcvm
Kl7hfk8fJMUGHrXhVb+MtQN3NKDPby/Ze1+m9pQlzpTE2Y1hbl9jgD5MadH6WqsGYf5L+i+cXNFa
ftXF2lYYbaZN7vNKJXUFNPZGMlJTttD4J6NbVv3zuTpqJgk7/vexMTGDEzWQYymqQOsJExWnMuFV
LPbHdoC2YsFlqJ41WbHWv4lpBxsCoT7X/Z7PmS77/dYMXxXvIy9waiZlIiGoKx/QlCQA88M5/uoJ
ATOB9MByplSXxyJv7Lu4GqCqVetDIDM1zt9Suu/2iCbNpkn6lxcFyE1wXBtcIb/zetJmGLc7SnKa
g9BDl6lnYrtt9WiiQJFzFh6vxu/Ck/TXzNpeGJLmwOUZyqTtDKVgF0DFgZu9XcqnGJKalN4V9Y36
ODUMveDVKoXAAjlkmE8YXwZsgmXy+lFBbiP/iK/39N8XNYwGx4xMOQqL1LNndXm2cxkdB6J+Obaq
AJ9XxoBZg2AanGl6KhSCnZa/WIo/6unJoGKHEbTTrd3e53IXvALX3aWHFc2t6K5QsqGfvJque7HS
BJYvZz0m9uuU6ZQWxafhwoA+8yT+M/WMG45MAlYXOs2dwMKqwtiafQPDmCzjzY1AflaEBI6tLqKz
qX8bcG/cLr+H8dKl7+ZlNsNDcmrzWOG0VHPS4CifKq+PA5cg7kN8jHRNYXzw4mL83To8xob+qr+b
KDglvfq6f5pwQdAjVRKfzOlwfqUqrAJ+UYKoRNsUUO0lzoIMGODRDROQWvAJfnhMrUSscCdfH5qS
Sqe8HbxFLcESpuSR9TBw5eFtX+QWWDb5vhIdOP0HNHZDoKXvaQ5GekPXK0RYSSFtYeUjYuqhhM+M
so2oOkOuieC9sLWd5fv7eNmTroZAIoQvCIgymOQI7dN4aUwy3H0aR0HkSX+YjriktnEv3DZTzz2V
YGSUf70TI3zknRI44LoS6LGITc/DZ+dFLuOeN8T0BvHCtSeucmHfSU06M1BLaqArQMe2RHDw3yEQ
2Itq7guZX3v+yyB1sYCOFiNfEVpGEnk7cxpu6a7QQSULk1fG281jda8EJZ8R670Tdyw5wmntTCBf
GrvIlzGGDPDbLXi9PajkrXXSwSyd8y+KVV8kv+KxTYmdxn5Hx/L2TXLXrX2B5mV/uyGJIR19fwNu
88cBKR4en3uw66oVGhdZnKoVipLQY6x9KrcgZLk9L0+vtH3O2z/UZ+97BG3kVJ/qFbZB3dXjamHm
BzpvkSnAZTW3TgMIRiOAXesaOYmzw0AV8EETf36VPeNzjrpG0wKB/KWTbT2Gfc/bzhX7k6YOKl8z
wG0mdTuHglV5oBjtCINT96yqRbfKaKR7E5X/xh4kdtSe92Kb2OL7mD0hjto8a25M8jRyrsZcPv07
jWXrd4MR/Mb9EfJCuiKbTxYBOVDpsIrkyZl0p/2Oc2AekKXPprb+7M/y8ummVxLmii4AS/G3Pkfm
z4sxUa5wecbUUhbkmwZwI59JYv1Eu6mFrRqR3suKxYIWir944c03/RwcTQg6HeFxaw4zh7+7UN8r
UH3cQR+6fB3I0+1OI5+ZQu0LqDgOS4K/IzpsSFwFHID7WvnZe2h4aTdMEgAc8Pn4BTOxGpQIj/3e
DVGTZjsl/54MPmvUemKKT+PeFl+qX8H+ECpYtpYCYOQyJyS06fJFX6aOpFWZJJBM/pPiaQyA11gX
fbXuFBfDGPNgThVdtwfsUjc7eUB/xVvwIC6XDLo+B5VGHhpboxHJS/+vv6XPsTqWQOi+2zGLQke4
rWbvooqoqnI6E8pame8MwaHLNZ6wv/6AI5wivfKhv9lGpW5ZThV3I5X/xikdLBetX650A4/tksoh
E5syn6jwm7ykvAkdYo38yfstq32bZ/Qj0iBiKZj0ZVmbnW9EShX5aDlmW5mmSqfxPCGZKXzg4h22
gI8P5rI810cNtfnY51KSOkjI6BQRWk4Q8fpJEyksBtB2npVtRveCXa7xSyEQDk8uDss+oFSWodU9
WJQHXgUNpdYCkV5/Ccxp3snOmZsshm+2oSaGEXR6q7rc6z9BVI3lruVIZSng/B38qoQn6/+vDXJ2
LS18SxrC5pndlt8GgPL5rXAprxm5NskA/x5ZHcJooW2XxJyDatvM3fmHu8AdqzVXVJXU+wMhqNkM
8hFe+r1yM06Q25bYPgkSnPep3OdmptD1jFM9BhFc/pqMMo904RB3X1/W8wyjdegpUGttpQu2AfhG
SXNzwVw+cpD30upUWdTWC74SgNKA4OVc4zL62BD6p9c1BR9XUZRorgL5jxP1H2oqJUBLmUgQNnnv
n/pQBzQq5L1SDKiEkiUc5VYbFHhIZ2nZchnXUPgq0jqB6H0+cG87OwFX4Ctm5VBYXv0odd/B9VsZ
V7lgHjxiuiSM4hX6uWKNlAJ60a2ckrt5JFQxjczGHLSlQTV3uJLL2CZ7Gzj728QnxV5PTH7r8LXd
4FYnEc3ZNksohyu9p9voX/9Qq1JzSZ5udPE47gdSiowZoeWMlUNQVyoTTue1NJjoMCmkiXZOi9zo
m+3/kH6PxOptLnwub7/YRS9Fe5IFM3dpavL89ftexuRIAqe/RRQjcbhZVHDSLtwIGNIdzUEaokWh
KF12lG+Dl7lmyqzeHPEEmUzJRI0lA1aTa81DsCByNbkUavD1NWvOfJtMIBlE9zJOUFwdzVW9fZJ4
k2pBj4qqlecosF0mhHyNd5CZuCITKG/gN43ngBMo22AHkiYoONzp+3mcRbZu/gR2hl1lT/cHT7Ed
PUQ34Wqgj1oHCjepQfj7QOnr3i/W7l6YXTpTXUAISXeJmcUK8YHFIe2Oo3QmeMN2tGGezuFXPI/a
WvKGRB2KjLMURF9Ez9qdqstJQYp+7PxOZXufSLPk6S+38r1H631auliEsf9KNRugoDQY2qI5jqxn
SIxkSaq9sFVpapvoHgaCgOPYgKJ772l+a18LFN8NLZTP+0st9R1CmP1XaGWtAL04ii8PnBcQRhjf
m7noRNIC37r+zxYkNzMNNPwDypCK9xHuNyiNJxME/mMBMPLrnf3Z/MeTJrUvmipgP0f6ehV5a96Q
KrZ36X1BUMrSEiTwKmadZATlaZZP/dnV4LRgBRwJT9q3GIzLRLD3PJuPce2KrvbBL+l69HN4MkF7
v7WlVqoOYw9Of58K6gcFAntnMmgnY7kvMT8p5pkB8UJiPWnOA98EfR2UYxLqaJrRRxNZgEg3NO+K
nFalO8RkpyjqtyC9XZIDa8FpxEdifXZ8EcUXKe2PjVtmrd3JbRiHZzQx3KLzu5aQ8hHSOWJxtPHm
bFeuYzeOtrj1HROnyVXBomUes2C1SCkModhdOqUw9yYxe/mwQMpFAectJXuLzCgB1wOt3Xk+kgi7
fslJ0rvFsy4EO1Mvok837VShwyMII2IghRuU0USdIRucnifvlf0lcTczUa2YMpD2Z2AxD+9oDaKo
8FdIp61O0JOT+VAnjgo19WdVjOr8UGz+dHysxPu4pQtLxr9YiHkIrS39YXt/9JLBdgVzay+1oInD
9ISpRRp5tcouid8r/2EUeKIRw32sHLWsfp0iAoj8PTxz2CKB3bABvdBhDGjriO/zTAmJ0vNOcszV
Rwu9fctnHisGFUmEXGS6q9uwtCa292igixfth7t41UUdIGH3QM1gGbvfxza1eAWmb4CkBjbnruOq
S/l+KncP3+NVR/tXMuXSweqUYbPpwQN5MdGCmt56QUBbmuThztXHQAgoxZDRFl9mUir6gZUqwDQ7
TnMNipnNCz8HFTYJ1IDMOkedqKgoyZ5mvabWI6CeO0hzfRgV7d8Z68yoSqO9bVldhhbd7FIlq4MK
W2B0mQuwdiqlpy0PC1Fl+Zi44M3EFmcq1YZxJFKfZf9Co0sPXOe11wIEP6U4q0BXmKQ+FSzQG1lQ
VhQALNN7ReTJZ9cyAva5h5CU5riZQKHPD7V6jw6OuaItu0TLlKuEakE378jLuzpp48SBDE/g4QXi
zAIQpO/anQNu47+NtZ7ImkEz5SM6k1HZgjGt+ULaL8Mg4LjzO22FH08oP2Qdh7Qgl7OC8uBUZmvP
I0NOldC8FmBQDVm1z5Is1F8ynzNzYOtiLG1iKTQZL6K7yrQ26obnyu7W/zrpGTUYOjoFK3uF0CMg
kC/go579ZstnW469mHwVAQtKaO3SWy176TsDJiBNc/u2oOL6qqK0XUbm2kOYKEyS+8PHs7KSC1mY
gm+5g/CaFxZ09P+iIj2uvPKH6CuwRQPtI3O1NJlbCAu0pXL1wDAppvy4cdaHzG9o8tP4ymKqSESH
nbGeQQTCetz7PFWVEgiklA1Xz8v8s2vFGwg1UOv0WBUkRf++twajlytQCpEb6cwJPzbeQTvzfzdt
6gg1nzmyQAA9FMaaiEO+B4q9lGQgLSA93/WMqM7tFG1TBtOALqq79P4vjL/RVKtJ4P3o2oqdNckB
0rh4oc1d56wuvtCHQ7BDujTDxy4tYniWA/c1XQGTnxosAAALmJWsCn9vHA+KwAiQgLr5lSmHaQ9B
gvqmvk/6USuEEGc/27AsjDjV090MO+OqpWstYemUzrv9SrfOUgrfME4mbkeQ3r0HTQoDFV+eXj/x
hxGA+bM3gKpKAMUsacn5HDaB0v4FJ7vBWtYvk4WylBXdp5J/q/OBh3DFs+kTQ982Rrdu0oPSWjPd
pttxLFEjmKcXWMu8691p4v33y0R/K37rBjnwd/AMZ3ylrN0iIm1dXnVN58o+aIyrVV2ve2dDmp8v
abgT3BvkapA+7xsEhAGeTO+AkbecoZ9o+OIofjxpvNpR2+K+wywML8hZbibX3L9U1M58p39x+8X8
Lw/W27s37wLLaBG27GgkIM+AYrAqa17s1oeS8SfVDS/16Fzrf6U82m78n9IX5AlmI5pgjzU5ZYW4
gtP8kEQ3Yk3oBARDw7VG+HgeVe1Opn5YpwI69wW5V6hx1n3dX5FeyGaSpZe+ghYotQCFtInOYA6W
2pZN4wNhR3THp3XJb5aF55IzZaDsXnC9mREzyslBJ3FB0K9TQ4K2JOkqqEznRyTHU2j9pmJyz8dt
vOC8X/4qXZZqARrxXuOzhLt1IKFFmQUDYOL3qtKSsoM8VTQJJWsvUzvGLwD10p2LUHDeA4PGu5qM
UU4S29X9VGfsFeOMcFHNSOYvhm5FuVIZDw5NsDknp6h42toRpd6OFh0II5DSO+LiaFiUQKkPTw97
189hpVe4S1sQejT0tayIkO9LNKIHMjC/DH4G3JpNBfwhZbb/E4ARbdeB6GCphqzCn14E7CFP9MWW
qgUQMULI2bhMQeg9HO6XKyxLwDK2UkGPZ93WiAkGxozfHAhTMumCna5w9GAWI6QKcRYQt+THKBsU
6Tz1VozWs5wpsLZ/490W/upTfxzczkowiFKABPzAeC5bXFjSjtht4NquU/6cwMlHDsRGp3gHbkeJ
tkTymamLWH6qauIW9544G7+4qeTl3sAnqQmvIeC+uM4QrB6SAfW5lW9Wzx1Gy9tabrZnG/ro5rPQ
XHt5VmKV4eYzLqTmqIDwPtcBrhBGdnbzMe9JwqYrMGqJNscZJd9zL4OjvpaCVObDJ89E1hczMXkc
UW1wkqFx84Wp5ZuaJJDLCNKayonyoL3Ik3QH75ABwbL+PNroVUxXBJUouGATHrhhuoVnbTz7g4v7
xw03wQqORIDQ2o2VwnUd64Q2Nwbv8uI0nUWlQ+x+HgZn/lqluB7FABCXRyZe9VcVhK44LG0b5eJm
qCdCIj4/8fa8KPjxaTI9PfwZeccQsWiqhtSZ+3jEoOMvr+2Ak3KNYDip/1zqZRP4Ni7EGIbfJ0R3
rUfA3Mga7nx4z4uLjBR1c40R4zIOx8fuejvVY5C5R4w6TxgxQJmiSfgcjQAW6kbZ0+tcVQh8YKQJ
FZqdWbCcTnY/L9x3RO3i42fa4VBCEFQYKGPJqN9/XUCiqZijFHAehlyns3747MymILsxRGwNFYxz
kwNot8KzkBAsUNP1YsK1KV/5PNC+WZj2M+3VH6m8ZGBzM6Q585Q7wlpErDrITDCIdLCdwQFdJXUg
vomOn8oxsp5jMxAj6Utc6+ofjuw7JQELGVOwrIicjtVK1Lj8dZg2g0ojd+8GNwxzmihE0sxas5sA
thggpPns0Hf5MRPSa4f/Ik+HLeJyatnrxfYgmzAwPMWBVD8SlPxeOeTn3WAYVlyS5nn7/0r0WP0v
jiZWcersC81+sMuglxZl00FQsW3qJA2P5taDFmpU3HKmEfmw/cY8z81qG4T0qOhqitBmcLd129HT
0Apj82vF7nWFyb+7GKlwsk+4Y9kCtCYAQxS0lPwpy92Ec3DAlcVMew8fswpvMGKNn4jjNtWMVNZ9
7TM5SmKpvMnMc3aw9D7V0mPCjuuqDydwBzHejR0YMWfM170tQeAx+jeXIxR2MCLy9KVc6UgDZggs
pL/y7AUJi8zWL+vbX62z63bNPL9hFSGYvVhvcM/DSnyWb8fFH/UGHoInD50zdO3dSMfQNhl/NlJh
+aUm3KGray+fUUOiA6/0Fz7U7Pgzae4LnC45wfE+kYFxrDS+YWcNclQ+Po30TXFzPT2CFpwonqs1
t2VbNnKbP/Q+7n3rf7tIQ5/MlVi6IELIIB5x9vfo3zqESdUGAtJcsLvVENCmCDV3wFVUsqfsaxYt
lJxlv7k3Rt7ypaJ1DQPqEZdO3JCWf4E0Ybaz/QTpwdYmdPX7r8WL/qvetwjUlKfhmxSDRmuz4AhM
1a9P3swMJsXLu4S+bForbeXjuurcg4DC7t3h6yTDnn7GD/MIWo++MQWbn59nwPNO4Sv6VhRlhnJ+
A1A7G00mwEwn7R63wc4KoDM6f0N3/GYcr2EK51Zh/4ugRX7NgoZ8sZDW72slgkXjbHW4T6OL8hQp
vFjzcoKABDhuL0YlZHZip8PGeYoaFYxcRS2mOMD04ek2ZSSdTmmTQZHyXo4o6hGyR3olH70FR/rq
XyfqM3PDGqSzpbONZu47+SIUdS6Eb+lUnWj/SExc80lvknpkbCdK9TQmWG8zTywI7HfJNYQVETAP
KIMoMBH1L0ORaSbRXZEcLVFNApO6HaJI9YoFBpLBGe8+r5eRVqlWTQfdjLhV7kw2lyEpgJeTZKxx
UjM1bNRbRO1/6QErppCb3BTlLe59ytEZK4Ja3Vu9rl0yZ/qw66Q/zBEJCpZlC1L6nGlSr+cEcSeR
JeWH5PDOOen+h0W146wqqkjjN65UieFw3916rKvdOApeOcUkaLGpHK6yhxQH+SyNqPWL+PYYzD4X
/S+7ay+IH3msaKPx/cTIxBF/RxggYMjzXmsGW108mcPSF5ujO9icKe7ezI6EMBfyuLt9UWOH4RmO
Sep4RWiBwHridsc/pROv8XawC+O9WQk0/irC9loyLVwDATTJHFfQmr5cl/1k6SHRPvqri5Z5mxRI
C/DdDu9tGgz4PYV3tocPc7uQ9tEJLcAfcf+zoNRgKcfAmzEpcpqHSlBdRCvI0cJ2MonIpPacDnSq
DGFkyqPMs2i8UN2cccbgIYevJe1Yv2tyczmFTqrktlmnVuPL2r2GuTwG1Sla/DEqronKMxIfrimE
zzRfqQeuD5GV9+0wv4eRsgn011/djAVIK9I9CGr9fEPqQbtYo05cfUur7JMKVoYFe7Sokviagg7y
MOKsWJJaZ9c9tQxuPh5kSeZ0xIwD+Xi8J5leAg/0gC4QpLUHqFfCNBLpoXX7o/Jo991vRHkigvxi
9c9Jba/CNsVOdjd4YGuVw2Nw+MtqOfZcecEI/z7Pj23XVubAgL8hhIjzULwDqmUvgZSVwdBU+wtw
PbaY/aC+mmcld/IoHvlFa7zq4Z+fbmdEWNJLCmLgNKdZA27GfHDXRXsOGBgw3sbTYVpHmbMC2wbG
2LECfDfk16vfHyTWxdgpVRHLPJEM1DpI2JNncqtOJcQbdJgIjSfVvZeAVkNAgEUKwoWx2kqVpmJL
ibGhN6z4UOWXHzP2alstJylCiHZcg3KWhXg+YqBRtyXWaIJ3d0DgsJjxQgPlGXp6OGGWZUEBEEaY
SAZ/WPjqDrcOpFMkXaGA/i3Mf5euAd+9HkdXAy08CY7ntzcmFmMgZfm40L4lv61H1hK6O3L9LYUV
RixTTlTru0UVhjwXK3XJzYC6OCgAW5UHrDAS4pSxfi/xr1jw5CmEQCMhqdbUJgm/smg5TlPn7Z1b
BcxWByji6ZwL6StEDvsBuPu6dXIKnR/fwLD3g1HQWVgYpBcDjBNaiXNYtop9uwZ7Ao32xi3H7VUq
aGWvUsT+IFaY+xM0YREdT/5kanBqBuUezgKexXxM9OU0Q89lUZRfCkJxiu44XJKO5oL3x0fQq2ic
6jc9GzBZC265CzW8/Z+S9eSWQctjTVJfe0WKejVtvtqSEs+lUPA/G0xIcOBEBJ0f1BVt9JWQwhEM
kz7IAHXaFNHU7A/h1BjJPk9p3qFf0SOMLJysupuRxXRMiAuXB+avE9t18s6fOEAdr8I1J0JA3xMU
+fM9gwo4XFkNyv8EuBgr+c6x1uTLxs2RJQIXCY3xC3v6HwK47efT4C7N7cB7hVQWPmDlAW8t+2dt
p5v68LhX2tNqbUNKjvVNCje4ToQBKuVG00YnhhMTTZ3SN8Gpr4C+mBfjkS76TcR+dARWxXwlLyzx
znydS1weHPAKoFGrht6ZlWYOrYTIyfYgsLqfE+y54iivzv6nk8kff1BeCsDChPcDRtNvYRaLm7uf
m0pe0nLmUhtW+JF5UPWi3ZAzF2MyiY3wAJxCXk8wUZiguSGpd9Elru43jLO4ohvytDKJOwLSTX2N
z/sKIxF99tSBhmcn7w6c4Ww5pfSsISe003kGYE8heqtorw6AXDUXALixkvYTo3rGrN48dtRTnJJZ
KgURU2stkh0mrFdR6xRiwJVE2gR3zQ5RNte/dmm7gg4LiGCn5XWH/PeP7LFZiDib7ptPpgtQ75MN
x+IYC28nDRwFeG+F/XNQYNcd5GoedKXuby9Q8YnZnGFHo1flZLFKMJlhXXNQ2TCt8fX1hNc7etdV
ddTzv924qS72bt80ybQHQZCKKNNUKyiUjQUTo5OcYGXdBWtvhFjTgdVyxPnC87U6om8CuD6wu+K4
IibQ5l+4HsFzW2+9otp1e9HUJywt6Nqam91/Cm5AKeJq8FqE6Av63azP5zr5SyGdYaiic25G1Ith
wLZyV4eYm1b6Z2EeAfdBifArimAM/oFwXi9GHklPl0O43Y/Sh7DpryjfDUVCKz+A9ADYrRbNXnym
KU1cRpqSfVuwAZJPFD1Ysg7Jjc6CnRFrZSBrvVz4Ha0GrOQ/m2EZAU/eJeM9fAXqcVVEo1Ym/uxJ
8LFssX6iUmlocgp0f5FHiZk2/blKdB+LQsQn/0Sa1XhvNLfMwna6U4RSsM3NSMtGt0tLaVKkaoRr
JB3uoAtSZDQi1e5VAxM2d0GYkapANekJzRHo5VgXLBo83Hz67LgTA4WGQrhV7CIaEJr8l02VAyMU
VsN++d4br99aGq5xxCDLD5AlF7cG/U1R7vSHni57ThD436C6MayVqU+w12SHSoG/JXCVbFVRcLeX
v1bBDS9hK3Q14Awiv0j8y8MGxGuruvqadJMWM73EWB9ATe2mv6DhiVX2dNcS9L18G603UVQlZ0U9
Uv8RAWGtP16r56iW8pWeCudsNEkaL4nN3as6naYYPWNWfhcLCFvHlwBQ15nkuHKXY+bV/K2nh3xf
bO13T7QW4DbtG0hXBBVnzJj5ombksmLc/hgix/1YZXCNUMztFteAkq1srUSbJ5CfOiEHiY4AiG60
nuDixlNk8IHES7SQ0NonBTL63VF4V8HQl9qsDmV6SvYBQ8u2VgIeOFaD+gVT5dKxLvfXB39BknKB
KxOPRNYpdi71rIMTDS98N6KsP6oOyF4Numz0Q3SpmsBQ6ZXmryC19vTUp02zcbQ3ZAZTXbv2esTy
5lXFgT7VAXsb9MmjECfVb7mZNeVkZp56hWrBL0x15WuRlzQem+tCFD74rYdE2TYSLNAFkUPcvXjy
oaTz0VXx3XXmIhiO58/7E//UNFC+CTf59IHsW4MCU3yJVN/8E+oHE4fjNOLu6mny/+Us0yK2xYkn
3lkj0Dlj1DXJQGVXY6kEeLISPqIK9nWkhLst+191Pl0wYu3cE+Z+mKTzlWHEK2FYE/JPvlNqxzVv
B/T4NVVzkTujbZjYCn5Sfa1GBebYwhXpq2HPdtogXX1soVsjAVOQ5Kv3Vw97mPqezjZE5eSZSIYT
w1eGcRjUYN8h4ykkAcjq0x1kZGcm+MY2AKquS4s9nPjQPjAuM0Z4nxKEO1Q8MOVSLUko79lF3f9w
y0oPu5z7UgVavj8VIKl+PVOG31r7vWepAminKZpknTg1GrTm6RnE4SRa1U6QV9sKBaw6JN0Y3FQN
q7xW2nzpz0alZMfqpjRBWLF9/s8lNOMNGIYWKbyr9W2nf3HnSkg5JkvgcrDQMDNepUxDl58y/lCY
WkVs9J5DSCcgYopslhM6CRWju1jniqLPfS3hf0DUTJlvYriU1DUMyL76ZahG2iVl3WWx3J06i6w1
n1RPYg4i2ioCUvcMyGmxsL4oIEix/KeVIHP1/W0i0wJfzVd+1LuINnvEfL8rYO8iqxe9Ys0+G6Uc
YnZZjS3Q21xi4WfPTMF5451C6TtB7NolF6EI1kFWDyjxcOxOaW5ao3754d6APXPFz5RyCH5XgGgs
TqEjKRMisnOMLpPqdev2TMjftzknfVRP5qDCam46KFEiR3epkaIVbhmOPtZIfw/hX1/c1VLiVhry
SL1eX18JKxgH7IOlz0jFsIQWVF+yi/KLfrBIhx42fGHcKtVYiXCcirGZ+0c84LZnKizOIA89Mo4a
MGm0JpP/iKe1mkcDKDMLDJHoDFIe1LIMER+LjRTxDXA7wvSLB4gxvGok7RnbUdeKefNOIoXyB2Hl
ePDElq0gbLCZuPEFUL/4NK7ZjnI7M8lZfrct3LA7/IW/obW9S1iY1Y0OB8t5QT7sq7qVX58+BKTv
wCax0e7J/b0v68i1jzT0ABUEiyZTzXfLBXLRP5B4Xk0KfiDXH1F4AuXwaQQt0VvNsIWDOF9oet8O
1/3XCaMVpjgh5xPN2B+xCu8YkW8oUE8T80C7m9sXJmpvguDwJM2VbfFadX5pTrHGLpHxD6kQF7GO
f3Wp3lQGcchetk8DMVO7u+kG0GdcCBCd7I+X4s+g+14GL1ojgA+txbRFrf6t8Dy8tT0RbUmJSLsd
tmkEdw2veV72QRHgIdohXaP3Q/FhY28gtcvkTZjUx+B3J08YyjE35P9hzX1pSKkU24cvz2goRWW7
D2bneOpKJSbC2MTbFBBgrcB1RtAAagwUDKndK3DueK3xMX8abR2U3uJ2P/HWN4HH1zc9rktEs+GL
hC4dq2GY/QOAIS+rivcA0008fuex6xi1WMpoM+ZXtIIpJfvUTOeNmN4DFCpgeuEz+SKssDsobGQh
nV8BKU8rqNUjIUh9exrs162MxMmbK6OC4RIH1ovI0xnsInYtjjMmyIFnnPk2oyTOaKXwRUbY/5RV
vIX3bV6qESz7V5ifSy0nVY2kKRKFT7Dne5ItdWW9Z3IYRhjDtNYEypkVh9ciKl6hqKgqJ/KlRwiM
VukvnPdaiCMLmVw7Fzn6MzbuA4wMijZQZZZ4af1misrwQl7+B83Fl5uYpPXNVlJA2kBPOuPtKlss
/qtSnjVs7ctqXepLeH0rUPqzE175wYPPamftdcJOoCwIWLzAaU53AC48CN6GLknzA1+5t2vscEDs
vT9NqemXeM8eALczdrgyd3sLkecO12y0t0ysZsLjF8LYjaE9iGg9Hq0PIWCJhnPBbYVGJEceTRoi
mHXGw/EX6XjExV1wikaGqfLOh46YyQIjRloHKSQfgmGqP/h0Tim92lZnFP8rMMGJ6WXY336inywR
6fmrZcnG3nvaFFrjnrg8i701h3V0BKi99J3Xbh6B6tlMBQJBgxQFXnYB0BWekGnmx2keNsJkbvHF
KbtgE+5AQhAGUhlVx9pZZ+NcwYR6LQ7TneZpBs6FJIGJroa/93fOXt7b10UTDWlEKjkPwTLNVarG
nFT3p9i4Yp9lADaRUHZE77sABTvgcOM6SMV1AI6+ipPOd66ey+bv9Q5qBOAf5v+no/Lr08RPNJKe
aLkyNxRma0z8XgJ3Q635zOrEsUZEbaOkMBsB00kIUhbrNtuumQefW1wGP8ZTkIvsKMnCrSOhuPwm
MxPv7uJCjth3kRdv5AGwu7QrDHrjBFKs/0ux9D4Ai2wNDKkLlIBt65xAwG7t8kdhIoyUu6YLb4t4
hAQJGInKs8XaRIVSAIs6rQtYPAgT5rvJrqAlEpLoF/gc9xwWz/bMZLgM8q0FsfvQhZqVCsWbPDeL
rHFuWDKISV79RPSQbiWNzXJ9P+2zbRvbbgyMZ9WDSOCyMSgLe27ByndJCFkORh+FCAR0S/oQUHAs
Yrf9d7bTA3Z0jRyY87hwumuYs8X9b+bVy6sM7fNUmRyOQnf3rmB8nc8BJ/YAJYE8qo2cuctNWtHb
+B26x3fmd+m8YO5mY8enPX3tUc0KgFH1dENIIn0AroHm6/QPR6wkq5i7CHUqAehbsETbXqC23j92
Gz/mQbf/ON7NTT+0dWtZzBt7CYVVz4bnDWa9W2kEuttnWHc1K8+4MjWPB66G6hUomYT0ALkPHg2F
QKbdqTbnasMzd60D33Xv818RuXxNbxCzqRDIruYVtWcNDSU/EtuJY5olCn/alQAsPLx77z+A9qNL
WR4nU6ElkbjuAah9/FvAoOE3ioCneQEYStTKbLWtIagHOoixqHHlVIc/Zrvbd0cbaKLl1GCOqNXg
/XhRty230+agyVIVGJibu9ZNQAEan4r2cZLXq5rUvAFtSFB0Pxk1HAbe3pxav+zTbtL8X7gLG4X3
ZSGZ23NTfGV3yotEL2FLixu4c3raiTXjn6rRtWTRiS0PpSzJ5PNen8Q9NuYv69+M3f+HwVxua/ed
pdT0j9mVaIaX0mwmw4k4e9w3fgB1YYdWnNO/mk+CC9OPnvghRoe2+5ro5R9c7Iov75201yAHdvkY
5fWwV2N4a0duGscA/b+b8uWrBATtB09C55ngc+qQMZ0dYFsuHAx5IuAXa9WgTava65A7b+ng7hbX
SXbaUHFthgo9bDgf6XB66J6ZzHHDgB6xNcD0nfSba1FMeeAxA126WAMzVfXwGHirPs9dw27WlpwG
OjirQxPgOnq+08CC/8qqVZj03nOQO7Xd3ZofMmDLEpUG+8eRlaYeIgRS6UJQHSPJD6eLxli18Wrp
kJv38CGlSYQrmGGad5xjT5GQzjPue8ru3Q+oPR2bgR8YZ2vp/d2PWQ4UA44e9laF5ilo2BeaZUNB
wZJ9pcW9oYYmIBWTouBuaQ52je3+20oag1LcIafEWaKolvF8Uu2CjYxA7j+YvyDFyJmNFqnGpFgP
qVvpmWvkqtkMlg7rXxv0rca96gJU2oFNFckHtV4FVxX6Rs8eZ32uRfZCRf7A6+wLQ5ph0Buvt2pL
ARCKj1RjuT0p10f5748GI4miWzxgRrNDEBcLP4ug+Y/MGcL7125Gt62PjSQk4SfSDuuIWhzHJfHZ
FNBpn8KQ92PMuMW7dnEK5xz9pZm6bD0H8KSFfrNtxRFekSpHLoQTZ/5deTVa5tKhyj/v7bL3wqPT
SKTUfQrSOjGSoASW1WsYWqgT6V8dWFzv3fmBl3PY1ltPLDoy2NxFLTZRMz29J2msfnrvFRJuyaB0
irFxPscCMoPbj2tfR6b5QYJud6WPgpPN9Dc7dny/s3HMAIm4Kh2dfI/bg02RTRFNYHzhShdWZFUB
J4CIA1pZt0pPs0CNlRsV2VrMHGoaHBqHWcG2NB5A8pqlKfCYRwcXXtrtkCmOt1dEmKbgErb0OGSi
GFsokP3I3W5ZMkXHbkPGtH/ttIl0Vsj66V6rZpFt418WIwz/ZLeF72pcNaeJCP7L4RzVRlkdbDM6
PDyaZkrM5W2zaH9KoXzx8GX/g845qwnPJfPIGM/mkfO2J26SM1u6d7qH55i2/oNanvNNWULWC4jy
Eh43+ObOik8vnUsqXJlLYKyUm62W9wKfX/nYSNxbu9bdb6msUteuCZtQIjV9xoxQwixtu1mNwQq4
VlvE0hmYNpCF6lq7RK6SXTsN1a5d249Ko3zc9PFjkHms7V7JbyuCKp+vR3ZHCFV4h/4hpkSDKEgl
DlbFi+odup+c0072VwacImFCK3tkIFD9WU6lVnOJRnoiIXJ/NeHiHwhed4hsBg3i+Od8n+LgXO0X
b9RZ1m2oml0P5evK16Rx7zgr/KcNOETTAUBcbvCIWosdtcYgWsWulYDQ+NXEPb4xLba0eV48slCU
xf3FLxJJYaCZdKiMWM/9E0D6GvypgJddRDfMFlOETVPBX8iwxH49CxfAiER10jmh9bpJaSAKYkQG
8mMSoMhXeMIfV8pQ1mPCVYi4dBecbbCCsBARDVrMnwebC26aY8Pjf4ezCqhrb1mNLSWGFyJkvJFT
zf6DCb6yCycB6im6C5ujqKKOm2GUocBzDUKBXU9WNCH5pn83oIY+wBYmqtpacB8BtJWjlaGXXb3R
FEOsJ5o9G4OGgNgEG4Ylp0Pm3m/OBMcKzip0lK1MelrKSoK/M9ni4rxJ5MblhiCOyGrOu+64fuwA
FZzcGP6hpWo+2lA7fKabjGwSAACuF8ZFpyA8rWU56zD679qhAidKGa4RHJUomdcTtK0TMiEgru7W
Cck2BDOEaqtaOcyjDdNSWQvNrLQKiO1OHqE7Ol+B+rcuG4pbSucYbFdc08N3cxi3lUPZ5OdO8Por
T0BhM4zAIx6TYO53NMsqn/7IvS+9K41pVJkGl2toC2H9ujivCzQhYKnf6pPIcXxJWuurcAAC0pmp
zdQPkMyflCAFgSxwMzQ9TgsCCgrhVnXVp7Ws+heTO9nAwRLz1BVQgmwA8V9T3XGGVMSVMjX6FQ6T
I6Nlqab2ad1PwMOYDdmVXjrhZaU/2iirb7xOC0djvbZakVEmBliFBA4ZUjFTSFBGjq0jjSJlIk5r
0xQmSeP11rQbhVW4zIXBwSNFWaCmhlJik9/br46XlJuGzWyUmimD9uyfJhWA5yjp7GU/dk/r3NsJ
K9j9GJh/SaffFZ8nLPE6rRRPtd+6FFJRlNUDtnbqbh59YbKeuEYY8EGvkZbiH7NCAdNMKsTYvodP
B1CPjULd//ouZNUsagNlk36XfsrD5uBANpKQkrK704cSbieDCr3c+nHhHl6TMJ8m6gExKu1uY17y
PFyneGstcPRD0ThCVpTtuPZCJ7UPGa2PQBiDPJEcs/1QVz8Dt2HAMI0Wc7lJniIXdFU6ozz+QOqF
nqsDRdLl5aVgzLUEKtiYufDvlNhWZ5qvfig4gnnWnym1+9RSx76Jro7Fr8tozvmCcqOckmaD8O8v
L+3B0cfmgP/92+M0RAFjkx1Ks5MuN2EoSs7De85WMWhj4TC47PY1PQg83egeiLkdQGjMwkKGPSBD
OuFENTGk09Y/oDdQrJeiReH1mNf882sk5r8JPAoTd2+4ZAJZjczuQlJ6ZpHlfCXl9ZX9xcTXBiUM
vDVd4WSz2S801okWRjGdEidYp+65iIwCKbAs4UWmbswQD/u1Gx2p4VHn+Aq0fhOWQQf8Gpl2oEE0
QVnxhY2rJRe/5srG6mkLTNc4XOG/szVVw1Bhw+XTUs07KTiPYYPLvjxd3jTrA9H7TgNWk+Vc8bfU
1XWzMAg+f7W5izYQS4ckDx0U4+pHCwWahImyTTMPF2/Qwnqq6wMk3QdL3+h6rHUK1R92IAZ7vIh9
3LsVMZcSIx2AlWQtncmaWg9Q3l2eU0vZ442p/Lcn7cGpnXhlFn6yy2OVE4zMReg+ntoZVnWWh44I
QInC/6Y+uIOkefsP93vsWanihRuk5MRA+/pCvbKqRuV5fvXicDj0pQbvM0YQknRTuttfmb5xooyt
BRzbxvf0HjKzQ77tg/mYVDfEF5UwZHd1ks1L0wsEZ+CLf+AZH7m3Gvrax0k0d6mxIfds4ktJ19U1
FqUu457qmMMxfIRzyIDD8ADg/YFgK5buAWCTP22J5JBFZq/BkOdTaBt3WV1DGMp7vh1Vik5FkcDk
xw45YFaKcmFqUyg14fLeJY2ZewJcEgBStAwZp+s2w3sjBKYYnrtRgoH1I4ghfVF36PaO3rAfRP4u
xOCzKXGzhDe5AdwcvZkADzq9s8goCH2hvyItGKFq8wvyAWxvaLwd2rlDwAl/4D25V6XYFyw+yW8j
2YmSfo4Y0486LxYF6KqHI5VH9f9MdbukL9NkseLb+SnpNcIsvFIKaIZdlKmAH0uv8r+NbjjJii58
nHBj8WhlQwO3XWtdEkVXcVpwxACEl4WS/qSsLdIbjZt226x/YW4TX4ye6AD2RGBByEY4ejBeg6MY
jNIrKUZRO57IZeaTllvrwP7Fi0FbHfEzEHASaBwrNetK6ts1KDbFPg5bb63KSK2iXqOtihu5a6Bf
cKJ/uQxJPZzJNQbWzVbAHxi35aLT/yD4/u29IuxHSGjWjqVYSC+FKx933h8wiFdFx59F0JdYS0jg
suQyBc3dHBAEYvw4ncvkz4oALSLRGrETc+RFcRlNyq0oMjMnHPpxsYybM62sNdmAZ94z6zMae7V1
YFblYQxW5DX+0Ge8zsQ1PcvU8D4vM5YRb29CulpTmtYpRhvFPaoPPJBHTV6UhB7kyJDrvc8uQWWb
h7AIwIpoG8isnqWftYjiEUImBkV6qMxZU4FZZYx9Xrhgg5UCaO1luZYXrw6jtzhSA4zogjqB8iqg
wdRAimjic79G9q1ZwGugxFs1BvsCgS4uvtxl3Ft8sei6nQAyQ5wzRWl75BjoM+vLQPCp5C7gKi+j
Ee6LK5u80WyvZTKd0b13VxENOWKIv2SdVAe4ZSYP1OrLdSB0ZSUmPFnKK+xH080JgtPGtojlso9v
7NVjy9cckL7YbUsxn3LPLntBbEtDduRMSI/vlnaVIuG37SLGl/T9DNfKFNvEuU3PM2OlKH9KGYu6
e9/EqwEBe1ZF1054Fxb/cR2FozCZK95f/a4zi7Rj2sASysQ40J3QlINWAotGkIjNQQuWZYubJFoV
xThVay+16qW5OsqYJRrfrQKFzIUHJgHTYR/8brfZKhrlYar2Jq0s4rYLk4usZXlbWBSovuMJQbPC
HfGgC7j3G2sRoSsOu4tfA33kzdEfzkMQ3/9lVUKGZIxBTifKNOGQ0pM6e8Q8fuY6gVdHPFSkc1O8
vAxNw1biI1OHgJz+PBqnCLKGJax8kdDQW2eXtqUXGvokMtZzxaVPcGCAjyG7/RAWIrsVNFnyayON
PZs0ht9vRuPsyA7zmvVfdX2UfLti64ssq6yuBo636u3MOwPvEsT3YHCOfkwfW0id8+R/nZxZ6RWz
OsptxQyyPF0qig2fRA0n9S6G3osiHKJIVOIR9EG6ZiuMTrWZ/9LKU5BQIcNQtuwh5nNR2/bx+w8r
QNBVqGqi6v6M9yXoLW7M8X9wFHSIuncoP5SyerTiOmEcND3xFx1VJBF3k6Yc7eJgnLjSIoaQ//Q4
HxMc1h5gUuFSL9S5GP4ua4pxSCg+/FEEnG4wY4gQjyrjya5yRbtDsSWErOrTZaERUpBEEqBOGoNH
KYWFI/WYiar5WF4084ahYQb/VDnLr6KE9VE3ygbQYDBAiJNFOt2GbchQAwUT/VwSha6m3J+BW+iM
FarBGSpdvdIClgQTREgntgkXqpls1k0xtMNY6Nw8ZizwrxosxFUp2bYNOID0+btWSnxlpB8Q5RgP
/neMjHQcbwHnhoqFHRvXXetyX7H+PzLCQOcdVmLObNLpHWoKiK1SKRZPuMzHt1OL1MGkzjj7uLDW
eE1pUZXR9rk6oE6jUjTkn/QRYfcOyPWUejaS0rtYIMZ19ocMB87TSkRP0489qtthJVFa0bLJ4ZMV
wZSDV+I0o6twNttbeQcRx6WiSyA4P8HpxwG4FKr7lU2OTg7lLmastLDL434KU9HNoLcgLg6Gil/5
WE1LQO2RZBmDvmvMow7wW79p6bR/178apyzmwgnNMpb6ai52KSVfUYRcC2/Bk6j+OZueZfRY4aWN
lph/YOqTn6KZiOQ6XFxkLbMMthWi5OJoDJIVCbwBBW7rBxhhJfJDgyjBinXO2/vchRmu4Y28g7B3
WDfC4Az9eSajzCQi3hGoUDutBlJzmiJ66lgXfCs8iWWt1qCbTEA/AxHH3MpXk7i7YY6yIAS1axCe
LrvZvRLaAFCVSwWnXEI2HVnevxNJ86VMQ3jAx6d6f+ndp598+UsUANkORz9SXXI5MeX+aHNRGCKO
qvRUiJCDDloNkuR9tMEg2wZW1qSub8fy6qM+Nw9AMW+XHliGgJgkg0wJ1HmSvwAca4O0cSd+vKcO
P7kT7eJhjas7dU3Bc9emwPMvfHZQQFbDCsDXJe70doFKLsrYdFEqr3n00/OGX6sWDJFJ8CwVozyM
yQWkka2gP8pxuQtyH+7BzaHiMf7VsSksSejhgvvi+EJ9W9GN2iEBAnFwMDn0PU94Kkrnv7RJyB+u
MKzMcnmNBX7kBTcioEe0dh0qBhYVZUWhnt0Ur6Vk04n2gFA/JeWlaBYV0/mnqFauKabaDm/mIt9u
u5iGFRlOZy04h9BSj4+S/LsHrXjuDaVPKI8JHYbcUD/n874knvQ2H9NIGzTK7c1kgcRZ3Oc5ErOW
NZQCo7lkzFBZob0EXN6GLZpEc89PUaSKv6E8uy+TT7fg5htaaMdUzd5e1bVbGJPEe2Ozxw3R1IOz
zT8OIy+yOAo6AzSiUgk2+Tqw4UI2qvqV0jca2dzthCLAatQlp4n2XqIqV09DcNUlHv67wXfo6PXu
ogTfJCknWDhG9XsrPNgh1MvabfCbLqRomG2LIS6pRPbPE/6NaTb36ndRlX20Nr2Roby4sSpRuUKV
vHtscQFW1y909Fz/QdXAs0K0eD93/B+Qotj/2HHPm5qQwJiaPs47Urxhd2TXIlmQ6e4QjhvDJt3y
SKMlVpZFmDBzOr4XY/oDdULXPBA/neqJ7Uq5XMr23uXI39yR0oW7M6DgXvTS1MX9z8c4q/yqDFgI
+jM5fKCZggch+ID1dlhvicAk/1+JGpZ0yMgc8qZ+xR/90C5YDH8EU130f/M+98+Q3UQSU2hZq+Ub
C/yt5Vh4UjLm7M3/U+azJuaNd4wAqW7aMn52RU5V7jWAaRfJv1PFJgAnr/a543D8JWhVOG2zQicL
v27G3xjbiteFhTYDiu3sqZFf99MaEC+iCaHiQ4QsFn9pfsqYeVQE+ZYdWx9ETxIaSg3CSRJPNoyI
SeQXZ5p3KdIXGNTBWLfgvjCwim2bmh6KDKhqpXKhNXYTPXGaci5XdbpquzsO7nTx8ggE97P+DVvU
/xw5rgahsAsyv3Gr836XH1eoq9TgFuhK5y2NotYoj3ZCgwYcUytYMHwqj7j2rBozmSY++XE22R0U
VtDd26kWb9Yv+Sv0xNJ4LMamFyPv+CnL3PTqqtkaqFiEEIr2LaJYCyYj4km4nnL15aw4hmY/zK9l
CVwWWV28tXEH1jT1PcMFJD9aIG3LAl7kQIOHRhgOUofmmmE+y/IyvRg0NDxeQW1pTeGK8qghZuWv
VEaA7Y1uy1kSve6Kbmv94uc3Nknpdoi5VIfU+a9OEWxhiJffVahfOrP9KWZbT9xYCtsqSJFwqfzj
cIDwTm16r2Lvwc5QidSR0b4Ou8TaXiPki/RzFqiyUJpIX1jV9RPns2GVO33a8HcMmvwjrI2Jw1FS
XUjbcmbj7t79c1cY85jC2krXRJHnhOmzN2nAvy6831ovKs4SV587NUM5klnpKk76FZ95B/KUavGu
ixv3cnQORGT9JMbt8KEH896mJZE9iAKOcgAsvGkQN7MYoheLFO0t3h0Oq0H02fPXy3K766uc47HF
585hmLdlfIhSFKhnrtFRPOZ260uzeza17WVvgIg7GPiU9ZAwvn/7lsVpb7tBIZjXOop4DrMGZfog
M7UhjhmmaERcfibGdwRr+16jr0nBJd4q+ZdHhHXEFqAI3VcjOiZ5aRaombvTe9y49cbJ0CHhzE1q
KFA5J1xKdG8zASisqF0sD728iqw+sACW2GdcnHGNdb7Pn0vz60T1WJ5v0Wjk1Re8vv/p67Ru+nSW
HT5detGMpwRD7V1gCUqz56W87xRUcF7POrsguxxpCjooc31hod7inYk0Fg/h5WzGu0Gp/XCUQREm
QCPOlOscl0hXn6k9LvfTCke5mLCrV9Sygk5JIzr68h7ZnOlIPDvbGjgvpvPkW0ZIKCKqH/JzanQR
I7+rhEdvYFd+2+LflWt7PMick4OW1rTfrcczHONfF6Lb1x8J0FgUOeFLl5NlsPjQzyW6lZRxuCAm
Tx+lnTI+PMb+tEH83hLkQR20aBQrhBfP/WpHjnf/KWmAFGMx3qSNDGmQjIvHj2U8PvgUDGKkxJpa
81O2zzB3q1euS263XJ1vMy+y8ZIhnmuWn9CzQUal8V9md5QDEzXEHs74359hTZCExtUMYPdN2s+d
cA3gDJroIgUxjYFFfYH+bU4i2GuNEXgVQmPWb3SFTXxeh3GEcPTb5huULo8xMMRXcwporc3zV6o3
zP5VbYYMfywQiZbLAdSohZSGn1AfL3rBKn5YgoNu9oWm+9aPHflJltej/fC4aIKyJOkiNLsRTYdH
GbCiPdab+diz5zKUPoq5fa90khUtLV/resrv9ro6WudiWf/pS7lqc069VyNGx6aunqQV8d9oUOjA
TM8/EsyqGbG6CSBdM2Wq/ue40f/CZZEcdtagJku/hRHoD/XgmXbQfZAo8YYkKf7XORoAmfoL5u3E
1nLcIJ0QOWnhh99LQZjakHNC2+o8V2nz4H8rUZToEdAke9DL4nj1t63hr61kKl3Kr6mYPEnAH6xF
EVgbF/4PhlN1g2dA/2vF0lQlV1rxbB4Q/CY4uf5YaJH7CJqqKyWszOWdnZE58aApOJ2gzoITptVz
qwi72IGUHANnOtPlyiazHM3mhd2nDM9TDQV9z/dUSdCrvonEBNlHO6ZXEw53X+IBoIrgkw/XfXtm
wBg8gccCNvx+cKSnK/39LIz+KSgNQbEpVBsXBT/kHn5ihSBd1zLcznZ1KN/ERpIGryi9WRaHV738
ezspQY5tViZB1KMGzGG5e2S3TkD4biNvisCa3hMDZbAw037a6o5Lxfir3JG2ySzDpev4NX41sHjO
/IvYFfexalWLEyly4ANxsFpY+F6ElbjmXhW1G7WLF2+1UC3NZF0ULKId2nDw//UfHVz3erJN1ZTR
axAbKIE/CpC6SOSdUaAg8xgnAIHxjOKf3YQGCTR1kKFzJnZhPbVn1xNzRJ1fyvyaqzNELomZluf2
euI6kU6HI9RjGHaKi7jpiiKk49PeD30zESKq0jKuENTZxREhAN7fJncG/XHEvFyk3l6jCQwJ8eVI
YOZ3ZGmjibCwANnyxzAMxs8BPh32ukI48IjiJ+z/9+eDre8yKNeCNPKLQvnrMJ7Ll3+T+1QpupNk
07qJ8wk6BUNhVWmVB5El+d7r+sDtTIL+Xb0pWjQ6molXk2g1+/2/LmNcDDDAssGzuw2s0KLAZc/c
o2n/Ego7IV8mZbQVQH0wCRgK5h1jhH127XtWUTBgAmpmr7GXMfE/d/NSFpwgjNQ8xYMThB045B9S
eE9unIRhbjo29wVR1/ST3NBkKOTHLC8zBglwC/EMy1xfAlK08sF1T9dVawzzrmJOdm1pAveDEtE6
oASPABwARy2v1ZQRrBrmZzj+2Ot69PYBntEmQUmOazujqiuGyQJw7lmufrN19Me5vGV00LtCbb8a
cMVAB+YbAgEsy+IkEJIOka35U+ggZlAZOmXqegq9qvvSUmZeyxR8AMukTEH4pxSAilpLlJcbDpij
H36AkfYtNLPruCXS2iXpX58LTPqu5PNc7k0CNEQGEOhwNmZhUjTewBevH9EJrD3XXeGeJY6+buqf
zGZwrWX0fZr5G41u3CxNjGub09FHfgPH0gLE4jvPGlGAdw+MbQaYwR41nLm5f/Yz+MbiKZe8Wcen
WLo0eAcryW0CTZQT4S9K/PdxCtqNjcxgJumltQl7jVzO4p+Jpj1ltBDrTyoDSIfKeW677QXPi9Ch
+R96WVfodjqy8ieiaKD4tQ8aOU3GtR0+/CHo5TBDF3upsSWTEHTKFFlofh3yTqyyA6z0meA58v13
AWRGeEUxCZLmlZbg8828QgEzxiZBfsNueFr21hsOFOqTwlFXvE/dkUqy56YM8MX2+U9RMikJRZDk
emc/uGrxWIXA5prYpzJUdg39rXD/ARFh7cRRUI6PBGK8GQ7V3Da6sAe22WeI/MrYf3wrAgCBw8RL
YYrrs6vaXfYV4DOw9SNVjFyrqKAORJLyI34XiRRDuudPFv4HWVoVdqo0jfRKjIinoHo1wyw3k451
zXimKT3n2x0LAYnnMzURD96KyZjpvabwJXpiMycZXQ8WxqT54oqNtDfgHPiHmY95tCHxuzUwbQ1Y
kB+9RNfCOmTcFMBAhzW/eoaaWmL+mAlsFNTRzwCLjXhjvOyy6fRMvCry91fvrtSt2l3wJU6e+mx+
LdBwLiomMOVDKfmBcHW4ci3W6kpKgQdDilQftt4Ds5Z7U+KeJRoUWdO1xIWekBMgQVml+m7k9M/r
4l2FTZ+pm+11uIM5nLSplUVFF2ETis6O5RHw1h/OFxFljJkI7hmrXnKq4773why5Iu7oN/V/mFpG
wX6SGz+eKpB7re/8jRW8Akw9s4U0Tb1QAVVryIPzxq76lkoKxdddB0b1wsSI+pryohmRA8E/1biQ
rloKV1/cAhUyXHtlAzLgaxDyQzm6N6lSsxALgTXPtTpCcfL5gHKV+0rZg7o0lkyfjhxxF86eRO31
HEV9ZJPm07QCzeuXidazEC2rJwj3sxKbec9MqmfS23fIy0lChhTE6gRqieh0ChjcatYAb8QR9814
fS1AvyG+Y6B7EuZ1DZRfvGfWWra6gxmM56HRPGw7TsCTVPkw8LHkOLXOMqSrKdG6T+dwLPFZBoac
7uWn0EC6NBPAvVEkDVsBYGsr+cFiqOin36X7O2IpiGLI26bAjSCRN99vWzVmgyhNVP8CsxQNDTQS
uQhiCigtWu+3OTWt3wCna5yp/sfnPog6W/O5oev+HH94RHk9WJeGt++mzrA+gbeL7qy+GJCWo4ZT
XHhGjB+sDEtn0kyBpdzsI6884Zl3MTAsroI/tp5Kfkb+igxYNTl41JBsdizGCtSb5xcM7ZHX6WUy
0Q5MtaIO9//bPHvD/i9A+2KQUMZSIlYVnBLw3Lxt2Gixr0CxkkvFTcQ0Nw93ryenC6lVUOoaQM5d
yQ8k0kUORg0Rej9tBnFc4H14CaSnTaDeFXlhgpDF+Y5NNYU06xSXWcwmU/zlpKJ4DlhV25GiWoE8
swDYefUcrLwVLLoH62xVAJrKG4qxJij0+3HfZyWgzBkgtxQTw2sKDqYRkmzV1YeDtolvlB/H3fwu
1pfEjacZC6imROiREB0g7/6uXkY/n7nlRIV4cbW/WbIj7WY3/8wBPbGHjcdiesEZqiilvRZVByOG
rBpx4OdZ1bjkoVFaXoBb/vu7oWJWmC7CnarmwyewRaA7My1oY+S2qBFBUtlPDmDlOczi4N/HhZxE
OlmHD2J8stx1RCYpZcWH2XPu8whg13HuK45ftwN8SsnWQV8H5e0Et+MgiViDR0nMdycLlDfsXokT
W2CMLyFBTJ1iNbsBvFhopAo3aRn4ojJShQ082193PHWgwzB+iULdyRCkRVHZbtFEZSHAR5ZIX1FX
c974rhNlW+cfYzGI5gtCzEt+XJdZHLpAuxPr6Z27sj/E/YmKuBFlxIhKHiVyoLgPxzdwVvEfQNQy
DHj+9SZqEMyrMYoa52G+AuH0zle3j+VLbkN7w7+leDuMyr2fZATvpRON09S4F8TBmMJVsZNavIor
CGx+h2YfJ1meI283V15URaLkOfneW04Zqc+v8G2AtstdM1Rokq1v2yBccuiRpxOn5cJ+pGHzJevV
rUJ7MGZK/I7JuTo8JY/076NqkORv72e1hIa2v2j1ITjxTyTvLPcOnm8q5EfIiZ4McGqdfrIFhu+3
rY97rriOTUJeStV0Ly3YpsHjPE3Y3HD1yvAFT/fLTHBiNenMITjh2P1w/HjLYOsZhhU4B9rnBHQi
vfNIVDZJp/BV1SssKw4wy4gpNEL919SkirBsb+y7PCVPC7Zxrh7WdJi+emFSC8U4CV+yrhrMSKih
JY4tR/ZEXf0Lq5JFAO8eCc1A0E5z8W+6FExdy0EyMdkmegmG1weEPFXqOe4ZjQTZjtX07gclIwiF
KOyq8IaTMLPy79ogObt39Evk1W98ovTa0R+zm5fhXT/KXRqABev/CtaIX+rVEcqFiio/0HST/4E4
I1jUfgWdpFyUaLQahUMIWbuSlUrXj0dRVZwwkqKonQ+Gwmu6lz8im87Lm3MRfl4+zIYmYjrg/6vS
NEptDzVfsNmD9X9sRqB5FDys1qAV3wKoCO7Ys7Im/5CrR1sNB7mtS9YAtuQUkDJ643StSDAM7x45
NQB0Bynji2PI/6Qwc4HrDKiiFE0QAzUWlmMNwkXOUsGcOjkOY78CdKHwDN7sP4Hiw2BkkWuVEakx
sLXxxVoW9qu+1H8Ftafoj71d8Lnn1l0vh7lrCgdGVj4s2tUJLUkDKEmChdpigDgIvStIzvU76QlO
11ePh51+YPNTnqKoqSEKclVh7Q194LxekT8XosZtAGzLouBfJjN5oNYjUb15uL6fRgQpWYffPaix
HFv/IN6BJqqv9xfbA0oAaPrFMPSfzQSUIlErhw6iAfES7Mk+18tUVQhvKZPNmmDHjhIF3oXxd5Qa
mRnOK+0hqjdhxggAqM8FpTfAVRmqTEQALdWSifPjbMXg5IRBTSBozxsKAy4de96Ch8pC/8dTQLsn
8Re3+aXdE1jZIV/7qZFrUY7TVuRB3K9ytbpHvxLnIVXIVRcIl/2Q525AvNXMtpQ35/IDSbXN14Xk
RrhhpbNCzcTrPxLGYDEFXEKemXrFURpfaZRQ+/r1vgZRoAKow8i/nSSDmQl/wNCLWPEvrsfvPnXU
VgE8lvcZf2jj4FiX0YxPA30M1CjCpIR/Im/vCYEGTbNMIxvmxm04cE6HAg03IKKElZJWxQMFUThN
0bL1u8ayb/GHnsYrXGvpOhaoAv95uQzUiIa9QFwQsUZzxEnKMCqKy1oBKP/9OKLsE1FXUVzzV1J7
J9XkMldk7ahR3pPN+wO07W1W95Iq84pm71GNyYLS/e6E8jXF5H9Kfcgoi29Vd1P+aB3FqrvnXwf7
Vec7+rbpL3idosdFzuE3m70iD7RCtZ2iz1BvKSAwA1EKD06QnDAeMnko4R/MhpVe8o7i2nGQ7d7A
sVtyOvnx0vKMBSowoXlqg5CebmbWiO7Tnkt8EsXoUkIy3/y/mCOUlfYlycFw6kbDdPqr5KUVclyg
t055vZVg87W0leFISn20Dk5X/SXbZEIM5EvYeVhshOVWLc7L0IcFU4Y2qLjXRNTgfM3f7PSYFwhe
8x+ATzjF0musY6/s52CapsLx508escXzSbslIEFge8oGrt1fJoVSRRBEieaSyL9QFuY3wNekIv7v
BBHU8P2qhpuubVbrgqj3Z54mPOpDDhaR3T3D/3WuUvVgeFJWGHlNmFJau9jnT888sTvKiUPKoDGt
YjconvkyW6PGZ9yQdfBTFLqH9kOxNDfnT9WThXVuMQtoT19vucU/caEHRnNRWCuzDy5EFdhI8Zoo
d9hD9WikqK6Z+OyfngxByxAS98s5YOG6Sn1Pm+bmFgNBI88zrOlbscykmlKZQnkxnbyh3uWpx2NO
LRxQXvKiyBYOxGxp5tRHA1UmdXMU2cy7EV5UOnjufRGjk/5WIJs/TFNVOI+jbAajZLXxucRWYzrL
AWdnUAXEi4SaFOWf3JFlK3M51qoaCyDscFk7b/ut0CzcI2Hg77k15jlnoBmm/kGjef1a2SjX1UP2
cdcA94/nS+9P1KuN+/cX1ZJdmzNjUKsjIYZOCRIiaWGIjr0nPDleyb9vYq0uvLIvcLdbmFM0twB0
knzhm8gIWDvrXZdPVKGW4Jcfw2z0g3dohCdKllRYPhXPkc4tk3rznqJoYVDZ2s/nVs+NEtDUoyG4
cPyWhbXOm3FdTSb+APxao5Ku4cxw+y7iWDqwpfY8c7QBZ1P0mkCqD6+WBh6E7BewhZ9pJ43mPReu
6W8gijmq5cQ0fSAqQTj/SxQVJDe54TRW0an/hA9EAVG/MMh5PImxmOK3umbevRmURzHJrRBpdZ6O
evvLaXvpzcbkvGdBHOXTZquKNtUael22RNwcN6pECY42Jg7TW+fNxy3+0ViTSybdyafBhrH6zdzr
nXdZjeEWc8SLzbm0t6lcme3SozLw3JIFNlFiYf5cITm/mNOjs/ZKeKnQ2ZMAG3ZXXSsmjBwS7ql8
cGI9Os4d3bv9S4xZhfXUz6/ioSCW0dN6qrGShUFzeIZmIrAWE/sl7qn2BcEdS/LecLpBOoqUkfx7
0K02W+w4ZwZUAf/OyyOhOT6a1UwMiVYaKi1bYScai3hdOgYnIIZeJkdp3pHZqyeno6S6EjH4h37y
YtAAb9BfOxeeACY31NE8Ep9PLwjtTbDYadj1cE793oegjYbdyhmtZXTzN+E9BY/4t2Z/1Se0t82G
eaADcnGkMU12wHFW3DMes/fL/n0bZlc50owkMGbgi090mdExlFcMuVxUFHbASjh/aPWuM7uNYAvy
0TuBAlYpR3Z+bEpRhq4XLXE8fQNMuCmR8E+b5Fd6z2S2d4GEdhj9/mSbOd0hg5mJ+WEvDp86gtE0
mrWAj1dq+L9tyXVri7PR7peY8nKQ63s/tuJzb6Ai/352B+MhnGda7F3VTwuOg64bZ1gFbqxFRFrt
jrc+msMQEmWkRPbykr1/aO29bbXNFwRtFdrEIm9Gb9+FDTb1lKvl3SLnwwtnRTd1X6w8o2uSZoxs
n4GSGY4quMYutqDNeI3dFIwtBT5R2948QlUcCPXnmomhxH2lbQbYVJTlk+nDF+CGc/6FvBtbfEkH
OiY+/DQP7l7jGTYKO1UqmI7HGYOxiFihTGeP8+5Xu+GVucMauL0b3Q1FC4HmS/Jm1U/eTs+EVGrU
rVKZThpD6tGgZx2+SMbx6BgQWrszb7RNckGOg7ezESi+DEvPcW0fE2AhGdL4kmaButMI9KF+bEZX
spmC7BpuQvhY+7ENHdGINPmmh5F2UZ14w8MNdKvLYpATC9BLpkFRI+XqmM0S6NIzTQq5HjDLLaW5
rXkF8HZkOQxft1dwzuag6sr7PRhOdhriZFtqIFRS8rcBtNDsKkrArliRZ0ExF8LR608UqGVcfK58
DWGYYFbdPaDN7CW/FI2a6UnFkM1ad6fcQCV8VkJiWh+t0H1QfPwyGPJHMMXNdqPvYQrZc2HXIMUK
PuXwkhPHvBMxwA65z6SqzElDE05OrG1+60ARpUrFLlxZlTh4x44+ZF/MyFiW1CXYfcY8pmIxFPOZ
4xyK1tT6rUitmnpfowNP6aabAf8P48e6xhHmwoACPcgW4m+VZGS/u8/C01PkN8Wgm7z13QAMetpE
q3MGssXbiJoDZA2ljZoCWZDVhQ1DwjHd3H+v9vZz2XJKfHHMAcarYmVlkykvWJQfdIgb30g8vuVq
onskjihc97yMEga4se20z3lLpzKzNpShNRwY8r28iz2w0P3VR9V8PbmSi48A5/ygw9k0/LXpuKsQ
3XlU/narbFi1CAxqp2qOjL3IfbKAz5HA/lnkfaz4QsK/EFPgvD1cstn+bm3wioo/TUvIL+m98LIs
fL8PlXsWlTT0hYVDb3x0mfdBL3GuimEVpKPDtN9G5V4Tb4LwRn5loP1scuAIqMEJ6+IN/rNuz4X8
ajjl6uaoYyo5CIMFxoV+00Lxa/aPHeTLP5SWA1qm54ZUcg2o00N33yG2WWb9JhoKuxd8F6fpIW3K
ryp6Y1yTgIhkQWIilfoU/Ta7akO0TZgClVLUjfJi1W4pcQfoBsrFpWRzXNIqmaIjyDtRSDfLGwGL
iNbrVHgCqf5pYGhMjLvHVnIWwMItPQquphz9SJxvgBNpqUUR7SVPFoqKp29JowYoPAclG/564CZX
Q8yAL65ELXUGxvvSLqb3bWdWrn800qIXNJu6GMCBLHDNXdjaxKDZKE0d81F0XBDV3fBQLa2ZNkXP
ZmiSva01Qpecw+85JsCnUKBcW6OZjgO+Zkn9Mdu+nX1NAD9w8qq5KtG4ThgZnHuvyiI4PrWm8Fe4
NpLFV/kPueNKKsIJMp39yGYQZ+p94RDvrpOwSxHi8FbRY7wWq4Cbp7/Xt8W5srNJXZiMnmupEXz3
U3A0iX69FMehqD873TWEcB8sYFIDZuXABTq+2tv/uOYHEJ/BCgbS9+Xhh+gL5bAuht+sQxL0RyMX
/RNSiRfEnswbBh9YbH3qLE0BwLwDor5Gd7VRmF9kGJvljq5P0bMcYT11XFILtwumsczCF4G84mk5
Uzelu9yT8xBrtq2txhkoIEf6dO1KuxOY8P8Q/AZL0wXJsFUO4hVe4C4kTblnwOEsLV3crLnEWD56
/WVSSmaoinnbMAG7B7jg0sOAkn0nffU+XpXvjLnx+3O77MKeUaOK6rO09pB8p7BUIlwFlIIXrCxk
67ctSpKHWMSimtj85Hvc8azmixlRuq8yhdzjxvz563fTc15bj6nG7WedoO97TZj1YTY7T/neCZEv
NH1n5NDC3Sj05fE2RiAukH8l+zX8iL3w1hoFwfo/XP8kd5wAskqqiDZas5Ec3tKSaq3knAoBMS9/
nk/FRrudt1srtTupH79KJWWRhdP60Zw7Jxdjsv+/Pfwm1tR1NbQ1wmV/8ugGC7zYhf8lVq19KLlg
LF2SKv2dtNPmmUG0IG52bguq3sk6zCyvqDpdLnONpOumK5qlmIZxEQcyqhdxlwt42O0N5TipEDAV
kdSJPHS7Zti59BiOM0vP7G8UfjlPpBu/mHseYSCiaeaegPNNeF2VubX7cn6HQKjfQApJX3ms6pSt
iUeHLtobacYdfdFUdotuxXVM0d/kZKbA6UtBAvR91knAK2fyNdwbb4TKNXvcTX7YpKIkRvBoegjy
2h2r4N3bPrUeRVXqddf4/apg2EVzWezc23p/Upmy1fVIaexSdL4EHn3XNPnlIpXKl1Ph57ih1p5Z
/QrnT/WbmIuXca3e94Wf0bUklPpJWpw2QEJDQmaJEeBtjEWKv+wNbup7TluzGoH1b2G5Gs+16SqT
kfDGfExd53Mu7okKMPindFHrUrI5P0qPwZXjR+R1DLHxLJkiNOj1VTJDtkBjln9QGnzfgZvJMwcU
JpNyz5M83dFJO1QA4Iyt3Tn/CNtEfcPxgG5IXjRjCShooEvG3hEylPFmldJtH1RU+BilRoSSYM2V
tZCtnQbtf94/hSHtbvycqUnN/bYa1DXl17h6REUbQaXW8S90+5ZXsj/cs2mDSHB9UIVyjvtZLFgd
xW7wA3t0UcjobirijG9JHCjRgrfHSRd1v3J6ymP3Jt0j/FkSUbmVmUHn/jfWDbX4NFpW8nBaW0zL
SSzcCahH8K/9bAbhq4yFfOtXTEsco70WR3JV9YweBNQ+BEAPArkZASXyCaDfayUKymMOEzPCYyXx
8/YlMDwPc6cKcwtBYy072E7KYVbRFcYHQ0S5Z8qlKN4auSvA1C75HAAbYgFoccTRVgKPBO8pfEoN
vuffSVfrrMKzeqRnx6CWR6FpCoo/zQe5chqfvJe2gHgPRGqaGyJFzNhpqsxu6JLE+KSo2dTNj9HD
qCxufbFrp13BEFV1egRS6A64Z7ume7WwcjT7oyyVAl2hnYitykrX57rMqFGTwhND27/fpUul8FyU
ziB8QoDa0WsikW1l0eqgfCn95qqzgyoJMYyp82AzF4PzwWM9d9kfsIdGuAHXYgqUAJ50OOfzOR3s
gGqXZmRgsAmEm6mwLFz1S6y9zWEISsP3qOjNQg9pqiv6vfQrzhfFpvBrpemWnH4hES/vQpYhrsYe
FN3gcy4xv16FOdi21pbMJWsYZxQ4UH4/S5RXqw1UVhV8x/oVZtaLQHpdkTlQ5yIKLE5DRDLqhM+R
ZH3sd/TCzkuYL2psiVlkk+ZbXewPfbTETHSzQohcHHZhrf7qnxbX4aC2QuaOptCpBP7WKNqk6XIg
dKQ6nSVVxWo1EWejkh3bTRxIMylZHQR10LGNloDeIL5MvvpP4/AtRsxRmXO+a6oDoqS+8C8X6qs/
pP2TaIq6y/ZGPL3oOdYNc0sEKSUIXA4t4UrPvF637OgruAqetVDpt6pA8BtsliN6m1mBcLPx3Szp
m+Xzw6VqcSR7RzChvpgARt3Q7II/lHcVYjVJ2fjGfqhcL2NauUlK3KN+dZ9lNJKwArzSW76kDhIy
vZx9y1vIdeTctE92mnn4YviMxDnWDX+2muWy2y0U+DPhHNc1rdzx7PbtOz/b7m5/TWG5gbIax8r5
NFPHvSG9NiuETRF/1C098Jr8v9j7MxMPF2V/x3sabVLsZiGqOc2+Jm7vFhetmQzkteTGiNY30oGT
phkxaeHn1VCgkA8vIPitPV6YWCmAF2cBtT0fRYP1eEYSBwaqqoJEq57LcYuZiKjk9NvnABxggC/5
6USiu15/m1GGvT3WTSk3wysXp1f6XAgybr6QTT3POQ0qoJaJVrCYFs849xamlSZKJ63ZezMqFFwD
nXkqA5V9P8hTScLwOMj2voqQl5N1cZRFi3Rr4sAkOuHQxGOnGaHEG8VEiSUeuEsnUtPDlUo2Zu68
35dfpYjXk6u9uTxHvzgFD9nmUTnNCtpScCkPckvt2tEu3iragljPugeCETlrNTkwN3KXvPfhACJx
qzq9L5Mr6ZIhkyn7mfYQm719640/u4RUKLrrTVTSQEdlv7HfvzTmsnohgOEqyvDlmALFusQ7iMDe
+E8aHkvWqaYziK+tkDao+QCwKfRu6GJ5WgItIKbv5W3SNhlRdXE5Ux63bp9xhj+PS//MLkx1X0i1
EdCWDY3DQs6MVTEZjrwV8SKyGN/FyaFLOYB23NqpYiqGrMPMySMuG5xaZSLPRUBDMmtxcFJfoSv/
uaOOWEiZt+ArtKrRS2QD0x8m2UVE5pH3bxO8BcZx/Oo8PaOonI+2VvGikStB/7RFE39LmC+n+LPx
GNUXkV7k56xEOQ0SMiTUyLozbuaV5ExNiBpmE2A9ZpKywas9H7QuU6dx0VdBN7UuzTDAoBdyZwmG
XVnTWH9zb+5HgOM2lJg3M7oCqnmi+91RgrZyuKxw+EG7w8DHN/jxIj4CiCOuDLZkAhB2VY7ZApp7
XMZKdxw15wuemA6HXBcw9z+/l0ob3dNcg8wdK6zqJAY3GjzCA+aOX7PtHXEQVelGt3VDE9PFURAo
4y3Psj78rDcdp2A1RGbKnEBOokPEG1KDzQcEacVL3HqsCQgfeSuWZgzoVkVTbmr4xfI9iLYdJGpj
QeA8qvx4IrFoPn9XWsfIqfPMMPy371HxSPO7KiI5F2XNOK1LTp5mBwUbHo5S8lBozEFZF+3W5Z0P
yHF794oJOTQ9iv1WmXmTQOcQ7IFhn5ICZfJ7LSbwHdhu39T1duPsxAgXV7G3y9uWznS7F4VpAkmg
ssQjqvMkN5bAVFKsJYeDIx3JurAdLCr495FmwPYueZY5ARhAgnVmjCSIv8PCTQCRatFyTf231VBz
5PvAjS8vo6rW8Ra7h6W9ZPuTRq5lbLxxJJSbi1EG3jjoYAgRpQ5sNAn8RGQMKswpLlG6EkThMHBW
5tx8XbUPrTUHRP9vMZyFNgKYj0qM8Vr3FuKAEP/wmY1VgXEbI2AX7BPZukhnjdL97o5CEfu08e8E
//j0Tc9QrNrB5LivUm2nVZv6AHjks9k0r0obddxrrHaBC6iwq88K3n2cEoAWv4OQowalb+YdCDuV
c8/ZZy8zXoBUzabzwu83K71ilE1aPk6tGu76HsqvZeE7j6fnN69YmkPALYvsQsgcAF/SmMwEca42
6Swqepz0V8oZUf8pGTXLem7DJ/d9bt14Ibmxi2k/DBHpEZ4KOGvE8C1FCpAoMEAIE99g6VHvC/1u
ODfgtjmcmKnGgSIctXbOgYwbY+4gD9TfjguT0DNt8hG+NEcj7FAgUxS2bLMzCXEMm8yTJg/XRvbc
JXUX7+JHVYAaMnI+zbbkXOj48cz1j1TtpsTV159yzQxDg8J2biO4+OU0gMD6NbvRcwHinOnfik1w
KhPOG8UCjya7vkQoZZOvkIM7K8oVPm3xv9UutJO1w5Ad9dMcCjMlSFhWqahfc8RpoDXCqViaqSMT
g7Dlsm7DpO4/jYz4/v9R9w/ko+AaUD+H5HQP7hyrrfR+6m8uKFJktwapH3T+9ARS059OqkEa7+qi
TdP1oguJMyM/lf3vCX5sdEuJ7V9JgG43t7UH9dxnptMR4HEFub185CxZW2O2AVmoXYSE3kBiqFo0
yH/mV6KIyDUDxbs7xXwFs65Sch1QS/87ODu92/kLiVp4Wps7gWmb5swrY0gTvdvqxlNAs5UCWCWS
q5L3AvCrMlT0I1f/QGqmuznRqt5PRhXvAyzMzGgKQc0DJzdh23bk9bax7D/TcBwg7XPQK05ipoiA
udIdTAqug/wouyxZzK1IYnKbt8IUWpShZDz5YZygKS2MMi1wW3b3yPZ21Z9Z8vm1g/Y/nchf+y+F
UpRE3qLZJ86vXmO35vm1OjdAmvCGPTNiZ1mSgkKb0yiVNEgpCOvsrAmEy16coIDL/ytYLXdyaR1N
sQzzzEP7/Cuuhr8Bs8POz8qqQ+rj9cXLo/a9Mfjme5igb1r49PStkWO9o3DN99Bn1vX2vdW/3Uqa
75zqEYG+k1ZIDNnQlZQxQXIlBzK1Vp7TtBJrc0vKSnr96CFWQ99dyKjWtwyFLnFu5Y+WwfUGl3n2
pEsz4m+hBU9jM0b0x5sCVxPqbbzut+sa/dYUM5USq7PS53q3IU3D6xnnS2bcX+H5bjtBYUQNhvmP
BIydQFrICF0lyF8SB/JS9JHaoiBCccdhnbd0ScxyXqsN6Rt/XF7tnfElGmOpcWqbTysbTaSGERqZ
ZP7ZB/4s9a89oMmzgGDQL5c0O52braffMvTVaIiCTKLjAYnJ8HsWCbeLUj/bkVRMF3R/bxIEi5cw
cgYCfjqls7aoM0NguTIeG3VIUlQeOMWmip9iZ3cJKovY0v1zxjGeDZWpoGtUKo+rNBaEW9GqJgZ4
+1CuiNtc/Te8JfuDsv7OOYCtHeQ5lvk9ZnBu7f+U1zbYLUOK/6kLueHVlnNXW+u5TeBGrxFF1RZ7
MUJc58lqn3zOChbBaCPRljdUMo5cjNq6OAofQFH/IkwFCdwhzTBJQ7ENIUg/6Mhp5j3Fjh/tJh6G
fR4hXEzY4mcSsCcXncMp782BuN0iXWOVAHIN6xIsGOGlhoE/ewwOPFPE+frCl5bBj5WqKZJl598V
e4QIRsYsumpRPYwPVPe8wLkRszpTfPsFi32XtpVE/rUBDDp36Um6AO/z/fn1Xp05l77EPLGfuWUh
e0sfTHkCKDHLqVyFxJfMxi7PlpBZp622LGkEzZX/9uYssueqmCNWTvU7DN+ctIv1B1Ia+8QS3EoY
mNSRNO/2xX8gtZcSCox7D1CIDSw1f2hciQmBoXG48IE799IgSP9bHHOK6FMN9g3tMwU1i5r5OgPj
YyUWAyd3HbLw3utEGEdmBt6CUX4JrfUSfLxF/Pw/LAO5I6fw7xnrDw5BHESKhtPS44OJbUd9JSk2
6+LqHg7XEzjd9wXz+Yodr5XNtv64nFwLmZMHf1ussUilBu4TVjM3EyNbJS+l3jmklw1uhtT26/cQ
I2LC+8M8a8fY0TAgQXsQSUYP0dtmio0APCWLWxHCcaFKfMA8T+nIl7rUs9GvSgcbges+8NZ2IQdr
XY5ZjZO5X5zZSF3QBvRELiPejoa4RsNgLEoEa6J6rR6YtPMy1YH8CL0PZ9akdNEFejZVy3fZjjL1
zcgnxpMTNnd//JQPjm61LU67Pm1nD9uV2LK+6tBO/yyJ1zVYoNH+gU5vW4hJQKdMa4Ye366D5oIz
vmi7R6okFdIlevl3K4aw9WX8TIQFrB0xDsOFWgCbcacfAPeMCKGtEwqEFIy5Svryb/585EyEK4ys
2tfmn1SKMLLEeaq+4ROCRLGiB+ck6SBch99yiDpKq3eBKn4cpYpXw27IRZKVuMrCOuMX5tkDHxKq
y+Cx1uFqdm8BdVSEuwp0+oHqSabNTsfumnWjxalguC8xx1SXxrRZF4e8zpUss4NFI0OFZwnsclRN
t3j1aNc4RXac8JhKuj9HXaz9KD4QM2hfDGoe4NOXVNm8axaS/afBFEVu4cjYXFlSY5WxLs78uj2u
L+/WTf/M2ImPPB1/1jSrvlCB3JrPHFl+j97IUDHQxp+QySoEnElQkULO0WGUEHIhBIH32txYXlq1
GIiwkjcWMDCPJJCj4jyLmAFmLxEmkde/nS1hlFdR8UR+SyqwgHgjBG0Zczfp4eWc1r1iqoZ37Gja
7u6e0qMOEv/jWZxffn8u25I+BDr8GU0AvoFSVfOWiYSFRd+s49tZnh8Fr+p8Pts6hl1pVVEoCQka
OHjD06sS9455dS1vWC667Rs1McTIdEbMZdkboBd6qv9e3JsYidYg+tRRkQeteQqcdi/tKTmu/k8T
25O9qhhEwyVU5N2Qq+DxfwNUD7toyZiKSe9oKlUr5FaHAyhbGRHqzfmqcRUb3kV7608FegM0N7a0
BHVV7HGLSMyYP4cFo+syQwf2XRXJ0i/sbWb0S4vVl7EjDNtwsJKD6/CZ6uCoD65ups/s0Pw5mFo3
vtcSwcigJqfSQi79bGo4KFaYR1zyPilwNQl+SXfxqS0jHcmUhk3dDmAMDOv9k7AdllmFUcHH0cQb
ZODgbUeAfcEtLm9tlRjdHengGbSUNARDod06FZAWkY7JY996gGImMulM6yHwDjDLQPPSwZ3NrEEX
4dEs0mHygm3kv1Tdans4wF5KjjNnltuy/J+uL3LYkhodWtmWL8ewRFXnT4BuK0NShnVPSVPbqbRB
hw+7fOCOYO8bq4KD7puIzHLqkaiY8JgIdpw91+4aspIVUIzFLPJG5pfvYN6AYqrBrkCCxxsN3dsu
BEjAfK9VZ/ki1nDb0soKiMcIZ2ajy7v+1g7d1wgFm596bFtN6VFQxkBgmMvAj2wUtiwNVoriZLg6
S/U95SNegVFdxETNMB0reDlqJnK/oqrmVMsaw7hpGhMRj/G9iugcBuGS4xRdTJufuqwnsaB+Cr4w
rypXrW0QNCkKTveaSxwmov86H5Xlp/gxjoVAtDMaIJk4+0Cr5d2C0aUzcPXF0dZ42qAuGwAVadX/
qNihLuVA8UkVFUBAMvsFrAFfpnWojl7Y2djC1qLP9+vcMDYpGz0iO4spYW9jnwefFR53lVHmunh4
jpMEVmvfU4EU/RLvlgHYai6gSXFEYbHCvQ9ZS44bTLgfz8uA1FAZAgVnd8x3fjNMq3Gy26A3C+DO
ncJbDNQZr09x7eAQbA+N/raJ1SVCHg52iZxKV1a7kG228D4jpDx1e7VI2sIIP8K6KenMfB6b44nN
uQ2bScBG0gEbkzoNXNPqTg9ef/muBWbNylxI8TINBMaEDsTlEVwF7oamSz87+2liB5fMGUBZpUlu
RCsJ2rv/HBuJloGBn9Yvm+XrTBYHwUkUe9cyLgKPkOZ6+O2Ht9+JD3k5n778zPuYBEiFpTk4J02R
4rH8mPbT3tImPFG7GCLNmeat3BSyL9Qw5r/QFGaOpn7yt5rHDBz1zsLbIxKyoJOO1M86jyirLCzH
McC9l5KVTwQcXfjp7zkpt7AkofwLWXFHAr8CvBzO08iuzbLKag54XtQjJT2YHnNL3qYI1Y/zJliH
B7BdXRUKpvLyboXKokV4RmMU/wPY8938MckyZiE2+B+XIo2d116QJewYQYIFsLrrEl6v0Jgl4U/N
R5vqak6TveuIdCZ0mwFvKcjKGRxtqz6q6HbQg1gQHqRgSg/bTnHkq5pDgx/cs4q0hT5f9m7oK7T6
ykF+KV6a9jqUP9QK3Po5F6io9eHevPnea+Ukp5e8ERROfFoYJsH+/eqGyo5QVaDh/NcZCyVmMsGf
4RALJPeqqATUjtL7KW+uj9b6vOtv4BpDv7sZ1wtpSu2v5CPWuBRrQtK88EYGiB4CB4kyx1qznLEo
pFbLedptlpCog3oiJw8H3fWizd1kvwurwz+nOz/AYRPZZ60dtp/SVCsCQIjJYOMT1PI5Srl2Zz4D
+oqs+NmeXmD4QPj5by52fKUEuiQhoD2kDi+JKWtkOHvhtCKT+O/gPcDtcFgsuZ7XJr59aA65+Hqp
G3paf5bM6MFWhiKQS9lu3c3mxJTKIkDhvYKNE+vj1jB9T8jlbRtxjXUOWaHpehM/Vy4Du8Ct+E8T
str8NWaUM2gDq6uxzSRuJHK2iFgDxGndcM9fnEWv4QHHC6RBgv188BBKYCFmGWxiMRNfQN9grioX
vCEWZb3M1sI0PVj1w+61N55s18ZeeRTHUXHrYq2h8R51jiM9dlQ7saCTQ+AY6IHAKE8EPgb8EIn6
ZTk/07hgiqCk9F0kGvLpFDG5lEDo1RZ9qVXJign0E1kJ3SQSubpNIdReBq/engw61Gk6k+LWjKAJ
lZOdfH3Gupc1bZdsL7m7H6Q4XJLRBbWYeHhImvtSUjkKShx6PmFDDrQiQsuxL33jDpLGUnFyANwt
LNjLRZHb81evJT9ia6CsAQMBXw5n+FfroNn451tq0bVbiw3zyoF/QIkPEIP9XcJr96VkeegI25Hj
6MQ4cfEScjdlI7bBHnoscJd4jqSUWCfyHuI2g/9pFwXZf3rWqYj9HXGWzXl3dSRnlf9vEggOaoz8
CyajuduL0XUMW5u91Oqh87CqHWC6rgQXT2YWNQPu54vb57X0zuSYiji5ymF5wuu1WqYcuAsYZFUs
aU/Ck4sLxt5psZKznXX2BArtHh/YXYBtripsfZF3bC0wWt22o6BmiZeBV/Tz4eBfEShlK/SSyVS7
Jji1eIgYpPtkVh7sBQEFaJ9C3kOzSevnGI85lZQ/t5sTRrMUlLdg1/tfRyD6kmREyhbVDpivpVwN
t3y5Ou+ZpDNNq2tUMdwGYI0dD7EsMQHpvY8Jz1j9x56ICwM46htA/MZDhr49I5e6vZvjFYLNP/yi
/vpUpUdjzkCqROHIuvKlXbUExmnpudVfe9LEoOcisE3R3zWQeH10e99B/xVPc6ApPA65NAfepaRu
tmU4AFhtmUvm91R0PPDywFx6HxDxLcNc0tNW5F72g5xrWrNc7i1WCEHuKT2uPox8MBq7+5NKBrVb
Ey3jU1vfFaytfL8619WPKabKrEUFceELBbgklHGAg8mls4/zkO5eEJ8I3XUQD0JIsJqCZURVqjEl
s6sctTlbSeeDtIUG90z8M55ADXkm3g5wd+C2NbHxyiDARl+1SaKee/tMPHYMmVTkxyWITUNEt02Z
XVOIV5ode35o4b/DRFvuHcot79hS/itJwU8b2wL7IxjJ3yUjL71sZDcRZqSGjlvTWXZginS0tIur
y5mPZ3UJn83erXluyUW6FuMzXdBU9OwWlXs/VsMNT/Rb38GBjEsxk5fCW5/FsOzU/If4xPPr2e5E
Yd1zZ7L1ZcVmzBnKwgrn2VHjDkytBG13QQsIFTbg0lsxDMMv8Ih7Dblys74ESi1wGyoHdalQxOEh
H20ZNxH86tW950HUNwU7veJikbenGPZ5aOmWiBK8kAzjftS4Y8jA1guQlw+h4D0fKxUjU/DwfKUb
fGrZuF7LLYrelCNUWwlC52/7BnfE3d7Mh3Hj145rVf4Lv/lpnleRzW5FuObcIshM3XwZ92Fk9tlW
tWL6puc2WRKoZKDPNRtfxHpF7bTien8ZrYfxQV8ShtKDv5sTT37TR9hSFksyDC0miaXrxpxyjZHv
89Pe2hXAZ2y3ZXcT1H39Nav6laHkRKYq9tycwNNy9ccfxaesgESdze6Zq9Mb6RosjvZdyAj7LGgU
wKQHOjzmPzUmuEiJFN/iJ9cc9GxYYiB1i3Z3vPy2R64wI5aq8qXkP0AXxMXQ7yeylS9EN8yRF3jX
kbDxBtDen4IpPncJ/YukpnXvkX+ET36a6csx5A0WKFfl+CbRu19ibaQ8xIyc9qWuao1ldPq9dfuF
vN4Nr9dtENDEdqGmZV7x9b6tB+zFy/JWQy2zlWR8EFozqPO8hKNyI1siBxtDg55NNdRjjoeBt3EL
Iv4An2YuTANp8yZG4DyVa1k7tKgYmE4flR6HbAyPPm3kqvCHc/cLtsx6emvGiJtkdiUvsP0gCYfz
1ZEiklPw5afAoBNi9Z4m+4nwBm1s0DEcuJ1HB9qmdUr6/gUyuoN3BBl3hndN5vCka4R56gqKNxg4
1G8ZQjDC2AejvygSV2ApGlBZ0dY5jLVO4KwZBcMSJN+O1nZ8FxPNl3d2UkeVz233OT7ipwgfcXiD
aXXXKf8f6TzHglPqL0bJeF1/OWBtSWePQeKttrcZGKSY17vV2ElpS5kncdz6oqdQOw8nCOgduLKU
JqL3hc1a04dWUWg1r0YcEvTop08ALNkt1ImoNDg40msG0Ud8i8MBG5p1hp60dEItwPrwKq5rrTnk
ogXXmF6HT+YMpAwr2Ft69T4nHJqj3gwMuAokNXZb8fgLzCUQ3VhQ4OBSU+xdsozklrMPl5zodsm+
+CY05F2hEsKVgOfagVtxHcGUo0aowBgXVKs6fQBwCepAen03vfyGy7XADK1pxTUhyQc4E8+vMbjh
ob0JeXKTrXCk6gsIlZl42A0LkXHbO1gt7AbFNWiXNVKwQQiOgFwzFh1rg4wuaZvFVU/HWUyTQkhx
/kVClt9s3/dieGV91bIHvF2qp1HncQBS5Td4Q0/sWRpze7s0eSQbMlAspkWc45x7vdBOZYdsXD+7
CpFVV5vgHGKLGmmqZv1qcB+rD5hhXXhRVSOg5uMW+R5pbYdHtKNU8jdPj4wMRgo59tpYGBeaq1XP
umsBtqKAy6c+ld3ocOJKPpbjWZ0zUOSwAjB+bpc8YVjnYf1/inZlTC+hmmLMiApKwmgVqsRTujus
qzTWtJjkjW0LN2g3TXyPppm8OqDaNrPlYWvEKA2q/sru0hpTdH+WoOb0AZjx9r/2Mc4UEG1o9C6f
y+6aKIvmKYocAmMkztQ3qhnzcHllIL13BP93BjUV/2/ocYPUM88F8mJNdQPDawlHHBJOFCXrJSc0
y7uxaxb1nyle8Pz0WdKbE3bmD4mjnikxzfrBhlPQdgGEjIEPaQ/VKW+5SLSONEHGYh3C1L6Br6kY
dUGo/5d/dfEfj4ryA+OhoSP6JjjY8QeD/xYKsvDP95xXD4XVqUvlkqgV3nVvxt9URpl+7CYARxFZ
OSneQ6NetcWRIbpVbodj3puyfrcRXkMO10/teYkDMzfS1UMaGzsB3LN8oG0ws49W354gLtWelgTI
7d0e1ygUIXb7raYnEEkonqAIYHx5lbQco+sX5hhO6b6Qbi7vpMm5HEqHVym0HUQ01o6b8LMnFT3c
qBpQm2tvk0OlKnwIitxVQKH53TZqLLdq7Wjo6/61DQM9N2yH+WvFuRlwDRy9L+azWHMtnU2UBN3R
8eoYHiZejL4r4cULVYhbfnowOydvTzxwTRAM1JTGqTA4D2kjwi05j/KXnaKes2kZ+eyG7t6Hp69K
FvN9r9Fp8Olk1TfcZ4WP7oqGrYHZB5kUyOSSbM7F1RWEBwXb/jI0URrK9CZqfiWZpFdrdL4KOZU/
aMdPfuzxFh6LXoKiaN65cVlLZd52YJZ32NGmnh71ioBzsWDbPEEaRHx3HOLpLO1CPekYIhMXGlAT
vXcG5PlPJzDRJF3F1hDJ/zJtzNCIKgnJoTML0pphixYfPbZW4zhu9NWD+ihsVhdbE8Noo+/xjktu
m52n+8SKZMrEU9HMJYnxYlvHuelBoqDzRgIB4lJCQv0VbQsjiNLWZqAVlEHORHzoOLrtVe3VLDni
ROFBVPd+OnBdwH4lq6Vn6bX4SHLl2OCP+MtItTmCVJzSFjpUbxS3ajktOk2ciQQZwmJLZKql+dIh
d8ZCkgDqEM8qZfrcwDLwD3femjvITqLUVfm78MvaoBj1QjFn8j5T2dsjybHOqxUIGQEpC6v7Bfn7
MOz47QkriVc9HUHXpfGDU+y0ok1BsBu1X0J70LEwqyrQtBeBIWUaXTeOC3OOcw4ADPKYKbjpy4Cv
9zcpXfXjcxeY+azIjewKAuti9xy9KeOeMJAKrDxPRGIbJDRJZ5iQgR8+OuuDHGoPmYoXrSVw+42L
ku7ziNrYV1UzCNzl1HV/fDCeB6oy8CWkScGLcOrhUCdoxehMeTFewVpy86+7iGAABV4DGZs/qzNz
UyvrGFHkNpbts2NTpmFQLvSxjh/PaiWgwVkjMH9ef7oP703AXiufupeEFfFlT1DOuJCscFpkJldh
nMalPKdPqz1uukHwe0FOm0PCRaUFTIeYEP7O2cf4kpyVugZ7V7oRMOArCY2fBHYC8utq4CChvxQ9
jaQ76GZIdzxZnTRKIHS/Zua+rL9UQ+CHhs2oZdHz6JwvLiYQuBHwhtLoWLVCNkEGHKWGBT87dU/o
xpuORBCiCMA+iEhryyBWqMn0X/jUXjHJoe2XBbP087Q2WTW7VSKpaSeEMDncatLnapSllQ99hwzH
2dmZhCAurf8ba94tTH0LcOoseQcz5u5x6tbU10dvLv9QWxjGOGkQiqxlPz9ViXsFARDt1+bjynPz
IQoG9L5JPGAGQp3GcUi2fK6Z0zbpAfX6nYaHDRuY44y9jg6UUXm9btA8oWVLt+2NVwH4naoXPHXM
bdAddtXizkvhiwi+ES1cT+jNYuRNWKd06ORogRNDSAb7lo07dItlBvLduPeLC/wT9MDvdr1fF2LZ
pTfzaGvgub/02kcbM8E1pgmUmhNe2OLjKR5YRGryQN/JFrY3ZZuzDeyYzyrTgw8Rwp0MqZoJcxgz
WsDR9+zuRQryBUiMWUrcV+WwJcRFKOaxps/8TVBr8L28sCBqsAHKHlWSKTrvbX1nQHFxiii6tlTx
L7An7yQkMUf5XuITkZWHNXkl2oRd/g9yK48oiJKYjzX+0V5cdkV2byaP47o5tufB/Zpm3ucAtsqk
7vHVeLF8nwM2TSuBpTflRjGRFXiNnup636jFTCYAQvDItBydcPRla7IT9gduScsVO/Ef/xbR/fX1
rEKrNq2ClWIw1ZCy3QJn5KErWJylDSI9WL0K1gJP10NUDziiPrnpF9wVmXecPlUaa0nS1ZbH1PMB
/GqNYzV8Jp7aEJYe97JCE2OJnem56pm/qwDL+sat5P/bQZcu5k/WX++w3/sEJYp49NcGER799Dbg
3ffChPOfADFKizIIE2GD1972sauQ6+bVTcf4B7J6Q4lPBVikQ9j4E27jvfqPX/TWPhvwPhUcDQbT
CYAoVY0GH8cdjXKvV0DbibGqnxE0Dqd6SN8ODBPRfONJwCifAJ6ZYSxoGVMgQa6s7KwDgYLa7arJ
XstilBodXnXycEwxJ6S5MUqwZyVTPj2a3J4F/ObFn/Vx+SzyKf+V9tLsXXERwpZdrUNEGnSzIOhZ
YJwT3eh4tShI2JuRViuowDLyfAoKvPI5zjg4yFTD/SiNg7+Yd708HMUB+0UKr5c5JsfQRtN4/dRf
q5M7iHCyecMKpDxbOKggbafI73B9cD5iSoA4V9xMJtPjzPoymOkVMITQ5ZPaP05L231lUTI6aZHu
EU7IADtbjqU+vkhnCH3fc1AnF5P+1UDBSVss0ANP+v8SXPGcU4brWg3JTe8oZ6DnPce41BOgH6aA
LStKtVMCqbgku15ZUVOl1SY3rjMLG9QLU6xNYOyVwvYCPlghdBp7m1oB9R4YVwyASC5F2L2RXDvY
y9tXo9vZFgwGQRRFo38T5naBdjksQSXXJn01qMKODXd3spQtzFw7nOVZQY3vlhzj0nbWILl9PpyI
Wil6mOQdfZAVumTtt5c4B60vYeOwWNazfKarruPesar+HWbfPqGYMISDxQiOB05lmtBXzg6jbYTO
rGfB20BqzpiMogl2qtBlvOq80f4bzUqvtWNYG1la5bfoNTgwB3HS8PBdKo91y1nyU/AWWdC17RBP
E6TcRzHfXip9QBDCoHaBYCu5bIX3TtEwFCT9Q1Ag/nGeo9NRB1kTqm9gSgOAa0G7+AEX9BXneHy/
RIDZcl8OvyyiCCv/sHzm6+SsqSWHhWupu9+BZ6CYRmBRghvqb8BSTlq0kIrfaO+hUzzS6GPGBIV/
CoELksuUSWmHU83evPA0vgFPushXlXxLrHblzqG4v1gTth8gk5KaMjN6firGg0l0/9VqghlxyyHP
J9bmfMAZKLgjAtPsA73lSO5XEPAbjAXt59Xd9dRlSePZJdHJ6rtpWurYk91m4Xb4ec9yUi6dvLfT
xhafsFAqC7koZKMGcpSFsPLBQuVTVMTY/7RFy3MOa8hgZBJOckZXnhiZUbV5+HQp81B9rguScaaT
jcaYNBGsgv1+8uv1CYxr9RrcIB6Kyuyhpt8RQYEpkD2lVzydiV8N2x/WhNcVncs8n6ZRdAYltPdt
uHmJZacoog+gyrvvziFozQZ5ltqrfCdD/hb0sFo9YJLmqYeiIjomwNnutKrYFLjrFDVSl2EMIVx1
bLkKi+I517ofJmZJwEploceYeHCBNOiRpAHsBYWrvWNN0seWhd0DnAxoD/ImGA3trasUGUrtJhFI
2nP//c7dthOBychgfQCN1y0Gc1qtKw1TDqa8yc0CSz65RSn0T1LLy8xziFiLLbD+OFO8ly7/sNlD
fORAD+pv1LIPDLq8QxkzmE04OUAhEyld/pKRVieUbEJ03bBmzRtpLmRJ9gAaFurV8fIQ4ogR55vo
iGty8xHq0jT0PM8nUuBXzw7AxWtt7rz1111OkXc5xVA24NCesCJmHid9kRdR+2n3ClFw6RycJ7Xy
M2HMGEKUdo9vdFWimOYt/F0fwyNPIoynyDDjYVXQRSLpjAp9ZcUqn01J6w8/vgy+IeQyjyr5Fnqs
64RxS+Nv74fzn1R/UVTKXNp4iTFhN/Vij75dCSrScwd+vcCGXleyGNKyC1+62ZBem/j0FvbAAhoW
iAPET7EsMWMHUz5aNeS2h+/YqRmZ924vTGoSvdtBWq3BTtF0qE5XrEgwAFCJaFsX93trcYK1v6sm
NQjqIehXKMkzMbp4P8QgHNMcfX2PgF5q+GkU+n6RIZ/7RDlrnx6HglYXnKDBMWFmTrNJVFlr1fMX
Nzi5ExweWn+MMbudTSkfgJUuiXhdvExWd4hK6k9rRhpxGxWjdzxn54C4VHB2nd0Ygd7yO5vEm8/4
PhFvtn+fp3UO2ZGy5h2ZbTTz2UhDgUQVA8+vBDD1tye5AgImzzf+rwRvYoOVekhyYlAIHxYF13pu
HIXcnQA3N4x8dE6jAf500n/9WIECPeUVzhUUS9+70fTIyv/Kh68TuKlkvm4ddf45z8scf/nIYiLx
c6DB1utW8n4US4zaV387sCK/q06OPXra4mSqlqMEgFUfihHxcFlcl5mId0AD7NdjPa0oPUedIPkp
GAgR3KnFnaCF2PkwRj3LAGLTN/EajkSrG68Fad+BbhUn0Z0Sf2BfE/S9jp36toQ/lpaIzKLx8gBN
JNbh+DqruKBZZ3kjBYNWrm9OWxJ2NEK88qwmXLtCh0OpMO+HdhpQFQ4yro96L5fB3xX/6T+l4haW
j0a8F+N3ZhdtFtc61CscizvATqxt6xHhJfNKAWgkCXpFUCZCuvvoragEgyto5hubd4ELEDfnS58Y
Do9mk+Ko7I+j1OM98rrk8rDEQrAeo9VXzwHQH29aiVmEz+HL2EP3FzUtFNDdQf3MeU6ucyu0ePt2
hsBLhsKfm6NAaX7eUUfYTs7IJ1TrtAinzko0HG/kqH8Dio7A4jYDB4F+gK6sZjgZpt/STKfwAqa5
3NDJufAdEhgcto8SA1SPbcu2fvWOzZ55k46O8zv+tBW+Gl4Fr+nOiFcBI+z8bApWJqdp36HullQK
QuYAivgsG4LMCkSFuiAkP0w6klz8oG2A2RZjSrXV9OgqsFyGg+8FwlzLeVIZrM4OkqU42Kqhx8ob
+ImHIgqZQWsTt7FDgn9Rz4HxC2J1d0/S8UkYbwRIEc7Z7fm+iOxQcQiUW2Qn+vdUjSNzAXfHDKRd
q+pNKm9rLHlZkbPKZk7j67N0CFI2C6NfbISPJFBqSj6Lm5tPP9GPGO8Irp7sn6v0+A7wqaXVKKHE
+RFw/KpSyy4XQj1qJp6PFZ7vxwBn4mst0/q3OMLRZnrLDBlgaQBXI96W9v2vo3iXCCUW2htXm8Zo
OwiatBuFsOP7f/rSw6FJ0FjGSc1nXDLlPRx3RNtF/nyyUMhdquULHThAnMFUZlUksVgbEikKkMLw
8TYeoh9cemUQQM6uvVjoOjFaOZRrgb14WswXLZPR2vdEmxwisttv2/SVeQl6l57HDs+u5aeA90aE
3EaC33SVq8/4gbK8eJTgJmhAlXuGY32CuSM62EAovBI4qubR2z6mRHY/4dvOq52jhjx90qBX+zlu
3Dc9Lkow+VmTuqiPYQjyFu5CwhPwGGMrAkjccbmDjlm9oQ1H0hO0e+EKtBkWZ7qMQddWkpOpR8rP
/6YPQGnhZQ/NmYTHX44yRepnqDZaGwgArNGWtfNYWAFqrUapnrIlgL3kcp/iPRGjptXxWlUAQRAV
g5eWKDuTmedIjvsdAwq/W0YvTyxTu4K4yU9/mWCQZK230KepHmCIieafJYR5JAlinmka3AuAMmld
bbQ6lIiCS8r+K9CUuIAZ8MJLZjQT1C95UCfKBw5C16oyI2V8Oo1OXQCc0n+L6Nsv3RM6p+ymaNvt
TQQoUH2bfeAHw9up+qz/+8vw/p3NBeMnANQmCVrwCUd5xoWe0jlq/uArg3z/o7isHJSldo97xoWm
+WFB9zV99AGutFP2NrcOsohXuaRP9Ry8RT4o7Wc+F9xLAWzKtwSIRa3bigORkH9Ls1oLGrA53cbX
yXlSxUMRaGJw/l262vwa7UqYvru14zE1/wdgGlEJpeYqsWwQFf8x0C1BGPtPfuqfUTSBEB9E+CLL
XJQaOHPlVyrzOqe0zyzuvwskxXcdqvG7CiKnic2KTAk9KTshM5w/Gun7bR4LJsN2FBW0iqTv5DGL
0kInckcsOuzYsbHDZaEPh6uwymw2KTazx7qcG0bh4kB4wE8bgXMNAbMfLDSXAJEvTHLCxcKU2ogT
qaRLeIwKoSDla/Ch/wZS+/bEjfYLpjKSZ+GpOrB+Sn5y2ONQrpyu0Dje7rPqmnD51C71M7TC0D5Q
awcBlpUfqIiD9oSQ6vYFCj4+7TwdLgf1ZjeBTUPjuKzD035vnSqeFPSh/Xbpkjda7tuSUsHdIc7H
LVzEY0jmwdYfL1j+YIwSXCQ0DrRtOrXTiDrPp/1yAxkVJ+j4ulBw5QOOOhN45fDVpONFRmMhgIML
vOvNTFR9PLub4TGdwSlsVdlxCAFWZCvNnpErtSAtpF+HyqscUJ0DR+lgxASxi8/QukFxoAJc2CtU
8FxfpeJ8G3m3ILYXGVp72+s4/5/MVoHVu8Bg17AaAw3BoEY5+DWVgR+hk7Zoz2poBlvvPlFDl/wy
8eKpclKqa4IIGcn0PrQ3osro+GMJ3mVaGWCYHkW3ShPCsb+u5OS6Lt4NEy/a6l2rGt8Mti+/DLIZ
goYV9uNU2u2cISEBflJfFp4mKcBruYD8cyLgVzZ4dxfzvGxufDr9Dfr6KN9sQ1qcWTDmsvolSvTw
9unbF/ZAw6N4EXh+jbcUzSWCTcVPydU7ndhNpQIcX9PjYzzlyGbHkvkPI+1a5CeszKdzMSiULIPf
y7mLFBWWXRPhKEm8RXTzjLbI5P/f2sF6ySjCw8xG3FLg1r8eNZ3KX/5dlcvREKg/+tV8X1mw71PR
W4RGQpZdlfA8j0ieQWftbxj+Y7kuKRg6IqFU40OxTMOGHQq7fJEko/+WR0khQk8JXhRLCjxapzrf
N6snhXODyhB/Zb40kXXZlt3UblD72kUXAYX/frA0Y9RPXLdP57hnuhyqr2mMsIXpC9IaKpo9TVkk
gx7AfbEFxyBfdDPyL5HVxO15jhV7y/LgMKxbI9bQsOSCzEYVH7rmTCYgvVm84h8kFgXe45hZaEYp
IWOMjvXH1QQBbtzgXREctvWql1gbhY0HHiX2hc834i6g+o39lhp0yuxlb2TU+NfR89XiNfUYiwyk
kyYeqAY93xImgXygOthjvoIQWlSlHn2R0TCZqXZRQAMQIgRqO01eyNi9MizJrTmX4JMHnVrb5COQ
w5QJ3VMQ+R2E5P5UqbqcIMVeKB+/A8b/YeI8jH2TlAREQSD/kTSsUAzgd0LVxIPMxUpoa8/mjPwJ
xsGP9VAzrd0/69JWzQact07LgFKmlPWMNnAeAzPNNStonbxMuu5c1NO9HZ0XwAy080KRpy6g9KFb
lZvaWSvGmu+Hu4Pyioe+XqUr8JDrIOt2appsF51+iJ1Cl/kBGcALvPrl6MVTvEfuVx8uaIKDu8/i
zjPojMUQ9CGntklQz7D1Tlp6aw9ZmvITCVh15Hcz5NZYE5H+GK4XDVfb6QWnQSJ+iHa8WICXuzAV
LZsYvVhZ5qqSpEo6k0Fvd3DukB2P0/4Nz2jHlQR2FXIm/CCfBT6tu8qZNgbmfLhoY70qcb8sQROp
xAWsK19WyCszLquunVb48+yu7Q6BlL5WP3UNZ6xjeimPY2KpgAd7p+SlkJ8j/UDk51pn9SO0P+hr
Vm3ec+w1nCud9Ea4CANM8j7nx8vvJNUBw7Q55bL6/aNa2JLE90S5qn04rCtnC7M5TzhY2blev4da
gmTE38sIA/Akyoi0haya1kqVOHFP34k6rpjpycgEaVkKrg9G5hmKR09xA4Cur56HODTO5hy8yU+j
0JyKBONc3eHty/bVGIxGyLR/g1Kv0LuWWE23NNQnrt/kpCPvSuOUSG9BYg6/doY3MKje9bgi00ff
ZFotyYHfASp2z5Y/KQZIKIERUBzWq99BWQ5FjqAzXbO9r/Fiuil12Pm5F7AC+SjO+AZrHJ/YXtJJ
84Tp7+ltvm+9UqdDrYlzfQKd/HCbJxGrlEzYLfMBO7bYjKrMMLTKwKDViAOhP3ItTU3dfLLLh9x/
tdt0fO2q+DCXVCx02GtW6WN8mfIFCgJ0+kK8EtEYV95bN3sLPBLHeRKOKeZqGaAQoE0lqBDfJfob
fS6nz2iFMtGcPtjEOKhzhzMNsLwQ3yFkAh6UlWiT2MMuhlGnXkDB+VqfG3PnIsJvZznX3bo6tnj6
r4OmwjLuDyUcUQtl7ecrX6nnRzAeVoU+obuew2+qtTtUG0Rg+wHYYIVI6gigB6nruNOqKEHY+9C+
dQCkdZhI86QBomwj41pvB4Q5C3MFh2uaaiFf0PHItuqJudd8Hx5zxws5CN8sUwnrnLwHtuBK+9Af
+tTV6/nK2uRevQVYedYiPy+5VopYKKXUyd9YoIe3gGByh7rydNnTWFp9j6G5NJp/SkEIbXUQhHaB
R046xY7hdxNt1AOX3jSVQq05VDqyeCnGtDZplycnYBvZx3LYQmbQdGn3KnGZjXB5RJJfXkaTic+Q
ccOiFYeWuAxxMJ7EBCU+K0UONpQxktjvIUUee6qqnGiyNgtv0xW5US2zHeREBEOnq8SeXue8x06x
5AfjvxWImq0QS/gqSjrFODEOYrMofg2X6ii72pRimW4J/gV9+JsWjQegOhPJA+/cgIUxNjzPDhZh
cMvx/qHYsXIAh8m7UPdo1DL1hRCNvvT8Z8cP6jlgDwt7j5bfPkFnxrKeFSIGd0oryXijao3hPqlX
ZAITpp35z+X5r9qXc+uUS03YSM0CtXTFKHjnaGB3PrW9igH4n6lERZv9QCaLZ6sW1yJxMZkdx4YV
aXjqTughAH/AYSeHmlnokqQLZ61TTN8eDAEAkQBH9qKVLxrz8J6BnhnOtCa7gq74kHlAtAoNgVyZ
2mGdK5Qn6PNh/ZP2Kff/TFu6zlfGGEklcz81/fHugJz59fmK3laea8J6FetxQ11jitT4xEHEWOo6
85L0RXsXRtPQFFtf6K9H6rLlpt3UINCFfswXBCSKee7+LZWp00PsTyUCkPTzF2rFoutIK3cX55e2
gRCgoA2KdAHYO1nrFTuV/XtDAKU2+yBZgoqot+ILfok4HaQnRWzODVP0x30gt1K8KD1fCJJiUIlT
4Ae2Ft108/qHDHvQvIcR04+RKVr6SSRbuBUQZJkLJUf1tuY9ebASDjj7ocEhn8+O5wQ0XjxFlJru
QRu4DWHF3CiAwElYS50ZCd2XedxKnHuvrfAeDsKKZv9v8BuTeTUTd6DIOPlU6Do6JVw6bm8W3kZf
lyH+26J1ovsCqMa0kW/ma09KnfGhMJ/twlF/XDAgqM+sLkMkMm8ST6egs5Z7vZUFgCf5ZEvku48Y
UMxKwKKhto1dVSmGoXV/Sr4485ELqpRdBg4M22R7Xz0qdVoE5XLQI9mWb6nJLcdyqRctKYvZjyg/
KVtboL4oUrEwQQFBhPEJyRtZjJlzDFtENqTojXj0OpzBXaLaDsF4CkI5lzbSJus6n/azr0YwZKk8
g6pmf8pnqoNSnPKtNm0RmAL8cjrV5Xn0qph3uEa1t06g0AKCU7x96CDk0H2xsbhE63UQYdjdSy1t
DQ85EWRMI4OOQMBlhz0fE+eFJKN1fKnMFz8RztVkllPZk/xd0CVAZLDxKvgXzrlMMomu0xjlFPLi
esQhUPqPZH47OpdvV4VsBaIJyZVAkw4nOFZEjUNBuNxBTj4Jq1bfzcYzSE0dVSfrdEF4XxbZ1gCs
dEh/DKPgzxjP4xsU2DCqHIl0uCmOqTXIvZenmCxuEFS1IpSn6NdDnfh2ITro7ihk2csLg33LzGGQ
SAsOMDytFcn+y5NyvAFU2cvXshQMYId8DBECseoI3HnGD8/9vdsShWefmMn5SBjc8/z4nAzWOU2Z
R5USf9ziiIkQmuVBHt9eMbqpsGVUYlkgoSui/qyyFMdtVRI/4pnxhyWz4fnxafIBMfmGdT7yKstc
hSskRNjEwLw4x1c88ZzgZcpGaam+dDtoO+FPh5o21sh3rzIDb16tkhE1q9ccJ6eAhZS7aZcrBACl
csq45IwLz1/1F/7BBxMUNRaSlQrNQGYr2dTUlDLOfPnxCb8jN/y216uWOhBYtLV1Jm1Hpn/cGyuK
bUDtTCD7dLM8kAjF5bBRPxWdGqacEaqjtu0EvVwbdeT68sAxzAi4v6pt57OihgSa7f1pEgjBst8B
lPxzJqx+ZReDp/2I5VjCV45exlFTp7VlyNK+OCnSKJEDUAZJTt5r3zKS638fNjmxdHh+njC8z5KL
yykYGWtgwqvJUqUWVqodER2/w8mBKdfNCv4n5uYK3hR3lrKEp2JzNMMLI2d8i/PikDmLHEBYanNY
HzgfCUbAuTrTlGwxSdWRwtMgW4NVnhFQZvo4/SEViUffCtngf1x+PXsUu5cnlHHKI7BXfQe/NVKX
9w4QbyamyU/WQbcE0vCD2RvTP+9DtY6hd8RvU45+6yyr75RnfsFKaFSpicrIc5SRQp4vbqfeXq/z
rYAHkJYGuPTeM7+FHO84pnad6Ft6WGh8YvgsQBQfWDjumVNJjhSt3HHDNqdJIszTegTPsMnmFWti
6IKy3Wn/NGBGnl0u0TkrdTFjRDSYJyFRcejXOlyuH8tfTo7Zfczq8zk+DQQ5NJ5rgECA4YHKzE3A
yrisAkfd/zmX+ExyfQZs7e4uM0Nkh+y+kHEJ0IukEqdIsKeQa6gr4Zm9NmiZDyx2yqqk1ebSk0D6
cDnrcyW6ersvrhaVeiIHcHWUt/R3og8PeQTWl0JzmEt3nhC1cbVnYYdEGhWaCexds5vpZ/ZLRJro
bVpAS8i8rS+Ed2fXctFdFiUQKVWAx8S+fdpqlXbPHncaA3XWoY/baCrz9o+hbdzYmzmrXXE9XA/w
rHREhteCxqKaqjL3fy0Sdgr7XcDmOknB0pWmg2Sn10GY+IAQCiogzdjsxQYeXdV2oO+f/Ipth9ZB
n5nDwdy4zIRVWkUy7A+T1xAeiTEdZD2DMI97E0RrpidKh3e8arBU2sI0OGDFVHx6YZ0NIgICdZMi
fSEQi2gzGybvPIXOka+LT+t6irwp30Ba/CFtj/jLEDZ3OO4eC3e9JE3gfXbFx1uh34830LaApz2h
kRpGHbNHCM1Kds9BuMOjE/lo8pxqbkNwdis4yohfXjXX9zQfJOWyHBAQb1sHJE9tyMVBioER7k92
vLJebf5VzvInd1SgANaooHunXVDbRLnl/zoBLrZaFxQ3AGvlLElyTG3MgHlH8BcMdXLl5myRbRjE
QfUyNTMiiu71Q8fCarw4M/Jh+2CgLv92+uxBgwqih6UNDawOmD443G1fve0O9x6YAUZrgGNjqAMS
u0T1My1zavisR0OE2kAQbs78ofoS4jXkx6f3wVpqCBK56e430tseWYJ136KNG7SE8ixeG4p0TQYZ
7pQow//94gLyv/AwlvenwurroMrkG6bXU89tihCVD+hjNQKGuSdnWGbMJ/BApTGuhud199bGeSo2
3N2GuuqVvnkk8AAwTpk/Sm7LC+DB6jlg6OWrf6HEAhsr1FI7bPhkUKP0PpBSgQl36l0wJ+6ano7B
pwsetnYM84eqq/WfbKgkBFal3zEmrtRl9NSuXnP4gNZQWcDHI9/tf82Xm/31wjXW5P3z7Zs7PLtI
BWIeDqP+0+yi8uJbouqNiwpWQxXJ6Hjm6IKvLaPr4b/QDaOjRl6NZHeF2NZU0/sz1qCvq4fw0GLR
PYp2JlsCyc9Tez6IZzED/gco/6uSsOb2vPUk7dQXWLJyAnXeIYQEqW18YKpR0eTvoqBwl5uaMyNn
PSGN+YCclXL4rTUtICEhYUzRZ1lify+katdj5y/Dmul4eHDrhzyZE9W+HWkfVs4JT/SPHXLyK93T
RlwTIVPM4TU1Q855tGNR5lCwm1u0JfJH1HCkVWNk6/cDMBkEJarxQDhATlPeZ7BXMiAcQxaHMH50
lcup6TAPxZZNNsloDB1J8S+12ctHM7pbA8ImYOKfof5PPsqK7o5SLAzeQebg2YE7C8+zBpPQabpm
KeU+SkDKkXmm1lKCKAoHnlQA8tQpoQWgqD3k+vgV00s9t1DnSi0ikiMmLQld0Ynv9F8mY8/zqw2C
CUAvq2pfyeQILu5fPtzdWHoeWP0hieytKiVnCwmc4bsYXALi5k/s26LwfBK1YzdzLgC548GI9+LF
itJzUv/NNoLbDqy7sFqFUCpjDusi8TxQQli86uoFJQYpK3Cf0HXpDbonceG/+yTT+fAyI0KUXCe2
GwcfuVFkKAFjC3KrtxWc3kefJTnywsOuOgG7D+4eUk4B1sFnhayNm5eDuZGK3yzUIur9/WOyDKGF
0RdgqEJn0b46hpa/lWa6CMnIJl+g0sHXZAKsQ6EBb0uF96ornAEJlRAsIJ6KxwHl55QJG0M+yrY7
j6sJj57MDwtEKrE1/DLNmopUxZW9itjRJqAJj/gk/QksGhdcC9zo7ChJyMVU/Pg/azVdGeAzYXi7
ZBrZXEhG3Qni8gPiRhebUZkPuCqXaW9h9LB2uWjo9XLQrRkzn9wMjV3/M1eC5zQ1nrUeooD1vZM6
YIeHucXjraoYYlli2WMaXYIkJGe9cF/6qffM7tNdRdjbQHpeKdFjBWIuoPDTtXQ7btLefqKdjSYJ
JxL9HF8TUQTP71QP1GJTsPXNXC6pYY/DRg++mW9BD8BvA4O6zYHg7ef10zSeyLILllmmpi6FYUGJ
PJA7wqief/S/ZDC5XyJm3qLd5Ihi0vOsyBS2V3ESgHQW0ZkrrM6ihUm8j4ll8rp4H5pHRJnl53oD
XbJZjjdYOxVgWm5ede8dtdMc4H0E2K3R6PNPsZNBV6FMECAkKF2Xcw5lUEvLp5zcAvOQFfGMpLhT
gGhlHFzcgEBx/gg2FjEQaQ90+2AvjpxeJn+k3OP6a4acjnqrub+0jVjr64XlKhxrwXX8RoD4hcfL
i7fiTmqClsJ0+vnXZA0dGVkvAi81ubIf4cSnB025SUEL02PIuMjzG7Dc+1vrirmx/yjpYbmjTcaq
8TY2gx7+d7bIcKeHSW2GSARycYguAs8zDwL0HskFzPGv7X8u46IR4Rc2ukDpNYLWSNSgcMs6mbiU
Ff8FXC1GHj1exFi3rxN0GNh2t3ENIdGXL2ADX8w5g3TcZm0fJn3rlg3QAoMYOOKiHlB4ChTjviKU
U/wDsjkcvd3C/y5VNGRQOoqrJ/Ut67WOhm9TSDGIxBLOS/q0q+tc6kqebN+HJ+U1CBtfuoq45gxX
+pIncXLO+9JUX8VPnQ0FWlS1TUoFt9VaBJr+RKoJQhs3G22oKJc31mwqr4S9WVMaYI5z6G/J9AfB
K1lLhGmSB+ft9QJIuGLyM286WaZ3SNK/CEoR6v9CramC9FEWswr7WiNCEN+XwjzPmz5GPGkAdk0q
FOX19/Bdq15tl2zlbxD0pvr2TJcSuQIMabemji1QeY67JQdkgb89Q9nOEvjOJOj1Tq99xwX0UXob
kMzjub7fHDToG1hi+yLuyqtEUeX4lxkAyZTLFrz1htlMh35iPvpQIJw5OicQvw03CrNRqdJnW71/
rQAI42Pg3jn9eoPw21Zghca8T9GNfQpN5/1fzRVDhxzFn+JXrjCuFcR4n5+SQiJDn6HLb9UyeNlU
8kAMVW5+Nw6kPXYvb7/pkvg7IdxcyyiKvqCn56xREnGT0L5GyzgQFQW5DXfewBHyoH7rLLntzv5I
CUAzXWkq0QIIdvFfXmfi++Iuic/gGT3yFXfUkBZvHlYOhhEGD16R0+PDtwxiIASC3vL/TC+LXhuW
bi02hemWIb3Ov5vm/NH/aWNcX4/bMxnpg2QIqQNMxI0vEc6Stic/nt0qXKlN16CqdWASsckPW27S
GGgDm880XarSnh3m9SRzlOPdyuxucpVmLiPNQzybWcFqNhQvOv170uJwsmYqQ/JxNMvYKo6YbAcv
nc2e0vmIPk4BWpxoWiii8fLYgNEkzFIK/FS6GiqoAHxHUK7M8zWBnhL8i+7iIcmPitnE1jR7mQvM
asbqON/M94ohHjpaJNS3P17deyCaUgUggFNr92llihhDsPBZte+4Z4UEskxucKEx1kN6YPK1bSLS
quc9I205ukomCdM4t9A8CJdHMtVC/IXpRu0CfM4cZvo8Vy81L6D61q7E0QwQgo5ZySUwayY3Sypm
psyVDYP1b0yLiKFTsOyQ1WK20LlgCnWtG5Yr7mQhfjL29HKCCjOq0IenuMk/RUh8YtGK1oEa3dpL
MExghGnGauHRrd9V1XSALdyG+M4Pg3p2qTr7WDMjLFHFJYwpDsZnKUz5iHfIXC8faGIG9vvQ49Ca
D2VbnE+/QfX2AFftPc119HFMbWmsj25mRanZMr+uagJVmHg1fYWR5dZIuAY6nv1Ql7gI7ZBGdJ8v
46IQNMwczVret1BFimBHJH6ZTFJLtIFa7KpY7Qc+3ON+tPBV6CNVv8CMEp8MqUShdwAy9IIUVtbo
IaWwiRRq8AvaX533HKu6EwORgh5QzS5bDenCzoiJRDGzpqxc8plplEhOHTggnmJySK0vmhdsr/iD
UPKvPAI9iyCohZ4nZ+v47a4ndzg+AXhX6o8NZtAnJsln2qdg/RGGpnfvf636kGz+14CyxgoWrJF4
qXCo7Uk5kpewGbZT4nXZ31UzIuPpUKOnaWMZ7bCjkqxcPW15/WSU3+8gkEyyXYBZc1IrCkuk0IAn
cJ3+5qLKOJjwYiS/QGKoau6hSCNJKUbta3x8Iu1JlkQkPkz9HfBWhg6S72HFGr6UBtfdwt4nO3gq
b/V/m0Z4h4vOh8f0qA9UVzXYzO9pHNhA0IH0Zqt65WJZvZxuuIvuMcsBF3ejs5NAywjNPNCjekHN
4ZI7fe7cVoVZIdRFlYh+ycmzzx93i4jiTll1QvelBcllUPRF7BqD6OzKbygtZSmKfb5XRG+U/yrI
5wiagQpVruU1QMzpl43dpnnxw2w1wLTMZVE0U0mtTHBO6LvmzcjsZhbZzRIBfBtyO/swfgX1MEHo
j1etpIw707FfXPz5FSsjxJM4JUeRy8qY+0e83W+/DDoVrKR1XVaaFy6CE2wMZrVBjPCgYRgzLmpj
aGQyubI3fka2l2TmhKeDC8VYvnhDTyY5p3jxJxMM8AXpY5Ygf/gyARzFs7BEDK1NqvmBYgH0BeUI
hwexxluQCN1P7znET+Qmt5PwlQJXPs590BnIRvFZDtwFyTt5foutjwEVCUNxmM3sR6/vhd+qu5Lf
owiUY+LeZyPX+eKyGTTD57om5gV/7JPio2eyM9R5Zt+J81osafZwzzmak+DdCjyoLmINc4xV8Agd
XExuHdJbJzO2eQIrOh+Wp/szp4h0hkNd3UFgG55xY3vwg63+EEHS6lwvtQyMxjTaww3Z/fXtnzOw
6MQo/L4B/lE1fMEC0URkGN+luUWtTCwq1F9Gs7fmdnHvucU26OiOhMjz7QBMjHo3SvZwGNA7oCS/
2GPZkTXLuA/TWEzCZeD+ZbWxrJuflqeJxmENPsZAFRlZObKotMVCE7e+mBdZFXUSRH6zkpjfyB/O
ZguGXf+BzgzjxiQX/umGQZD39m4bqU5Mnjsy2lxOjCjAVunc3z71bDV/DEuKY3KQu29KWCH7d3T7
F93V4qJ06a6pq3iqImFknx3JIdxdDVH1tPf+RhfxSPr2IHL5bL70W36fyTrqcVDACwE8V6fxmeH9
lNlaucDQ5UQpUYtfxHn11gQm0ueJ7L2Cb9OTvUnSascrpPKVK6bzrArwewtdsuLboqbwmVYbcefC
CNjwC8o7qE/8PbaqdV/VrwDcJeMKP1mTSTNQSfXm+I15sOWcZDF8R2cKSnv/N/oOgxOys8HLSrmt
kI3f8N5JQlv0Ala2FPbKSl6nyO5RRgfHAHk6RVdYvNmS9cC0lI9pF36r3W8eWJT0I84IFnEc715M
OW7n/MSXq2R00OFg8Fr2o2OF9F17GGPL3O2PLyx7Kwly8L16wQ1p0oJ6z+QYp+eplwaNhWgu/JT8
4dRFT0OpCx6ViGrQTyplfKq5pv95kdkqyKrO2bwE+WIQqTIN8610oB5V+RoUYSyLajt/RRI8GguO
XZ5aM/FM5/uuNPXnRIMhmJj8OfprWFUPujR+vbZqF0NRmNyE8k1WEKtWZ9hW2/b8m06I16rFY3Nf
+tOIFR3WSlEQDbrPsQtp5u/k66tYrtIGuCQLy/wXp+4LLldP7yxi0CzCSB0lV6zUm/CnfqH3qhix
nfUK4d6aP3G+dvaqMA00SbuFMRURM8YQTlefW7+fbt+iatS+8ZQbaS6/nn5I235pRdu3RjQ67HVQ
fgfJUZc44ZHfIqD3dCT3pRqBn4c9wCQo5suJfmv9CBrhr0TAJFKuszbMfd0B6zpaoN9VNhsFWT4V
f7fI/D+gKEy1YnUVv2l5ch3SpZtSKq/l4cOV8XCFR5uDgDYnUk2/qWaTkge721mOmT3GfWDXLuFL
vg6cK0ed8943k4PJqN3WUJOxIPJVRSWTdDP/cp3HapGI4twsBQSsZ/HH3f4jVKqfuAiSYW3ngWbD
ocvEBKYNIPN5rG1Ud/8tdnByJ0osmWdWwXCUFpaq5+oX7d1OIcu8Ps8G43UO9Cbd8bEP3+U5ytmi
3YIq4TM4hx0+2dzK3fduNbZylS1AHSWojkEzdsj3KY03rUox6SYyx5ttC9Si8aDDujjlbIil8CYH
Ikm2V84jK8U0PCdbolz4xwyJjSRsN2NQ5Jxc6CpfjDTswoKdht4SYVA4gWhiDP7IFLmE6+rb9yUL
nQP29Np8wmZOd3/LhKVqO+/RTsyMTxwwI1pZCFSNX4flqwcLP6gLCzrPIqRqsOSDIS8gWhj7vt2/
sjCadffw+6l8XWaRDDaODOrtftZffkyoxj9YXvkoicv8k0XxWtReFt37sDcfIoov4uOymkTg6OSG
gh0RTsnSXRdwpmOqH9QrEmqjTpY9TndoLSF44SoHx0yzoxnEx8ocAzHTgxaDLPT9n2R5XHL7xphZ
reTSwg9TbYXUWymhmGssUDsNnIozMKaTCUIEh0nMsT9vL1YrdmG/hfAMIZGCm/KMjf8xNE5XRsyQ
hZi7thUCBsOru82nlS1GPtGuVhfLvDkAyU6R6Y5lIKdRrStBLC87jC2KP6nwmYyGMowkfVObxCw3
M9acYrWmqfRtj8ya5VuNGMGckWWbCx76aNzX40+xqyYMNYXghTMt/3ItApa49mq4F0rYBFuoZWG2
OQp7DumkVtALoNc5Jzsf3ogLtvLF6lnZXBnkDxhDG1Us9kzyQIQv0hYz6R582qriPn8MNUKQ8DP1
rWLJi6B20WqXw6OHkO0bfCKr0yfeRjHXTjoxJVeACAfW+JGZGDdhNh1aa4wlHHNxHRaoVv5xhsMV
3vyh04bju/4XVOe0MVs/LWKzGhbs2ccZhylDT09DXJ4jwZiPXX/gHF+otHY+yil7xr8rdSeF6+hB
x01d/9cN3Ym4kZc0D6aN+lWbQwES9Whez1Lcn0MtRiDb2vSNDJtitEKR/svY0ZdokIQg/5FtMTqE
V1QrZnhlq4kX1tv2eNAcxGU7rSWlc6QNZkD5+NzsUQzqIdxF2dbyhtK1VLlCzMMSB50x1mVWpjOK
Btbp9zxa8CgprsgTwuYDu4GzO0lnBdbESQDB2U9PHhe83ys7zDwmLjdeyR34wTdJRZHGft5fJNTX
dnpKX4RO6/ItfY21RErcPAVYNsL7q4UF9og4BD9GyOwEpTBQLnZaPVncBKUs+qOffUJWr0y2f4VY
GBlgZ4l//uCcq11uF+fO5yeAq4pXgyDJKnU9w1/kFCx74usckz5TWX+ZbkbsnzF+v1PKMtPwd2Fr
m4wisE65W4RpIzs5nqjff7qq3Sc5Lwn+QG0cXbGvUrIN7j/MK2ZKGJ4qYUJsPVr9/T6yaldj9R9v
K6HesVQyovc//9d2m/kRrzsMCfNENnGyBb2OOZ+2g1Fbh8GhvZtDwGBpNyAGGTPDo+BVJIfBXyMG
EcPz7yqluCaFNUchsU0UciCawe8ddSOpw0spzIYy7GEkuMzCrX18VfXRIoSdFd0OefqitSChV+Qc
JwSBRIfXUxwWNKpK3tBFbxX9mKp+Mt9kPY8UbIlNj4u3Fq7oy299rCRV2BaX68IaR7wgshQHNtfc
v6HnPiyO1Ufx85e/oa/RNMhZNFZUziKtejScTMWHziZzkmkTlMU0hl/ft45jkksk70frYqtEpfTY
zkq7lf0/AJpQaywQkdYiybJ1mkC4Qh3WrJ6mw8maPP+Hq5JLOI97wLOqWEKoBljbmWvXNhD9tTq3
beoHic/+tz99dvXoPT0GvzCUJkMjlVzLy95/ylL56dZkd4pQD3g8wguQVjsg4V5DXtVQnobmdFwn
HP3H870JMl0FtywGfDDAWBxs87chDRZUvciF1ffZGcFM0gDxW402X/0Ygj5EGQm1A9hb1iN0e3n/
r4y+4w5zDHnkiHsfYBlsaT0QLpDs1/wtbwJ9FFxhZPmT2LeyAL6JNAveOV0hjjaP4/WT3P7MMj6H
hVOsNBb/OylWcZvSc9uFOHq6xLI4HLkQdVhfu8R27b1ienLiEddWJJOlMxEOCrtojGhNLz2d6TcJ
yMGMJDzS4Q0mhy6MxpYqQ5aDeDlWd0gvpl5THCEwFRnRqanqBDMyueufKbjZfpM9cAZ03roAil8E
mWOfI1kZ7USJpxxpIFngEHAjvcmQCKcD3BEX2GbcNXsPYDGU5uSCkTWNy/ERXEW8ydXn9NL1KTE6
87losmcpXSBl4NPc9LGaVOmFGK2LgmWWrxrkLCGnFlsr21Dd5p/eXOcEprbBwwFyuT7I+6qjrLMa
AdC9WniEM9Mq7gU0/NZU3eeRkmE2zUJZpVsomhEZH1Il/K7/LZBtP2vT6NTpYTvrGInJQjej3/G2
BiQQxaEZYyT84bEql40Yzb5UN9unieWEAuv43+Ha/Z/I16L7cIcn6i4Czc5yCPRelkoocpS5twMF
ZH8HaKGXZ9brw1/lwyojrwMFQzIrNR2FOhE9UTAabraZlkYyYz8IwW8O+EC2GMtv0mJayRWEj4hA
MsRkdtJxgzze1HdgsOPPlUNSWl6qV3y48TlClVrTmBb+A3FryO9lfif7Ohk+XAqbcdkqYPHMJXc0
jUxt6tkm0qYNCHPP58LblW+SDvvQbPjLb8KFTvlfHTEaU2lpE0iqHIW2NfCnTH3ZvTW2Q80KfYgN
HGVw0LPEneevWgUjelBtsoOEEC174OEvkew3rrU4BRT6QUVz4okEY59UHniwEToSti3nli54grWp
tGZPm/vIiEUit/3jw6Xhyf8UjGJcUkTehdTNOWKudEe8emeJuZfibMfva38ejrDLL6k1YnBn1a6b
MrteFkaNSgnTQ9QsCwHcK5XVH21/Ck2gWpWBleY/amTqHCVx6gNMXHu3kEIZDCJYtGla+wmfYYFj
E9vZVLjTgIxim/jshf81/uo+f1QMOrWgNYq95ZxxwksDjzFoqvDLySieyW+wvMQTJHtxNM7VocBn
zMs0EUijnvdS+3L1AId1venvai9/fIk7I7eLt5HGO/ll1ioy+fbhoutAfyiiQK7gxM+8Ogu/9JE3
v7sNyOazQZg8Sfr5/nm1Lab4Rd7dXZA5HsPDiYzzBo5u1UclTjga8ueBlXBP09WeYMwoNY9zxqrX
kWexrsUzuBGj+lf2gJYjNhtWVLctRW/k3GL2Osq6k6CODmk2DJXgCWVei5uRkLdVBC7T4t6IBx7P
z9qJt07/ZjDbe+wMOiys+MCfxf5dycLDp3nqERv8lmGFC6j9RsTCSL6A9D8hYBav1b49oS9epC4s
I/H+BjZrURq/7R+f/+SiLHYeRADgjm/xkr7omhwlbnGK2nXI/5Q6eJpZu4HWKvC3kCyBplWyYSh9
Q2bx+2VEkDmv88bokflBsevhLFg26PY/1ax+HqIL2k1YRDf81Nq6t0UUxP2dhbXsm8NHPGBTCM4J
wQ+V9Ie8Xceqd3LAO3+wiaM6L2Yu6wXix9u1RAgSQPIEat3fxle8nyHNqoQzo8dVD/Znk+84v1x0
QEYGcGumcINN+ibwhs/zs72UNl1+nMBcmqRtZzaw61VSiZoF0T9BqUBmxs7yQrrOcRrd5RqRgVgV
d+tl+8E5D6+7D25J+ecgrLThZdEjOiguCFmAw6Y0EaZsl34x8eMUkuMTZaoKz8uAH3DOi4aTBhWl
rGTqikDSV+KscYyEc2FJOPS/CrEv+Ez6XmRrJ6wxkNf97XO+7nK9c5NoAK++7Gpk2M7qyAb91ftZ
zSgvJGP3ri9BGaaZdj6noKpgZehqehwordMROem6amT+1t3qE5th5wGo58Ux2DRMSX53/nD9Mzjg
jT2BuBRYy9l9qJ6zYdBMa6shdRajWNv00IKZTupb2g1IpTszFSoYjff8zV5EKoNCuNio6TPdqMyx
DhyaJEX39xj/M4p/0JOVODTYx26z0Om99uztmHkQhsk5qRcJFXHpMZJFk16TTUkhMCVzWMh1RuxH
XJuAI9bo+uCQWfe/YYGDerIKICFXD1nkqnlsfZPLgFvjIyDZbVsRKvNKviCwp7vOJiBKqQAqAJV4
mTteeROPf7ImiCD4a/bdlf0QTxuSm6FUUvT0rG2HqXYrOz/wpz0oTCUysB8AehJNwzU5EBFRg1vt
zoP6E5xItsGOyerg9xrW8IM/VkJYGWLlBkU3J4pOKg42oL9XTBqtX3qz7AZohTEV9oh40+RXyKGG
xms1WBt7Rc5WzHKPhBQpN8iziSG3rNHGMHO8HluniVW9Kt0ByLn/pH8/thY6OJXp1O2U/+QFtxLZ
Ac6Ukq83nnV9ObzGOcZZxG8D4K0pDxnIHoZMWl77z5ON+dAjVZVA6Kz6mM77HSbjajgwtmo+a+6R
IqS2kvNrwrDbUQAmQW/dTwL/Xz+HEQafWg75nhi20kak+P8gAKp46wm4tklzbQheLdj4alzGNj0d
O1IBhOqSlxfEalGubLoN/qBhSQuWFONzjYAbz9Optfi5xwDfsA1iE/NwXKBX8bs5HaT0luj1d34D
cC7zNTBsRMLPixcg1tMWKzgJcEk6W2BL/scmwcFcQpuvlwcrUV4H1vfRxXRXVP4MN4pamk7x8c6J
H5iYQjjj8/iNhSpoCOdf6ojVDza8QhcMmJhfwPRw83MQhL7K7F98jT4klTppRLk0FLL/FMHTG5Kt
3kOx0vB4ZRXOawL3GcgiMk/9L2cRoxK3EDp57OkCG7ZcYY4BAFcdu+QasB17m1R0O9HTVPgEReX3
cHgvMDXHolvGgrJKqGFgfLPP18urJo4cpcNDbD/QpWqAJs8kd930k11qiNBKM2i/ykYMZpBege7b
6XWzb22CwAJNScpSzMPyoCEjrCHN5S1x6Stgib3v4VsmufFjl9T/VzwWJJ2213JuIyEQmIlXIP7R
jQ7GQwFqzVyknLnNW8sZ7IDHfu4eKS1d5yojS0MSp6/icNs3GBkeC2CpO0St2LNdTqEK++5JNGUp
GXrTqr2jancd2dOW+5bvcQNYyjY19rXDEsU7egap93WLEA7mvpV95Y9EP3r85dG77SRyzk1X8HeW
W/qhBwEqRw1rQ84CdgBu9DaOwaNlM6mb1Rr29TRHNqQmYYL8tK2RgXbbaLW4daMDomho9SOKCFzs
l8fqh1SekyQazWgxfmUz9tAWMBA+7fZXBFVRbTOK4LCmfNGJOm7OB4ewjoR8wEyvcBv5cLd7Ildo
+eJz6s9rEOXBQi2vYgZ2rO9EM7opgSaFk22Qw7eLf5xlUDvXiOoshKlABCOF90m/2m38p8Ib9t+E
bHya0dzpZX7FuxvbS27GxOiRQ22RMPrmmQ5l9NIAo1UWtDeN66RTHxOe+w3wgDHkIfkp1Ai5Mpv3
7FquMzVnfbLR3qrzyN1+Nr/9QZn17B9SXnnM/JADDWOdY78mm2CjyvTEPyDosAvJIncwkMMKOUBK
83myGa8VesuZhZ4a8oRtDgw2d+HRgzHvlEGkO+9ai6A/FqgIwp5CxiYCgS3LbbGotqSa7GFuZIB5
sJG6E4Lzk2GF7e0/xLjmEkCdPGlBa4/1pRpETwiHNam+GQ/z5I/8uqAKdaQlfodHMKEZcrksG9Lm
FwV2VuNjjs0GliGlJHJy7bagqXuqrSVOwz2Z98NtCUEqhP4bkB6t6uHAW8NiIVmz9uCNwR1hK9Zj
/Scf/g3+JcKlI8GXDA3kAqrX7e0+j854Xr4cqZJ/P78k/AkiJl2kcDL3InfNf3mxG7Gni09+3AG+
0GtixUtvRy2l1u3tW3JEFSVMSTzXn0umkvsJ3Gmh7L7NWJiCE4tVrYPTOXglljLG7yK+ncslAR38
UnZj8faM++13cc2jfb2+wBw914igPdDAzHGRcLsFU/6APXQuEiS8ONaE/sJzIqLL/Yn0MV1WON76
a+POJHgUQ6zZ/tSzVjF3BsyWo3UkWvXA+MBgVDHgSb1StlRFudi2YYkLCQXogQEJNYl278MYl44d
GCAnanu07khU2qhK+Ap1pJRaSKVmr4bodA0xqlEnQFkHaiKg0J8oGfnscVBjdkvo6dfrAaqiGIIq
RNEn6+5ObG0Udu/5a5A/Vxm9maeVBjCrKrTxIEgReuIu7u9hNJtZJcXI1DTlczUQRFFyUKGWnC8b
M0sW8oc3qw9TXOQjUWLfQzmEcCknQBkHwtSR8Q5RHnb3OaKqBqs7S+FFr3kGIQ0GQD6dOssrN3qn
NefLEp4/P0JhR8d5/ZtgmppHVT/6vW49hcjJaMX4hHTqDN8DhpfNUmjoN55Txz2UURlllVaBwkoI
qChwGMMbBERNv6Ddp9Sb4e6dZs6qlR0ZLKazbV0q3ICRydpExiYe725Ku8cDUec1wzad/n+v37s1
HBl10LRrWIk3gGgHjI1LjRosOlrEWVhX2XT7p50KmkLM2IHld/5o1JWTHS3SmW72F0GFJgYWhLRE
XSA95cpaBJRA5StIHbYWuCa6FhxDCkHNAAbQGxZR3UjTewb+9bV4Qe7mdlxCMljvNJYeFVHlcUuu
QIpnGJ5/B3SvOPiWEG/ozEVFiT0F9BuFESXJhx5KRAOOCt4d0XvDSGHIcsLpm3XdMLkTIyX51y/N
4XXwRM8YMZ3KGkHPdYq7b3jSxMonwuEMlPI5bNP34wjhNj/3vBWDk5WCz4M16Y26dGF1vu1HlAxl
eYzpu8NG9+Ruiwb/H9bDUfcLTPFXT87C1aShVUdREQb+zHCS1COujAzbgmmwI9INTo2muJdwohHL
lrqAhyhJB1ThRFqyTQDgD+Iu9JRxuj0KwlHoJhb4Hj7oNTifJ+CTind/wuLEM1nl8ZlecoVx7c7P
Kr43FPIX9HegizrX6hojp+6BsKh/dxmbxOZECM9rEoABMNID4i6+7kRkst3jSa2swtSa6Zsxv0dW
1G8t6ml1iFsry789q58Hzj1FaWx7lMfYsnH9t/FpjewboV0OaGyGkzNHK1GxbCgzQFTf+cKElzkS
lur59M0rWRuiAWtzSD4AWtKOT1dGOH2Fixkj372gOA0bCO1Jwy24Af9WhdvHk5/sTCWf/unjLrzw
4GkVb695GSC7BGGzUK6UXHtKX0/L1srMO7n0xFGfgY390SaWRU3c5Fn7gE+/8rzg2pWee+WIUwwq
BRP6p4DKQjh0CuVDl8eUUOt8biiFKx9wDGwLVugrU8GfUaJiAYm99IpykBEGd0FAVgkpZZ0LIYL/
sTG8jqKDigy6cU5bn+Du7YB6p+ehXQdQQ4pr2DV6hD9mAFV+e9TwD4NiF8IG9x67HKaIWmsfOb2L
sWGaLcccsU0kV6HR5SFjduqt/k1yjc/E7Eli604awFC+tLLJ7/cRIVS/aVn79VL4I/4fgu4JyJkR
GFkUa03R51JFwo0x46mjWvCnegZDW3F6YM+6TKJN+QhnI8fFjGkBUJzTki8AyZaowlfBk84gWxO6
Oy/2pU6ApGVmUds/jMFEQOEHhz/W/tgwxTXlPYcbz78cEULdNarV2skEMi9OS09Hv9BRVcHx63Q9
t0t1WIvffbbDH+hTIRH80CGqA3R+mrvoB3pXISm2q4e41fRL0zkVOLVQ/r5WadAN78rX/DBfSIWt
J5po8Db1qOpIqdu2thxaZ1WZeZxBIwyapDwqRaTjQ1YK2YT61EuXThn07rrlo/+1nXLQspV/GnMZ
xNa0zBLQi2TfEnyNtEG3UTbvy2AF3poJjKipO4D8nx7KJA0m5LP9AddYz9YbMss2NsVNx0tbBRRg
fq60WyGr9B0vNJTgY5RFYdwV6MoFO8pQWjcvCBfsND6O/DKiE8l6q1ZYtvtliFExounwpS8bGMFf
yX4BgvgBNFMLuPH6EZZru+yW83zxWerYHIkLz1ad5SrHWWk0ShsYG8lwFQswdo1m+Po1mBxZ20ig
4NQBr8LxTnHWVSnZR7Cop0M46aiRMLYU2vTbxXjDoOAcXZlTUs0yu/do2ihes8uTwUUYXApJCjCg
weadQ10Dy6GkA7wh1npq1pNovIrXWFrmqiMCbNxaWRM6u4Miz1ettt4WAU6CTtoHtYjna2V5bX/O
2rbvJfQ3nSs60Hvqi31bRGmAFnQeKRM4wge6dgetkFtZxrYOcpI2TJwEUT6PMdculdkLaSnND/g8
p3GE6cLWC61Z/0d8QQTFjsxXYkpM96oAVjRao0Ws9Nl/GBCLHBPSk3Cp0iNI+KX8DfpagMK1MjsE
pe+qx4qBJHHY5kqd7OHehKazC3yzbQUzFLbtnDAKBqp+KpyKERKltB54pwEHxtjL+L15Op5jGuna
ayEh2GeUJdCsyVuv1ykqYLeGoAxVvKsctog2EJw8tXTCTsmlZbojbSWeIHoxfXKnvw64Zwgmim8i
2dtk7941qM7qzVlqM0/Ejwx+etxvT6ofF6Wj2bDP4zgIuprJlwtlIfYka9YpE/qVZCORfTwBbAMA
uHcMUM8R/H2gGJOUlPCayY+eal2vOlP/BeBANWEzEuwffDeWdn74wm29T7RhE2PbBWZi1oFkUNzB
g1130pfcPajcuyKIq6NUGvOdq5VlmbppWPKw1BsAJde5ewFTlokGi1tQsD39TLv3afJaUZpZ6unk
xozMVKPhIzfRYpSfrCSw84YjzJK0Mu+dTZtDFJi6dMTcm31F1YNnAL9bxTdI7YJ7zPUhKm49yc/f
boPmf8nNHgt8ZhzGb/Qjzc15bjsrGOdictwY/G+IB/Dgb/BMzKAeWeykh00tH9p+omgQBAjbfJh/
R55y9reICd9Z8ETMRQSvm/lMLwTC9rO0u0Qv53+U6swrWam5MbylpdXI8LWRAjkZWXhfaqKEiKZx
SfGFmxZTVKNdRNDP1KNWh3IcWE/taJ33t183mAHXwp0i59s8ubz34rT8iR3VziqLgBbpVX9WT90w
vEUkCJnt6/benI/CP66oedBJ8gU5dd4rCNqL5CwimIG3HW9XXH/G+9IhsXQpl3cosxNDmdm6/c15
SXWtebFMpVIMeTJwBbyE033qP2yoo7h3PhDlSWqGLY/cZBSWtlD8DHXrhIs2eoUCs885/Cu/7Swo
dSVa9cRgyj8XPy0AwpcVJQ+PmZLZGT0K2ZlzUDHjwNN827dfo4p4JufgDgNvl+XokUBiA00y1p2M
AZmrxSgM4OH6atj+t85+zaVpB3322dUZvuunIuyerqWPLf8E8vrsoTECz5T8BHXXCb1lDkzbZvfw
fXb3jlE+Kky3jGVrWNCmw9i9QwYqeA0/G/PefevqgVuoQkZDydzBH4A3UgLoK0tX3/gyfdf3QNIU
nnLYs1PNxufqCcxSj62sAbOV1aTkuxi6blJ2+EVqM02NRNT4WIHccfUdxGcDPkaG5HjKfgmKNb/t
J/2HO/VWxWhUhiyH3hO1wezv6CbAuahv8g34/lADR6HQC1MkRToOTe4yoNpwdmolZN73uq6AYEtR
rpYJ9bi9Lw0neM1sEUCOHSMqsgLNlugRfu+elBn8EHJk9k7/SAhBa3oQ35qMJRO54CSJuYFPLTh5
NZRVwYKYiqTgfpU25cOC0XcyoBBBSyzT7tOyIwM2vI4XQzqwZFT8m+Oyc8WP1lKQ1I9AVftiDl8q
MPpObUGzS2KqtM84c6+cZ12avvORccvanI3FLo2wLNhgM2WDDky4oFsjj+hl41rkHOuU5JbJGD2i
Co+mnr/LAhDjPku0s1n1lKb5eVf/4mdVlXIGfJZ+vUJ+/UUYxHCDnJ3RzUfFgfSw3ejP459RKjwB
m8VaTmVrY/8Fod2K018JYSYycWcUO0zVeACuR7ucW2e/FVqesWKxD1y3seLfco0aZY+6JVtnJt9W
Kfh7eo3ADK59iV53X6J4wCznr5Bds5Ov9uTa2EeLyl84lUGbH5DF7NixN3GndcfxGHPT9564CJGi
63tH+050epF11BpaJAiuOSPYHLaEXbLfmKTIoBzQTYDC8j/PU4Sl3rZxHYcq6g75UEekBsEAuvWR
OHFNQjI5LSoxnj+bUI5KgqcHpcoxobzdeEhrP+XpxGKChDKQBIiLlBYlxRnLA+xTtM3Ncmh5D6z8
Uzqmp4mId/8N27UGL0VcixfBNeVcl/QnAKsKOuCPMSA0alxzMJ523iorAFCGgOX7hQVvgh3ZvTAW
PSIr5pstLs0dyY0AdYtPwoH9wx+ZXqBcsJ32rK/1PahK8wjNcX1qilagSLZOztkpNGTgEy/auAhR
zwjdpmxi5q0H5snU0HXLY/2YLhAqURvux6GjgRvu2buNisaWwlZFfdrV4vq3YIZI6OfsQVoRqWCO
hhLNcSoRHvuzjo362CjAX0Y2m15GDBkj9d23YgpIKZnAIZ5UbgKa3Wkdesk9r8ReDWdxU1E6Ur1f
8yhDigAve/tGLrj4ahk5Xpcj4cvSjWHtZPKt7I+fEKfBmrdCBEc8OwJOuaiBpCaNBWDwMTt1YfDn
wbzLqQyCNqBLJh5Id93CpNSJzQyBYa2nr//smGtnM8F8KSw4GllmM8IT/AHlxa/JiZwA0m5MAeTZ
yTUrsrg6OHvhmfndoI2L8uahHjbZfTXX1ayXXXfTzsS+0RMFh8dlBgY4UNlKbC+ydaSsOBVN4qsa
YYgYGHVd4n7viDl8QYFvdIR2w8y89GpxGC1/XbWJKtblEsMPhsmFlI04850o3Irk6gLCRbKilvKl
vYGKhcSFUkma/oln9YJhQCOk1ExRYdwYjIflUdQ9b6xjCQk7/T2BtVw2XYvM1UdbB+SxYDIGpO0v
GSI6CchFsOQ8JCrUogB2eRbaqx3ce8e49cHlMpJkjp3w+GD0/wgB9QT4718a0JIQIGAmy4ahnbcK
HPEpcAdmbA7iiaUxHwBJ28VH77Oe4JlpxLyYNwEJhuLRDJEseIb90xzmSqLkWuThfVNc0dEiEexy
99OzTzQF9GKnVNYgmv8pWDSXT40TjaF//m9FMq5my8qVKnmcPRAKDKttDhuxpNwSpoxRorG0c7ck
/QiQ0Z0wubGAbaYoUW97xWqAmcwWuN+EVLJXDHJ3wEin/RkY+hhC1aROVLOBfJfri+KByaxlkakp
3ee2ClYv7MHCu4ec0dAisDXf+q2wStiT08k/HNi7EsMMb/R+3JGbWPXpOeUjBpE4jJLWUi7DxGG7
6Vuo6TT0Dc1LVbnXr9HCLY+3kg9wqisnGAOVA26cYL8NQ4Y34jzS0KFGLxPj+ICyBi/+No9rqbVT
WdjObDD8WUSn7zKHlowKu87/ZmznPmRw9pkbAh7IcDMMOdVzEvbzl9W/lJ8vJwQe00wGsljoEsVp
Ely8bZBc58NHwJZf4Az1Aotth7oGWQLnX5rxdeDCqMM9fhZw+MPa5KzqspS6SpnwkpNhE/6tou8p
ymqqUJhDjIukISg9maiPXV8yTvGC+/sifINM3Ucecs7Y36H4eb4Z41gqDyvyWrx3cd6WhpKlzmbZ
HaNI2J1rks4uFt2z3IYYimFseraWOTjmuElTZq82glxU/rKa+oomFvvaEKIVyLLKaInMgiwJ4fE5
nzjkFHU0Tl0jau+UMiXAJP8emiv186kwKTxJDDB/vjD3b1Z2/QTPZLnyRbhFw//L5LjcPz0v4BNt
P6+5vAqO11x359BU+h1YTg9Fe7WSCVqqcSHsEvdrYn/ikX8Hl8/X5zcwPWmEXGq9KiH3drJqHbhb
yOD23HVax3WSflgcoDtUvuOpOUXvHNPwDqSMRo9HvyJk8mKTDRD+f/zva577LfL5yx6xPHEaBal9
DOQjWSPvK2XpuzUm0qao7dKm73lDetfgHfn9X9O4cm6Jt/u3jgEyVvLvCPsHy6TmDlwVvxt9rdSW
0DRloN/3dMg3d48V3ARIADfygJ6BsnVfI2/Mvprr+OkKBuR6SPy2SECLSB8HGqKGXcpFwLnFvuAb
eEtK4aodODwFqd0J3gE78cTyiPgoh7+bEclUFzmf5TPS+opzq0QmSJscvCuVLCJl9Nrz8TrO/0Yt
a1cMn7tQpWdtSZHx2hMCLcp2C+rSgWzU+goaaXrs2O2baXtASH1WBMtjV3sCePobWH38Ea1uFNgr
ORSDF8yOsh6/Pl2LfUt3VZTCLgOf7cWgRtXeklBOdpWCfLVWs3zlcSVkA5FRWWVNYr1pBdtPcnjg
VxHGszoAcbrjZ8hYPvEYFUoQ4dUkQ3vcH24cTSmD87L4AkNwYX3225EjXpLUTnHeNmSpGT4V5YNQ
NnOYZ8GYzyWhp0yiqaobNeh46j6QIgcUPeh4BuDLiTKLQDaygrFGgjY4CIRN0AKcTe3Jhf7rNknh
hBBDocwPQwm3Gc3oj7e8sQCgXOrFsP08p5OZ519/AT7dEMk4ytyUUuHeIJOu6QDkwQyVyqAFPEvF
k/uCyYzlKXdUqjAlgM7DhSD7OXmEiy/sz5LpEFrqLm1lDcvEdbT8TkvrecRpmBmq1tqpMmzejux+
eDJ1T0+4p2lLVlMOpEEXpPDfwui57NQ1nhecgjWLWEPa+oVPKZuq50F8u99DCdxWW0k3fgp8jxun
QFtgK4pVMXa5vwpBxXy43E7Y72WusapIr7+wr9NU9HIoPWkEvW7TPKNeaEr/Zm+rZUAF8kJjuHno
uersOObqOq5ZRkbxvEKFHn7eCbJ8x8UAKvayK255fnIqnIE43/5iHNjWlz92+03v+iIqfqqacryp
ajgWb/TjSsSiM2B0uB7jnpOV7PsMOvUzSroflWJEcn8523xjOSkz4D0OKIo9mbuvvd7b6x6fDZLl
gBsvSESMcJM9yx2tQV+3li+zQbnsD1XcBOe0sqadIKcATMs6K4hdglODqcewjZ+hV5aD7RPFgu4e
IfkK4DoT+8gDwTRu6/7yqqARYAL7fG9PXcb76GI8kX/CwZSP9FKsXiDtwdckiAtk7pKL2EHa1ugv
5UP8GwKQqhmikoXzVCBQI0wiNS+TSVM6NgaCpj/QJkUzqnfJerkOdDDm3WpuNT1QEGc+OV8xzbrc
Ks2hVwpYxS2UvSLG7fLwdMa1h8A5vDgSIUA8rpqrkjqRE4db57I4SwjSB6h3Vgt7//hzGqKV1DmB
4wW+hbCZiigT/M8FOwmboSDaHhT6f7EMkv0bQh1BITUJj1O3JjliZdFP/mSHByBT0TbHvlOQ6xCk
TNwAINga/jbBK3OtEFspy100rlwjsl5KCCz3V3iOIwxkRjQif4uVNKk40V3EVjJNHLiomvYWscDq
Iz0T4Gtx/FA+oe/3HRk8hThfsdB9aV6GCMwQFDq5hlytP95YJIgawaHrbz8TuGhbzOSKBl2dZWN3
o1LBMsLayo/l+Euxipo140SOokYnL0UX0MfTkb11FDRV2VH3e+6EXMfCNbX+0eqthi0U8zPNmtSY
VR13F6VCwb30CHSuAv9F5LlOrBgPokSqJMwp8z4I6Dszk0eOgn7bY/7MAnrnxeCRsd4+0mqA6TY9
p70Wr4enIxVvGiDXe5d7b62oi2qofCrWxFEk0P/mkcV9INlOegYbTAfwJkSaOaHNHvevDax5KmxE
7DW16QMkcbeapTDlbgmpcYBMryaNIUjLQKgjEyI3Pzdr5BarlPJnPBMuZ3lb4jhV/NZ9t2mkHCn2
Ph5MkPJ8JnziDnPN4KaBhpBxM/jwxOxmX9a3PULPc0r83s3tIE3FMoTaLB17BE9XDaFsUeFOU+rV
hVRuDwzjaTQVJawxJbpjxhWwnaIvyjspQQ/tTHMnS7DtzVT4kw6YuizeinZy3yI5UWQMC9lPhgMm
qlc8KEX8tVekgITzWQ1G0E4LMKFSH/uTPO3qSMHJysH0X3fz+REVx9iiJuLv8+2jz4p79moOAG01
3U22ogz+5wMXWQyD3ezaWel381R1SuPHxBJk6QYMO12HOVPbVvrp1NRJt+1GBen5uf7Ft4TNRWLn
xXK5UhSSbtYZ9xa+kIbj3uO1mqcXaJsieTUNMcnn7zybAWCwJYkULW2YAcnrDyqELR0qv1vr9sLY
mkt2UwgH3Rp7fcyTaL/88RlLQajRVgXEdHfkZliUpfIm0Pg4TPQQWyGcQ22U8KreDGVtDtnvi2+M
+jHcN8meqkIVFHpiEkkkQXqkj9YbDBdMVKcbpJFtAN2ZwuCPw3dKVVNCZVmxMFYGT0QeptnM8jAu
rNLHMYWpZ8Ku8/hgowWdRYG4zKadwFrRURW0CNjxb7aVMVd60KW13FNItyHXqMNdkedmxDLV7VKW
VXJ7aDUVOmL9fB1f/3KB7/CActLmwviJEwZw75E3vahTe62Kc/KG2Sbp/Ccv2GXdQsIgZGLmSwDO
PxMrl6BNRWdV7v7Om8d9gGjwojPTQX6+o99YolXXkj6qE/SCq/nG9KeuTR6cDxhyTGgSjCH59fDO
nG2zGWgUpiMJc9/v0YbXlTr80n7Khqh0AlFihcrjM4mGTJuVUGyExDwXk0m5hmFyy8YLxetOOipf
c5zxIElvuiuABPMsSJROnicjOkauwFazW3LKeBprwSb0qitAEHMFQz3P9jJ/6dUGI+slu2yH4VyX
eevfWkZB0PtPzTkGa9MxrECAuj1lZx6sobR6S4B3SGmllZWM7F+I13mHOvVnB39IWab0CvQqJiCJ
0aW0tti6LoUXeL6+FPw9Jfpj4Om893JEp7+ujoyQ9vBElH57/j4pkx0RCBoDiv64Ni6jp6vsmR53
0tIvqvvU7FzPtrM4AV6vA9FB8JxYzsJjHE4q/TGjPzhtJrUYDZ8p1QiqcQRt4WSqZx6/dvZcOEU3
WLVUyEOQb9QcowSEp5VA/VWbDknK5YRnkh7pZ1Kb1GXMneoXslfM3VVE/tA/vXFksGoz85WOMAtA
96XDM2jDP1HkqkvoMED0ahna26R4ypBB8Gw2+sS1Dw48iuP+tC/4xDKKWnHjdiSXGzl4tFcVhlFN
CZm2PgUcvQRw+AVgQHkAMj3gu46LP01jkT5bCvPKl190MDLCTvczJPwjliGP4cqfBn85W5SQ+2LX
VR9/LGrjKVaB7jLHAOtS5fD/q3ODstG76H9zKbsVGUgf2DyaeeGIgfKrzPaKG36HUG0ZHhhcQo4y
FU78r/Nx4LmW5ZeJx1zO7ABh8HBn+jCfRuhOOuataX68iMHf9ZLruPIZnRcqtkI86YLzDDo2L7uR
PQ/tWZUKlGfV8AjKxZFtAbYnQw09c86t0+wvh3RCc2lxzUnVKMglyx+GKNvlGPZ15MXmgd6KEbSG
Iq33DZ71zZY2ok8B6XKD1BWvz3qPgPk+VOBxXpqTclha9h42bvowHJuKhLWmLI9fer9XivE4Dvz3
6qFtRiR/mLskM0Yml/p9TbLENUUmRcoX/QwWKnf2a9c3BT11L2yro0YFqxXJGhhUA5PSfdBdgDJM
MDLKsEO7Lp9uI5a026GckYmC/2NGzlJcb0ozElDMvHZBsLBFYzO07OHsARn/ok1KTt9r0gAApjr5
akBmgAUyQ6UD67gCzRQCE+yhWDlyGD/2ngRkgBze54jb13ru50fshUmytpFL6qGHNRLepsEhts+n
QXIJQonOdCA/7uYI6pQT5bJblxLcR+SCQOuhmK2GUO4VLgz+hvxQJanikn93atNJxCiAhEf59ePv
+Y9qdPruP6dCYv2lw28jpNDpkY/whO/DbPZs4YE4lNkGwBxTW27I5MuFAiZnUiKOTApzhGoHi4Qx
UYIlad8oD64JYfd4ca/mGOqXzfUTBR/UwnnsUEG8SHd08qH1iDA/SUckp5jy1V5RcAtVFgEif6gQ
Nh9UUxTQBAdps+KmH/PL6Mf8zOCYC/NRdvT/WfhJIZ7pW9LPeDXVGsHggbGl/yCxf54yUmU6bbIp
o9q+1xwIcpepLz+YhvzCuJvw+MUkUKx33TqrFSYu6l3JAkY1xcPgAtiTaaOuX36g/3oUtBMG9/QO
uJzkOJdlA5OG6zx5YCn8aVJXWr3Mho70ugORh4wtxxMp7tcEnf5bjs3mJmaY3oy3VkgcHvG2r5y3
FD/ihjkFGHZDSFl28zcvb2agXz1S1BGMjTm6LUBeb6CvSntvveYZ6jIW0mKlCem6uLCa+mKKUeKj
F6UTHY5g/93p3RCroaNxpwIrJgnNV9z8iBQDTRjcsHBGrgZz9BmzfGas6HIjTz7/Zn9vEIc+DKFo
SjZJNxj+74DqTuXyt4mRP4ZJD+U/PEQ4LaWQXk2xBtTr0ho8Gxl54Iko8QoShZLIxTwFEWgzB7fr
L0qunOsBCws3oUQbfmysjycEIsaQBc8HeQuXkLw/VIjfDt0NaH8cHou3lDUnGBeauHwSiKHzva5a
UQanyUn0AxQ5dPaVfHB8O3xJdb/y3l8rPtO0IoVrv/gi3acvX//I2Jle03pvGP1DS9o0PDa+tfE2
A0npahTsjKIaJgxzoBcYAPocV8HunTbmZ0b8XCik2vdybbMZ7kU8gIQUwBrde1a0z4VezM3qSAz1
JYOR0rFZ0psIUKwn6dAoGHFfZ6B+Moq80lGQfgrSSgQje4M2BdSYCSIU59R1Swj4v4I8l+WIk7Oj
pxwiBHrhDA639acoPvTUZqigtOGL9CUl+wLGmA8yxn8FxEE9w3gTXGE/LESmJEqKrecmJCMYaHuJ
ei3oXSoGQKQst7Tk9PdiT2zgdE6nNZTy9e+EEFpmZQ4qTEL2JQ8rhVObQYuOHV4rS04bEzAk48Wo
0qBKB2S97F7XjmGb8NyAMXTrssSwQHXu+kOOofoilMz6gwcBEQBLhE15LlNpoV+0wo6PVGUQ7w3J
GT64VYaqWTV4Ee+TF5TSL0bWj2ZQUXp1NMyB6do62GCGn3UAh9xNkMAjiOCejs5lKRq5Iio+O7ha
t8QCQ1fIvlrkIi/B9CudkmUuPjMceVGtl6LQAbQRbTbbS4s3/rRxV+LrNrblh3AShitoUasrN+37
vIAsRjmjlZXr8+umii4D6D3bc7XIkLc/7mYxsEl0VrjDmaMQFv0Tx2FsUyr70nQ7lID3FCXi6xD4
hhZ0VUsPIRlx0/HUAK8l+/LskG27R7qmDQP5oBfhBqRfDTqizQW40L8IKCaxkmL28jkkjCx3dvk+
2RkqRdebKH/dcC9111J3BKcO6gEot6HutezCnX/qSUmJHtL4ejtFbfqYY1Y4i9ETd0vKBOIPVp53
j2BqW/RyWChmw4agCpQdby/enwTHGd8VShB/83MveRzZTzB/3sc7OaSY1Qdr51XWytTrAd7zWWFf
9O0MTRtTOCc2XA+bIZKqeDCcNv6sg4YnQNTmERReYjzzDsw6Pe/lUBVuOPEo3+RGOfL/aRnNZJS+
yOtT05EfaKXhipezfaXPfAVV0OO/CXK5Saq1Kw1/9IrmtusrWsDwYuJrhvf8V74preIQ2vguTR+X
0IqmKxZD5+0Vj7k7duJjgNfFk6tEuBVlr9GDn8CfUOb+umZMCIK8bpynWB2uVnRoyosy5Od5D+Yl
PKx5RVH5p/Bo1dinNnie0OmpbeMt2J7H7Vs5onA7TJ2fe5uM45uRk3tc+7T5SY4Tw6Tf/It+dhir
cg7QPTJKul3jyT+284xi8RLWVL3XvMRG9DNJcOBOJmPxSpn3uxmA+S3t6rT4HyB3y9fZkjfEsw9i
72x/o6xRDAba3ibjLNA54CCZViu+H2mlMDq3tZTnaNoTbw6UTCu8T0oOt88ZFq9NZRA1YSMA5fuw
kDdTp+A7MfLYsKq0IggzW8EAq6jYP+2/p3Cmz/PKIAy7y8zCP2+vkd8YpBoskHGMvsqEbin8z+J1
mKlv7eZHv11hEOYOXrNB+33L5utzNwRPUZUq0iXSDM05HQqTeYsrE3Ejq7pIJbdscjaV+58doyDn
HPkTcARsg136GwjMQr26jbcmsIS2iKZtT8ONAPoVHiXoK//ONi4MQPyO/wLWPsc6HHsHrDzaOHl4
8i1lKg43+srIT6HBbWdFhaYdvfDrc/26RFWRVIJYazJbOKn0WqyfkFHuaHoTyKYIqgoN9dXHJ2eb
5LJZznqHzItdqqIXOlpeDRN+9gRfeqPaBrn7vP9b8Yb1VAvkwOj/UzO+aIL268A/GU970XesdazE
HePQejZcB1++gbOyHUGfIzSw9En2WpevY1TRxPWxL86v4tm43T4r7P/0BsorW6TvW1bWt8X0dUD0
f7dkE+RNfr+StO7Y7AtTyTDqS65ndMEzxYesgLihaaWGJ6EbCs/oPJw9FlZ+TxVnBqhfnUB1RxFv
zAdRb4c7Hhsyb2WUq6kZ8Fi4Guz3nJtc8h1cfE0FLNkvi38iwNRhndNcJbm92gFk2NEvwER3tlTR
P1j6UX+xatGjiM4P6dBGuGqzzsMJ6RiOR7wHq6g1chqERozgAXIZIVxvsFxbBXFzUC15zhhFAkqp
RHY/QqAabK5akOfznT3haa9hLIJn1b1QDl89LewstwRBNL1VxeWUOzNM9XeAr5WQM6YU0MEGe5Mo
Vh9HCaNfuOxnEVzsV2egJmsf7SrIFYU9Wyxtdie6D0jqWpeVjImcfK/qtoRSQLUUqABN3YapRJGa
jfx5ZA8PF4IR9i8oC1YOQ7zNpGVXnCQRmE1p7G6nauVY/TNvB9s2OAEa1wiJfOUriyZHFo3mPSys
U4c2zsDOa4tObN9llNp+UNLEWatw3lkjKxZFqny0rH+cHdJFUAHwpfKxXpjwoShJuy0Azx4VdedV
bTtrzA8rAJ2FqwmIQIAOoyVJGmSyyOqbjtemtwecNbENluy8hSL6MW6AH0rMD7hZYpXMwMf5g0BT
G3rMAHb/T2l+SqvcbiLa+Zh+s2VVv3qXyuBDhzFW+AkCVWGhhp1jKIEIugJNLrLDE7Po/zXQKNWS
9RX3CU0E7L8elSSWCsB7AS7Q+yRmieRGI5mQcr9TAIlzpXHh06dr6DfwaEKrRAg8N6WcIVd/2nLj
bXPSU/mB3SneXfpkgPa/X9XpDoHvutWxn2484YfDXLH+48++ZblNZ/AV9lPA/zBUBzrmxbrCqJru
fO3f4x8gwGSeH/K0hbzsKcPO6wQg5Qw5FMg7GNBv2edboPBCVBn2WChPLO3cMLrjHlKnnJ+E+0EF
GJHdDEKAfB2uv8lkX2wrkei0c2PfbtnpLWKlBvXvFmqCiXk20WfkHrb5oT9WxNdba0S+ZRG/SiVO
2x7GAPBhBHh8K3rz8yilBC1F5swkTSw28k3V62FwRvAoEb1+94yUdzUB41mj04nRC1jasBzpOp7i
p9r9ll0BPqbj5O8pEYx9tBmY5hrXEnhcR0h1NTaJGPI4cc3kGY4Gf3Wmg4y14Usc62xuXbm+waTM
N0Xp7N85KYICBr63VTA2dxOMkNgr550jGsJgrZQcXT7TdWHAdPb+4i6cLrp6LiOnmDwb42ue/QL7
Plv4FDLuOw+3A9gncGaplWU3xfD6w4M8Bl1piFTtf/rZryqopTUjyDImkwoiDyuAQmDq5rZt9Dli
MsMozX2xIqtJDgTcvEojcvltYo3ShZTWmepWFQQdeiVX1I6m7JvSyHZ/2A8uNxFokUM0dRQ6csSF
utOMPdnYJhk7fbNl+4OxDpnjPgHMUfZzPiD/5S23NMZwsIjveXDrICG0Y6xXMfETLKXR5SrPwDLn
ID8VO+Y1Z//IMXPx8esv+foabOo0h7hWo4fS4ePAby3OEJwMzU5ymcuKpkNBUfSOBuMn037CV22V
3utjkhTx4kP5emndPNlyTUjLggW5XwnwyjBm/Gzm2gKA1MXL3E5d8fK7xhSqc0saqU0a79Dbtxtq
vbsHzYl1ZKIx6vYr6RSlOEpKLI/7zThczh1RBbnuH7OotpuVp6pbUrFBuOWFQacdxYmFIUPj8bl8
9YW36qmWM1cJAsfOSPqR9JGzmCYHxs4UN1jh5u+yr5+xWTHg6VsXXjSYVUMieaDSQov/VllA8EyY
XgLR8E6QqJuCrqhkA3mxcO5AsOJo6lb2+A7ZlZZljiV6OpYVp/D0kVP0mb8IvXTxg+OSl7ahvWEH
Lw9CHztGlC3fCYlMGwXG4vYkooSFHa3f9hTtSaWUiWhe/UyBIxDQfhEQZuqZeNQVw0YA1cPlY92P
MuiHH0mp2+BQb2umG9wbTGPPRbTtbx4I6moMPD8UID/0r6hZ+wjlrFFvK5QDVLdQ9XxHFEigX2HA
6L0DxesT3dVMhbJc/32mpBaJ7tnlSYjb8dvBWzIxkiJEiBrW+aeOvhC3aZUuR9UGqg1PjzqXvQHj
LdAfMpiik5v7dfCtgNyTo6+xiO7MaWnl7gZ3iWt1jVUoi3r1pDVbJTYmM7m+OOcAhYbr3eLNw722
qlcj9e9yw08nexxeAX3WKVKsnH9kIAAdLdYKUjqQBbP74ouR3iZmkYcX5sFqVRAjZYjRrP3npfq1
PU31TWfaTbe66+VdybIv0MufHBKK6/22wm+iVSKfeRa7ic9CrVgV6PdL1ry0QdVKFleRZN1wcIsW
WunExtbzEHj7oLXg6uMrIj647P7XZaCTzW/3WYrunBpYKV5UPAxW5opFvy+kF5XHk1X7at7Vuo4W
g0BIBYpPpCi8Dp9naVQARQ4TpVq/ioJ2DvU+Z4bZTX+nifvNDyclmNmPGIrCpFXalvS918/NQWWM
eBtTSWWH2e0jb718rEkzRr1jOnUzb2oJf1mZI3QweWdqfhsnVegX0IG1Lj/pyOk7/bKKJ8+6HXQv
sChYXUiF+MrOANGyiRa2lXzdX0HLE+WeAsfTiTP4781yLjF31+YOerApUPG5CYBOeN56xiIkeLy6
FydMxojA0wcM0hcFu2aLNujR/UvZrkdXXHDzu0+1c92FvWQGbTLvlxRNXuH9NI+jSihz9M3I6o66
XyWKrUP0x8Jv1dyWBNorlehoxw1iTS6AOqRbf45H6pLlhi1Kge7K5wx5TzkTdpl3TxP4MoO/kAdS
I43N/Xe3787l1fynpDrLztadbrBkK/FQhUBkCqghBiwQfsSEpp7L1x/yQLgbQGcHowx9X3+gSsim
qaIeenlypSP2r979TTC7xE6Y0o3I+p144eopiLsr5K4ZHnu4quuyAgjiklC29N6GLahkqdu1jBIx
0Ab5XSyT9YwyF8nLI8BbOw/SkbKMyFEmeEltqMJA571aajtxqBmSQ9ZQPBxo+RH7cbXU51eCSNo2
3Vorwl6JLN5Dsx3uUZuuwOZNECTNgrma8gR2kbxdgZfeNA1TzmUGcIazL83P44ssu8y1A3XJRuO8
Z1SZfscimd1cM1NiwO3z9AAnagGuFIG8gS5FANyh4qE2dYZNN7CaVUG7iIV4GmYKx4JB2mfhSU1O
5bZNsgvcm++lEeDM7/40nAjiqpLgFWZUWNkfSTn0cIf0CmHeY0a0H1sn6wMZvy/WDdzw0UxiCl68
MI8ffxC5RxKgSnhOsDXX03Uqns3Oi0j43/Fhw94jbexN98oTShU5xvoWVpKrpo2OK8UJYT8/Im6t
beQyej0m/yed9QcvLT+slSCVW0+IuXJKDKUsyp/yxxMXVepEZ7A9hKqgLIopglHX990U5Cvcw678
5H5fwA/mCQrhJ6kRVgQDNethyc2s3b6pznQVbbmkr5xq2y1jOgP+0UWSwMQCbbvAcf02ckhWqz7k
zIl3k3vgT9GHgZwuGTN4eHevb3VGjF0m4fSpBZ8AMaXNd+IrOwhRko1XO9xxwMm5SxnIUxFjYjCm
vfkKnf5qjo4eMtYBGYzsof5hS4vOAIhIGFNNGU11CaehTKPdpaopp3yrejD8+bgncAcbnOxy8KrE
W5d3Tz6YxhmV4ggdFne924Poe0JVyixlfa4wfRPjkUKyKbDVFV3yYZLPGLGvXLvG69coihrBi6sR
7Eggxc6LXcWfWma1R1QLQO/5QRng9VQimLn+4JRfss7rzCLYOXB0aLQR7QH5be75BVvZUWs3jX9M
lt7Md4FMWtDjJoxHN02/thdlTALk9R2fLha5cZDTETnhecBI4jYA0Bp29npkaUuhOfulLpb2Ab9z
Kacl4wpAp0HXYUSKkcl1nbsjjaJ4xuCi8d8mRaVRKTy7IN7m1ZPuoL4VzGtbqSZ/z/FDmOXIvUI8
NpB9uWJaUU3MM3tV5um1WNAdoWJhTTZviHUmUBzSGFnVGjPaALeYcZRKrY3IUl1zkuZRzaXVr0qO
4e7IahEz6Jtjgfk49zmYoE8qsD23DWll6p4TO093iZwBCBP3ESb42lpquj9IyFSsSZ2mnQvuW7s8
O31YvP/l18k99oa6cLA2xc82Kz47ByHpmVRUGI/S6C5DtXCkS+cLbtUONJoh5sWM0fzrEklLAL3L
Py+fhxZ7TzcJsB93uJNdaq9Gia34FYwiWSBjMsmCP7AWxZbRGp/K4Q9L9HAscLGLHnUVUKNqck0o
tlmKV4N1PwCq4ddBO4M0Cc7SiRa6X7GTYCGrLJaBxUTT4yD8QHxwEf6x7j4Cpm67IEFGRuZif6Sb
c+OoQ2FKat0evL2+wY5UC/rdGDnsqsVU6MVaEcWTI30oc94TnUi1PIxRAqZFmxentB8Yp6liZs8S
cimVQIbMHtf+mdtMi0j4M0mQVtIu903pbIlk0UAqsDCG+oN+UkmCzFotGH78GcPGBjZ/L9hEO1aO
ONn/2dvNbr8KVfduhfuoDuWVVQhOH+z9enVBbAbvafd9UJbE2ETd89D0w3ylfhDj0TDj2Cx2GmV8
98P+n2UDRsWC9d9zCR4JTeqVDA5JmbPZEA4z4cKvdDyyCNzRCVE1pbBmTXjkf2dgrO1syu5wnHvS
lN3+V1erC3qJpCcxOvRhveEy+DU2zm9Zkyce2pGhCU5B9wy1naGTH2sfFCK8t3vlZqNl3WnFFZ0n
mJd9pLs8WytBHLcRreBQHc3VJ9Ds+Lv1/+IAxKzpBPXN+AY7wiLmQZ1dRNE1/e2PMPkHlhOlB0Bz
jhphUda4MYOQUvKgD8Nt7xPEJTttzw0cAsuvGob/80j6UIQbm6JCxsGudHND6y8/h0jF1nA/QQyV
55GoSNPWBsgvPO/Y0PrFW0Rd0DSNWoOoe61Xlrh5o6ahL5Y4sQw+q393a2UjFZQpcRrFolkPM3Pk
WdeHMYhvLOcQCB81y/iIwOyZ/WaZsd998SYpELVJNg+TQyZzNQNXmojv+HKU2nDoApamC3TSqPFw
6x15wp1Bghq/35QCAdi97scHhXzA2nIzXkK5RwzZ2niOR2Ii+CqRHTPZtqa8FrIBz3bF1lsclumM
JUt8ZbggcQHxO0J3LEwhqHyJYo9Ija614TmL23upioLYAzzjGq4aFn+KTYxsunhfsEd3BalBTbOM
Uw5JQszNtbDueo63BB4+nL7ytVyrTuyRfOX93GnBJl1tLFjbI0/SqnmOkqj7vC4BGats9ICv3TMf
3/R9e1wWdyqLrbqTlJphfrVV2rfY83R4X3pBTE1dFL8HtJPo7OGg8m1V/qK/GcpYD2zCM4lmCint
wcMcjdISzu1Cd71JpiffKBCNKPtct+diPSI9sKVfuDPEzmle/vWC+fdKiP+skH2kAZ68Tfxbp1lV
zc+/lA2qsHf9Fbm2519lbYGjqMFnEe69T1Y15/1FwkRwMLPZZnhSoPzB84M1zXDKZUqNaaKI31rv
55Xep40BUnA+m6ANz2MqukV6vBN5NxlfuE7GYLRUav3qvgnoKez/zC1sw/B5XBOo6b0UU9IOF3nI
5moLxHAbt1bqGQWfTtNcMqafqUBv6e2pTUSDEY3BeB+qnqrV6u4ezDesNx81kkWmsGjQKxAs89IL
kYnef1bl93J9UbfG1xipMHRnpoXZ7wo32YQhmm/B6le/aiDyM4SpnbloLAKZQkSCeCTSS0BEbLHe
bHq/TIBpxZ0FJg+KPJYZpTtJJcJEN4Emuj+AW0imL5EY/HTPI4YrHkZZiKqf59tAEKcHWtDT7491
AD3C4bRC5SB2iiDKOEOGAQ5f80yHZh6ef8Lazl6ABVmHS1ts2MVgW7U4L0SI8fxJW7b5sHwmoMQ8
/8tFCnTriJWSyC0dg2vnCEpn5lz3jX2w6tQg6r9q3S/KiGGtNGjZyPgcvmj3Bv2Z/LeZFZx9BnkF
0zjzEDqYRqjA+QRvDWv+bABVeEbRCpPIVImGU3k0Z2SD6v1cQq5sDFVFIiPXmuC0DxRz7E67VihO
phWiPPCPeJz0SLyMvoUHk6pJ8O7+0M6q5PZU529QaG2hQUclb0PaeaJKUo5cvv+Hhbrky3Sjtliz
N7LnR9dL7o366mVuJ9kputf6mKW1JgefsRmwrfY55a5aB55UQN4x6a6Nd3t/+Xbxi7Vgn96GTzF6
zJ9XEorPkygubI/H+x0A28DJbT8PPQRVb+BGwbvs8sV2Od24jsyu2c7dsK+/BHAKwuu8vp4kYikD
KOvWD3PdfO0XQphWLlWQsU06lAnd2d/smv4pmyset+miwsSXN0sTUDAusbIdKUsSJYx4mRKPlxtq
uqAK+zDoCpNWQcwlA8QPiLWcNMFhj/H8fX3wZa81MrrZZ4tRqMFk0g+F+YbZf7/WtI3IDRlLQ0Kt
ouDLDgxnsSNZTUJO3HPkyf75LeMW/0ajzmitB6MznsB8iVN6rOLxebs2bGUaANmND20uBDwsRopr
TyLF8hcT0OKLMmdt+TQoJSGnb09TA9mMr4IKlNWjdXp7CyL5/fltVli4HvH8gbLsnwc5FoSex0Ht
rovWlpntFE4PXYEYmpO81zBsPWUZ/yQv/nIUSJz9dtqEU8zs1Q71uxLSJHSY9dUM2H9eyl9HcvhD
yGVh75nt4M9kPKLcsdb/mRL+9FFHi8gRMvqyoPDpuXDyVPxpiSYWK1rTgqhlo2SrdDBD0byfRvW2
6e/nnH+U2PxKMUxrABXsslK0+98P+oV1QB4/tS4OPmXoLCLLttlLmxGhMjUcW+Xv8Ovb7m47E9tr
pQ6DYrN5spFjVuplMbfSyjnJDi+lZ5LmilrkcPs+t62/AeGJsE7cFDdqfy9uIIsUbbd65wfDiNPJ
mBc2wfFDsgiB0GdQ2wxLgq4cUJjUoBVarnfhn+WqMZ5P4iyIMjrf6TbrpEwEO55bIm0mDY85zbRm
0oxmhVNR8NPKGqCxg+MYuJSXUrNQaQoaNQVXI1mrXiAVCDBBcQ4AqKHaBayN4kZXBaQFh3/jvooI
CT9iHRaQKbB+od/xNSRcOTufNnjajzOWynycPOi7FUNom70zDEa7AqTIkyY5nga1A5+WEykV8kbg
ndhjz6UVB9n5dVjOlHsQkPrdKMEgTCeKveu/puUU5WK6kcqwNESsptHFHgIuYN0iUukj7IqoJ00N
6UQwbPosI+HNcv3LHZ+LKyZ+taO1yOuKxsjAXCG/mNMj0kBYiiatWCdRnU0eFducaLlC+IrOkwFz
Io6Iriz5vIerm+zWSyjZphYrC6lcx5Arj0zjoeC6KOG04+boGmC5P8TeZ0Q9z29MliP090JdYxHW
F1T6IX69xn9VE9KYrYIif1x5iESSGNgbHtVJweA9aBHM8zULiWoRERZHkfjJfedNcU/PXP35lPJ3
qoptCMCpydn9CzGBX18lGKaG6Hchf6pdO/I+XsQsBjjp5RHGTf6B/Qpwmab9nU3k2Cy4iVYGbxZ7
A/G7nIZyUR+Y/jf64e7WFaZgrAHQMfNHl2mHRTgwHJSXNx30+/U4WGBixLfoG+ix4PrrzUihv0aG
YRNSScD2/RslImf70bAqk1e8TxQAwOK7xhXD3TdfmwnPlsHpS7HW/OdtzTQRdqplWkrOdRYVRaY3
neUO6N+LFZ6Ev+JVTke9W97WoEoxkc5q7rbgT9sRMZDLYk1PN6t7xB5OV6CxROMz1fBjVqNZYx8r
zV3qfOA3hu8Z5SHvZZmbTQtRwWSf358HTmy9JsJVouwLFGhXBeUdHcMpd+cD6xMTnpoIBisCu1Ef
4s80jF9ME7T0XawBPyhwjfef2v1zk0I7hJKEAv34KALUiH+ipuOdmhiurP1/ArcHCJX32ItIzGBn
VeQ04wtqG8+wJoLSpy8Zsg2BV64KVi2OKUMtcnqg1Xm/ZCHVSCv7jXcae6bHgUzUd1jJ2AJ80U9f
z4qtNc7xDSOOjQ1gzTSGoTeQ1Op/68XlupRwT2JzcNipv7rDiiDAmEnytYSms0SdymqJ5wLXgTzL
eI2nbuWcc/3SIGBoHyLBIWm2sfqVaXSYsEZP4n2gCrgx4tMjIrhOWQq4zeI2rMPvsit9Kyx4eI8y
nEIw+rpAuipgbH1dJ6P8lkzRyPItAgZQAHLlqCg85OLSn0tP8LGAQuwpC6bDDejrqB9GawGmkmWH
x9GL/4Co9nRDJ04rCiGkspzL7RV15Po2de/4N+XCkc+1CRXEsX2Hj87nVvZdEnMuexJHjXXG8wFA
0M8jOQ7p6lHSgh791UP8AeJc9ToA9b2ASjYrAzvaDVO832cTNrt8IaJROrUixApMn4xhN25WapL5
0eD3hBnO2acnYGfJZykr+dWnhEO9tNj3OimcFk1MyQAZqNiqvoB5zaSPqze7pr6Z8JJR6UFNy2d1
O0rSGm29usD/PRPJqHJoC/ScUEl8Wagfg982mxT4TLVNjh0RM9YHFiim1MChU12zyhPCTDfrW+QF
+HqUKmtw4g/zqMDNqbfn36qsAqEsGGyk+hk65kVL3vnpdDlwJZHomOF0wOCY9qxz4G5pzFbL+xgZ
wp95nkNkpD6lITX5EgPFm/ycYNB3HVVZuiZTydYpkkEtp7jC+CJS3QSpZkJ03Tr0GOXFi7tLaTof
WAAhbdBIw18j8yWuPLqYolV+7Xgyj5QD7oPxMxZKTetN2/MWgudayGiKg6UHfqKC3gthop9L/uY/
IwHA8AsS9Vj5VndloLkhdjFJ5x7YXyWFGm7TPc9irsRuI31fL9qs1Q/RTGXqe49Bv/NcLdiDNJpq
fXE8p52Mojj2uPCy+XV3iGumWGoGBeE7ngGt5YF7c+cLJxgsd/65/BRzCZnJLWgXRw9txEPt7hz4
B4Lm4bCW4WTKDhMc8ECun+Z4++E0EYvxYr0mrlqg0HGJm0wOo1zbkWrhf3wpusryQSLzBvBK7YyT
8vGT/faMNSMAgPLvAPogufSDxH4d1WLWX2j3LNoC5ylheOiOqa9G8mDM5h9MBvakh2G1sTi8BJ7x
wiqtVaSHmrT7z4lkWjy3P4KhbJ8eXfMIn/6/33XIozJBTnTU4XG+p3CZFGek7iHghSkd9WyfGeGw
cDxrpzs+AC73SxXSIZUTYhabZRPIeDVes0pyzkQRFwjqPShq/Zlcqy62bREa5Nlul17uKnWgphCP
vcsZvX/tBzc4g2pwDaDj8/MwzcflLzx3EZ8YHqJwitx/0GwulDN201/BDJPSU/nV3t07yeI0ZoTN
dE7RDYrBfO6EhInTFdbI8YfdoHc1FtxrfpWkMcK42ECt+I/0PhWc8qfTkCrMdPiJQwF3xpblcU2F
ahvJIJycaVCkK0qk2yFY5d3tE9vYssD+N7rb+AQk2oLOg/kjiWzNDpsrWPc8a84F0gS3p67lN2yV
XlTBTB3rvr2kT86D7YIZrl4eGSyeEZYyGHR1fx7Vl5tPETRVqj+QAryp3860dFqOwbTFEptPeNN+
4JZvu5Yvn/D8OKomVkrtrQVNVfnDdrzrNE9sZ1yCvfhd9EzOFltIn8/DfypkTiAuw7I1mDElpK5K
mXC6YjxDiPf5depiwDTk8j/WD69VJwx/WkjSF3Me97MGIsiPmeewPFNeLEnxrPOVUTGLxDdlLCVd
P+aNnWd47i01qvy+5cplD1YXFoTdhLz2Gh7pgJTaUykJdOclLx7xscU4PajH8AOi0ASVz+hhfEUM
QTPUrGIuYskq3qpeP5lwUThEKwIgB1T9U+LZH2f1pb3wXJ/MuliveomvXP7EXSlTON9yRI9Uxr89
1xKunB1lPYuygG+OvGjfJLP5qLDyZBotfjYpt1hSED2TdoAZZnjWgxK1cxWl3D3wWeGW28qGSlxK
7T+zeLgbwxxtpBgYwbF2L3AT9909EIYqxgtAI/AHfg5ZH9+AWjbGeQ+S4F9ySU/3P4BEU1aKSGVO
YubVc2C6MdJjDlPMsi1sXVOrNFu14Wmzxe85s5RP8dyAtEw9eqBaCOiTEXeCKou2nM+rKxt53UvL
VKUQIklmItCyL0U6qjuJt6Y+mOLWwz3R+3P8ZGEsZQp4HJ//H2e8p7otNru1D92czWIlklLWGhnS
gST9BZFhlYx2u3uxsN6AyneLB1rJaX/Y8NnBn7vdOrkQev9tiwVaaqYkE7WFGyI/wfU9++XGFvFe
2M1RWbWcqyPH5A3E8oOzdCBJE8Yw4Ku11JWSGEesCwv51qMGsOM5UZVKL6uMhW4vQYYkmqx87/ee
ObqJ7tyqvsZhNAN2+4T4EOv4un1uKfoJF5pPfYVtdYTOGzmlLd41GSe7kuWs8RdcizNrk7O8Dwp0
/dkEijUrDneu80i6juIme8HIgPS/zW/BRbjI4QWIN7GWY2TY8ee2zZVG7zgK+bbZvg5V3+7V1IA6
E9uAw83poM7ervO2RMyaSZWanyLe0Rrl9gle6p7lvovLKIWptJAREsDILP1lXyelumxPxQL/wT9G
MkwsoZk3Y4zcUPEIS0zWr0TswWq7yD40l3agEsencV8+iD45oEno2OCcqPU/uAuc5lMhb4+XCukB
UVbQYv2acTmGdZe+3CCClbMql75MsuElGkVA/U5O/RoTXX96f7Jz2Dlohk+KZm7N5fkESltS164l
ZXt+Q0nyLtLhbyJZTQHD2gPaaM+DPL1SWThyuvGKdNC8AIziFN8AhXpYXsmY81bKQvx8uMRixV/M
pOwq49KvjvPWKIFhnN/kI8GPXcqQxK0zfjRtMbdKvqMKiuxEo057wE3s/jbFWwBqId57p+pqS3kN
6PgPIkjUM7XKtfXR/MeWmFc0s/LdgOgZ5nV7Z4QfLork7DGsLh7EuxR+rqhcd8f4G/XGnjCgeDxU
s1UhMV4kWWI2/7f9UsOYza62zQ0E79srpMWRRgYZ0VB/F0Yph0BYRrOJOxH8j7DT5pxWsCjKemph
MiQpRmtixI+lA0J4W9CE1cy0OZx04mcd49ar0VsnOnTkG5Dinpl03jnlRr/LgCYZ5VbObsc18c69
nZ5JouUZn0bxCDjEiKG0Epi3zFYWApZ2OZgi+8XCDT/iCzi6c+h3dSic85EUsf7w6C5aJ9eMSirK
Mggv1rypI64yAEWHeszQhZQehVi6CStOO9gT4lp2D9Qois3wgTNNfF3G8Aq6UUcCU7T82SJex7u/
l/ysp2Rj066NABb9bG04+H4L9ACzbbOkj0sSDGLTkF92I1U899R552QRKDtcc5MUdjMjl3Rs2lAK
wQRHfy1Wv2Y7t9fNHw5E6Qr6BuXRgV3CUn3qdwoYBTfHsa5tzDAI6wrCuPCj8rZw6VYQYNT83B9W
RL6JuZv1RpFEHbxcc3gU3WHRfqR6ARaVDw0ssvkaXGAyw7NzyDtDhQZFcYpU/Z5vdr7PX+MCZrMy
HtmPtlQumefY+mOacerBxTx6yMbFyoI0fw6WdEgv5VsoOwmNCOCD5/PjOeHIYoi9uUiqrDliNKu3
17UpnjRHqNfWm/oQhjZLAbmPtWim9bigDhPdbmg1Jw2CdUjCOq177FSL9i9RZt1Arj3Szx+ccnbF
2f+QWtbKO6qlbP/blRxybYEftdk2klcmetEbqAbhQGPeYNHH7o7RgPdCHXNbSrD1MXhh0wGez47t
nz9CmFif3mvydpqmcEvmZrX1exNVzlsj21sJowm4jtrtmFD/pvzkJbkbf0sqrpMptdI4pHNbYN6V
Zz4Y9mZyyi97NhradHHvElEA8WD9A3Z5JG447ohw5KZ0W6nuVsdZ1k/7B1Q7m2aijuyO/q9TYms2
h1ltzaaaolXZgP0J/VXwPP0wawQWrR8lPFdIKo7YezxsqG7PFwvZtheLO99itbXnD4KFvQFxmz6C
0DCaSk/pFbkGYIY61LPo0rUCI3369mQwUPLzIpBWS0mCoNB/QDUCw2es6IPf4tUFuTTEiC2vC4Vl
HADfSwUEp2j1D1Q03+BKQgD6NFuTAWjZ6o2Q65NLAoIo6HCrYfAy+NImAdvZ3HEBF+Z9iM1i3wl+
jteMjDVHyoZhBzNYOyl55XNY3q+D1MOAYlAAYkY3ehsedcQe/R3xFu73dXRSje3g/EKE02YK7KG8
I5NsWbMFBNWYRpx88ER7SqXodV/mMw7T4z6OKJw/ZfsjOi7W7a6cfl5oPYKgVpYrhpzxnBDQOxvg
HvIaM65dCfPZ0RQ0KXcdWs0cPCPpmzB1gBn+zTfqQy+KOQSomeIMEgI0KuSjLmu/8nLO7LNuRv9P
BDYo5vh4W4B9ujGsrGsol2/kZxsix/CRLXQOH5nXUFfS4T+qBjgJUXsDfXbd3x46bfx5K8ToYl/h
9we8Demh6k3xXjijJHWlX1xFVQvGJ00HgmUl6Q9M8lVAd9XjLv450W8xCtLVaWPHP5odbhOoY+R7
RuCnZSZJ6KYwSVW7ijTbkM0D2WlUAlnbfS+hsb1F+6Ai0fJRz5HoeVoVp3MLHvoUKtJKi2JSlhUF
QYiTWGhS7q85qjpmkQsw+q8TADgNgDrU1yKEtMkjg/HLL/iwjtO99+7drm18I7dP/RMzWIE5ExtS
jqC2hRtWKzBcSNd2t1KKJ/8y8eO5Y5EyUaKDr5wI9zqo7MD/UTPBuZpixjGpHaLQBdP6sMWU5tEl
3YCM9MshaDIiNFIZbhLjnBk6ai5Lqk8KUaDrO1PFSQnV73dl4Mqhqz88FOW3tUH6gNdT4XE+6gCN
NqjPzI2pzkbkLCNqbyD697QWlgZbZuWlwZdksEM3knF1jfdCklsQPk/XcloTWmFBMNJc7/3dTtrl
7fjNPygfDB3OGlErWu9XOYO7FmnJ4D7Y0KomMfRZzPoCkN8dsKiE/82iKFQUkCTcCDblevXWELYi
MLE1gDtaNxZoL95QTrE8kvOhKRfpzC27q7T6uWx45D7BS+R/9CxH2o/IFyKU+qcQosTj5HIgIaEI
e1mIRyKMS4ta2T8jVcUTV/edlOzj6GDIw7Vq0KbThf663gPGlr/hFyo4YxgjPdfaIcE5BkWTksU4
1BGMham7UOx8cKDfY4OJz7u+AG6NTwO+R0x9o+nuhQrJ/hg5/GuCwG2zdQAryXxNnwBbkAGoO1PU
Zr1K6LgYFDx6TLKm4jitumSOYxklyMYLBnEhzvZCC7S0bjxodXFEKnOq6j0deawkIiCwX912j8Vc
9gpyQqJxhqU9mrrKic9DgywjIGTQrt9nqYGv2plb1gbdCnu6ueQdWaHzoQHjAS3+CKoxpR2975s6
zYrJbnUqRAR5rP30uAU3Xx3h0MAq1aei4F4Z9ZawzCKmzFD8mw8I9KgvGkqaSXU7H7npx5h6jwHj
sbZbeIIHwkLTf73wszGqYilRPvq4VuC1/ZwIYv4YlvUqjhRs1n1dEotW1/DwieNtH+Cy1j0otLhM
w1tR1TucFYJPMSXknXlK7q4m8qkeRNYxeCgsgTztkdFjb6uyXax6moRXdlIAcwYMVfnCI6SGK+mQ
nZmleEXjfVrGV63lUx6PX8fMPbjsDN9xFrBWY5k79mmRffi6eyCF2y/sDoHFJEaNk9NyaWjDn9pT
M9oTnXjEPl48X3XR6trEJWHlDtzIeR0kWQgvjQEsd1jj+pdlgBzsRPD8ftybVrlY9YeTXVRtD9oF
CG+LZd+63zSUr/bNGKmaFVOlcNoVmF2KodfGjBz8NERF4/oq4ZgiTbv9hL0BhE6ZI5r+RepUA80L
q2ChutaRZSdOpc84SY8HQkGyh2EcuACntdLXiEpKC3mPvtLpVQ1YrryLV+ULmjVJj7GkULGibDbh
oe35uOKeqylDXVX/pCDTSTF4DX/gY56KsN/7grhoaKQ0BtGhknBJJSxShqwezONT7dm8S2Q3Aknw
KaDQcYljlBaj+HRIpeflJ4f7N4I+WvrCqSW89+H3G1ZuUbIpv9AVtLpeSWVgKpUv6yNyMtJQvzYD
YbKZIOzjkFTWboNYzxv91btUb301RgWj9rlJy6akXKNOzcZTAPg2p/WdfQRcHpTLTgnc5nIvlG9m
Us9177xtQCzleHp7otFpsCufSNNnCSHZ98GoXO0L6jPj7M7gHJrKfJzHTmxMiggM6yYcC4qRBNSx
c9MKNIJjhoSAGnWc44FTsMDHIte1oCKln1fuAA9ryIytUh3oDZf5TGqYwgqeSyx/v/ClHOKjkeAJ
fVvoJc/tahk45guz4Wpkj3d3hJefnTyEkCExC8QgshpyST5KNM+NfAl0N2DwvS4zhK+RG0eX9/mh
GLEyljaXe5hz99ckW8Xze3gdkJBoj5JWT/MF/M8/hEMV41NPJAJkyK+0AJmjJ0orRgnBnGRsDpQh
SgiTOgHBpurc5g9dkwxJWR8KRnIUwGbSibR0b/N1hB1m/DzhAp5m+lWuMYi0AVC/2c7KgtvPbMyD
MAqEV6uEbi1jjJSi5vXb7GOj3WeaCuA9XNldYN/RLNWI9pUgwY5niYLrgh+Uvr9bGsVRwXwCru0F
d71akCYvVllBMu1v/RYmzDoZLf4cMPpSIeXAV2jF1Fq89W7H0U1htP1+9XOI1IjeSlFG/Wjm7R7k
fQKA//G36PGQ1cV8OsjuzNsfaRxH9j5h4Y5anWMd7jFoh0DI90peq0+9USTNypuGhtIv3QfkYXfl
wfDw8/Aqq1CkdAD2yiycRY4deoSyH5wOMNDJ6mDHvCwbAzjX1jDYAmKEgMZv6IMD67uLY+eBPopK
sS5xZyAYQLTkTArrSCiHJS/krtV0FvmqkHmeVxOBQUbSdIc9lFdP1F8FA8wYuicfAP7Y2ovs9Zg9
Gk/0NaZ7ZQ0AucrcXHs1G8C17uoFJGu7VfduC2AQvfizXPPy/Jrk10jJDyD3I0p80gm/XRw6rw1u
IbfPLlpj7pB2PWIGSGC2oh/aw8UDKin51xHTgnKTxv6pkN0VUfsCpDAo6Fdtfy8lbzgy3BxxcKRF
uydvw3iuScFrvYn06BBtaM53T8W56QOxwvTV0DpA2FiBeV3k+dm7kOs+Zc1vdVEfd/KWfWV3QctZ
/NBj4uD1CBB9eG9lTNJgzvm+BmUHNTFPh1y0zHGVXkXO9ggUztDRfRLUSIzQNZN/8CK3wGqj5xYa
YLHojpk6U0ZE1U+mUhwzheXRFFbFkH+nrbqAE2xhR1c7uEPwcOR6J0MdiU7vmi5GG1iPYsc4dAwQ
YCseJXAffHbefFsVUjcOylbjPWJh8xz2gyLNlVpykPelr/isiHiGVveXUnSHj5kZEfRI+gzj1cRY
PaghE+BnYCBbprunWUU4L/EZcF1bfO0Z1pzxgedDxXBnjFd6jCqyoZAVI/kwwUvqqmZMjEV5zAKo
wmjoNM9pCC6SHqBvCUPnkYVX1g9IKt2yqkjOz9txm3JSe/hzyUQWtIhUIiWMhW8EchvjKZsY04wa
PrkwPA7R3Op3M8CeLa4v6Xl7kr90keneb83jkxvbtp0nrS65WFCYmv1aDk9Uaysa57VGQi1Kllb8
/JRhVmH5vPG+nEyf2RL2rP1Lh1mJ66jz1hzjB2+qhpk4vQBHbs4Jw5VfiH0J+DfxI2db4RiSBv32
2j/goLqmDqbH/LszJVPzp+lQgrZNLEJkgRX7Q3pGVLClNeO93lWfiSSgBgsr/1UVI1nmXAYffpkE
yULEVmLXE3qPWvfrKUviwH+1t5Cdd77p+HSmswR8GbOL7sYkORU6TjwHsdon/bnZ18fMEi/w//cC
ERDUs+0wpcCV8unjXCMhfhjWrBuk1fIXPvq1kpSBSAT1YijLIYXh2+FA0LuAIvO3BshmN73CoINt
XYaGIOgeBhD7f444vOhH0oXvPBPjm4gCHrgNzvqDsXneMdkn8JdoscvIfN/H3YbYz3Nl7LXKklUT
sMLyYbGlakrTWieNPDkru0NtRoI7fkoFmTmyQB1XCBtpE2xSs0AtnvVKCLd7Ft4lWMRfC+sD9aqh
9EyerHz25PRfL7Dm2b6iFzflESm5pAJiZOOsRhyBiO0/esN9s6fpoUq6zaXUta/3nuGS1c+0CM4I
8n4Rzy5DvKNPuDrwrBC8HR3PgAFUXJ3g5Vmfz36W74aifdXwt2K0N29+Ach4MteBOstDupfAtL1B
ZQfjI3X6DphSE8at0qRnNWiFGvHm3pTTvlEinw+yUcxkK0TOvZ//O8FHDtrJPSIgdvBtu6iUfQYT
Gfk5omAeiXmw8L70SKcMbGaTDtJrjFAmsepLzhExuEniTiKGdJu1n0LJU4sT7/K96mzvAi8Nnfal
wmyxxh77e3W+TT2SCvx0qQ9Pw89qqegKaQ2oXjPCzhCdOY373p19wPGjpfu0oU9a2LLlhCOIMU9z
wRSO2Bs3AOlai1tppKm9ZUCtDawv5BMYC8Ul8JwpVWKaNqzRC1mwIDsxXeFjLkV9J5cBf8DxNrhO
chKg9koo/I/YFUifPo5DECsLvLE0hJ3l42zxpxU50PO/59YCCaASVtN3xrIug0GCnGSRdPMioY1i
mu2Y4Gr+xM65j++doKgr4zfsogrl28TJxbg1fPNOIyKIIkWFDynxl136Yq0ApixDRb32L4BN8NK9
wRhHxbX7D5t/8iQppA/h89q0LgOWswQfB/nE7w3vrUixL6Vj9QX2xTigl67DIJbep2cL9KDOCXS4
fGA4+f/SjMGQpcN0IRV/zJpunAdAY7cKoOM2oq2ZLwfjiA4+1ux5mRLrA5jO/P6uqRKCUsa8iBjt
5kugJ2BJg5yB+pP0xTMUHtHrlM/J7ovlu77ZkDTCP/vnsytq65qvymU+jEt3cw0WMsry+nmNLo0N
wYP53n8FfbWhr42xOqkkCmBEbdHvt2Pji1QO/sW7BP2fjNC8lGuOPfUZ2Nft7TukGgCcP677vI93
ElQf3q0H6VHSfxV2+RTgL1cuRrrmhb/doi3N2Qmx516ONXsAaAqB7ZF6OluTx6tm+Ge4SF0AkXOH
7H9rmvWnZ1MslLRJ/jToAFWWUhO4qKc0NBx5W2cP7xkd5Gp1yc5z6tmaJy1TCn2VgBd3GUvyaizE
VNfkEUJWJjtlZAhhvm4PI0WrJajGk3/j5Il5sl49xeDJkxM4ZugjK504+J1jsbUdX9R3pnCs8Q6x
3B1PPop+uw/afR5EjqhdKeexwrFYxB1YLJnzL/oBbGkNQz54/nnvp7JVuz2SiRSfhB8/xeV5lnNI
bwaEy9NUM8JQpNGzaJ7peKDano4J1pDC2F3sNYVwLnPXV96LuC7avmLHAwbsUmzNBlUjpDhcRhFI
BwpwZyLRuArL6p3dLk/mE8p82ZJHbSFLjos9YSgjuDas5QHwI0yff469Go9/BfDHNzd318FFOFRG
ne3AbGEoi7CTjaVkPs4wj9vlofFtXqQOEIswPIGac8RvlTqPPqszlyBz7BItcB25wqHPpjQ/rJtt
uLF+4tCDqTVr1ws2akCpuH9zQzeQ1/Mh2LU2F7pRuA5UTuq6rSaZC6qW5w6GxOkbnu/5714b0i6z
cQJqYjDrZtVonmLIKO1cOLgN4b23i6QxCU38f94K1GNWdZJsilExfBP41FsvnsUqLvFKEl55y2mN
GYFBO7ZlJ/PzMGumvFf+D5auIZ7SskHW3DvYvubuqrV4tylKn6zgU8s5Th7B3vX1B6MbAibSmUhp
nihORowRc53L5RmOLnaDu2rH6B7Z11kKyqVyBEmlAlbcG063hrK/+HqTJT8/Bede8UUa6KH9d0kI
ANU7KdOdwDLA/1phPIBoN3msDojKY+oH8jr8BbTHvrLA2ccOKPw6fBkVkXFoU/qnacnVNqiJ6UpT
C+dfPXGBXiIHYcRo/A37HcKRv1nY/gt/Qsc+GFJ+StIix7lXMiqEuppAnT3oDqr+0zFEWF+9RxwX
tTFPpMu06WsOjgUPrDM71zlX6NGdd/QSLNHh7sQFqwXscpGRIN9yUTy56De0tsNujm8z6dykE340
8DaTUJEssWCr498L8QVwd511CeZyzguNNd4zF5Uxdb52rkuf9C5AHBR26plKMwMMIjutccBzAx5a
M73Z72WsTwRrdDNLqAWdsXqV8X1BkHgVviPO9vEQx0A9ATEea6IxVt6ap/mShBa3Tmhxz5wyyoNG
2XEG4XKldPnKbdttnmdj9xRvRa8h0NUmtRoE+Ez37xwr+p3sGETkbwwlZs9nfNEKMvfEmaCaRZr9
twmqcJhl+mj2zMbu8HYDxHPQ3ErB0kraqnux+eUxrYAdhT3yYwnuYpCjI60UsMd3FpKhD8zEEphw
mbkrz5w0oBZxHKKNasJIr3l/i/jFdbSeP0sCX7KPfgiTr7RUJ4JpQ2vrmtznaZpn1kZ+4YqsKpCa
0IHOiCgsbVUJTtEAY/z88YRfI/RMwZ14GKwPqdpkrHIK2th6XKo+nE2lY2jiTriEhG6SfthgeNfL
AzycyDGL45PrHGO++JMA/MpL6Z1NDiO0snvr2vmEObPmLj44gKY6yFMmvhCoOJuhnNbwKQzIX7sA
s3Zfa71TgEjTPbqYrLa6+rHmC7jmkP3xFgxRsj8i/X4Nhxd2TPvr6j3Bl4D7TnTj2GHhjbOau/ga
G/UfahNH+SSLVef8TLJzDXjD0HuMBUHbB7RFxXdVNNvTo1jPn16tAhCcN871PTuqoKZNLQpjQLZx
1n7eY/5ZuvDQO9gu9vGimOYnIgrhWDVp5idMtkMpCMQsHLe9q9pytFNZfDvHUq3JOlIH2k4sLUEx
WSM+hkyXT0LLFCxIDg2tPYqVYPAnEh3+gkRiw3Gq5fY3ty+sCE++lFZtjRzwfQhhArqFF1lzEplY
wEFCuSgBu2Bp4I3IlbSuJqI21/cP0ybc7pB8Z0F2vt+2LXLbcSCvFuVikCtCPbgtsfsoTrq1qedP
B4rTXTSaFdNmgXEkW7SR3EIX49GEozgqMnfLHJ3sxobWh0lc02xUJC2KP/REpy3druSmwk2eCG4+
JJw3pqAhhxPWSiZBG/K2Co1bjQolwZ1z3DyjAxOzlAPXRrEcQbuaeWJ1jKVh7ti8lZvdmFzz/he1
Voypqkbewj2/bmZIN2AmLnbf0RE4wPJTv+bMamFo8CYhxf0uzBZrqq9oSNbccUDumOBZ7pXKGyTU
CvQSpyp7cuXZgLWDEVVkjU4CFOBrHIllwuICZ8ReC6+CW0NCdr+7QTZfSe8sR40Aj1ayNk6kg5jY
g0uSK4K5iSz93jmf6kcvq/dX05vfO3cXcdi0gPF2JkVMjSsoG9V07Uf10scpICStOsqRo1IsVBJw
T/Ded6fN+zPTox5Ne3VEz9L/+baIXLdQ+SknA1Iel76A1pJ/Na7cGVvUCHifRy/UCl1JosAXqBCw
S7r8oG4umBKC6e/4c1E9gQGesjMQv7K/RmoYuiuuZyBVQpWzg/5+ga5hXK9XzmRpdtwohSlkJRvN
glztPnr3g5rVCYjckomiKfLqgxKCwe/JhMCJCQOSmdiWZP00/xUxxREDLaRVnNjl327RQfEbnjfS
ADgt+dTEdpy/KKArtgbmFjIci0bN6G/CWo5JI/bKJHcs7RYYJJ/ur9Mf9SePYPsfOexqTYCKmzFq
4TdvPjxgznk6CV6WbPbGmuoPU5Z65XN7bEcizCYpQZhFfYVUNloxexBgGNaQ5h6fcFAMe9kXp4mb
qqOiYxBIJ9SIZ1mhGCnPfvKri9Tk8gUwyTvLhJGRZl9P2l+CaO4C1Gk7HaNq9mwJ5vK/BOsJcefP
F+XGCSAmDqIdCYHu9bx9nk3tLzYDJRKYYZ8grJYfzFWMpg9uluoeUvt6R66BC+A/5rt95b7IMevT
dGV0ijebm0Y4PqqyZKNN+sEbHrbP0MyUE6m5oH8QLZCjo9qgQ+Ma4wUeVJk1AvsVwTnbPY751LMh
9CsZPLrRce0CuJ/9VuLfTZQxm0W0MJjMUuax7kOlT/jybEhQ+337Ypl0hGmiBWay/VLdMF47SksO
NWOF/r+kIeD+Jp4xVlVK8xmFggOEE/9u8M6Gj2xfGq5fp/Js8am6k8kIh/0ALDhBszaY+dSxeGee
xFb6iyBPxB2cRz+LrGRhjwju0hDzgg+L2d+c/3oieuZU0VpJZO4uSRvIGEuWGacluw+XekdhJyqC
OrdsEfOK+rLiUFmBSieI2ihsP4gDp5VdNS40xoe9nRqQXiHdDIbs3NqQ2dR3HT6LSmzv/GIU7nUr
5GYcM6RjTQPWKFWl7067wV+UXDLIXRzQ1BNrH04tBWoYhsN7e9zGm7IIt24K2Ts3BOPYyAAsMrRB
U++dQz8r01c2Er+REXaBO4YjKrpE2lvPc7DFogE0VcU/aUOUdRcXuWidxU/YwX/xhRXhJosuhlrH
0lLlAqRWQErIuu3JeCwVdKDzOmr0wkgnxV5lTf+QHUEwZ/5s6F06hJVRLzaoPqJkpNIRxA/B2mYE
zybQmxKbfdVGMb7FS3WN8hSShOp9H5l7mRUBdGICAYA4CHkmOMr56WrIrqnRJYr6wW0J5Md+HPuS
pd/6GoJ1fkLCraOhXhx5Ba0XMv4fxU9hnhME7HH2nRDSXdIH8o9T9uxoOVb4bRmyfG4EuUpVhKsW
EhlRVdvbA75o+xAnH/KZob4c997CKMuFXmWqQ8Wte55Ri//Y/g8MuJFOnsxGpuoyxL9RY/X9CH/5
LqvM9ex6MLpsZYO9uhdRQmhaNNHMqzwT/Da7M1/R7/NADmwelB+i+3YkLf61hmJ6uumiC9L7BGMA
gsV2V0naC6foVE7GWIBPJ3IOBNXF6JWqzKiVXCBLrASS0elWEZis0t1sFx5pOOQIDdPAZUu09PO4
B/GTTqkhA9xD5Rz6+eYBTAtqrY6dYFyjwC3PY7SVbq/5VidiLfslG1Zl2M6ZuJAAU6QEci2zN+vI
xJuaK5M5dWpWtcHqC5Lsvbv9NuzmYt4LIoFQkGbPF47NWLDZVxtu/dxFsdQagrYBaLzRm2ksRQbI
kAdUieJQQc2wYYfaLQal0tJT1O3NmaAFTCodxoJ/A6/ytT1L7bfyhlsxhDsIuAk2fYqMcZmqlGOX
ifVHAgNL3/06gBRx3xV5QKabT5Mmn1LowAx4wpE7pauQB9LI4dZ6MP/l1C5q2yQexRVs3K2iUeSZ
SoW/B+kZO75BvOtZuzZqcvrozRdWmNWOKg3IAn+Gx3BkEPL8QM9KOz2UHVvzojZcp+FAZ7fvLC5M
OlYYk0D7dssn79zzDV7oZx9w+Q9sM/+Ey2qJSGlsxZ+vBA14E3PkHOCMqHdMaKgpmhxn1bD2lCUH
AkM7mAf6wf0cPDAmy3Nhop3nsmaneeRBBXqKX0EiZvLFY8oYDZibNUjPW8Ftkt4XHy+78mF42RpP
+0vZ/POQBSDJGOd/oKy75WYbxPYsABxMfVL8V3intYvnWTHANHcqqVs98iAU68/M69QhAUQOqjNN
wHK9A/meU2VGmPMHWFGXRMqR6DsjmKpQJ0ge6OjMobU7i6DUbLVn89DT1W4egbtfnVblpDGgQXUB
t8l0vKWezbv1hBysF2u6uxJe/RAS7FRK72wP/g3CfKZnGP9riwljuXVjHOvydiTx5OYjGNovIz5u
xVrJoNVIwRyWP2pNIEYbEup6BA9IGcnVIFCGQ7VdRqSShaX2dtaTjnPlvNXP7qq2sz1QInMcgSGy
bHL2fZXdQW4iFjtQPLjGmXeGc+4RDN/QjX0S3yzXBAz/xAtVNP1b1G+G32FmGAekQbg8WpoBJxfH
0MJQiN6VRmNmIYA52xpkUoUYGpIxzA9TRKXZf8pJLIMQHLmfkAm5dLeKDCo2xNRNztHnnstC9KOq
0FGkjdD5gB5mf7ZokfPy0y0MIwb9qLA/QnnGLObIDkAUUI0GkLyj9j0/3VgVl98maM46mAVX2ILp
X4zswTgrvGFSp3jbAFUWSNySysIRjF1FABVRzBcwtHNM4t/PJwkGIDhu/BDv1cPmRUU8B2dl+25a
1SefAPOVNx67h0vthgVGbO45sOvRIDN/XpDcYJC0N7ygrGO8fghxHZ0fpmPec44O+Jnwz8z6BHYO
2LJFIchF8cf6TKehnXf9D1zFMT1371ggg9MRUjNtN13ZyNxgX1pW2CVz2eRs94CIRjnm3Cp5VV/w
cT4vczbvFMoBpxrClM7BcpOL4o55hvcR0PJqw8J51Vq6kziVVTi79V9MNq/h/P6DabG2Q62kL3qB
iXiCpBiHXqJHOwPSEAKbtjx4VjCFIw/DY/np15Arswcvs4CtLsepot4xlxHqGczCBfIiLmroe37H
J+06sVLHaEbhcq/+yWqiJ8BMujDafrT5aBdNPAuCF6g/xeMJn3dlXA2LsvIWwXhCA1hcZPjcrq+X
Kg+UwFSF0i8A5rkDhE3BQiq4I3cJcH9O6Yb8N1oXBQ5Le2z8fKI9u/UxSWmMYkZrugJRYzQpKcPg
BMNOVYigGI20vdmy5ujBANnPZ11lSE+8E4MEPwfmQFv1pLEzi/gdI60PlzJ0CGJjWDr6iFSwKGng
pqOazYluYWUqG0HhZ8OXWBzLlvzaReSb07WfGie3oEmwFSWutGMGtXZOeRm1qWBc+m6dDNXkLb+6
Ndoa3Iog7Ct9cWSu5HSZUpmxgqKsW1AQej3QCTHOD53IsXUMDJ9gDgeAz836WKwcKCbrbyFgqWAT
g25C414g8pHCy9MXm/f0bmp9VJ/hHdgZsO9DCPW34F2d+zUDrYHqhU3pWac+A0bj/2IqG/52Md+2
lbgi5n6T0C7GfYbjUkN5gtYPR5spnVMPeFKSf2LUtqSkHRw2QTxHuYBe9sI0TyB9NADP1DMkVwGb
tn5k/BqC/qI7yOObamZE+UPy4r5MDIUpnnhuidiTfoYxoZqBV+VCg51ahBWvM4S+PUip8ZU0R6rK
C9m1FB3cIaQi/ZBCl1nwA4i0AzvJWcitRYaQpW15CsP7ctcixqSG8XKnlPBgX86XU0wyoVPlNLNl
aV2hlfYh9wG4w/oRd9pZ5dSOZIPaTVmt2Mk/tkYZ1nfD1HUeEsLmXD/BIRq5J2xf35bK1PFkUsds
sxu+wrXimRSgonnsXjMoem6iCzfHJoGZuU2Zs14ABjKTX743sr76wN6ZJ5KthdS0/O7skW4EorCK
KSGX3aDTm8pPuH3wZH9y8Y6jZ+8UBtt7bAbYcaeCgb0pK6RmnlXXkj+CCpo5d8miotZnjHssPhk5
DECtUn7XD9j7d0cCSprzSQb/2bJPAo6+0ikngYFFpFnWpoyFCh6YOegLShjp3qNjrc8FTkJDvmhH
Ls3mM9fE/gtv/sKou5OHk4RDbaQr5+io5Bah3iIZyFsJ+iV7UntUGJlIDzwEz0EHWQv3KWZeCFPQ
Ej+vSMTwa2abeOsaZQqcP9LVkj0DyQdBhCktDXza50wqORl3MWGd1FJQrLOqnUr+f1MEEBMyTQKx
bTUm8r80dtv2BGREVkrLlMpzIb8BpCIBpSu5EQwPNozOhzDDKek7hdoLU+XqBqNF6RxqGixgWe7t
jBUfWYdfD4RE37nRbpHW5gXuQPD3PyWk4wKUWv9rDeidBFDmMLSz5dfC3CQ/CpbzEDde39yNFYT8
gFyzm0H8fXNZ4WcfYp1BHoWQ5o7aC73yK/oaQH+vjiQ+aNGTwKERNnesuOxMCTn3vgKaDNskjO0q
1qw6rq+LgiIuD9de5Z6ZIYl05nXUkt/DICPs+m7JpkRskx3Yn/QdiI97SB2Ir+eXAf7zaXfHmIs6
pBEpqQmAKXM3Gh6GZ9fwcqJwRanOKjdhPxRKK9z3qV5GYlD6O+XYI18D4uGDyqCmmN+hqaRSDEMG
unQAXzndDmUa4kWfFSWqMoNclJpMU1sct4Xm60CTyPSog4PMMOZIVQ8v4vLmFNCdB1+d/VktsM0L
7CRCNMNU+cfSBoAM/HZtl5u4bv0k9XkM10jW2+KT6Qq15yJB8XDLGMjW8NvoSrEyS/9hOIkuGgpv
h19vkdPEM03JIThC438S73E4mUwSmEaqASM/VKFhsj/IV31Q2O7NjU3T3P1mO7S3fjc1NjKMw/lU
3E/mEX/SRIAKblFH50en0E8UkRUdhw51SY+Gp5pzyTRB8rNBwj7ZkuifSoxiTBjIHnmZukH9TmN0
wq+fGQzgcfuKDa1G33u21QpWAUfAvv20qvd5O7Sm74n/oF5A2iBODpJ3nKT2TMGBH1x61S8mO1tM
N1VZfdvNQ5qRuW2QtZvTWsg/oOoB5lgAf+UNsfbE6sBH0ocCoSVtR3mKVt7rzw7aTZyws8s5la5y
MctTvdxqneOAHxoVn5EuzSC209Rgo5lqlMpTzeRt5fAmAplloud17XTlFsLL1WUVwNGqGgVr9asP
SnI9ZaElV5SEbKj59VUtYuOZUP5Bbgap3Zleh0pgSuAa+nvPzmyRALVWD51q5mr15xJdOKf2Nucn
s3p5uCbEVVXhjBQZNhP9Xi5YS1lqwNUKPqBX2EHQtoYMswyLhbNT5hVUF8RXNBFInC2shx8OG9+t
H7uEUO8rxgGKSOD8ogs5qMxstekOz89N9U1z5MgPIcuYB9blqfUj5QPO3eYf2FsJRWwNJ/ndlVR1
fHY5H3NNpoW7Gn5+5I9/sVxqwgIw2Q871Jww6pNURTqBtJDxF6AYQgsNczg+6ro8Caqr0z9p2Gck
60JD/l4yybKtqscBR7j6aVuyBqw/S04UB4lHsNAgMaYGN8sYdsx3eHSImwGQT1Ip4b8q6akkRVf+
OBQPe9Dh02FiiKw6MZBAaNH9iBEnJjBAw3lR2/5DhWHmSwJ/U6By2FFG11G4KgBk58BBdczlAE/C
wqSZIHg0/10Rr5ADQ1m1T/E76EYq7tZCuFte5/S3nodENuy6CkkReygtaJXi7vUmx/g37aHD/t3m
Z4t+exsSsQrRq2CXshwCVS/wk2sW2SSopUAuvINnFjXWFPBgtz+3q6mG5dg2BhjmCF2C4RyU6yUS
6ZCnrdW22TaCO3Y4jphEhDde522+Tg/IAMD6hNXB6y5xGO5JKyneXJ9eGsjY5XQvG7Hd+W8FteJF
l3LKKq2887TqPDtzzqhCkCkBDl/pboNUed4LxZPHf7JPAShSclB5nbJTiq4+F13z5tUIRRCDlHN5
yho3fE194smqtyzhQbEL5LN3BZZ5tmi3tOCbTFMVEPmCbJURrpCFgeCWIfU58H+5rSqHNaxrIgP9
mIczekusp2c56pS3tIvZAg3XzKZP+3yIyYm974HeI8BjeF06D6PpGtF3VHxm/pad5lFmJU+KsLej
pWRvQpr8NWvd9ypvhZGQB4akB3HcwwCKeTZQ5L9Ps4vlGjRrWJ41REoOSFcVRNen8AgnNiDAly+R
DAhWbquQGH2q745Pkzluj2uV13CCRH6MpRxUxK1T3K0DRUcmfr6J3/6QXuLt+uirHfGBgqzXzsdF
4Cajlni1Ke9aB8pZU0oSIq2L8qE1FhyZo4Na7YSl/42GudVaemYtwt3A8x/LGb5nextyXSkSD3dZ
hcsBBRxQphGUP9Z6kwuXEq3E9iCii6lut50AQ0FUw6EFYR4KZk6hFg4z9kdckFx33cm3q7DYd8Lj
wdO+r1qzmpHz51Rx4kh9o/w1chsZsut4QH46XOMw2U7jxwfIKOgBD4Ybz5sN+JkUjQfViEMlgW6P
7pNH+cPvlr8ZfTcMRBgE9yFzrdFLof7MU+a+q2uYJ6y+KeMn9kvjLNsWYJEBWX6PZKtbcNe6mB3l
bqm19ae6/psSPv6jShBsy6Ydr0rHkazElTp+rEmHbAQ2lKq4MI0PznXqcpebOD00w89FqCdKilld
/iW56IqcBmc+PWVpXFPmP4KLmE7r2MxXrqq2DePSDN9pTG2uApvn6tuYQyKF0UqiwTmxzgCYq2r0
zIZk5GM8slOZXDtKG26of5ogfgCiOeC/uQzqR+p7gQvUwHjQ7SzDwjHczXzU47EM94+9+WK1DSRk
a/3GGud77nvt4VdTgtKyqg0E3xhZA8i2Z+rvTPjh6TQWi7u9YmlDkWB9OBWZ9Yd5/on+GL9gSejZ
V5l/8AognD44YbSOFrBIivgDvG00/218OlqigwQh3oDCZb2higKZKr9th6rXhQDfKSRGgRbUrb0L
xrsrZDB9zcUKBtsqelRtY7ANDoquXQe74PnlPEQD3NkXfpBgV4D9qFRA3sydo/tfY3X5pb6cQCKO
KVIARrC4ThJt7d0ainweKLRhjF7lAi9gl0PwoGgytNHmgA7QZBS5LOVTaGMWYS+BuA6ZcNStshaG
8OmQMpg8UQ+Z9pLGVUFXpMC2Gh/4jXG80ZuE/0/BIsjugnktcm39YcX1JFEhSS8sAetT5mHsgieh
0FGNhyV4f2aN69h3cQUx0/3txbzJIbcwbnvcFb3E3PdiENe4H1KLVBJ1yzWd9DtxsL8yDugaGvzs
tBPIJ76CX3juIS/Ni9Dnxtq06kHKHhlr80zyRxvSBNNyMu5jOM7UyFZcH5g7Yp2KW/cM4HPZmAuH
Tl4MEtWf7kI8Z4OGfa7So2HP4vfjiS7aJgZv6kK0Axr3/RF/u1v162fJJtnHySPJTzpakt8uwJLP
ltf80yGu6tGmJMIrYkql0NYJXkHOCQUEoPEp2zeziVJ31IJNYHlSFfMv1JGZP6B5R2GLqUka4B9F
f5sCV0iWJ5xWs48/jPklZwbdRZDdFSpjeGvCPd4KJSJauZGejLMU6hw4EwqYpxjy7nAxMxWkpxzE
1DxrHssn5QJpvfnAeg50Ty7+bRdBM4oTmz63FItwYBp345C3zUqEbZiUnWMbjL4g2zFYH0yArY6b
P2VP4AQJXA5onVTGqIv4VkleJ93CrmI9Br/5cGJU+Zjzl6ZyImqn5Rx4K71POAyjGm6sPym1FKth
YHG7PQsTYAmqUiYnGzNb5mNsREXCNnAp1NYD5daeQyovtn2WnVo/9UToMlpB4irk5gLNwxiw1KjM
u5+1n1/9ias8IuJenSsSCfTIYW1iWliQqKV+nrFjgbpWZmXMWduD0vdaSSoQ6Bi5chZQDqqA18PD
w8g6Za81m/4AHj+LUZ6kqjZNKtnwg6rb3z6Zjw8f5w75XLZVpamm3OOWICHsrVJ4FJrE70puEqd+
cDFjLUT2ljlR7MCJ7fzz4gwYtmNizs+sV9+4gAwrYizbMQIu5IxSMzyXtGktBpCZwvjG/dyQN+GO
nzB6F263MmlZdUHcyqN6g2f30vYPFaW8HiTyyxJKu4ffD/TZBXqrOfNQ6FN0c7nhuCnji5hdi0Nx
wsTkH8i+qT8xmCYncV/0/VdLI8CWxGGV8riAMrtFLFCNp/wYlrD/5GgAuOrJkjCCWfFdhvXmySMY
GxqFn/iLqvJKyPoH0BGcDCky5XTnQqW/k8pTPZh/7Pfvj15ZoJPpkOB7cGOuN8A8xxgp2qNsCn01
ox7bXSXbN4sWkH9PYFLaPvm7jYgHZzCfzfi3w4N3IGFcvvBuj2mnEaxyMr8EsvMjg2frSK88zY8y
kafcK3fmWk8mbLGqRclroSuW+xGcTCItIrIBTZFIcpRdmq4ozduYiduHRawZ88+4hVyfMKKADD1E
DaNqtwDCSLc+Zlnk/xca+Loq9qsYAdDjbxDGk24lRvE7PREabelCy47E1CyyvrG9wI7xrFfQl/1B
UJ13FswORyeXPGcGlq2UiLBV549J1+G0ZCk/YFEbhFXyTmHkSY4K7aK+OTsdlQrZv9mm47xNcWkb
R8rFqqYFzs65JK3bNwCqmvDbnJ/4prL29JuVV2t+01r6oGyniR8fkT/hoFh+ZSArW082+p5UwWmh
GGbn9W4dbaTyPPOEQOtZaXkgueNvkoNVcz9xf6gUGFCx21+O9cofJxwQg2cB92iH2j1mid9VWfjF
ZPAUHSsmmp9M0AJxJZsj2rITLJZFllmiNAedqD6R4oRJTkvlkulkxZvrt8hHcHbbcCLBS6pZGSjn
KIeZ65ty6heEqjeXdOplN/WIdWAw97+B/0jyWkeKfhMwCZs6hK6JqBZxsumiwRyBMpl5mn6fSdwb
mIxpW0xP84/+9CFg5KttHrGOTm4ZaMnBTTfI1kKAFOxsah38Db6aTmn5AQufDDsteGoT1t26nU2O
U5cO+XddshTfw2FrBgaKlEzY3E3O+opccNxb/6d78eHzS2+Mf0XGctNfT5vlQL7K7hgpODQ67Sfh
uVeWfXl/sWPma090WlCyzRkJ/SZXOamwvMlfMWABbaC461iupoaGoPhRcVzgJpex3xnxOfg2hkZk
tT3eEesSea3Yc45vMtojIGGdntaEHlnWb2kpoGJmYv83u3zi8Mh08iDo1fDUycK6tSl4vfrCwVXK
1PreU2agVK6u2cKmHFfX/4ZA1KJSBvPE9l2oWOWE8X+EAIVEWEeM11ETKaBEbSIDjJz6E03V8JBj
xfduK+/R6avhzFoUj40OWrJjWsTPwVsu1WKg5F9WKaLhDWphMOlTuBQxLib1nH8WQOhqjgxt0vgf
uC6vctKruENx24pV+S2Pj8W9Kfe0WfkTy/SERGajFTl9SDF2PM6vu8uVF+0HXjc20eWXKOPGjA0b
f/w40yCof0lbUSywsdBEUjmsrnbVN8CWNVRDBHDrOCCCEzpHxEBR+Tp3+rCEpJiD69VUM2W/RKw5
+GY7WC+DOiNGFa9gVeB3cxAfL+0LNqmtXWqx664AADGsdT15cZhTlBBzOGz6plVtIdt3ahM5I1RZ
ftz2krkfP7/YdTT/INrW0knI3/tC7bpG7331pcFoPt4h1N+rhPkLq4U9QWUCxmtHi0JOFlE55Kvj
lWfpQ6vCFLxE1jQHCZEAEQqjS6CgcY6F5rBRul4cOtU6xsSAnIk+iW5GAjxAngVAKDZc8uH77J0+
JPiVauxSkwgjZP9FP0PpMsNJJX/NkIwfbLt5JQ9XCqhlncxEfnbOqGXDreq5ftUeXU1xDC0O43uu
iZzqAN1shx4BzleBdDRZehzULdcN06ob6V5vgpXURVt0FLmpnbifNoTpaY4GCPT079YCBbDzKr+6
MElh8lHUaVUAv90XwqFIEj5NOkfERsOff/p/logyV84fsbJ5A9jSik/taFkMJxH47nOe7lWPheW+
YmDs9urMZgK24g51hBHT+opDReawVTGAB280UYPzDmMZOtSVW5AeVBLbqH0EpC1dLcqE6c2HKHGc
tiZ5FQy6Cbx6FXSv4bRG0GqUlvtLL2kk0CYYRPxdiJN4LVI0F3TMSitGB7jL3bScVelrvgXKzSc4
xBUh/ARSaO1gaNrZAensaoR97jEj4VVAO9UDy0rFqsOsgTnMBo0j0QE02O5P/7VAdlORe4ck4cNc
K6S4MWHHbCfiduwTroehW4r/TSnq39VoUMTkkPAZ3V1OADL2avF1Q6OQTswZtVHsw03cjC0Ll1uE
2FNr783q4+kt3b5XHhQhByW0zjBzL9OEF9zRzyQ1u+/UcMlI5YTzXk7RCohxiZY/ir+wbnc7XuNw
bVrjxb0DGDRMoKMVa/VDq/W4eLKlNcr4pmmNIMlMfBHohnOYKgju8eAVe6LVqa/xoKeD95ur6rB2
Fhe8t/C51yOEjzlLp85JLPUGp83PpZQ5HID/zEiMit0RRE8w1CQpbQHn5utizLbbyhsV7LPT6nL0
vhc9+Ak5hzY7S4/z6Ro60C1gHBVztQmOzG76qBU5YcJQow2iOsUvASEDXgRNma+gUW++IqgQl/8Y
DP1iU4/vpjsGtyM84ThUxxgQjM83aM4S14aASDDrANOYYbFZQlHQ5AtCIJP9iNNn4ayi0BLOK0oW
npgJGu/kEOHlUhPWuLT33qMLXHnKWwy2Pz5n7ENinYnH/smGONdt7/dFcpt5GepZRN5mq64qt0wd
TPYiwhExfwMn8hwBD7onBNGG2IMTsAfkUtVNi10vCqDTu8gs3HIpQrg6dyJ+rqTL9Pg6kFR2tPib
BCAR6DXx+ZyZts1DGc8Vk7kfvCZYrcvwNFkTOz1XqgknvX8mTvWTVBjlDl50yHkktrt0AkJs3XuT
Z8w8d1F/be3CFLMpYiD5bCsM9rlSGGPkqrZa9eAep9uGTGb8NkqEhLxERbtmZDKphAxT1cBxs0yt
ANXe/Vf82uVUrZgUtM6ZPmeyLSXgEJk3IsbSB3wxO8pCl6w5SzfFQz0n9zwS7WnzQBz4hGycGo22
dQSwHZaZzVOHFS9ZKeArlOkoeKZ5KAzzU9JAWAQnRVAWlXTCeiCmu8AKd0L7eVh7KLsbaPS/zhMa
uzYwriAiOWGJ7qmUWte/NZPZ/1C3RBcKptyv3y3t98UyHpXggI/Ej0Z7RfeOXM8flOFsxwSMuen+
/KKnTFSBrFNp8izJNGt7xFhYNAYXrD3IUOeRmjqLXEiD4wV1FALWAFbpXvYsmuh7f23VJvhDecMX
Hgyld4BccPcI3mBSF7wMSmCH+RJ5yOREpH1+a//zhxEuA9MiaI9DYOCTUcngKb3dEFR6WHW8QCEe
vy9yX1YPB2HdpiAm+rYTCXd9H9gTSH5uPrAEb4GN1Kul7EXIma5jRaJAlnaXKJeoNEoVKJRzBOCI
z6NKUntVac1E4nSnHG2Pt/xRZJlW+GA38NKBKt2DXNBGi/cSwsmggLdt2JVDgul9nwtsAJeFH3ud
Ub5Gmo3mbfdFPxOSnhv58WTQFgRN3eWCIPh4aPQYwMHQdKn7xT78VWO62/j7kGVzfiYzO1bbyQEt
ejuvDfFwsLevPscQF3c7lEO7RgEJ/I5d44fVwN/2diBvm78z0YeSqCOGcl6y/FG+E4GD/r9sltBA
E1ZQPjMuu2zAS9utk7Ni/GM3GuGdOmO8qWT7rrnSDoHTL/o53JhY2FeKBJwJwhd2hT4o0mP1n0gh
nRkeF8190aB+01gYPXsAjiQcfWGk1jQ0gwQS4Fj0uGByc55ZkNNpJyVCf48qv5nYtEjyFUZzXSr+
V2HxJydYFr9QB7J8nWnYdhAclP+BCjxpEW+yxusEw1fbLGS8fs2NONefN2a48Gssaxf8XZcxvL8V
m/X8Qo6tXdp/DQt5r9iKBVtOU7CcwHxyDBeXUVfHqobdfQvUBJ+HyLzEOVrFXcFothuapqivlVhv
t+FhiqBCVWLx6pJSPDb325NfF6E3vbCwSvp4d3Aq8paLD/tYp3BMfSP40TcQ3IHyk8OLhV+PJc8p
OyRJ+bYXijnjBfZOyaSfAZw3Vv+MtQALmS5mkfe+QQhr4mwW5vKT7aR8ARFBR+BkRcOynKJ7vQxL
2B8qnuD4jY1exUaiMIKOfe2kMwb5lRCq/9eEXP1nMDWe2FJOiy1fHk+E5wHvCgl9i5ktTRsjx8R5
fVQ4ZagjSk+5he0DPj4BuIZNmIzZpd9UXzyQCCncMHyMio2dVZmar/9/s9rqIE12hL/ay9wz7Wsv
H3eOHhhLDrCytkiVpkfy+n5UNJFGnLrSCgfmw9YTRlN2RIVeQHnjX4Ge81s6Gpn6YcaGjh5911wb
5mLwz+qrR9ri0ATPuPqDgwScQANvli+RDFbawFceIpvYjFThS5xg5yNvtRp/Go+jKvibzeXwaHUI
0ozsJC7DEQsup66s2lWlDnoXSrTPdwmf8os95rSLl7LV0DdRXskoeW1vpXUeKYBmpQBLZ+FXNCPI
EPYkSbdqE/tGxRMn+HHOXjd1jYvgsEgN3pljzQZqVIL4Q1aWqsgK460mAW0nm2RQBZpWX2aXLEL/
zLxqkLjMF07DgAoJ8X/U827CAStQs81sR3wh/HpeFCbwqNIHS02F1SLQL0mBmUHOoknAxDH9qHvX
96kBIIfaKDcVDcJG4wS1+RO22zjT7HXqDTYhwIoIGjgk1Gg+AKqEg5Qw5PzZCHBhiZF+EDNnWxLN
dKScZws8Ee+oGX1n2kBNlMGYHlcXOOzWotK2Ksr656VyI5KJv1aru5acVmCwhjJQPV7cd8Gqs9Va
rQ4QEQB6OMswi5xpCLaBzFyqiQ6qs5kK2q/A1UfNClnWhWg46Meo8x8ME3SaPijPuJW6RjEHPYEA
1J8FOSqv/Yeyl3K1BOzJ/eUQPuy5B7Fz0angT7vXO10VNw12PXT3wM2T+sxDeYl/bfKoKIQaBx+P
/dDySc5YYaW4Ahl6E960qW+yiE3sDesE1QtnCXpH8vXWWEK6Uj6tctnSQZX32+lqi4wqU5Hv/k5a
VfDWqxd3cNNnK/XP6Qk/2cZSiWHYpBng3JYyT7f5UAlsO/pQAklAAdZyN0g78z9VhMyX5uAxhFk7
sSo80R+YolGTjaiCUiL4tGt3fkei2GXIKND4mfjdo0XA4n65q1B3TmoZpe672QloPSuyh8VBBqC5
XthlSGD2zBzqCTT+hPTLV+m6zvkmhBcwoOzdJbdZ0ZbFipKZoXwl2YRdU6Lb5OAma5Khbw3deHHF
oKhtBWZ0rnRz9EQE/YMamgiP8lfNeJnHl9ruTk/g/8U2b7op9i9yrdkeSZ9c3SN/ABSSJd3/AnPA
qa4KH6CMlbRYvzLSp+HSr90FB05/GXsYk/x1uAzQLGi6iWgCwSR+hNxPmtlpC/NSOUTDk2JqDVYa
vNDKQqoebvTCdAr89q2dqedcg/RYseRhlpLmrTsw0o3pkGI/uXwJ7FwNur+jKJbsrkqFbAfEgSmM
A83tId4O0L+A7fPmn5QOM4qTSf1DkH3Zabycaw7ZdKeSgH41UjmNXCD2knCd4eF2R3QCDOYfaiSV
BTIlFNxNhCPgcbQixt42Jsl3eEOr+hNYJpynfNSZ6Ydy4Fa7wx7JD2MSRHlZM6/I+q20QZtcNidw
T5mjtRgdUa0sRTaxWBLpTZQRjkcVmSwd+MYT+lZiFzVQoxpt14Uka9feUMcQVSlzKJSCgbhhJEp0
rXyxnysCPnHPRztckAzEbj7p4ARtjFeZcic5LrmGkZ9lMkwglXtXwUC9ZF8/7jPxk85heW6WScgr
ribTcKc9vbZf+tPMuzbrTTO/+cUnhVPlwcxeOahfusCIVYoMK7gi05gzUtoFh3Rt9aGEIYu0KXnZ
8cENbToBdzTj3Bb+rjutIp9V1hee1NpVlqPI6BWHwK2oCb7whuEyZ4DMO1YQehzmfpC3Mt7nbWtY
Um0GdyqEKMIvXbf/pebN+tECxd2aTniCgDiSlwix33tSVKIqRvFWPPjl2EHi0K7QBHSK01b8xR63
4sWj6l4SiOVgNZxP8mkrMR02C7D7aJH+OHmfz4H7nKYStF9MOfDJnyGtu8MX2/MN+4UpHsfyl260
RXwYYntfNqgf1TMZtZaBSrYbKt7v/O48knNt5UDAvyIScMQywvzpLSb7yFZgAlpGjVoN1GunP9T9
cb4rc7XlCgNsLhv4rxJ2S9vtagHeQGmf143n9aCNKNdyg44LoQXfPdG2fOFJMsYh+Kb05QmkcPNv
S0HGuS0D3aWDRy/ZSqk6fJ5YlB5Un7RpkKy09Kj2A+2PBRdRIJdfwvRJz5Tfy02G0Vp4iaxWajc+
zHlkJOy9gGtyXkVea1b4c2tQY0SRzjfAvst6IgI+/BH1tVu5tkEfjGmD8FV2Y6eHlFOqYJfnCGGR
dTgua1tWg+alEECs2ZXinoTB51Yn8/LWwMnRsKDpLfHDA+UhBIRA6+tWTnNCBPDoewTy4uXTchow
wwDOt4A2HZgRySJxomxTUQZ4LK4myX5JeabvDYoFYex1yy/js8zU5CycavWXAxV+2tAQ/gbkEUXx
ivbuhjtGu14xI6zuoAqtbWTLDJgGImzqtwvRswPPaX85hI4XApfAUXYu2cG3p9IUxpxN0DMWrJlM
Ow1u71iBC8cXelrnfb84d12YrVXrpoRWtf61EJXHOCEPDmMBlUjVuaEkHI7iAb/VXyKn33j5cu51
FZo8qqg9ApoDWAeqs848ozXBF1vcxj2av6lT8nLQDEHxA5PDByKIaAH2JbcTZJaZg3fpK9IuMfZm
3S4GgZ68dnokyZibxpdvWOdh7UeY71kxGazw3KNoOqQmlvUbLijumji6BLV9djZ5aj5ivoF6kild
vTP73r/Z6Wl1eAPzB06EQZatDxS3x00ncd7Qdrih63wkHT46S9WAjkWgi3NVpkECSqdMr4hNZ1dh
GO1zoPl/0jSXhDwID5LdT0fXEB33ZDvtVcBUEb9lOqMZcFsRYQOrjZbuMSaYDa9ND1qG6sFEc1Yy
pgXArMwkZolOf7Rqs9sG6WW+LtHIvkXV/zhn9JYJuEWB3xW2BeUnj/mEfnv8vWOCLa65gmBUIMsh
ZHDD//PWHuuGuWPipCR096K0+VVd83F1tBVlFsdFSmamVFfW0hiMo8iBzg9io+mmwPM9mBf4HT/h
Tbd7Pzem+N2+ZZrRxlrZJi8xsh6JlYJuR0ae4FYUD5fo0lLDkQ/SOApED0mzaqcAve+A8fVk8ZUN
r1pRt7BBETpa4yDE+si0PlLI5/Y12Hixf2efx4rC8mIp4KraJThZkJ8OqoFjMG/BUdhB+qhUxJo6
udbHcYTMsD3YZSx218DhL0jBHvdIr2p6/FC+edKRlvnbbxWNv/5Bvnz/Cp4AQ2oG02BtQ1CF7cjp
A1/ThuL+v74KOIt2dE+Jr/ZrOhY9dovXmCfX9SxkxKnCOZD8xqtwSmCmcaONYucj+Zx6QoQX4GCa
z5yxpV9dq+QD4ZpjlzUZNB8e0b84Nj+Aw1YfVGxvAZ1YPk5CYH7GE3yh+whhfk1GRDBkGnBhAaDa
xXXMSdWOhYE55IWM+9TeUjRs6Sv/gi3PyEcohG5XgypVuBVHTuxAPfaPmgU/afcrkhdNs9Ey7xeo
JmBB7+WqmCU15O7Ofc8ytTwz0M6oGxzeTWAMsjWU5Zglnlqwo7gWZspgc2DpjqenQzH1VP5oZXPt
59SwhFKUBxdE29qdXpYce7HbT4R5u95D/rGlR0SQAgPyD62/OC+xt5fLnNN4wD0jDQSYa87lD6TD
SJMF53i8U+ZBmEf3sCZWGcohrUVHCkr882iNtYXFF8UqWGO72WSjnFH+sxFR0GQ1VM9JL9eKm55D
ehqdgenwUxpTNQ80HYShf+zQsTLYohWdOhb41mXBSNKUCFgV/xGvxHAbfOcOhpdLNdTSeO/w5qsT
BJ1vTFGAbKuRRKxX5GyCV3QCHHkh4SyV2s48EGzhL5LaX5srSvGzf/mCRWoSdsim0gtwo7z+aAkK
Gz3d4/M2M58Cjfxkpuqvk9Xfz2BSKnWPl/ip6Er8AyQgzWMWzz+xswtX5euWJoaAjgMcVR7zCG3g
2z2hr6bQgavY7C8pO0M5z+3T0c4LtFcHgw0byWb4U2F1j6dVZCbAJwRL7Sd9XUXYri5seppZ1hiI
BKYt5e9FJrOXgiuXNesP5iiS0Y1G0uvOdghwB9qu4dkzhEKT9VZDsxpqhYppxx20LoUQ7xtL5UNx
+WFJkTpEYEvX9EQR9rj+4HL32PP3ma0KsLK7NUBiUKTnZgw8iLGn2WKRkkwZyjHf5bwMTyp8iV7v
y4qAcQ1pre+nzYMLVzQC/niNSmo2Nms/1daobaTLcTwyIaWCo2QfC65bVTEOCWlp6DxSGCkl9HHF
JACXQWeWBi8BeyjgNxbhcZqJxndSBP6d7Zu8YQvxoY+1zCbAe06212/EMTFCWFPIARsrmX1GKZIP
Tm1Xboz4rqrAHwwZ9xot6pjcrSsM8sXCwZ5F1emS7i2N+BGpfbGHAPnpFb6RJKbreRRY/Dh01k0F
jXNeiH+a2BaJNJv/yb3dnIxPX9SAroEzO7Os84DBUGskdVQlAPDgaUqEnMThQfIjVbDTdmX9nwig
9sXvJ7tXz8QUf39ZOLC2uNiYbNHk22xYReR5XXKjNYcr/O1/y56l1XdJKNwMsHOQtjWwy8zaZbyw
xhIGoWjvuggvRNkMCyHuIQL19CeonDmhR4/xJgQPA1lW8iUbNzvWeROwQ2haQ2AkJM2LNld0Ig5G
5RR42Y9pI6rVfdz4ZN8mVoWo/gXPNrL1EH1mnoK6HzUhrHX04B9otbOslN55Ctj5uMYTPU/DDaGs
DxI+yg/4Le2mGqw7pdnpLNj/p/7lj/hMPcwPo72q668buw/XYZTriDEh9+6HMMk6X6KaxZRYaned
qxRm7acS6PWZoGefaBLYj9MT2Gbh5W+IvkXQB1U6ZQI28eKPbo1BOMs2BXnpN+h5xeeMf/p7rjWn
4lkrJ3mEebKqtbh9vS68qQodZ60LRgLz5yLNPMDmZo4tQJlelwRcE4V+zGHCI10vZmRUM7aJMGgl
o16br5F/K00iOitFLnO6W5NaVZWRO78Ix3YtbS/0/uu85ws95Jtd1+aYX8OFjoSRHhUASvfeW08K
wsK3EetWDOt6cOR7qVOn8PZIL2iRm+uXTBac5y7Xvcj2Kp91Uj2Elc57K6PnxIQ+EPI5gWbJ8cXl
9l67oMPyRY2M7r3x7QkinYafeW2L5/5FxhfKgl55NAPTy+q2DczQrzB63GZq0ccq55LJkqbmojLR
YuF2IYQCI+LfIyU+HbPesQob345mxwx9VhIzWtBwUk/uV5iI4BJF2P2WtPpIGh7hymIkg4NPkpCj
sP2P2/Lbr0sXVl5TEUT7DcdR0CasfRrCjLHbaP++HxZtL3pQj+6WkojlwKlRhKsefF0jY2Wtcwe6
fpMJWd2myhTnrNH2lzZAOpafO9e3f6ErI5OfVYbnNQxfF8mkSzuTXi1I5zv9DU4Z7kAi/EpLWZ9k
mjLE3vWKqzL8ESgVKB27bbtW45Fp9YQXLQtT4wYYFyHmXDrX+EADdl5GAIoOvOpcQaZT8y6wMT2x
TyqzhhYHlb2MhiXCVMMgLRSk93zqCgNBXe2oVOIVyH9AKG/nD5RcMvGZ0YJvLkKJKxvVfJYZnANK
QnuAitb7Bbgz4lUzb00JTtPZTZwSJx601HSeR5XY9fSSlCSh+dCqbJvMIVFyUfiTyG+sQXQXuNDs
kK8DQ5qzW+CNTD7i+h/plteH8mkGaR4IthPEKMZ/GVOsldQuAMTnv7lzHJyNdX/nrx0P3u8yPE86
Hze63P2T40JyrR81AiHN7R5SiDShG1HDDrE+LFSLLBZmLaCZBYisGpFBjCKjTCfH64ozjuXthl0Y
4klAxd51SytwLOZP3J+4zs/X1TGXaEnyMl7XCn6Xm8O25/Enl993F2n1qp+44J3uq6mk3cZpA+IA
gAgIuGprBrkgdu/QAmUQ6nZfOxFq6APko4gGTuP5Ff2loK5CrMhmRMWuGK2XZGdSSzJVYDDPc40K
CYwo9GYm23/TJ571P257iUplqR1Sa78bsstHX5uR2tMSlIkeZqhqRgiiPDc92Qg2ewGReu7MbAGE
We8N14JCzTuN4OmFWvwG/3ziTykB9NtU6tal+RmYJhcdxUXizhZTLuEchEuOKtlPhbGbYq3wq64s
I8xWn13wK88HZxPBhtLTmilGd4KQI84gTU1QRfhKG2FGinPR3tVO7f7+Cw3JiyOaFAp845liiKD6
TWYmkCJ3GDfdcV0SpoYGHPKTW3vN0dVufJHqdeHdZ0kZoY/Hil0Ev2+sfCNFKdCgjIVNnVEGQtjg
TxLNmEnV/gZJrASWR9FlYPt9lpw6MGviCDEoZJQj0ysLqX0QewR9By3e5MZ6yC6cPWM7ErNvGUGP
TDKus+Sw1kHC9de4K7RU27Qt7VqTAYNy0BfYpa6mUBhvUJSRA3EsmDbOsS3uOzqR8iamJjfNNyVc
yuoXH+OMhHLJ9kndAZ/3aizi2NuMJ76loxfpgX0P76caiRnJtEfz/M2mcY10Ukriokl7RC9t2F8a
wA7X47UKHULpgy6xbQn4TcBBfKIDRP33Mo7tMD/EZ1xt5sThrgip4twoiF3bwBVOK+yd/yP8eFUH
CBztnoHefd4HZ2kJeLNQ2dzsJqMuP2PVoppeYj691zouBnfsMOD9FQgPZitdHFNRiEeeCeZYi+bJ
Lpr4DF43wYrd8JpATFkbx/FlZ0uLB6pRUcxJwUX4E4TwA+YvLRp3UUsM25j1sNZY1kCWUZroMvIE
sR7IpCxiO1vVoeNMED8GCRfwPpEIpgfpPU751DPjol9HejUB0Ml+D+NrDySOoImy3g3TcUGW4leU
AVE9hSX0p79U0aNOYdbAGR57rgogPTHvBUGNbQ02V2MbGuVqwqJ3qteWTubN7ZTQ0JSQ1uPIdq23
/ffYNAr+iMT2A7qA9miDZvnNTvhLCeD9wEb/U8oN6L6OAkLk5xwqwgZ+kjQKDakybU6NSa3pjDMB
X5es5miuulq4LaDoRpD98pSTYCHSkqE8DbNBdynDVeT0MaKqbkNLbSZrFQkntpC7W59EhSNyX8Yy
+t75Y/+DDJwARtz1ZCTprDJ2XeTvIOkA0yVRG2uRN2hpV938qpw6jXFzzdVq5zTkGiToFe59NAsM
IZI+tDqTeRADslv+KiWy9E4ftbM3k+SXZPiweSA4eEBSvUMFNshMPEhR8u+zyPyn7GmHksrwiOvy
w32rEFHoRsJxRbm5QEOKd3CcxND5uVPT0BdjwurPk2V6tahjvqQBuFHgDGbG+0lJdEkq4dVkOJ53
nThHjDuNDs0mphCOq2mumzujVeSPiBX6pUuOOr3RByjXqD3UY7Pq6EuLIv9gBfhzhpIxVw0JYkzJ
tbvSZ0iUmeKvzWo5WpzHKD21xDGOATp5KfAGXh/1kfeVhvMNVR1Ni7VIW80rnBMcxkngjx6yR0ny
1l+JuMJ18lV9ScBCBN8EeGJ5O/12t5fNYNRKx8rAjZZQQlVJ9C52JjAoIfPwQT/cBAyKpY2FdX+c
JbYHqxGfUH4CpO/Rl0eEUyyGMcQMBRHe3Fm2gqLUi8350K1JgLwBRdLXouP0NvodG3K27RDKiOy0
DQ/uE5Zann5itGceR8J5w9AVyd6xxb4xIUP738YRIg6Y5DAZYDYdjirBSGoMb3CK/XcqLAbyK37u
w/UhCMjs1eUkPlAYQyHbVrjXp4QrJFUL85ssRS4C/2Olsx61hG3jKNyqfnAgKPsYdkJgIUNdxcnd
hJLOJcELVDI7BwBbStvhwsq2vkdvTiDOfgoQji1O73BJVJxxcOu8nLHs4TwARnbkXhbkZHkgcrVO
ZRauZJuHeMT0ZmdBNMB3ifg0tjABfbGWP9snwKZp6x37dsd4F5YNy229LgIpJsvhja3frjES3Z2z
YTZ0yuuGX2QH6MCz8ie3TckMXCzpgVvjZrxZa9FfCWPHLoI86ZnjFf+MNeifnAg+ADWzQPlMWq2I
ig/P5zZi+6chI2UsGRdMMpwbIArvU857+kU9+prKzXN9+duTswYAFLPeJg+lA+IMlRSsq/vivE9K
h3BXwWLraERMUl6qRsc2yB3ni6wCM4RijiMen6XwUcWVhTB4CK0QCb1/B8tYHczLASD2vZAlfDHS
FW1ACGzFgydEgQJXLlOh7Hreuo2zT5nvFOmt7VqxYJEL44xjsQUiKs1Ul2++wFy1iZgWE8Xp72NP
mN5N2goIYGTKSqIlkc3dQeRMnZW3RD2rXQmrXu53YlErHlRbFD2flxD3U1+tgOd2cVOedjRym3nc
PLaHb/AJQAAn/vZfLynDogrdXehXMHLv3cKSfgEL482yvgV39qkU8ws858xCnXUzOqqlNRvuQZtH
tuWk+hHn26q+98MoY6VlsCgoK+HsKDOVOOq0gMBjEftEmhfcbzEwXgzHN1rl3+5evmEBfTeUIcEe
KT+AgOnbCRBOL2M9iGnhxILmk62AMs+Mh6+Ya8LkNfogNLk9SDLVCYiEyjgXsAcrjXLbhCHlnmN3
yhgB6/HixRld4MCwS1sbT1YjUBbycNN44QpEy9wY31uN3YgESTIizXHmQ477mM4ypSEmTDumDlM9
QQLpI5YqwUncSDOE8GCjAZPc+NiA2Bg/MfqjWEC82IVBZFGxkj57SoezE792crlKyex8DJIiXSr2
i3P/uiu6RuAVLTEcCw6iVTv7kC2q8mZod6WTrAjhVbXtwROXmsTSupBzEUcDZa4gVrjPhMSSH8UP
lshAXW3SBPIcHObOvtlex38TafGYminhy6t2Ho5Di7jTOkR8AHsBIXImoBUsmT5OTfY82wua0GJi
LYlRRiWfHwSrmqxmNHPsg0xGSJsn8liE0N9HoYFYcm9KCVv8H9tE2Pp1+fZUXeb3ywSXOPA3Ed+z
n9rsgPT+1KKDG/ucH23T0aHbNlIchQ+nlbOrIkc79Y+7Alj2zrhqZo5bPpqejwdt97feU2AAIDvL
J0NW9fAZQc93I4OhpDsp79DkkBKttOtz7PCCygK6XAJl1enrw50Qe0DjjI6ypPS6qQzkFqdtHZDu
UHT2V99keSJxYROH8G8KFOhVunApz12h0xFr9Gajz20fdEzb3ExuxTyys7HXXsl2kF0vSiIjTxWP
PQ/zcSggDsnLMzbG4jsmEGnpYifcDxFGnxr6BfyAMG9Iu8m4PTIVy+k7CgKJlDcmx6Xdefyn7Xnc
9G/UF4QZqLu/Z7RRi9odDiKMNqJnduO7iX/0shdWsKciUIIuS7R1WA+N5FkPZPAz9QPVcVPUyoMM
vOEmKSpqueLaJqEVYOeexLR2tG4E9vUIxQ7H7d6Y8BjXkz1kAFg9etwtK00wNfGARnVB4NGFC7UC
YU0GcZ4FpwpD0/qfYWwNO7G+m/wn5EktH4DxCtAtYNW+w61uV8BEcdKyTXZnQcMyxM+5OI1rnsom
2qCOZN7i/FccqMQtHh3Q6Qujju+Q5pzh/9fhi3CdLbyWUTD+rficsT7K17JjyTHPVlcmCdH8m/ES
OX9j3/nLd2F4NEg1sV0ub9y/xMKMhnPSnrTChQexrslDUL/uC4iANGJQeDimHvuxgPWaurfs9MG5
YVSUrLz6BOo1w2Lx/0P9WkGtKIXAREtzcPMBmtJPJlogMJ50k4DaqrxSFJjT4WW2H2m1F8cFW04s
rjPlcp/csCe4aOOaVBc9WosDRSfmE1JJddpXQgZ1c7RnP1/6zT8VTdWqe6Kgw42Q/YMHFr7yFeiw
Ry2oDapVW7Ee9eqq4MTDgsxPmZ7oP/Z9zXRz3Z+TFjZ6qcNTBmNPkU8jSiuncRdGe4Vo4JFMmwie
Tdb8fRYjCzybhil5Y5PBAlhHL5WDDmSdHF9o6rjX7kD2soB5vyDpkPdhvEEG9jsirBsI7s5ri6na
1H6fLk1hy/9C0SvoTXHpIpohI8Vr2ZrXdXb8oJK8AQhUgwlwzTol//bjtkPfcS9IXFybGPzqJx2p
DLvMIVZlAiIAg+Wy9zhH/RODVmoBw7mypSpCsH0Dawe7sU+c/ZN77l+hMjiXTQ8TQCM4YhqSpTMU
EESief/4o8HyQfnLoA2xzX2RNzqZfHPEKHzCz2j7MFwYPumSo68SQS9Xwg8UINsJ7TmwYo+v+iDd
FF0q4ehNFHnd62LKisfCDMaATpWng6awwK88tP15Fgw2skic7EXhEPYMsvFBFJueVZmjDznOL1vv
0INuBeu/D+9svnplQxRfLGxHu9OBUwzhDrZ/NEnZroVBgEjgoqcu7/oiNgkFJCbExuSnTmnLU7EO
vsTr0UK6+HRxJZZimaz0cnOZd/y237JOdEVI4HdHDAMQ7U2cMR77fNHgmON06zUZbUWMvqFpjsDj
2g86+paC3w4Fuc7YaJ57NTAT6I29bz62gIDJ9B4rQ0WjGrLZnz7RgZH87dDgTkLe/OvrRu3V1Dqv
jBdAaevZGK5YGziH/9wqF6NvrDZ417xTx9SPpMIEewbjUkySCL+qG8zIm4titJPe5UYxUeIcstB2
oES9d6tWyMchOxPHTG9ZP31Ca8wYrRSe9MnkqFPVFaJFjFekvAsevtyx1UksBQG8OQyQFF1difw7
qqc0RlVhKw0aqUJqd34H3Htpq6qzyJY2ZgcqukdhH+7bj+bx91xZOSHop82CMaXTYYsGoGuLZIbl
pr7twAgj0I6iRhzpMxGBoUY7tH4qvOxpz3xZMlQUjl+dXXpEoCRVYWzzSUjKDaDHdv12aQo9E8r4
zyZwgQIcARmFYypRl7KYJvQ/IKSwOCMs73lCpkzM9sea4qWhsDVavqTgccrk6UACT5pdbmZNv4xQ
/cSor+qzWzUqEDlP9QMQ11QBU4RP5Ft1P7Edt9MCP697npLGVKKW9B8b+9e7SIzcd3lRBupZKX8M
7omwBRZQp412UkO38lFS7C/9WLHGjCkqw/7mrxyWBAQgr+3PpPLnO0Th79cVucCR8j1cHSUaYWij
k2Ya65pkWB4BSuzm0n3xegJ0J5FNhKBg4ldVBArsDzi2I+L0/QWI+fz9oVBbFy9RxltjooRGclWd
d24CX0VQZL/5OPRrYqERb0fPoswZNoQyOtsAM6dWzEgrPm1eOBmw5CKIkbG+sMKrW8LONVReRcfp
lfSiJSyE7qzzC35QibmFXHPYd5c1ZoeX1eJDjnAojIvmwinkmpmq/pCVMjSVG+ER3geRVdksXHTW
QuOL4yn5DBEPc04hilDQWV8C/gGtjzJekJe+yDHDQ2wyEgWgFLLQFjvTJQWVY32hlzsD2F9R5YVK
BVKmYCj6aSUUulgApmzZkjr8xkMwIQT8l4uJxfsB+jN8uoGFZR28vQIP4GSQ6it0Qwd64JaictkA
ZvTvm/9JUoHRJ2Xz2KVs8KxBCqOIXydwV7KdQOcmeE4Iu2sSa+CCv8yOfVEF1D6g9o/1HkpTjRa8
uyr+5sgSntCFUlNkb0FgTF9VCyT4pMzHFdrXh+onNvL19cc9ZNwjFmrIJZosn1xKsNr3iI+VYt6T
dPVlj1+pcFFK90SMa3HmdQYx2QXhdAkkIgwM0AQ0JcCRtUE/EwyFH10NzWSrWHiffEaSQf3Fn8at
bDO+5B0yDBXE2GIJVoRWXkkhinbPK92eQGV4Yt2JKyNvhWQL/V6+HQyZ4xj88a1kWf3OXTHf77qz
hSZzMrjxKC6YgLI1HQaEE2yyWVKpjE2Aq8OlhPcMIMyOvo2DSWIH5qoWQZguNyzG2m3ZCOEl7Nny
NJ+ltcbB/24GTuDXjv249LeLwYV7xKv0ajRl2T8hEAp49liS3sein3Hsvbpli2zLXvKW2L9Q8Vgr
J2CPw7Nq715ocNH0q2wdpCT7/RIljGBzgLCeWRZ5dercomOQgGPli0GsLEazKeb8DEJHD/ShecrQ
hlfa8UWQ0FfBRJT1khle2qwVCLk98fOQ2wQDedMDAhXBQALqFftRV/zX7ibvQIEsed9n1mDQP95F
Jh6StiZxDfHQGFW2RlInd5Etdo6ou6wr3fw2fjBr5O7gRPM9cipViW5lMYrl2c9VAJAmmni1jYHY
4UvixRStZfHQnIcv9ZdiDIFYT0p3YnNvyQ34NRcgcQjkvpGFa39fexlb7Oc54j+w11PzAoSqkV7W
MkEbrwnJLAw87wP4dgVbgOmWfVaBsU15ibn86bMlAzG3zRAZAvZ6AaJnORmuRmvam97dI3X/113B
5Z1qM5VswLdbrZrCgrkqVXL1sTb8J6RF1CcIiZMmCuTXXfpGgpuBFGtxTTIBbJYlDhRs4DIkfZsL
2r0j6s+oGJhfWk9bCikqLnLcjzTkmrQ/WT92/itNAsTys+FciG3haEMeVbUJshakKptmsaTYXiNY
5oY/fPuTEzUQzUeZLYWT1o3wM+DZfsx+poVoeDBbshVTZtcQ/2oHRWhj+yxxEbSKmFY5NW3nUbcM
8fSWqyJNmtgmGq/Pm02tQliqS5/GkevvsMxuNOUqNw8zSQKqeKgfhfX2GctQTlkQiTQYxgcjJRPG
IJdmdSDvStx+5v+TdKfZch+AhjXew3ijUj1NGwLlHxeihAOrUTlEvXwkLj9LMl11a0k6maJinofD
QtyED6OVotWLYMm7Gi2acEuRfbouzIs6WqZUR+tqt5ws5B0qMP73i/YxgI8jnaDQpAyw7cgCsng8
dpMwAw5uAGkpTnJuif/mjfJ8OfwlcCNNnHr7ST/Lzv4nvteBvJ3xH2QHWx8Q41sS127OXN1AjQUk
spG2kXxp1Vjaux78AyOLOB8M1Txf3T0+R9VSOz8GdpWHbnw5tIT+yU7zRRO9/BlctzcAAwdWu7CQ
a6guMGKX1NaFgyQuMawYkX2bGBegxuV+DnLHSfiChZJ/BLenaU1yxJSkjVkAcSj3zQA14K7dIvRy
YOjEts6t/KEXuraoxih172sutppldvoAetisEvUnioA/2RKW86PCUd/QpSLZQGELYpePw9uQUM6w
A/6aFi21mMc6ZE4dDCU4zTi7uzHue10LSFc6SMiR3f81kaiyB2djX367xS6zNSv5tJUx4J7YpGmE
WOil1eSy0CfF2xt5fOAd8/xQc7k4JuROtzeKxKibxRZbTKJY5hi7cnIcAtMpaXh53XriHisFh/lq
CkBLSlTEssI1imHh32rilEJOC6NPLdBhYXaSfSfg7lgIY69UtQ6X2B9r5yIYdCZm+cL+DPeMS61z
7M56Wuy4Iga2SOLkKvJxt6aayn5zIEl9a2z2ZVgjxTZI8tckRGhR8b1sO3vEm4QVwvrI9F+Hf40D
VZYEj7D1Vfni6Bum8LXYpUC9/9ZC15y18TfOpQ67Rfkw2QC0/7zBsVHqaPUHgg7cwgOyTk+jLjpP
s0HTe4Fr8x95zTpCGQ6GriGwWEBE7HVGdtWsKUmhLmqJVPvu7bUXBYtzxQ/qtOFhATsxFvH8jkd8
wHAqJvzdGWrbitZUAuk3EbiCkv5636EHFSZxB8ITv8Ous9DfoZ4i89Q4tRHCvVMiewUPvGybue7T
v7qScVoke2qpnRCE2TJOUWWWQSeWpXoMKJswiPzY8PgDpeecDmABFYiEsvBmv6XQQdXTNAHTXPhi
U5oGOGZuKRatpPZ7v/stmWHB+WwfjtXwqbzs8Po8uY5WvzVGbvth/RLVocv+fSKtijMxHLSQ/kyX
IsjXS9m2k/xdrnIAVlzvFf/UUQa+ing9zFvvpfJ8V9odHpZlNIgJAFt+ufgqbEnoO0h4wqCCrMTD
kHINyBo0tjhdSlV9w5x8TERHidV7ZO8EfmPBiMdqJCBusYkS5IxdjGRUVS4X0DWvesmmoZ9umBEH
SNzITMTpukI6KWi8eTHH1ItXbsBgyiO1JRZBuPbjo3pyt/dSeEcrPcYmo4D12kC/rYqzpD+QeqM3
n805JxifQDojyXovFA5rpqHGqsYs5r/Z2SXW9xrILfWdEqs7hPydhyFYApQAZRs0BJ1QaWJVqIE5
oA2J8VNEkm2uUODXuZai7G7QefAd4OKBKh1ONafQ21zIkhZCD4VOHXlSIldugvkbcxR60YkE2Wtp
lTLTNr9zt/dvqHSDz0PhpSpg8NUcKPv22TECSTNnR9B0aqb9xbMuDSeGj3cSFgkzcMO+eGFdZqmX
xV9alT0l2oJiHaOv2CAlsl3SB2tKJuN8yOP7e38gFINM07mnhMcg7dy83VyagDIkvV43HsuSVhSr
6ok6qQQegtNZFv7n9NF76oR5ogviAThjBDUwz3yvjpPtplbJbgzRaLmD4mAw1IssR0zYslVDUAy2
gpiTi8Au/6usvVbUusuXUKkENTOZIJJV9SSM9nY0ONaSL99dY/xKxFT4ca3YaXM+DuNhltsQfSXp
0I7TZiRYKCP5EsIe6Nqwi0qwIWNjA0RnfhgHcWafSdFjTvpNabtSEyttgkicLJseZdx0st9Ye7dK
OAtqXytHwLaoLPptp1pxqLleEgI8SVVjc65XTQfVvDwkcewsYlhCP8oWBTEoNcy6TxwBZ4xEVJOP
RUeckM9ZcGEwaDY+P476bnOvClUdVYoLBXXP4jjYM4lYDKIarsx7Dnzbqz0nhfxt7TStE5FwoQqO
CK1XpgELQ8cRkL+3JwhsVZpoSeFmkeEmdIueIXHvEO0Nfl/QfBhjyFK4ItGH6Hn0xEDdmaf/KCtf
WUOJX4h/XDcQY9+RxNlant7fN4uvctSv1Ao4+pMu7zELdcKX3whGS40GHSjHAL16FLahPvNG19mp
+guR12aK4Hx2AbBK+gwps+X9CrdhuE5T1BOD5LCwix8RE5qPF7DqMz89gmsRwdPBEUceqmYn6fyf
eRsNEZl9W+MZUqweZKkCDFIW94GpMCxxzDSAwk0dinb0biIEbN8VU6MdUD8K4pDxwUIKF1W22zIW
3TjvXFSibpdW4xif4Kf9c9gHc54e7gVVNlbx3Rh9JieTLclUqYBbfKOuNJquC6EV2WICvYv6UV8u
uqGRWS55zhnxFlG1fKG9dXiVdL4aW2L2LvKDjDfs+/G6iPKDkKoDqy6yVOx/CWK4QEu/c37ZkpbQ
m+V1FCvFwYCxV9sZCToTGDGDeO0SrTnmSY2nfRgmvWWQQNvHLnPTu4j039F3G1UjvT+3VESIyVsB
KRU0KK70mRY4RvryKWaXV4SIvgmfrhHiNyi31sCI16oeDfhj847atU7C++cUQrnFD/KmuRsCHu85
oETDxFD+IPS2cSDDEuVcRb6hWYpPk9KZb02RosYFGrRAH5wz0byVWTMVYATp9DRR5USQ4+MITOka
vjszb1cn3TkOMR/KYL1cZvINWAafDRxcDCK3jkkCIH5CAVCcNS9RqSmtp5/RhrB0sDNX9WWaZNYI
Xn8WCE85sFwZBeTJ6aMAmW9xu2RBt7eUmrp2fYhmdiUw64xp44N4Bl/HWmNRn6XVyuZ5jvBcawWT
ThPr/ZJn8fEFN9tOHot+IASyxxi/ylHxtQg7kXwR6OFT1825x/WzO+Gj52s65vwjW9J2bgmMPvbQ
5uYUFVXM4gVu3OvyQXWPVKO5YDwaoG/L/JsrymH2Al6mO7Q9OM87Of/D0qPlXkMLkzJqR+vM0JXK
a8+JaE4EueaTphzpLVencqU04gikmnZA0mTallfKdof/0XyY8LZVwIADj8vuN23pf499dETs5HoZ
eCt7OHzko8fYQ94Kh8fHsRT+lsWP3zv91UF69Puz4QfkBGKK0b2sQ+bMakuIxKThst5GJbvuqn4C
/WTKiSKc93pBoT9G8ifboXCQvJRDbTciLLYIXh/1gPme6B47nrOFtKizSEFYBnK+M0WfeeAQucZ0
kQ8shYnXMZ6EdUAXgAKA33V40DHJFkULXwBbRbRMz3D6YmLUjaXOE5W94uWPsIcy+ADlNMYMTgqO
b95UAw5I821GdDNNvJ5s8GqhhEdnZCGF2P0neMMellg3PsTkuoP3F6gXHjuaYX7R9XJj0Bw97K74
x8mL9YpaTbQh1qUOMx0J9QJ3NJl5+ca3HlHsIhNjlUCdc5hSwqE3wsJydC+wD17XPWwJ3NZGu8bV
m2ncGuzShhY/VW0hdQGDV7TIYJwHIWl1dDSp1sBuicf74+jwPQLH6TOrBpCrb/zxPFfltfzwlebM
R3fP7hq/u8gmE5pOD1Ynkd1A+CuTT6MoBfydYg56ADZ0dTQkY5UdKxR5J7ZVMrhBdUB3VzU8D+VY
LDyohHy/4HYVLZWHnhm5kYkr7ceVZeFSTeiW8sHqtuLNmOxfP1GDdKglW4xTJU/rYNrvqnrYnW41
/oBcfwFbzlioMvg3Gx9DjSENcLjWaUGHEZAA5y+/LXy4rON19hs5YAHCE1/+BPRdfz82UjPPh8dC
pVciDBTx0oROLlTTQm9fU63Fxh7c4qHLFBNVh/cOwhtd7W+kZd1cCgPLs5IV+qr/UjFig/f71ip2
9loTkAKmEMU12mzpRWn1FcvTSBmym4+N0mFZskeD+WUfjzM+pEpVD89ZrZz/ODXgOCvAbbc3xM6y
D/rjzTvgM0XX5mCRUz8P9TS+yMfjP9vXdDdksm/6vjurnTzjfmu9kieTij+bqYCiukIdL4Pgqn8D
z8QigYCv/9B5JUBFivO4ucVXPWwgAO3AaaVk3ylC9SHzzVqKsxWsuPNbRgZu6wuM/npSzQ9jIUsJ
8yOeBEPrTUypdyzRaldhHVSPbNt0Pk6uszFQNQ7xE/QKvb7wLtABk8VQTiNHCPYcKG0AVNSEOtcL
nNX98ugoD4wiI8+nOADhq44IS0EMr1jD6yNh9ZKDcVPh+VOTpeIzH4BGvGoctQwQ2dVDr7W2hFIS
51DthS0L6rBsvQy8xRSJqvOp1owsmqny8/uKAPF2ctUXzqUG0AAk2fbdt1g/0QziAajreByPOe5r
DgfW6hjiAk2hd5EQc6CIfyP+gkUHHV18amP3Q8wpMw3TCgWHtl9vxeyvdtR/bcRh0xaJTAWfDWbI
FxPhOxQkS8DXwrTV4gPGe9XcmcZuB5JvymB0iaml2vyLfDzHZDBe0tgmZaM+clbgZcCTj1IP43VA
wmTqQPfA4INVB1pCISXnNNZA98EpkCR12qC5ZHvTU5aiNAMxVe15YnFab4evfk/up67jTgB9Kf6O
Qz6fqiawe2zG952XlTYRAji24QFNxyxGQaLg8+mOw6eWxFFeclUxNAbk+YiFY1ykohRE8Qrapwae
rBgHL2O6snFzR2d2RS7ojvDrXImPvaETCkQxTP4L2MDn5bjV2iaILtlHsRrnyi7pNOW0Z/EbgBCC
87hkI1FnhmrdEtAbZLqD3ATowva9L2PFb4+UZJ6rJCDfA0/p3Dvrv1Nv8bPGawqXr8t/lZjRF1lo
g92asy3Xjo5PDpi15gZOQqD89DGMzNGPhaBP2EFdZs8cTWwfMlcyRARgQ/Vr4/au3q5bzdtckdJ/
DWs26hf58Kgl8udYD8BDNLFi6Fp5p5Tmf/2DROoqlKSvxS0ewl4EROfeggW18c5/B7yQx2E0MW1A
bo6RQxbNl/GpJ3M+dFjbMOGma7ws31BXKXtconuNn3eCgM4Su8MNB7MB4FikBCW8jt9usxrxDzSg
/ruYzvtNukAMpsZdigXmA5et2D1etUlZPyOEBVcqJ5oJjflx/EGy4phrd3fDXlgnDJtG7TM4+rZK
3HJwU+HPflCOg2r4n/7aX7vQ2WZOkg4UbNdD/gR7nLuyEtqLUf2bobdx3Zsbyr05ibhWulzIBZgo
laGCabrvJXoyibLXgl3J76ClQwJjnnMVQ1/KA9LRYp30i2B8SJuvp7IUtrMzzqrwSC1TqVynr0LY
IthByQ8Pkl5GgbGBueSNureaOBiuvL4gwQZi9vNpruYMuois+hwCHFdLCarnAx+VRlt6S31kECVv
k3LMzWIOHlV9jybfPy8SqsqrEcacpqa9jKeK9vpKbhl5SMga8ftRmwSUDZpqM88nZGW595KcaodV
gYwAyyahcMQswuRbuPQzcndhJYc24NPLCPRRoUO4p1NU04vwNzQezDRpJn4j+97aIELb7RnB/qtq
23/vH/RQJQH1Co995zPuVl/hSgxZSgIsjDt/PVk2LJVSAUVSCSGpXqQ68mrx5IjxDR6hYoySFXuj
sTTozMAXsZuy7BxUW+Uz9Bjwpfjm7qPffSpPfLuZsLY7Y/4elMD3ho6SqmNACFbjeTs6Zetnd5sM
qCTtJBxFHb/Fcr64xyXfBevu2sGEJ2ABNR3Xx+HSf9Pvj1s9DOYqkmWDlhtRfDCLRFqUJoOO1NFX
RjUlD3IKVfekdSUS1V5j+oQW896CFLsTKomvg29a9Pfs1T1V7/2/sr7EJKCItqyWqZzTFRTd+6dy
xQV1rLIdt5rqosdSZAfRrFYEO5c5sOV5Fee2ls14ViurpN8uBIS+O9bF6lTkm/yC0sk73oCBlxLK
ztmjhJZNB0GJ9hbHCR62etkVQMmtCECwZQ8qoYZc5AeSEYxQnGK167LCvQYaLNBLnaaBKtFiuK8c
ID++5XUCn00dt24CgSPKUMly0F15YVU51dFp2BW5D9noc+hAqxRbEl0ALY4R3gBg/tfr+SQVZvBt
hymzSg3JjL/+vDCAReFVLD8jFt01iqhHfWpY3tp6QEVv8K83gEYafAl9YGKTb25Et6pqgeHwrdo4
crYistxH37b1BQ/mI7ioLMGxliV3dHw0YUSfccO8ZK0BuLP6eQo1qzRWOljmFMNaxC48fQPzSF2Y
+YLCnTKbKBbyg4BuYFSijrWt8pY4AUez1LOFckgoXNxxak+IczG99tK/ntWWuBcnwCpsSTb2J0nr
0UglzOItdTycF8sRarIVOl5YdrUdnI48ITfljPP10Z6MHSu0N/E/CI7252y/M2/lkkc9M84YEG9w
P+uY12onaUi4MBJ5W7w5E/Km9zK4CLALz1kVXPObc7qdBTNsyPjubiKaL13oDjBdWmdzLKBpPzqz
pUvrUeFCrnSSEXR8XHbq1HZiUIGSCdfvxUUPk6CEocc4HiGfStM3YRw460KDK/oKJYKVo+zfUy+z
mdZchxdLRiyKcRFORUEHrh+V/lQKw1XAZu+UrHIHbbUp2QkWHLWM9x/YIyg1wGIS3RU4+2kw2BUy
W3uZf3VY/qdEZqT8/bNo2ZP+QCW1POWpfZ3bf09gD0jjgpZB3kA4/pZbAkg04UeuhnG0jogFocEJ
vvQ2LWc392qUVBcnrrKfJWqvthUNoJp8ftuPggK1ZJ8HN7h+Q9azV9sycIZQSbT8WeuUQm2konCy
3ykVzC46x+rMNEq+486ks+/6CpNt4ANzFuNEGp9fnerlIrdbhfcQkYjHL2TyTVplgGuDRTUF4TnM
CBWlS1dWHoSRd00hofyyAXU6rRG1jQNb+kpo165RBEnpzmHJNn9ghTjYWg+2d3RnnoBjqEjlMJyN
5+qhTj/n1UrD22+mCpMQ+Af6YRDUbyfyKgeqnA5zmRZkZL/TwNEAfCk+Pje4xNaFr/MAO8Hf1t4b
6ER4piz4aCb+IJCrlv8DLDqMjJFdsr3gIQN8YPImxbp4Wwkdf/YcxYZBEoVA5p3Xk0eaNwzCSMd7
4t0iR+H6MEowMr1sQEcpKxJAC8cSMu9yYOoFp0Q1OAnEYwXhKvMLlW8gs4B+RFyRgwsHSHgQnK0R
Eov+S3BorxEK8oxTXpVk8EJ03GoJ5ecAIeb6s6h+5dEwi+381hr6mDX+3qaRjZr8OZKmMBNRgGRc
eOILQd2J4hU7gkRSTsR7waS6TUifRxphuhxKOP0V1j3+PjfyzFAe8DF9zksTL8BTpd1i2mqJPQyX
vrNtRk9qVwnyp7d+IsHVOG9VSZBQWke+JAV7xOJkG2EuA5F1XoY08z1TnKyuvncN0fFa6dHoQKJw
tphwS6ApeH+XtljqMGzCW3N5uB7pbXri+1qFs1TwjllFwmwLBXeEbfv8MfT7Xd7MV8LxVuPgEuGD
nK/NMINijMv1WkLBU3psgPThXVnwQgAlfY831fArgiqfUcGJ+amse1eObI+C+sWAhl9kfpXAs0EJ
g7nd9B9CPtT09tZ9ojUEey3ELgaBZ3MbvOmGPWk+NY1i5HZDF4RlGsMljnlW7i6u6o87IZ9EoXLN
y6m5a7OvE0H3FnjvCCrfaTd3ZjfoU4F40MVs8XPCeMQUFwsCuvHzZp9U0H4IaQQROAjiM6fi15+e
CQ+eGdr/HGW0LVNv+oQwRDl55uy5vTTiEp+Sdwbpn4uCbWirKlv/p6jb1SrQrGT98O36ezPtuBos
R6bozL+TL3UjfVYNFaHG6Zq2zvdIjF3h+ZvCycgrc/xJ2VNqiFbT7u0hZY+kN6OKAJ0DPveGjcYF
7lMk/8kTEoChN8CeiU1f8PWelH9WQYHzz6TF3mjtq9CndI/bVzA77TcWGnojYifffLKYAuVzPv/j
wknFojFrXdRbaAyRJ3tLvgdOZu9bDVUmvBPLKdiiACwHjVMO2h5oN7RvELhqWmRkMM+YsTMbVFSN
vSdyGLCJ9jd75VMvsK/R1RN11fnRlhFbbzrKTgxbucdS6uyOID8+amyCUNodbxTm6GDd3v+NY980
yasSDbp++9i/h1VbuE2Syj0iAU3i/Kgf9ia9gxIV4xfwlL2HeZmbG0B9G1/a7lS6g3bPdpO4rPRp
OISnrc3jf//4rF0vea3XAZ0NU8JorAihFefZzc8r1z/uXtLFaS5voLFuvzFTsDzFa3JgHpEiHHTa
syiGGt/m7Qx/Lrg02j1bD1baaKnAreydjMtluQP9rUIZupkMmAtJCv+nenAVVyf0j25DCFL1nceq
lC8Jy3HFShrIKan7l9pYEsmkhk5f+6tPv6glzCqfK/3xB/d3XwUk7h7bi/rsq+rFhbS+6iGpV+or
jljI0NY7zlE1SbggbJ7d7remgbZOW1Zb6zfcjCCJLAgpHJPq3HPYPFklubfbAdnQ/16RRncLF/3N
2bdPdDe1hYdrXxyOgcRs3FWS5/bwlAEAOGhJ3Fkb4a8x/DA8MdgcEeyDARfTYIhRDHVUxUj0kBCa
PnKvh8ZP0Qo7/wh01FK2+vGdwr5GMp9xKa5zvcbXznJM1JwtsCEDMQvGwpeQg7rfGkVemnIkw1OL
RCKsx3d5Y+ePJqHeYtfUn6XD+n3pscan69sZm2ubn35MJnKdteMLm+7/GCMizrFh+zx+sZqm0IlO
ZiAURdNOwKrzVSsJPUKXm2mJLQ+v38ZPPwWxlCgsFs56cOaOvXuMYdwSL1dyPQj0jI7KiQxHKajx
jPfAScGzAzZpNC0LS2gLIxKfRKsnaf0YFKMfMqBzDDtnCnwfqC+xmrqPZpjo1zo751wcB0+JVApG
7w6HFog499gWmWdx7MZVgm6mzknn2IFMZvCS1bt/Z8aX+XHRCKYNnKzOIthvLL2kZl7AgI8dgAgi
e6N0dZPR+3cU2xtQSUlnbx1mm2AI8WYxBHAiudrZbI1PIPoCGiJLfOZQz4B/VH8Mafx43cSUreDW
ps6dzXMXeY74DBGR1i0JqOHTD8yW7tAuKHc7jDs/4vKRzemagfOxwy+l7IDfVNxUF9/B50B13kwT
UU82hJOFPZwL3ptpKDvUdmCBwHwwLnfN9TmIvATPo44fsS7DRUti3P7hTUXleTdOFEitA5ZjU/JI
txaKFBaw0WodArZfCM8lPexDGgm+TD2IDLygSSI3yhoTDTw/iqIOhddJBL9wGZP/kGwm8NLAGFmf
jgREi95V53fhZirVWW28Yu9Uk1Ix9T9+pd9zlAbUnmgJ0szA05Vxfszq4hwQBXqQ4Kzn2Tjl8hOB
Df2Ot2bx0HKnkqYYGZZMCE8GftgA4weZJpe/2lNrz5GPKxnAC9w2obGJhEn1hyp5sqIG0FsZReN0
Lxk37guzNK6R6kf5U1bm96tcvgwkHJNMO7HTSFyWwDltdv4wkMBeXggDmFmdjK4IgTYkLd34Bfuf
SX98A6ZQFXRo7CCtboRQtrDgpUP8/glyrQsygYaWQmAiia4B5pXACtQ/Tm0J1VvKCmhA52Cr+cpl
lux77nkKfw2A7zKwSR5Os57QpQOiZmJ8Pa8qxBqm6RrRgqDlj3EQN84u+IZZYXNCRKtdmgs6tEPK
hKOjmSxBdWR+PGaIw3IBKsMKkwKgG8JJLq3uyxTTF2cYbrM7aj43MNWNCQ/wPQyCnrq/Mm2en0BZ
ccZMAZBeAbakdZWUb/or72bXAHpNV1bjSS+TiQ6wug2EqD4vB6qs2Eocprjfi9YJpIJJgaInh6pr
LMQZi6uLnv1jN1pxYPnLvI8i4gIp72Tk36wkfErbyy+JlQD/mUqfQbW8Fr9YYmsUpn7z7Yft65uu
xoeFkYsQ5ddfe/L98E+7bXTMtT/cwZiNt2MzC+YXvqsBVjm92ZFRvEd9i75lKEeInRju+lxFhqxm
i6Q7FcipfELQXTDcLJlgF+tM3XEGbxOsIgkmM+qMa16R2U0jcHN6F9egHVCCqi+KEJ8uRjBcAqj5
sQXJn5qu2E+VT+qp8xOwsr2rRE3iN9fWWV02m9JECP3enzvRYXshvuNWYHRdIXjDszUL4a5JfBVM
r/l0ItW/IdnqXMBW+wkq71hMeYq+vza98sVtSOkVlLgEfZkTzMwrQRoFszeJPI7dgnYhcXZ+Bh7P
KIKtAt1K1NqtPYN3tRzpKMEoIi+Y4Yt6smR9S6f7v+KzvQSHk/u5HyhhGa+Bsxny185xV7x9ScSs
oT1+BvfvZDjYK/dkWeCAhZdH0dmcJvr5SUq79gpbPOht5oV0oqqShb39PLzXMuDaqIhGqHQX5hmJ
wBYt+0F0m13bozz91Iga0fHpyg5KqvCJnBhT5ESsNWyrEufOOnTNYnTn4Hb0Igsh1dYhny0XmKy2
+h23Uan4c8Dnab8oe2XWsOAM+jSbNbDQf/oNxAsZyGpbrBDHyVXLk0S4gZjrrlMoEi4wbWK500LQ
4CtTSL8i7ZqXPPtaOc/bfWSnoXAL9tmv7MfPNPUk0hBwWoMM5kDUf8pUmgnkePvgpksOAtSU+9Td
qi+QHNurQPTVZCE66pD1hnvnSt99MI+/bEykYnBLwjtBPEEs//AsHXX2Ppe218wE9KT3IJeMZuj6
3ZK9opTOVud03dULLLHhLvHyLC5kHNgHlyLUTxFjwMZce/eRfGxcWoKwzHQsop5EAWg7MC1DWse6
pyqjyrHJfkDArKRmdI7se5OUBd78S01ZPowMGaJ/Zd8TUGJ4DpPhbMWa9DfaOyHsJBGjS1S9Htee
9bGk0pbDYWqXIk3VRfjBDgoD9LdMdgArLhRhx9lT7BihH8D1j23vFiOzAxqBRMLht1cV8vXd0ieo
YiLvaphuVCAGqAlzntrSZNgjh/F/1nkWUw+dFg81WqAsl9Z/ZReL9TQqoBNvGf2Jllqn8pLdEZPZ
NLr6mxmeqd8ZyQODcCQZRRPlPodadsGbRX82o0Wk7TBuSHgYhtEQT79zSlHZKNhBRJhKPNdHYfHD
U3Ede7UZBXXCUvdkBuB6Xb9b/kLxcRcw36CMUu+PsxNfzvNieEOYut4B2tWrXoCMSHEYCKng1lHo
e/oXf/YCOqptHfDwu1RZ00jv/g254wO71lsnK/T0y6TWPND0p5F0jkkhFxzSz5eigCmLURf/ro6d
vjsmR+liiZZZGgJfqD131RpVDgEgmcsJJBEV9yIqe4wn98Uhd9Hgwib8rBwC/EN+0n7wyjOfGg5j
mqh1ba1s00BUA/cVWc1eqQODXl2iQCW76seh5ymS0Vp62NqI+2jPsvkOtY85I6LQd3FVlQkRBvLu
5cP54C+8u9emaUdtMoTcl2EdzH3P8CrG3YarhH3BChX7ZqrRuMPD6eDrgBnDlr+qc5dDbiTF9/Xi
SB2y78k9qmq62hFHzS0yKoZnc9MkW8fTyRILgXgbvI1M49UC9hjTOUlSXlXom96jkAl8GqC3ZEnc
9rgRHXHRhnamGb+bhzr1DfXsmLGYHMO8+sxtMa5tejILO3+A1jToEbJ8c9pxKlzf5xeXFnepd+uu
psObVI4h80jTqT9sCfalAM/UhAaR5Jf/D/ZFP17sJ+SehPK+8JMtGL+D7I3dbH2aPA1i2GgzFb6I
oxcTMfmGfkluu2VFbpM1IA4BJ2syLlQ8FP12NiraHoLhfX3XcVUqc1W3PfJNdmLXM1jw/4TCqE69
ak8/lv2xvdD70EhiNIFoAKHKZRzlPyyP5/J0eiYBDrMNb42zUlKIkOebJ9j+vVIfvxyrCXQM9Er8
s2+bUq4kASExKGTOP761Mf+FtOSAW7WtKqwADtFfqn7rMvAY5E/sisG/hRhS8YZGDg7qi2S/NRal
WTx+puLPiXNevCUY3il3pFby0fmuspE0pMWgGIbQYh3U0hTMD5TVZ/RdkuRCo3VBvnwavBVb51ot
n+s7Y9ZYbs+bb7FuYNaJbirsN9OQ9qFpsXk3yYA+qIv/SdusgD0Zz0RqZ1Qu+u3z0eC1U5MwZcCa
0zx/vixxDPClN6jraB8NRSqGexrslz3ZCr3e5sr1Daopod6s02xKsbuAtX2Lb3joTpqAv4icTnEF
nPSUE/k45If9AO51mRZKE4zaB+WV3tOdIaWVHWMlTshAiunx+m3Q4x73cMweIHdD3mKSDe8G7b/Z
cUDOx0vqqjOu6ye1dKQ4syC9ecwT7usx2RrsyH+NC5gas5dwq4bT7fOX+cMyGPf+DUv2Nhy50Wly
HzkCJuLiwWzDHqCUsQ+p8AWjmZF05cZZ2R1XlVnx/W1eUA8T8Urw3RmZ43bgKnamXuArUAqLBFva
gCipL4FN5tVS0r01RvhkUP6thXlMVNBkgJghnptbFkIdFQMg+zDjkbSn0I93il1l4v2vrsZMUw4Z
XHo79/017SEwkyrQrj8F5jVrUa20Ot7ID964Uh7eK2TXdhxbjvZ9lr132p78p7qS3z94n842U6Ov
2UU07vcx0ZQdQ3HnntyIKAkDPEz66tYccJ73W9JeZv5UYwNpk25Et+c2gNZT3pI7uKp0wmay6uoi
WmaCYJJMSWpsJWxSVjp7dAHu/7wZyCHFR2tvNOKgGUUoNe5x5RxefiJ7aVlc4LY442PewGYeJ409
xI9qC6PE5oXnCfrVSYavSEdWkoiKusisruRCpTWSp07AMbe+iY/Ur02+gBBk0fwF9FzhivlHPjij
ViwOi2md7oSSxA9rg9KN0W+Qzx3QfqykqnBzdofxGtFNShW6VONR03ctsnsn9QYoBph46EYVHKpI
NQUBy5F0L23X4qCFaoJpqHkoudc3mZmeTEYHUTqNqpXOFjHY9W43G1wwlYLIAgMtPNiVK3nyZHQ/
+YbqM7z+2w83CXusSjkVj8FxU6GaJHnrOHjzXKLjhwaF4yZDJUGx1njCJeF+GHxNP99HXqzB+Fsc
qLvN5ui5FwLnz+bTnWC4W9Nj3iSKUkAdRM/9prc/dgrqmRkeRJyRHL7HQO9EV6v+hKnAU35M5CxS
c9w/QSY/z+0AKfPiyHZESkQK0dCpe650dkdal8a5GB4e+NYTOH4MZ2smcX/EwxeC7/K/A+InuaeC
gWPHmjRg2Kz43dwWeEq4ymFjwmJy/O7N4TrIy2hGOglY3RQoIqaChhETnvxpDdvQ6BsfDFkG7ifw
ggfMxWmNalVmqcqyWZ2omVKQvwuR7OGKOU3yZhC4+ngPr8qwjpDOBJKXeXJRaX21qfbsI3LqzBTp
5PGfCsJwEg7r4V0e/wI+TBY+JBcyVPPQWlyywwYE668JpSpeUBsOgK94RkCUtPmIGK+oJiaIA5dz
5M5HOpn11R/UprHHGgrMh4pXAfpUm2ybbTGgpjMW+chHFM3ZCijvAuGfC9DiU4+0bqVlvD+CIwYG
PppG548/keuLh+fHXwKoUWs7pn+uG6q5UN018rOTceyUllH61lGxnI8tVSIk5TvfxJchjqxkG4/U
1lZe6GOx88xdgJp2S97N0LF4+DGhKkuALKcknmYqGNXUa+LVoBVdu9sPL3VvP0oIgGA0bucbj+fc
Koo4hxY5zHBgWPgwdrJcixLZrBedDrRvW7UgllFZciaG21UFbZ7WFZ3joCbV8vNCpdYSNpVQgwk+
vvt3aSRJPDjiXvTBKKdOogEzmCo7NF0eH+WKQ1yB3t7hrpXeg3HBOSOBKvMLO90+XnQjBvbj+v+M
Fx6FQzDnDeE+bcV3hl2I3Jqpt5zWeXuvs6aCKuNa2HqLhn2YAfhkK1jq093pCTSGfnhIpqyPOeRv
9avkINCoNqiit9/N/wLDHuBgGSoYNhzrKGjt5FjsjKaVC/87ZCpfTwNpdUBWfBSE8IN4lTp2CsTp
ftr2Z1UTGFkr7RETU36Pg3z025+oOzasE9VB8f1Ht+r+tbCul2dBLDujX0296PE1VfwXzcjNUkQF
M7lCQW1AlzZCTPw9vYIRFzzW/VvAzGOwnPZT7eBxlprnF3Pz9Y4rW4dTtHGWzjkXbK7KlmlEr9hA
qpYWj43XCJ3q6ekrUj189y4PcD6QN/d8XOYjYnNZBG81zkSd7y57Qxe6Y660eOtDDL0RcZIsQNCY
EAjbKeBi5eIH8yzQL8GRATeJyzyUiYMPHAI91U2B74SNF2I30NfgyFhCcWmLFppQhTACNk39W5Tu
pWLIGCFxBkz26OiQLmUBn2H+JcWocsW8nBDE45uq9MW9gGcfHbxV5vk8lIaXRM2xGbEFvcdABE9f
8N2jLOKP6rxSsUiTN4hyj5YME5Zr+AfyQHAeW84yAav/ki8lkeBh4ZhmTV6AicfvgNm6///5Am8M
LJpdKyGzk+7s+HK0qye/WYReUW7HsZWeU4Wl1RtKVT98xMC1UvQz7HuUAgzMaJVrJoPCRfLMAvPq
xTkybHm+gmVC9Ki03j2p9qDtAsReIF8/WBMrcmKtbMyTFCDb+zg90/6QxAIyIDLbD/fx1MVJGDHC
9//YAWYuz+eyMNGXLpgZRM43u0qtSI5zFSZNI92MYOpt0iThtB/DwmOiYblKnqoOnE4pnWA0xaAX
cm0FaMYhCc+YWOUMWCoTTp04b6s8HXvPvznaoAj/SLaK+g7mERDOAFqCsm2nnN1cDMeVyg00Tdsv
9tFVVHk8DFKSh7V82Ut9FQOvxUvw5XO9G55eCOBCTu1h2o9GLZBxCDRywNK4Pb4zzKLM4mgK3o82
/x3Rwj5wLxyK2565J0ogKnjba4c6nP39xSNFiCx07DAN9vzFUXUWejYUZYZFcrNmVewcmqZEplDN
v/zuWgs4G/K/UlAqJwSyA3Ez2R8U3SioVldTeLZwLQbAnMed9AEFLkceBXwPMd3pSSLCLpOW3FDd
g6hlUzXWK4p4+CVrUpdsATXEQIP2+l6FzDhXryj53Gl25zJfRehXUZzGxBoHb5OhcfsK4JmiesHM
Umx1bg3EigThHC2F0a1VwMUNTW28lN7KCjI3fmQRRsjDxt7sOPZlgCQ1WOU6FiEhzt2DARanYsn3
wptPPTtXNJqCJmAKfsYSnhCT+3oaOZMQLI65yycEHBqqC1GQzBb+8p9MabswZHfQ+9SxAUmQe76D
LUL0bYZVgE8HgsyMQQfrdF4o/H2RRULTz/ivZsU9CjvqI1vjvZQ3N+JdyO3Vjxnacp18I0E6ZC/f
GFgzg5z4jlLUOWR2TixoRBYbTl/FOG8IOFwfVowcH+XqB2muFvM5uGr9qF7PBsZriWjX5QHiE90R
qTU3Q5hTKMfJxtrY8ly6SfZOo7rItwEF/vwjVH8pvZvND8MDPNVnl0L/y88/erFlrQkWWEKpgJ9p
mHnwT3EQtbXum2WuQ12EpqWh4r0EXa1udhlTNskycpbOT3CyFiSu0ChOLNg3egwCli3mHM47MStr
6mLOBqTYpuYCxic5nvNe/IN77vKN8aq2EwIpIt0m3+xW/yoLDtutEsEQ+U2okTiTzN+xrJHMqFIN
lMhzOPEvFKzgPpG8jSBlvBbzJDWbqCUyw+TbYZ0M+dEcLZkF8QOSeVXiGGEpAP7zz3d71fLFMA9q
lADixekf6d2EZjcxqPez6HtM3AI/sRBwwyKAl27RAxzzgEDbNhRtlIkN0GqSmR6UOd2cDHwqmRf5
n62BRZuX3QCQomit7UqPCT+WEc7onKzCsHw07Zjxw7BoJuJAOdkoDZdA8Al0a8fBrYxUZAIy8+1S
SBzn141DZqII1FqFAmvoMKbzpts6yosOVvDVM5FrooQMjwjMfZ6tvvkPd2CZ2/vvre8n/6haOklG
Hc8FsyCr4VoRzO/6sJN12E/qKaaXKgKwfKZ+KSXumhQJVJZnVudF4d0V8vf3F0Wn+x6zt42HWNE8
1N2b0/B5rxQQoF8GfrXG4K+ND6uEZPIAIZ5umz72vlcZXkPMWURadNwMY7W0C2ymg09oUhg70gYl
hw1QE6mHlEtGTKZ1XbqW/kBiuYVd0VQJ3vj4KL2rJnJUgOvjofUD24FQiXUV6DVuPqcjQvgH07So
/S/KZ2PRYNicgChGQCXVW4KZFX4rU3cOrgpyx8D5gXw4mjtIdWSAkKfDx6MGM5isFzI1320GlO9I
xQkNJBHsDSJbj7YzJqPB7e49BwqPArzYaZ08vVSpzAhoDR/FYE9hE86TMr0F9JV/nLUsboodv98x
OWkU6ebNtkgAyqwLA+J1bBtI0TogcXFB4plRj6gd+q740KUyBFERjoJA4L/UtIga9VbefDzhbRJN
UT2Q3ZjdM6EO0vdyDRcJTZ/976er/rY2iAeJhgnOyOJeioVpqBekrid51jo7ALo9ovOBJua9hwcP
ivIsFElZ5tA4frGjV1EnovJIdZIZFcJ8Z/TvxY+LBxnmtN1c8FQqMLIHXsCDb6KNCHvnsrTVhq8X
YDYAupl7oFnxE2ccayL5RYHKlt69ftEfRN1UTL+eFNJJtfmd8ByDMJgFAHuoqYlIGt1bW9k1xglZ
JN5uLg9YSJ25bRlXuRInN3xEHaRt6bmLUmz/AdiV53rCKBK4HeKmSgiw777edg4Z5eECq10Vt36o
etvELVctnhUBuN87zR5AgAV2lO7R52084RiSr7SMZgZ8kI+kBEMKFS5HDk8zWsmuZcFY61XDw0np
xczLu+6t31ZHvG+l7x1TBJTaEq0HhHHkKqkDPiNcshVQaPtRMhymyCLo8f7DB8tWDwDBp7rrxt4+
dFgm8FimM/2U56J2aBUw7RsYsniILn4JK8qxZzlWIRKQzppuFi8BlYl1VhhAZq7+Kc6y8oDBvEBV
T66IjVzdGoT2xcnF1zL/B4wMSkvmriPYEZDcZ07IWKdB04olb2mLxTZ17mwCzd+1NhHS4sx69l/9
4AaN8pnjd4y3b6JKuSu0JLfe1c015NMQZx3JvnUFI1Clvsnsfk0M60CBfld+GHxwl3QVBwf8beI3
0TAmvlkX+ZGBK4Tw/iCVdz8DOiVFI5GN+sBiqbSUs3T0iME/s3pogE0ui0BmbVkmHD3lNy6azHZa
B+t2cAc5p4/dA7uSmMYdP1tUHenIImPZKPJ4Nsmv1a8xSxsmVYcw6FO1Sbup0NSIRdrCRLGPRgOX
EGYbEoHtP9lGSt+ALE6YkwEEExQ6mvx9nlbbymEUjIEUBQ+ySlqfYY5LFlYzxOtPm/fUO3/Y1q9V
aTj/s+/lBBdPdqYBdUCqliMBA4YGIjJXE99GlHWNVyhGumU+zQg/eCfRbugvvlyQrR8ruC4BywhU
l6cX6koB0EcX5GUGQwGSdbIRuy4z2K5ugpmxSl3Yz61MUxv5cp6MLx9H6YY0DY9r4kfLPWvb7vqm
q0Z8TvP/OekJM2pGjk+QchHEuDi/omN7X4tJH4Ua25vvziK1y+SrGnpRfWpdSAn/4bpB3SaV/8p5
18+5redoMBBpxi8nmMl3WyPuv9DFXx77cRj6xs3ktS1DKt0q3W8F4FkOUXAzrXTOYsoRINO197ih
uZnUvTKskpVOYtJZ0yoR6oP7c+BwdQwqVHczkvHZCsobEAuWkLUhbYsomr+/ekuKDHbfcU6/2pp0
61IPY7geun4f0L8cJij/uOo71JCLpTj+WNHk0F8apqKsoKv62JDQBwTT5Nf/uNrnt+fY5t8vj4KH
tjYIm2yzatrgtY8uGIP3S0p1oXAgnKi/c89fmzo1CI+SStEIm1Da3/7uEHFnDbPaxl5Lp9vDm8sy
o3wPgOhdHauhRoNKlvFMxF0+5/Z1Laz9jvhm+23jsdBDy/F4x/F/VeYHIUOk9iRpZaXz0A0ZUpZN
XOQfiFd/UsvnhAAC27QQf0gnJFzII31P6vZEfTm1tvH+UuCoqwLX99v+NuqexrtMlsffeuCkpXM4
bDKsVnsDOVNPBiQfokRN/AaPUzSbe8vLYw/WMHUUt3Tb8omEzgAMKJCQniTWngHvX9vcLmb+XSOT
h+4/2jRo0yTpssCy03ZoIozUW0nUkkg7lFs4nhUxeIDSctc9ft4v1i9lfeZsGnKlRv9vOju+Za8x
UxkbMV/Ohf5Ym+TrzUWNYj0qN12i44x9CZfaLY/FRa1m2e/nRYrQmXwufVyrVP0qPSAhL+SnS+TG
3CUtD5i5PRFZVoSDbpXuX54bxWF5NYL/rZZAtJguXYFJjcgBlBY7JXOGvhB8WTqF99EAro4uu686
4+gYy/oXNQRgYgwyyLUNaiWMDhOq7mxA4Ymo1roWM5NeEEKR81g7MO+e0ulPR83pqA8+RAY4uE7L
RbGjpDnARaTZYPqA5vBIDFhLChqIayuTlSk5sfDAt0a6FykMvHgfNHr1i8DowHeEcsPQmoXtb7BK
N/obgWwaPp9OvrjL5twir3wfKCqo+JnNi1KWz1uLK2eycXYtjcOFlA05vZJzMHL8QwatQBzKmEbi
NdXrHeJa381AUy/Zy2RC1/eDfcw3BUw/UTXj+CGf1PJTfjKJeR7ne5deI9lTvOiKl4C4tDwA12o7
BuZR2dt/aD7TrJy1JUkUsmrWk4mTKDzuffhQLUcU3wH3GeRtELt1csa5rIXkHd0JNKiX2moQ8oN/
UEE12BRtgSMsliBEsmhH1NfQ2+i0SUYQCFahWnQi01vDWFomSC/fbyQM+UhK1L9qoaP482UeviFO
TyfLhCZxGFeplQ5HPQbrHjhuq4Mi9jpJ8Cm2HRdXvTYMYo1XvWmtdv5KChseUv2JPqPWrWCjTlZH
0KvKJJx2LGMixSCJbWFR3NNQdUv//TfE4lquGmjmjmMOG+CnAQW7GEbdQjnwCvw89zyU2RewN+IY
0+MVIb8hOF146uVSTlEo04CJuTk0bDxyKyRwQ2G3op2tjZfQ6PtQRAoaNYknsvcSsrnN615EQhsD
gBWo8hfLSxTQ6wLpJge7O/8GbIBfYyODQIfh2n8MIdBPAMJ8bOckKRnS+x3ZLPFpJXgpzzL7hmMA
pMQoYz/hzjoCc+vciY92DTBznaHtxLfkJoymBW1IafZPjiJQQXIfop0Qs22YD9f/qR6NQ3U9Iikg
5eNr2W+GySb0VkMoV2VDgw/LrocA4cR2wXgQ5Big0kNdbcGkD7ETtXijJdYcbDclXM2Om7BJ3Mal
u9ZjAIXwZAIVaVZQWAvIzmMbCU6iijM2fIRSh0trQeLb91dIZYIcYEWbBfjWWjPO3EqgtNTfvgl7
VADzD+jpjl38VWenUZ3gN/OlGgvXcp1oTK/ZUoBx4bzj/mmpeh64oGVTmALp1Iu7SB7gsEgBMxzg
uZdieRRuntCXL/YqcvBgA51ZER3QW5fyCHzdzomqjng2c4sbvhrl0qWdkntEP8kTvG7bbDZy4jJQ
NjkCqoJmSb1B19UEBTQm9LBWjRYKjEDCYMVZnqyLE/is5OXMCxXoTv775SWt0dmFx/SeEjakCsxR
NsqPkl388r82yO9wbM/WC+Afztjz4TEDEXSJwfMr6P11efSCxqGYcO2vdHASDrUqR0kXMuv3uxFQ
g0Hq8wSA37gez971n+z2IH6PBaaIu3Lf8GUHUwuP8NA7EncT70RC2f3jHtQaB68orlbRDdPg5PRp
J7Y3FSMKydcQc+JSGjDAPhH7WNL/ZzGO3qXojHKalfU81biynHAcxk/rCH3FQ2+pcs+DsTKV0UGv
gkv8zM14vDUkNyGMH3OnmrD0XmD2WSx26m2dr34fI1d3hi7SupZuCV5rKPfkXAaG5GfMQsmV2rwj
2Kxe/+hP7ujGczQW4ACcecgMFgMgw40h9j9hfefANYdf3BzThgMrBeJukUl4zBaxYZZxgPq8zRdd
73NOTUUQ2+rmHYFwM0bWhuYmEVX6Y+u6KYJcfjWSjmGzs5SeUu/sd0cumy0eD6G7WgRBzMjx03Yo
S9Dtln4zlDxjQgiMeqbrVpBKZfTkqZLoRJLR65PUD3wEKmyGBLnf/AmNPRjfeuh5B8YkyW008jQr
/0dcxlDIFRySZ79njE32jMgb5FgKN3gEPyscB5ZaMKsIXith7deGQRkosOsWUIk3r/zW/q6IXCiz
P6RrsSQt0HLO/R6qmDAuDBKYzmyY/EN9jLdIBdf2SU9p2I9+vLJH3kuYaOaJTVKYWjaujHi8UsZz
FYG0od4Tr260w+GtYOnLfAfigyMV8IIXlrLjmI+D4qtibVojGkdjlLSz2FtAcx/6k4xRR7MdrLz2
del419StDhwqI0CS5NxzFc3cjEuPf6aW+IKwvYrF021KPglScsV3nlnRLOBx3JqEmPnT+GJcjVe6
HhKQn+kzvx1A+77+RNWwVQikGSZglH+vF4jptGIa19KuzbEQ5xZ/Bja+awlz48DYFpo6QaBEHL0P
jIv2KcbJdWVZEC0AxpL0Np+y83QdAKwWvZP2cQnKkz94LYAUIcMD9ozNqAxwy0aeRlq/99qsklg1
8lTbZUkZS/dTNozoQtc7iNakGC6frXKNfJpBPoYOdmtfcZiywkKUkWLy29CwcS/9AlAyoLCAzVS7
g+Zx5Sc4N6e/oFEcxZIeB03DRbLYBYbxjh5yqC8WFglG9zAl8zatUdJt3aKXCv94DulNJ4tVDQYD
TyUoudAw0jRNQoBl8CP4zxUwVmY4eVrQty44mLBngfAUVmV9kes9nkpgBrBN32WpZ5BW3w13237F
+pE61ZjcpHDOWCTuBWZtaWoH8g54N3Io/vtPHS1N7heDzmL8ldrQHBgq5uT1H20eN7sA+Y9EffjY
CPWgdSrwaQRhguukgPZ01GFbbuxzslY0Y+dzjJ7ZiErtzWTpgu7akovMPdiwupxjWbPAQqN01r1S
+GTMB3DhCwSNFed+OCfux3jJ/2FOQ4xWrxR3sy3McbjcXJxAjGcdZKBw7kytrqbmttZq0btu95zo
jlPF/iicBXYx+WW0OYYyxhUAosM6IT+4H1TmXNtfwIWGV5odvlc7zyG0PuIGARtm8IM3vaWophQY
ogQ8BfW2sNJOZqwxQbyrnaJQrrQn8ypzJ62xuql1fsFrUF9kYKlcWynfkwQ15Q3nnAk1ik1l4iGm
Ks6TtVTNezKij4DO+EFLDUwjkyUs94pfcX4fUwFK/53/TN7W+ckDj2ElCUMdsZv/Ld4o/pzj/lb8
TsqTxaYU4zjz7gf8nZh+tSkeqRXDHbq55O8escexZWOGBU9bUN+LOe8I2u1NqjEsttReN1a09vqA
xDK/RmTJNmf0a1rMJu++mL0CKcWT/Cr50dUY+pJRstHQ7crvMlrcNCHNWZkS/0PhHFPOLF9vv/Wf
ls6rDgwRca3Hkq/Vpj8JGqdszP1GYxES7TGWo6ur3eFPJxjtSN08s9UHsv22JbbwbjvY1vSU9H8G
DMh3Zj/dNTuwQZPEgQoXD3nfHyKg8oywK0oHk1KqabThC4vdj9Fi7+yQM++hLRV7vQFWrlPumxzt
uwcLzUnj9YJY7Zc5mOAm/xxaAbaK2bT14YNTCXlTr0AI9ZJkaxypYPG9cBZXFXf4xC5LBOQBezmA
dQcXp8bW82w4CQMCszsW4YCE7/e3g5AYSckWTo8L0iXkVbVVk+SnDm0AjAHn8f84GRy2tVgRioTb
fCrEVGMAcYokND+3z4Ogs9lR0LGfOWYVkuuc5AfeRfaOlCAVB2M+uW2k3vcOPphTlO4kAn6XdHrY
PcB5+OMY5Y1g3Rz+NItqkjV9GLkzX4iW9dQoBYEVf/0+2r/1pb72MnthYvBYPYhtHIFl2Iha419q
9tG47c9O4No+duSs9g6hy10N3FCnzzyZR/vz6Lbz1Om/8ItoirSbtDxOPh+iFept4csGusrhg2f5
n6baXmL3OOOvxQABIln3LBBM+U+YFtdR5RekGPphDlzYB1ibB1l8UWFbSA1Y+T12JYdObsRgOBWd
dl3upQbW2JfRZpORUC3oG+BghOagtFWnkZ73MeLe/fBJGVJnzB0VCzDISP9IvhfHxWwea8oMthD7
ucHo77qID3IzmEKV3k39OtAIrK1Y1E3bp/liTrIJ5JAB+vCuEQqJHAyGT/c9sSQOQZm/cOWQgBAe
W1HTSy1BcorAdXuubHW1QY+1khDr7eRPEvQBb9mTEZEy6n9j0o4wqGWqDZgSybvnC8qhPZPEahpZ
9+BLLZXcD/PYyG1S8KemM8MP3wOiz3jCwAeaTB7LZ4IyL3SDXBSgK94iJ01zCuIuL7NUaxznKDVv
n4ll5YdlFh1Q1VAj9l9ZqoNzAtuWmIN8ELFSZ7GesNgg4T57M7Eju5rzlQ/6aGz73C9L8TfTl3X8
EsFfVz/bL7h7PG/qjp5y3z9azZDbyalIIKuE3ikHfRCwftlY8IgVe47ZFWYg6WehDMBsGXnGwBUG
twGYjXqQ/JvxfQgpnqw3j98xvKaBXUTStbHqltpGbijOdquAIAtSeeMatrPBRjow07/uj94n0sUj
XZFNn1cAvjSIMR92bCiStuqqQryNwZS8RmwS+6Z0q9U/dwZVWK7dDbDsM2qQuJfGKvnQHtlMxwvm
XmPnbTIzc+voU+AepZfMswNsopkio9IzDD1WZYxwlfgQajPlfwpKW5DVMZ7uGih0V1eoB53Nr1li
5Et3gYw0DGcMhC21TVuh8ejUP9HL5QPdGwldRW1j35NsZuJodTkm4AoHRG1ipcHvGQdEtaVMr7l7
XzxwWGQ/zxV9zRMiSPVvDYtnBLKi3zlbsDDee3NxwA/UnQJrgXPjJEvWDslyCBVspWqHM/2DKF88
O0SGShaOK9+14uSxAai+zKH7six+ZlMMSwgNqPChyn0a9ohUyutXGp6T3L2/kom4pLX4ySpOfG7o
T5YDrzYuv/HkMAiy7okqbl6EX8Vzj9L6d8s4OASk+927ltiayIn8JtIILgSwAFPtFPJ3RWFjq2h9
RjjSP+jawku8oKgXfpOiAUdYqUWK6eJyYSjCXIyswJRhz1ICgwIaMDy/nPNGNLojyn+7JDMPRO14
JVyZf2WsiRCJt420GuLNrU6JVqKkQ2v1cDcKYqcG5LqZBwaQH9PzouC1yk7lMuX2I2LOfDHdnZm/
kk1TxjEWWcauIztLm3LpeLKvGvmefMxntEqMtbjtdmFbn61g6MTAJb7ZhqfU/Xn7X3dYvlzT/9Zo
03llffjqO29Q5/GSaMvZnBBjWZCe4NbPpxCwGbvxboNM3Xxlzue4akPngbmxrh34TfJb4QMRzsM3
zeuKBiRltOCpeaVu2+1P2yOyfHXqv2rg/mh3sxTZ1V1vWfdouCMN7CyWAArmkygEzglQYIBMeKMS
O2YeBGCxIj9mis3tFOpeuPiJ+CJNmdzLQtsrfQPiSvHncf+Y31EMrxKE8hnHksa6orSJhWLkoTso
bB21XU8IKe6v15eSn4ioBCBhos7cq8bZiPtlWjCt8UfsDg7AMN6Kd4LA4bceRyf80NY0nBxBQA3s
WB2GrxBgFxjDPYjojt0h83PlO+iQdr0qxPjmxnY8TtESr8GnY8T7Asa0UBS0NS0Kdg6eIN77+MRf
5RTQCYln6ziXNLfCys/7WZnaf+TmDnBNXOR9lunt665fsEnz3f7P7TyvxxNq74jZ1k0cPAkVx/Ly
KughSm/BbHFYxRhtquVDaJQ/dr3C7FS8Y91NJGSfUG9PS5XR1zymSdZpEjAI7JVlV5VkUfWYjhjo
+HdnplxVIYNcfFAfe6uB+AwaFiQXEYasWbZeVGNhwAF8GlZkpqfFJuvYVc5Q6b5YxSVrF82N+5Ux
6p9HLJQD1mLAftygSsQ0Qaz5eemIzHl8iy/aM/jmcRLGaAQxzemMdJ+BqqSWegAhgfE9iEFO4deB
dU9l0L9D+oIbfERWJR6q8Csq0qQdWeQBixsfAOLk3WuJmxgbuLAs52vAvgD1Qim/LjILQax1wUj7
Yzubof/5xl4PuTGBGGxNb/IAeiK4LgVZOlhEQ/UVP+/NhQ/zjoTqNkoJ5BqUBvy3cUdnnd2TLMwi
Cn93INGbCe9nkZCAf1Dx0aiVemR+KlZ3ZJagbJZL+RuLpvZxUysbSTO7TKGkzYS2visnVrNC9pXM
5iytVNQp3LZs0cPgYHyvnMj9ferk57l0XmGj32SyCXEU3NyX09APL0bT+9BeU8EGTvNzt/gYokl4
/+uJf9Ab1zo1z6OlTyhtPRTbfWhYFljauwa7VKAlx6TE2Ue1YPQkBHt1ShY13wpXu+6M7eYilExc
crUWg2n6ZSfxfEkyEQCe6g5eDpXR1Iq/FwIzR7V8Vj5Rbggr/RynAhbUKyFdoatXZ/4kOpE7v0qG
gUjQlyAUFTR5LBonOQihlFL9pwVOQnsdHOyaVt28+hZKcnCAF7D0kTFT0cMkSYvLeDgAxm4j4pgF
ioLh/cCWris1myCJKwudx1lx6mTOw79XPpR8nZ7lEKxIPZ0smkOLVTXwMP9/txbIjhjSGSjRVbXO
l6armUdXZhURJFPK89CsAg0p2AO335cdWnaQ6qiy8Z66QcocbXyGeMvdzSsb3f76n9xy+4DBPsUd
jWOtXqYwLgxJ5Q7RC6PEl1U6Te6Yy1Xp2VFjnCDvt6CuI1jJ1Qjk+eGrqtZO8q940FkLyxXIeE1m
Sgs5GT4ZgIEshG+DWsbqFrjfich2gC38Mf/e9tVsHT0i1Q1Ryc6PVCz5lq9APKDgdu53Lje6Dfri
lmydIHmIg6N++ommf6BOIU5wffcRU3T/gdVsb0Q5lUNFUS6NAseNr/DjOpeim6vPImTkc78RA3sp
yPos0Oq7Shr4e/eCBwFNg0yG5sQ7nCt2WWuw+7KMjaf6SOGFspqceoliH5UnDCpooRY1HeYYeNK8
fKuefMelr+25a/y2O1b7YJp0YdDrzd1iCpDIjqLEvg08wBC2dFd5kUmrmSMkEwch7rQhUU/zdU8B
KRfmupUQP2r4IxwZYQzhE+sQfzOrPyCV33qd8BSl6cY4V8HHoiti7c9p6A8vz/7di6qfdIBvwgvm
iAvo2OpZIXIzhEakr3XGGR8KzX0JX/Q+yr+DGZXWR8WutV27m+/N0HVfLZKhNnX6V//jJ+EL00bJ
8MKcGoMyGelKSIQW+AyA5/4sTaNDaoo2X2Qdp3pn1ZfyK6EZ9a/826Wfbud/p1/TQdSBtjm6S8fk
oxNJ/U9gwiTMYHplVXNoYuQ9ufu4xZZiCbjM0UuVeEOOOQkRGhtFW10xXUNe4WWwO/+uxZpSnjxe
R8WyNNHl7FYhcEMkbOzf7Q1rcDq7eCCzDzWYTEIHoQGi5mSCYUEiVUZ2+wbCpEv52zqML4CZPDmE
j8xTOSwmOkQZg25liBoZFiu3T+aCW0owVLQXN6cne72jMFleDB6zPcsqyp1g2MEpiiyvXujRajXC
gf+KXxBaOW9E1Gm5CND+8cYck/HG49iOVdp8HWV5kYKnnssAzTdfyKhrWWMHtUYayQwQUJkM3Eay
uta8C5mYrtFO+Zlyf4adJ36S2Wlpr7UCDylYcITJBV6YY3PBGcqT9gA7pJwdERRfDCZ7JjkprgZY
P0w62iHyXNOftluR3+IixLuQ8NQcaG23oZZwzDjTq6yvoatchvnhEQ99bGU1Ple7CSuzCVqyVdJl
esxNmDuikSSlsqEKBNht1OlS/s8clRvajhfyyeziV3Q9EqqBkdwG0y0j7uPWFtB2GNdOP2EIC/6F
+6n3yXc3cbMu8w6WgHoyNoy6tJp3/jBxLZcSo6VIwrapnYEjwzhpyoZG/kE2Wp/ejNbTLGzKqXhI
XmxNflhpF2OPKlbtaIRa32daM2OjUwE6TSuAlw13wmnI+kIzzd0qmH1Fqp5/r2lfZNRKCbOwV/Xw
gpImVpkGViR26Kvlv0kWIM7/tl4iNxzoir2+m01iRjLJFk0XbkY8b9HmGU1vrB6SrSrvnvCswLZA
Nnbhm74WmdTyYNILtbHDnWzrj1zIntFL/lHRrGeAFIoIX6pfE/ayeqSQPcYGSRs3lFRJZKdXwOD6
ltdC4OyKGnxo+pkJTuzw/hEUGQVXTkcz2fN9eckEbGIf36bgzEWm7E0pOKcU/JyL2WhSQX2abXDt
5SzaqOe7/D+53GTktKGBGcfovECO/FOIMl19Dl4oc4Ymh/BRFlE8oD94QeCdK1MdueAN6TtdS7xb
4AUd4rwK6meWmiVF8gr7B9PnQ0X6azOX3ltIVzEKCrd7ycoteLY6NG0Q1iMHsi+kKjdH7r+D5bVI
Db5eWC5eFjXzcSubCYw6y0ZW4W9FksAIe6+r5NIcMAIbe7V8fIWb5NHkawfO/Lp7s40Wbw+PJqm0
rYtBDMozGwzruw0tPCLsRkNskanGX+ftXiMEuOUV1YvU9Fp+jK1FE++wR8ZSYhFdE2SkMSpAnAef
8n8mwlKmovuNJ4Qr2D1QmjRh6g1AhQMqzHBSR5ZEM2ZYtJkRbPTA6RBMyg32Nme0DxfYijYE6Lx5
m/nrLDT/A2QBea9Q0vq85TeOuGbN5E+52Mzp0oIBtZxRsLYBqCKwtABQAJFiNQWIlstdmlHm+Unj
y97woVVLBciSOwnhCBvB8uvvGrTOnV1r/t1H3ENzZaVyHPBpxHALpkMhyiAk2qrY06O20yHiValN
x/2Rnvbk1j0JAdw3MvXa4rAKMZL2YfczFxv8F1KnH/GfMdXLPD2YRj6qIQSUQEBhgQ2WG0P4XKbf
bUf7LX4taS4UcMST48SG2uVW08AOXoaBd3QJvOx0iVgikrbNBjRwKbdaD6s9sisFZPQKZXU3IMO0
TEUFGUbMF8uac8jPNpZcD0uYrVsF3NrzvN1YzFnfh5gpZzdBfdinLsSY1IxY0G39hDH0n3nGNs8b
ck2jLum6ZD/b98bghYIc51Q5WZdrrf7P8lXPngSWjqAleHq7if/vlGKofbFdnvjEk+mlZRRmNeUc
C0HsA/ZRfYqpuBdTKjmNPuN/2iUVoIEzOMXPphMVQ3YKoaboXjwrL6JBgWjAlzq3TKrlWniT9y5O
HTAmzF7RxmPg3MREI6cRMSSCDzm/MnXZ4cRKcYpvdv+BfFWh4SDb21Ra5VGLlNeMyHTRhmeoHrkc
ajQEuAKY6+3uvupHEqCMiNm88/n3MAM5xS9hrwIs4zYPId6+V6Lco7SFwUB0OezIvdlF9x7oj1Ub
EBXzHT2jXn3TU+eS/8DOLdywNOfHlv4qx4p9RMMH8C9Du8BMFW4gt0tqSUlKmFuE4mjhmctkKO3o
sYwjP8RurWt2kLSqS/ilQTYzlYI5fkcR85KMW/qYbqXV50QOJmdVRB//kpOAF2i1wP0e6pA61vTx
yI2xtJRmqZgSq96zkTpYwlLaDkHAhPZV6NjirqzylNGwXOdoQjoRHY7iNE3J4CcyLmlNYuLjPsE6
JrZ/bXhBgtbl7qLEJfqfulNXz3qTP39wWsK4Vwjwz2He5kW6n61ayNSDrDa5ua1gVAxGwM3RDSmP
W6Tmm1btmzetnsqRh1ZR975RL3E1QbIf8HUKO03rigZcRB2TF+VF5F8PR+yxNeCaJJqqpxeM3ACK
tPFDi8H4atifMCi2bQ6TKRyA1JnlLGeplY6soUzZR2OSWfazCeIDor7jebw3AKQ9gd/uzUfDSZun
vqAtAIsMW504fAO7Tpal9TuRZnMA76dagV2JXa461XF15dP9WbjLfVSNVYtdB80j2yNid1TnAQMw
K8S600lTkDvWjQYVlV4YbLC14vf2vWmr8QwD+A1jWyfDxMNX0KMlMuyBfKhuxP7GWZCREkt9LO+g
BCVV83urNnCPxai2fy+R/nU4w+EsuljJrPU42qEmclsbOQCZwsHgLIuP0k7xSGn/9ZiZRPJicvzM
/KaMmEPIhb39nOYwOf+bKUT2NXZvA2+VhLdppNWHgQRlPwYigrsp3KxZNo37NF2Iwgn6riOwFpnY
GaJBzMoKYA/aSITyg0rzOcfEnlFG+w2EUqR394omAnL6pEoQuvxUIPO8Q5xWl+/vZc4ffV6e5FsO
q+A0dnWhgRGAZSj1UeAymlXg1kcnv9XqwjJXoGqvMkWYKlJgCWBeIinePOGJBXJrfkymhUVrckAg
SrQ0ZRQKrDCi9WesBdFAEzwGuOYOhupn/r3PncH1UlY8B/CPpMvErQ2lL3FuNpzEBe1F6SFmuW73
Sk5K2qsfnG37XGxCTrIKOHkhmrjufIqhFu36Ebzq7PMuzO0ouBajekukt1++34OKqF1Qt6BjTe8M
o4yVV8ob9pJIIkIEOCOub3TXgBF9kScbkoRJ895Z22PUIMbqB1ZObfyaY/GATTizO4Xq69oRXTas
xgQkQ4Ywuw/2U3WZxICKBxJCJxkuByKfReNutbBaEgtGvK4/s/ozT4RQkX0NevlSDHYlFcTLRLtJ
qfrLWTTfzzcnWgiMYfyGCnv7nrAAsr1vhWLu6oV3pkAu4QNqYdrPPeGVQUCIvEiP/6c35slObuqX
XLcVThf0QhYe1jvYlJ0CXtPYtOLAxSaSVMZZu1LzQuPzM9xqaK++ojpF1D1lApdaiLFRSdW25O1D
0Q2J4QKck7cdj1heD/KrlYKMG0otEBTERJDyB7R6dYa3nbcwTzN/zVRcPUd9VxHnwUwou5kl48XW
GFLg8ZTPirj+CEes1RSrrYScepSmP6XNLSpQERZx+Y9UAdE5IbYmlF1ai5AXgLXb0qeLpck1fyle
bbWwzwr56QWZMYSuK+uopz9MlkqYQmptwgh4TBN53ZhKB5AGqvU43aKOZCT21LXqG6ew1CMI2F4r
z96T9q4DsYafGrlWT4onQ42HBjenycszf1h7WuRrqBZQ0N2npAdSI7C+I5iJ3HnxJ367QEitxUE/
94DtUV7P21Qaq3xGU4OR6cidOxPDYGA8jtKIku1F1Tr/X33SRDEDbgbjFCXCuSXlKO6oH5wXTnB2
px2ThfYbRtNDJNZZ7rrzbKiMPSvzvQTMeX4ws78TuoG+TnTQgodw9Y3MAHYpQIlon5wyAeD+A4hb
B9+lNSeERVxo0kZ3Ig0MZSqMoBJTRnQD8aJNb2CEEbevMEh2Cy8gBJMV47LCAGT/a4HKPLVzoG6p
R/h2mWcD2Kvxp3A1x8dWpF4eK9offsBmhkZJoy7tbP2/r9Wm+UB1jLKLy6WZXVw3wIjgG2pPoX5Q
xFiFf0wAlNyzzro9yURseItsNYs5VCvSqoQtDPYixHBhu7H9KJYSKRThJ1tomeLmmodWpQkBsiWq
crtY/6BDEk/o1JZI9BCaOS4qrfDcI1vD77rkH4rOeEigt23u4zBjt5y6wdppP4b+EzXKJl3pKI2d
ltX86mClVVTQvZb8NS/cKzarbOxoO7sp2TQYak+AjqwlW0c1KpTKhaoeyjMp+Z+warFE9XHf6wKb
EJk8OUh/rPGLYYApyoKkvqSC/Q5PbMwfm8kuZhdAnrznH4NNdSgwVVWzW3j5SaTWhRwaHou+IrRM
wIN3sBz/NLDjhuXEnvVACH5LANwoCxGtY3j90jnRYiqjj+FF77FvX47W44VlXF1qlft+SRjszowJ
P8L0AkGblJpcH5JUvTIOgW4lshF70gcw8HVYWVv6Oiu3yL4mzS0LblTL85Ls9UfAr4GY7LVkLLYC
9KN1RXJKJ5Vx+EBn6pWVxjFHys7t/5CtiG/WrBTuQSN8cvGaas3rb4H/IAO9nJtZ4kbl69SNh6SG
3p3pBBNUSXn0eXU/IXyV78JvRN/VbRL9mdfUO42iIOVDs7B8fozhMZk3ZtsxcVxyDZZ/uRE2foge
wZbpFoH6k2Udcb75TuariaBA6SWcjGGLPtGRqpA1KVMeiZumdWvaIH/Sq4ffrpwd5siDjRfiuTCN
UlnAmETSyc4IbxxyGNwCHMjL53QV0zDMd/C2kZAdIPVgCyyn9F6Plw2fcgyJgUGfN2sJ8g9qSz1R
kicex3UIaotdLhRWkvKjMLIxxQ8XUqBLqLoeIiuQNLOJL2g3WVNYKaWN+CEGcAZCipoVLj18d2Sf
eV7Vh2H4I4+NE4egUyM8oHBpWjjWv+QaJSxkHROw7PXMxLMAphw3pjs3JoNtR3unj2069oLniYa3
lbEw5oW9y+yO1jBo62nQsVNKNM4l9nd3kdNYAUyxSYLARWG6kgolfgYuiJSWnhAl2mxk+K41rnqY
cPi8HInJKkHRi4T8NyQlGtYHw/7DyYo6rPx8S4LeY3F64+N4lxiduHJ5wLqAn7+G1P4OzoV5/kvz
368KpycQS9yjbSHEKxS38Gq061FT2pweEYl7Xuw77kw8mThr8CVrF8e8BSKy5Ia+SIQg6Y2Dy5Ui
T93Wcw/r7GBzdQBA7NLXgyDW3t67OHttN4n6vbOcbpiT+9Xu6Rz07aTKhJMHBLvbd08kym7J+BzG
YmJXGcJBLpCwCkwJ22hCd+nFIwh8MlifvcWUuckreLD8dzRlp2grMcYjJWNckYCeyyTUKj8vASia
7CmAK88DPhlYkjNtW+gn/ZZV686QULC8VKwsGoL6EejdWxOclyIl6KSTmo8RvLr+1J575WAg32Ch
oA+ixBDjmsj2Ud2w6Pl1uGxm5o5+dgxagDPK2MGef5rHAG0mj16lX8WSGvHIp194Tl9BDb0EJRhM
b1xlSjDgaqB4MQE8pUsyf9zwtNzH+2enmniosHJtdpyqvv20J4Wzq8p68BazmN6vnG3huk7G2Lch
m0KoWrDQocAZ7SJknIax7mEDjD8O17BvW16+nZrX5cicOpUDYW55U1/1Pb3BQ48aAPWFxj3vcvOw
MhbvyFL8PJvmeUqyAjNsJbkFrxoJlVnI4MJHMzNRzeXTcWUTREtMvEth3al7eOJRMGCVdYYUbERK
bd3fYZXaA7dlwQouVINUEekP6xXUjueHgI4aFbb0o0kdYf/yEnHnBtJe8njKehMjczyp1j8Ws3py
HMffa+vdv3RpzB7nfHLjVH4Kt06vsLtJ/zlUwBN5dQiXcDLlB+Nnzujn9HJPoMl7axQoWKisDI1U
/tgb1rTQelicSsi8KAqgleE1q3b6ZUUNAQvOR/UTvH2RJCtDsvsnlKbIpkSIcn0WDR0oolUOs/l5
wKu+5BX0bwdyJak+MqzbGhytGJ1EU3pb84lip3yDrmqJgpi37iaE7PcIRta1CGzoS5uFHJn+0VOy
/vtOjJRH6OOo/H+lOT9JBtqDfkqJXEEC9JUQVqK/CJmDoj/Cq338Y9L2hS2yVC1/dbwYgeZvAhx/
iLaen70dLZp5MjANqaHo1r/8oGHx/oaiM5Hv2lfHNcSHfGv1QvDhTeS089OkzQdVsYB3C89K8ejb
6qEFALsAw5ZM5PBnb2Sti6ejAIyBc5LWl1E8M6hsAxuEtHGd7CVcDHay0Lxh2z7MII2Y6tiUEJTN
8R4o0A/8iiqVfW46ym7j8042zR+sv2kGeicEUqwfK56N7/kOD8de7gs/fvWxNdk4bteoMKQDEfWu
EerChMu1piacFuAk6EfHHmYagpXNBsU6ljP1Q4jPFM5ULvCYNq1RIXQWeyn2H8lwhFPbNfSXgB5i
A+8kQKImZOSumPPWEt5tYLiNx/XeyThqXAVTxoktYwY5PxfC3AiqzaAWhPcdF4Mz/i4IeQrGe4cY
wZL/5SG/5wJFcxgGDrnT6hcn3fz5nD8rGByK09RoZ2kZPQzy0f5uRbRTS7OnArvNd9kOBgO33MXn
f2m3qsBFDonS44+XxfZbpknf73/K2msGwVwZV+jLLOjWXavfX/R0wa2Twd+fIXY6qZo+xYYG6gIT
AOcWJXIo1vP1un4Ub5QkJHybjRt1mVraVC/cRkEYBCNFSVvQMXNcewdv8YhGTWPhLWs1148wSvAy
U/5cYbfF80qEr6PrTSA+MpPxv5H9gqaqF4V2lf/c9REnNklZzGbwdK0q3UhqwECm8lfTmkbuEN1U
ZQCfWZcWPHclPVHqtyo9vajPbRUIf6+Jbx541/DzpnauqaQ40KzFreQnAX22cBBV5cX6nUPjq1Xu
bBI4nNK7tT1zKS6iDph/KdM7vo12AN9/I2fp9hoyNIu92PztzwwMCdpwQ7k/KSO880YYxxix7y/j
lwxIqObSFwjBAWsWmsxq2+qNOTaUvS3nDf4yyEEIHOLjIVMopcIFej0tI6odGuT9B992FNTGljv3
hCHckJTDkX6MJVgHoYdQeDNTsfBz2kLgAUyE1FiV3xnHLZjXO7HDqmQ0cYwjHfbdUjUQTZGNMnUX
bNFivrB05nizRq58jUr4e6HtdDrNqjXMl+SuNAfSu+LRGzaVBoStffD78pKhvq1DR7aN+FJ1hey/
KvsxnHU03fY+QXM6OcTGK2/09b6M6+LfUoekRUppLF3yD8OaUL3NdWzv60G4xptdtj/INfUlMRjy
Wg1xNWgB68xH68+/ZOVGCtjhZPeWRrg8JGZCbbKajoxPNpCpcmJ9yAkm9TYE6w4X/ljF8IA0F+8R
xtsko0ccmW0s/5ziv/HVThXyjZ2pbIewWtzzdIB13Z6OrCrBIzLVbp8ua2DTfNYQFU+uA8ibmOri
rVa6tdyHG3xLRGnB7osoktfMZctpvPt4MBxEDHmBUPd8ZAwurLwNW0Qs5fhOcbKi72nO9fI/yUii
ZjCdyv8Ni0/HfDqU6XTGBn0N1qDqsAV9lUbJT8AW+GO5VlmJSsDByMz/sUoGhtsgkUjPbbkWZPOn
SZm3E46jUlmJSdPoEqxg/P38SZDMPya6BIpR39Npjymkt5APCoSTplw60iAdtb39JFHndt0F0q6p
P87VZlzA/qQqNKwf8he+XxvttdNkk/NkLzWs+zGr6Ew3iH3EB4uGzDHp2Ccz89pfavyYxBTzwEon
SCJgySx8081FoYBR16rBRXqn3f9V/Bh9w458YuMdf6dWBEtPCoUoyNNasNSNqr4xbs7x5Z7KGygr
uRM5202OhZPietLFmbb3Ns2lZoGCWfMNmbBc4bmQwJYM6KgbO3blUWckXwLJdd7pFa699JGXbx+Q
cG1IumzjwfuVA6coPSuOGjaMXXSWmITxBCwnL4DDOkVQkBKb7/u3th+it3JJ2gOw5GJF5n1sF9CB
T4SgLAsJ7wNWN4I45JAvqqi+w43HZE+qMvpUP+y2n651E27ubmJm9z13RSmbcZr5syy4ZAJPqUSo
PwqxsWDdAyz9JBvEXfmqMmvDdHVc0WI7GwNf//Rx4mZ/8xNznIcx5RRnKLyG1TVwbGpCLMMpSdLM
rPft8zjjwXyh+kMqWRW10jvzHaf2Du+v1s+RQOFmkIsmMic0ExeFvyorUp+226xk6flblhet5AZ3
2L926a8dPyZkNNwYCNaGuno90EBCT5RopVVuTlLqaqb3vrXQ+B7bVEwEDw+W8q0xqg3bCAz1Fyyp
Vi/FHQ/HpbfMIRhFhDaARXTDGd3nmR3vcvC7BqnRqRDGLp+iH3BdC4DmoXBLl53o3S18zix51EJV
pyICHnlkdeM+h2lXY2K7H+/PW4TpzIxmTxGZRnSlkQpo/1nAlIoLDkJ+GO2yCeDMK7qIZ6FRD4wS
dg39OnMqZ1tNdvuxRZ5jPVSFFa9LU/CVt01oyWXghd9CaEMwHhkUxIaxqES/zGwuUYvLb5qMxK5x
8tuoco+QDXJSESVBFZpT4XTVwusdmDZhNtg6uqrM3LldbZf/wAZ2IRn3LMlIzHv9Eq7X3APxLDqP
6FN1Zr69gjzmMaRwBUPsGgkpEe62CWvGQmmF1IrSnuQnQ+iWCvxYMELIkluGblTL+j7uFWiN6b58
BfUua24cvJej5hdbRpbWTEEMaKRohf6yID2f3R0I3PUCnZBSgr+BtXYwPidNv8XQ24H9oclIBpfi
TgFB1J722Y77p13kSK9fDEYGLn5pSNOUHMZwV87OTH3tq1F1n/bBQqOGaPOuAPOBLQLhd6eW/rON
H/U3AADIZewVOmMFETXxRxO+3nqRX9J65AjVG7/81LCmQxTtHf3qLrKhRMHF1VFTtarGoTsL+05M
XID2CDx3OlOF0D2rSb4ZxVYDTBA0bK2pEhsDAuIJOokLwlusCsGdvXAt74Wpgkj0HQFX3XinTqww
nsj0cfscc71nti/PKZfe+cj/3GdaAuihNCpuwaAdnOwOzj37ifGlp3qbhgHa68wS8MfKQz0XQ1In
kfuoV3IY3YlwKAEZOwakxiiucBnOYiG3QS+yXm4NCuUZPsZCGj8GMb61LgPoxd71H5Ac/EuvSun4
cbwE/c85yOrTgp5kUz/TnMHcK1D1EGecq5/rrzoIk5gGwPWe73L9DLI46LPxVCA1uqc4EEjOl1tm
Vg0/WQDdoC+mLnI9YBw3GR2phw0HAYLHRtAQgNbUj3K/OTUKM/7Lf0dBhnOq0AhYD3YDeMnqjBO6
+eLK1TOtfmcqJch/A0/LJn9KRpY+5BypFwqKW6e31FpnhUBUKedtaBdmbSWe9/mFKlJSbJbxZgAT
yaskGt5GqbEfMYjIReUg/OPYokwq37TK4bka39YjizMbj8pzeiPNhVIwX1yEJFR3LwCYgEBzmUfP
Yfokj/sk2ZwpDdMvgUX6L/G9GuUyYV7kDReUmb9Et6uOokyjxNa7Bi9MlT+TLd14emOEUW61LKgj
mirLZbp6ne7xFVKJOB5y88AYxHX7p0YzVA012aIc0XLxANsNcw+XDX6JemkhyexpFyxc1S5qIyos
2YlvXHUhPfVmaYvdSsEeP6EBig/+k6GPX4pfpqPx4EVWbkX9tNsUoquhdvnTmawQTnedvSmkfrWk
bOoPT1QWb+T12+P+yhkEsI3Cc/3uG92F6edOE5pSzc0eR6yXNu8u4mGJ9vKVl6TWDi/YL0g+4CV+
wxKYmlz9Kxpy1bmRQm5UyPtxkaFxN27rBmRWP3JQGwWEaWFMNe/zZwvbdgDP6NcuU6l3ju7I+eEa
1YaZe0SgM9LnvZRN7QnzYZZrprXVtmzZ/Oir71CC75ONPgiyiuU7lYjJ3XVyC8IAfDZ+r2RDMYGh
pUij9rE0Fu+U9rrbX3ukETuldvcyjVgakychhKmuk/KR/Y+23ATkLq115sdOEEpjfNUFLdfDDToy
Scr0FRlIGQmEmceQ918Ud+zhFNn6v0yiNP+eG/IywlM4MC4iw3g/5OxwIoQMWnE3hMO4lwrFUXzJ
+bGE+qIljXgREzFckhds31dbO2OPUM/tO+SdlJtwcwSeQO92gUvZaD4tAP3qE/KrUNxnP27Ktu/m
SZ8Zt+ZBwY3WP6qoAvb7zmhKHkE/Q82CbyJuZvxgJIWL9SGMEktrAhk0bVc/jCdMHmmtZz2Zpky5
QP0ENZD74EvQ1SjdkZdBOlFbPSNNRAKhXXYw7+cAdGD6vLYrbB4WfWkpM8F60UmWTyVDsYhDy18d
lQR3OIk2u6vWgc+cUv27174ckdT7GVseNjovvfcsEI9NSuEVmWGrFli1JAmBFa6pmeKNAcwQ4Usy
yhupurqtEE6CmGimfO63SmBr0vSDKJ+O2+PxM4nkkfdzFZt0ceq9Hcn+W9BymtGFTIFnheMfsCOs
QEzPlstqbp4N2hvrb/z5SE4pWbj7HPSq4WDxz9SwLQ+CvDn8Oe62uW/fYmgEnknW3uPSz9YNPcKt
55GjKN7i6s++NP5DyIMaL3mb7A9aIo3w7m/L6umrhlndGLI0fR8A/D2CeLDR/nUEJ3Il0CWNOLSI
wK4fRWst9Hljsy1GcMEeftRbT8/1ZFGz/gXVG5Z55NfErVnf88AJiX1CBINmCOAUs3trl+koM2LG
ZaOHH+5efSgTQGsu9YKQUivdiBYNLohWbjC2NiXyn2TgCJJ1WpPU/6fZe1qBFg/HstvukUoKSx1e
4rl0CeLeXjTPefy1xQUJyBAGfLRuQw653ckhD2x2etF82E3Md06CceuZoRHM55MTX9KlHxL0/ffo
DhJuXew3CiEih+cAhORPu0TvR+S0e6uo33K+72GC+DeznkRIyAaKG4rtB9xwkmuy8xaOaSZ+DZRZ
m2WEM0yFDpuz7kAzzz+9itmXrvWkndwdymMgCeCz/U9bm7ZQOOHwUygVEq8yoYINGvPtaxKFc0Dp
glkCun5bV4OveWcQcfeqZc9xyd8dtWicOoBJM0TplUG9A6UQfvk4fxAtnvxLPEzXD90elCiGgGzy
81rgxJWAazfQAXcJ4uIVazKTUpgPwjzvPZRhzXjw1DMTH7ON+eL+nZ6A9h/OgQXqz8cUgb0mRvvk
ujxq8JeG1TqnuOROv3RG+UwlHIIYijqZFiY9/z7C3z0xmLSoVGFifNaFjQ5ujjOJ4zouwH5gfOQ7
mpbJD4oq49HYYnAunZ100nqNCpiCiYYzAX6KFAcwNTZv4r66P/dfe9edNj2lxYuXvEYmTmmFZey4
WVNiFbt1yxOgQfJlPuSzmgVUMdoZSzOwiVFIxh9bKrcxvsxiLgXh7V8KO//0IoPmOJNSSMXZpjUN
FdiE2iE5pJx2AdoEsJ2BRwAacJa3Ghfs8sidheqGCRicN2JP0vo1DkRUxcADbuVoAmwEf+aiMILo
f3zbwabROjpZU82U4XzxvGga7UG5owTAOxKynQs4cOoBrpiBihYq1PNiDp5hKqN27Yd4tXmnPfX6
s6MuOf9PNw5FQ3gz9c0jU/bbgQ6tbIyPxIVLyP7NZp6hqjbkshMhxC2d+XDCjAfg2wTxvOSi9Xpn
BTULnwKpiT9k6czkNWrecAWzqn1Azxcr1h+9H0GRp6gSt1czbRBxJU9KmI/deWILZd+xxk3TDiiW
blq5O2pNegR/fHLI1WyqQ/rQsyXZdFmzbMUBQTEjHty1Pyw/Qsdbc3ZU888QQRpbzCnj3oEfTPbN
U7a5pdBcQlFMFmnbDIvckYVxjIOBk0TLprFohoh0WR34E8o+ONEj9YEpmAnjbMsqaBuAaIxZY5s8
5N/2q+tjq+KDkK3EYdisW24qcV7Y8lTr4z4vpAxWfaPaCm/8Uv1VmiI9E85iXkVOrG/KkmnlFJXe
MC0eZUNS23CXqzwdy54iLAPmL2YaV+/+Sr/r2kPmKd1gM8PGWtLfI/Z0x/jq82+laZj2C6vKjDCz
kBoWNpaB4BP0iWEmfr63GSoCXNvYgiTIRenRVg3if3nUn/kzr5b5OuJzhgavWBi6QNlMD65znJSx
BXZK/70yUry/WEbVzauD4xEJRrNheh6yRq/w8bG+O313U9Kvbj38K15GNYdUnV7YB3ccMw4NNF7e
ugPqJXm+mbv61Y7FilaCo60lUYpxjRKbZsWYGngRCsXawwY4bL3DKYA/wltYIsmD3f5F1qa6NPra
na2xxGzjzbE8pp99JvGuNjAmsOhpHEK14Nc66pxEdz38q/p76E4u1nVIoaZYDuUIQdFvXrNu8aAt
CgyAWSqPXsN2N9HVs98eP7P6BZ7WZmyxz9bQxGrj/Er+RY7tW925p+n6WxudJHsExTP6iy9pjbGD
jdZzujWoyebpBwtLmwpc28ecsM9VpOYX2vu1weWwDrYr/Cqla78HWSNxUAdmybnBSLzcmMZ31Hct
yVre06qdIp0F9S8G3KysVF9aMhholmRbfv39kT9XBSSwj1+mZJoop4bTcmwzofMHPdzfqXesKTds
c53jQR8sQ5ZFxE7bDxRqAOhjkB7NpLwEEarL1QkFsm0C/n8qZL90zXRgSyb/1BaO7ailShSM8UKB
vWEre40ELXyU6IMg5Y/Jc4KSLjRyi/NBwI0mwxvh36CFTTs3nE3GhQHbyG87D0yhZAPOYFJeVtuq
ydHUL1M+ZRGEksVo6PFYf197iNvWSBmhO/85B2RgXT+vVaz+rNi60z5wdVke4TIpsrwUtlWO8/0/
rhaYESYr7VvNxuBQPdGghJceFXV7sdok/Z4fgEBoTHrtz/h3keRaoUu8kdysiiooDEUm1+2ZMbq2
BvlwFGexjveuTuWek543qU1uZysnIAMqMv1yQMZiSpAAVVXGNVMw5CY1624m7w89JgRF4PD+23gD
r1FolsnpTwKippWJbgUW8b05JHTDDbsJN2ocH9M0EAXRSu2I84AOJDCGVuHrgob9Q2W0dfFOT3o6
r5vjHd4OYkKdB3yQU/g8EGP3ShggDQq9lgKqkWnE6Z+Dos4tM9Q2LBff3jgq8eNdV4FPlJ5fPxaY
63JbPYCMcFsenW6h4A3gEt1Cl0a8PTTCThppszF4GzFSgUqyKv1QnX8uW8jqZdu0CzhWl35c1qm1
xfqqIRIm3Zf3RlT1ULLCtgpj5siPM06hZcArb2l8vbqBpKLUAmoTCTp8NeQp24DB3j+CP3xuxE2K
CnHHcAQOl95sBoVEJyAttXfDF4xki3m1ktPKyWTibrR0ciXVTk1PeZVAT56hCS/1S+rJIOEMZ2nk
EmW3U+fUAsFwtQEBnvLVl1Axq09ERuGRVxweoRkuslWxFIh5qgzRzpHCFNOihanNh6Q/sGvwcIez
AxhDMYI0yeRByCb5GlsQrKtszBQoJE9fw8D7VNEkOloLhpMoqZZQYW9hPNYLtgqGFgcp09ea3Aof
ZtGBYhpnFKz8gLTgcEbFMtZ/pmoO0MtO1C8uyRZCR7wylr9I4egtyR32EgWED7hDgBZaEv8Xoo/7
zL3ePVzF6JApOLOJXoffeCUb3SnTupfVUTfQAluwA655sk8KNVEqUImb08I02Zb5GU/ATbxAZ7RH
02ehgGcI5CcNO/P3g/7fl+Rs+9baM8I0ivX93/4ym4FKMxpZ236EkHNNYP1LwalpUbZs48Rn7oUK
P6B9ptY9chPTQHMJJgQTMs2vZAvsenMXS+Ztk+Kftj5szgN2D6MGAnL5P2Vs7uL21JeNQtbLouUX
igi/0lN9o+351R5WcYju12mdxzenCNQ95KaFvk4N4Zdox2ch+eX11FRMDPaswEt+dBbtb/me4vgo
4vng9G4M0Brd9u1ipbEIhloLE2cJISb5EKvx68tI7k0AT4/kcjcG0ow5xnLsEZwfCfoBc2yn+oQd
zZL8uWWY1Wh7lseX78yqE5wTAiC+/Ac7YnZBf6kI9vacW7U090JPvMkMN7cxO/x2u86K2wKxCp4s
vDwhhW3EfCj6tNt5nIk8s8hTMa8D4clblKcyxlR7fnVNOSFQrDpPsbj51leEsVH2SVL4DaaQ62cZ
ezVt3HJwnBRB8xyB6prx5y01kRFtLIm851suMyLTHUNUqSWjohXw8m66NMjjZvxEccDn/xvGELxI
+6MOrKYNtP43JmS/Y9TpSMwb8BPFvUQmIuXWlr3cheg3nUZpMPQZDu+Al7aQIG6KZATZUtWJoYVi
wgLjbXBJSC2V6Jzh4nJrzMnrLSnBD+286UALg1q6dMd8AFrmAy8wmRZofRLRqVdPEYld0Rg8y3AM
ekV3ZRzvSjmk33yUqM+VQjZmNpJyITbOlA1fPj0NUdxBdyubi0yLXcbwJPdyK0OqRkBj1SiVgpk8
+XuIAGl5ftBMMXR6/j9ny2wpzOSqeqUecUwBaLDX+eWEjohMI4UeTtZMMqCGIsnfNy+mXn53hook
VXD4bN5YHbX7lEVpSXcvZSUWPTDgWbWh8v4gETvOW9xOiGC/I3/8Whm9qGxmtWcn+gAVl5/TQ7PZ
QDHQXnrs+W/RHITmGD8Rnixl1aSmCBxK+D4NYGU5HTjO0xrmYpw+HXYMEbFqygFjTTj3ZTiJH0+m
fDniVq/NHBdXGAlb8v6AmmRlBx/ZA5P5TSTloRdpTsItTQcj8x/ZHaVqF5eymdqCo0mo4lXr8YvS
+yhq2LHL5CLm1M24ZPR+vgR+B2qWb6E5/7SnWUlzVoaMMcYcREwMBB5CApuThCqNG8WMoxcILYhf
ZKukHSb16QYR0Rqjc/9aMTYBdQvJgu1U9wQ4BX0kpCviB4v9SQ3PnIRufWhEbXamvZPyIwz3DXpP
cUNs4GAY2u/TaetQ0ArfZe0PYPetziq6eCgnvgLrIUmvCQT82HE9pr/E7LfmCwpSFjEzzhNE47Dk
Z+F2jrOlz7t+ZokAo/blUbYLSVAIB9OfayrFdtoP9f9s2Z/MeIoIMMUcERgKZELaml5EdyF2Ajls
kztRItyv1uW8+s9wLFix65CIQEwm3sKisJAFHvwWmVz3KDMyxekbNBuGnoqkrc41J0wuLfBUnvLk
ulM578yzqGRjGF51ON4l17QRggE3jWqxRjAiItn+1mHtYsXagTcCrjWH9xGsrHTS+XuJTbTdPMCH
lot13Xcep1TmYxISIPgD3GG3FZxIC+/jNVc12nzlL4/GgPUnACtxPgfda4zZUgB1dZvOBEBaoLmX
Po7zu9/kA20yXIGTXXP1fiPIG4tLjN2oo/Q2IYpdyq2WV4bFfMw7fjeiHOZd+W/FwlNkchmJL6Bl
SfqkwloMY6gr5pQKPxVtTQ5Xn3f2BE6aY2eNRSuHYrUS2kRt9y9vBFYs0svY+NMuCpaEUWDSKBE2
3QLcBE3WC54DGp6kQgrKMwkXIjG9Acd+6Di57hML7EvwbPuVcVf99RAcPPw4wYIkcSR+y85oYyCH
W036SfGCzHm5+iNWzedIyjb6nK/M3H/R3zdqiaCE6eG59NV9ryuS81n4oTzVYpZEYYFOQQEsl1ee
47/3fHekDJlpWDCtXoExO+kyzFS53gx2jrmySFNkcDfBFpbmZVc/CQlElyhU+x6eBewMChSU+6Ob
jldbvNffRoo6bttSTwFDDfpRjTgU0exQd3L2WfBCoFzy9TIIjISJ+nUF1oYlYe1I9PHuqjMfhuOD
p94dZmK4IBd/CkyjBWWoXThwg1QnXG/wLM/Ipbi0jLtB8Yg8wE3t9DCtlID1jCzp7KE5BMRNDjYQ
k5HAfuDsGeSpna4KxCbVaCkVsUhxU2LeMhoRwiV5nhtfliSgJnG2eO9kXphlThbwNK3OxW74Q4Ux
0+TqfMBP+Z8+W6HBN8o94x3FRMXorxaAtL/SP9M+ETYpy0+yRML3gCv8UMBa4pdeJVFDJJsE/mu6
nElg8n9dxynoOuBM5HYgVfjBjySOn/8LijPYPOryNGDa8dwVTB8lhl9dojgCshwCtUN6DS2zbOpw
fyAwpIAIxYpny8hlXDxwSlX1ICeVPnxDMq0u/RKsenia5cvzGwU4kCqNPn2oydl4xa8ELF+0+peN
FjDkBdecJ3j/OQUeklXOXlkp8Fno2ARb6p3uIHU5zh/Ewi7oIV7a5gvOuMdXPqiE0waFz3pyEoVB
cbrymd5nfgO/K5JRglUb+0WuGQJ9BGYfOmoyAqjvi8SiS7v6IjfuXHiRqSvr2KDqHFgICN4Pz0BU
1GlWW60IaZzQ9Ha46zFTGno+Ld58qfr8HCavJRhRgH52DckxQUKjiBWo7cdLniQY/pNvjB5lsxvN
U0GdrcaHPPSzjGMmP2o5LZ5QF5heSlCK5f66HaxOMMDLuHz30wfJccgUAHUNJlf6XEGa77MJvsVF
CYU4T7XTT/n6XLEf3Z/cCJ1a1gE3dWIjt4W3LvIscClP2EPrHwoVC1ntW6o9zxwJfYBv5lb8giF0
9tcrpIYj1beZvvkuLMxqpA8meOR6v2H+HHRuN6hmm6NkKdQHojAESqhLCui6RbbP4+NMjS4n113s
zjTx0zQMdhQn1mHrLWiiiUN639LrmgnB6vONpjW4ebgIhgn8mf5VzojOnvCod3hABHOwl7TtkHxE
+IQW22//CSMTnwwAJ4Hfg/oePT06eLQU4Ox3qW45dyyBx/smhRs+W+WQV1lQWLVelYFEWZYtUxoG
OyiGHVyjlzZTHFwlDgJs2EZew1Rj7i3XE7QanKFVjv+Yq5HPEMFrIetuiFEZbyslWn8ZG5SxhiqN
XdmNwP5GhRxE6SAf47gGca+HUkzlPVKL76WSAd4gOM5v6gmqCgGX7NGoAFOiTgst/BTAAxeNYwxl
18+J68Nvla1ue3gPZ6hKXVCT0CLBoIlrfZTMCT/gmnRjkj9ZLvh2iZw6IaALJtzt/ykfqkeiraFw
B7qz6bAXfUYuH/uTptLoTsgnRCtEdZLAVIRb3DpTkimp5LN8gdmQSefLd1LYb5S1pfQPWYJsJdRb
Qnxr/3bBi6628R/jN5WBKM/YhjoTK5/DbgKVUIDtGLkqVOVQpay3YMWqRlZB18tCeAkIYn7wi25S
u6gAfLRXuZ43kqkmkEBFs8eKINQ704vZFSiNX/7cmiZLcdkh6Blu+fMUed4dq6JrjsvjzppiaV+U
J0TJ30TVTvoLP+SMNcnx0XQjGU5/y2NzwlkWrRlwOim7E2u4dqm0za/QW92ynwfPFGca5d5iUY0+
2D3hWJOE5RpQpjgGAn6FIeImley0iSYc/nbNTArRh+sWvqz2nIpKPowe0KlvMyKYisXqKEPQCvO9
y9qwWZRGMW3fKn9MCOTWBEdTUcT20NFGwBcYxBYD9uV6Jf/Iy3oAWXaJw4eqph+mst9H+P3aJtuF
aozpt62AGSXBpLOCD2Y9/1FLPtrI5Y1nQ7FsDW0+6ke4JHdVj+xmTNHpPN2i5NgFIq8CzD2PDKMN
bmg4T1r0GUVOAyZgfjDyTskvTiWLil6ABcbpyTjdMH/X/drHK/GsfdZQ2fH3LjRvsfVMHnWxFRpR
HRIiAIeAYZ5EIFirei3IZyaJBES0lMUrhF5B88yRpW7mTkPBHsWPYyePwEcF5jcr3uD26fVlCNm5
Rtxi3HAXeUYnAR6PdY/Hdsqt9V4QP0VSpmB6t2cVPwz1nMCUzQhRIh9a6vsYmmWB/6TYfgjSVGCr
2kBsG3j9I8eWMoeBigQKjDW3N7dQ8rKLdo4uK3B29Bw5zaISESJpAuesAF/+cIgPJQti4ujGMkBd
04g0tnZD9fiSU8GpIIJxRLOO4xwTfAHIVK7rEsX6kx4nV5lbURNhEb6eDN5Ohh7CJo7PlqnFAh2s
BJu7xGJtPwQPCJYQKwvsQTGHOUnUD+3IllZSVcwKa6Rc7ErEMZc594xtt1RQG9sWmIkxsVdAoawx
1Xx8LbS9FDKChJSpoUwR2SvxfSPMW5ACmY6jRYkl7TPX1GkI3OMeRiIDdwYeXofJ5Wr4PMLkNf3R
M3Lyt/WURO1O+7K2Vk9ASZ71hZswLoN3o9wggKW3pF4ZrqkbikrAgXAhzkdEv1lRDq90c3Ep08Fm
SP+JSSqL90q+IzVuE3Ah6B5P3QVA7gAlR35DNiaahWz544+yEXdAbVRiGX6YFubVPuzHSD/lNC90
vDQI6453yU4eZ2J+n0H6fnYsj0bXsBT6f1OA2cl6kSmAqhEdLqD9B2FddCu2ZnvYtCoSIV6150Zl
2bsBQuGyvVdrDPEgu6keANzRKfcATjrld/ND+Hk8fHmJyBMZvnGX0yaEIF7HR/VadJXMTHV+oJvD
/67kHZtAH7wiNGyZuDsG4OVWuRXB8y6xe4qpPsbdGSkW0hxSPMFvR3/hwTnd+8OiKPwhACpjwC08
kGuzHei9NQtvNUNyaNhp4QYiXVeZiIFUYbrNtnEs6/3IJ2BynAQuOT1mt3/F2RhcQ4PAclUxDdcH
ZZQGZkIiy9VtoSKAeEjrFTWP6NNW+J8HZPwbutG/ztiobENgez6LEBeU4w5DvcPkRFI26RV8AxTe
tVD7c+qN+O0Hg3XL+vbJHv1VxT6UuDqiAsnHenxCyhP62B6/50aCnjNMCf48UPYSW5h0NHbv4VRK
OTChSXoc4l8r8WjpsI9/8GjWd/kors9+fOz+pf86ps3PiRaCpKZGTRCGLutNlTKrVPesNE1L9pJg
PGefY6zwoD3KYWr9B4pGMe1xLybZANCrPVz1pua5T8slBktScUdZsx05k0y0hTqhNq++U/ziHP3t
kPBZ+iSh4VxeXV+N56kIoOrJBECKfldlSdi2/grqE9alZX6IdQEDDx0Dx+b5hsdYXWzrzdJ0SgzM
bSX6AIQPy+wGmu9HPFUkc+KqzlCjJgb+FoajCN2ebOG2lES13PhoGOs9kq/MAHKuqu958yiljL6Q
R7bidd+1OKXHvRFmL62/+UFZkDT/5yKF7DpcBCFCxEMwpDfKkzty5FtHdq1hvT9t40lyokzY2RSZ
hHPufb4szekff1jBaplB6TduFXErIt6ZUsyRhUad+qizdSrGQsGwJJOUsbzsSXpGlFnpy19L/ZCR
3E5jQ/uYddCVIGhcZ08kOWb3iNNFivy7Hx/oluqs20beTLUulQe1VNJ4bOwmolKPzCsaL+Ap42fp
Z/PRhFsMvf21FcSRInPtZbaDXPL1/GOTwaUqKifQ4mKjsvU0NKosaq/HpNKH8F6MbKS6GfQ/osN9
THB+i7S5THTTZIb4x7sYsM+gWswskUlcskmyuF6JqZyGEd7hAkrGB8loSrvmd39mVBedl6hXAJd7
ZWtEBrfarj4SdRxUKeKs2u+dK2QFiAxFccIhIsY4sRqSDLCarLqck58n+ASipNDUVkqW79yJjSaj
7xhlwLF3o3iSwNiYM4TZvkdlKeA8Hd8AGhH6uRbLoGB8lm4f9uCyCDfGJw1T/SIuM2g0uyTNC41A
YM4zXOj6E5xIAoUV1qEBiGc5Ld/r5rvai/LnJUfK66MwHm5bPqB4TWVwINFrnR80bhpDO4/IaYcy
IHFQ8GFpCT9VjgIgLxzMu5BX5eYTKizdd0BfGq+t+6q/UfbHCaYiZRTaEmPF5W3pLJdGv7PGwV6Z
P35/7YKH45GDQ2BT6zhHth2+V2NST0P7uhaiinfF4OBpOfClFKDIwdeBcSkS34MQdAGZ+kCl0MRM
G5gVvnqMu0dpEhFuRFgJNT1VgElZ9l6mAaWelECZxJXinZvxTHwNvSrP9KtXg4FQNW3z96/zsru1
pe2RRWYxoDm8wlsd06E7oOpdVglApALcZqqNyRQowgovkhzny4cnQSRBDvE7hZ0H8DrDoEvHvT9w
5qA3qNSGa5W0z+D2Pc7Eo+H2UTcwdRJOsdvxP3+e4LrV4OCk+It4NazWpquOVUZwowZFQ+EbzeZ+
woBR5prARUrJ9YENVTEmpj+9Xzw+Vl/BCy/pJuWhRxDrZ7/y5rzkIdDX5rqDSjxJOgkcL0dOO5ai
XzC/JsUSDjd4pt6JXuwtjtWLFSiQao1ljUafs55wHYMdFs34aA+HdXDB0r+slpnJwyPXbVjuoyJ/
13eQQ4UGIKp2/P4AFA2PFR/KJi0rLNyPIdM9uX9zite7bGyaseyfwJkxjQ9bX/kyrSqJVVAEYtzn
ANVLC6eBq5bisoa3GgT295MrGd46TfDbEOTxBhH05GCnkt/WVKqOq2xy1i8bzJFBkXp58SdWlWvg
URdcMmUl4CE/RdeVJPeeFnYY1OWYXKvnkaAJpCSrB49gkKvh6tcrsOSwWwryWadEFWap8vLf1yjY
a1PxxicVVnOMluSSv/rLsHkXlYMAUvL/cjQQOic2Q6oE1MJ3QfOlyPT3/4Tn9JsHp3Ax870hfL/e
OJNb4yxrJ8HFejUuCkcndNVN3yH27Z9908W0X9KsNZZBGYPjTuufeto6nlAClOOdjD16AVvmHksA
2Ftve4zRjU77lWw/ouUcDNi3gEdI9YjqTVk0L2lSDIHgnIkVb5noh9+k1jyphhchNy66WSyzf9DQ
no2RKc+K7Ku8PJAWWXl3DrtCRgzBygBmAN+xmbRdSqZjOKWOxCQeO+WKsrrczLaWgn+GlHFUrDfR
2k1KOMGJIsmRnvs4XDUqWnVAlS2cPrzDTZRindCIW6o/pHTF71iOKKbGRjFINjeLLp4pS0DOEvUm
eZ/jK/sFIFWEBmTJaOD7lc7mNJhzNFFx4ImE7ACK+Skmy4DMrL4SlQ//2i6+lGdnuCyxd+BRmhQx
HgtFDDKuv2JwbL8jiSe3OT30MDqeFanWi18m5Y+mLXrXZ+z1CxbDQQ2UbaSqWUqE+I69XobWWbnb
SUIuACHW49raXD6qMKzi3LiZ4W+wZDe7kJlgI0Y5DavL1jyj0LORotDBBXo5q6VymZ4HR0A1iTTr
lTXZhWgfs1D6t/q2+4V2w3Dp4BUfdgHlPUfHtxYY3nAn2VQjjjoERKWS38HzHsYq8EGJpP4/Y+R6
WDWuwY2+tGOjLUqf5cFOeWNSFNHVO4N/z0QHAIyHl0HrAhbOwe9StI9nWD/oOjf7o4jkd3AFQE15
S+BBcy4NbvfuH/8RlzYuXNnDkjBXbN/lJh4V4GCzzfB62eDW6onUD7jojZ1fpL16tCH9wjRqQjaA
03nLYS2Iv2zUZ6CkpBqKyrU0s8WrPlzwlPjHs0U0zMzHFXPUcSU27+Xd9PBVUTtPcuNudbMvueJp
3jlsz1lOzSalJnqVC9HR0iP5hCefgtp8VDXWKwscy0JsZu0KV4iNTq+6yQNRT0FQ02PO9Y8KDi86
FlHyvx3YzC906Xts06QCi8tphZjQHnjUceN9sPCoo8aYT/n+DG+bb93WadyC7V47zsfxBGA1zt0N
+lvGuC2MvwLZSoLPPxigEqo6VFYlLtwL9WbEHu+UpKEIn0tS645n59MJl1ZmZGWWaMOkWKKT48eE
8wY22uLkzMV5TYneMLuOrNPSL8vIh34z7yXSqmXNgJFS9h428/KyqOFTnBlK1vIb5j6LUs5ybD7J
CgHKAWphuC2101pim93d4zL6F+Qpj8jTL0649YXfG/pC3M9GXLpYKE7eDS8d8+wjmBpqILo49qSm
8lP5HUii4P7CgWVbCIYIU4vw6J7JCqND2jaXqdRPUzxolvD3qFyagEem4zvXWfqlGQF+fDiM1yYc
kQbYz4BVnSedareNs9Qht2e4lv8hzVFx0QwWqVosRtoLh2AzVKkXR4GsFb7lCmqH+9LQCzPbinVZ
5xwoLDGxilrtzcYKiySJID4QxOQwO7j4ZsOkpyF7zwNThVPzTDOZ25xvOUegWMuCgT1umvzsq32q
6pS1YreGyXtzj4MVpBR0MOnYujDNM/Mrvp9ycAbFrmMB5tu+F5P6lsfoM0DZjZ2lrSYWqSKq7mic
bWn3o7CFs3THWmLG8PrIHwtkw6M5n8UHDqWP0mVK7N9XTRBM9wpqVV2+B8+JLew/cuzWsaoihnpJ
sx4L7/beSZIctuFYAgclnyoVbq7dkf8Ig2A3cs6RaktfFJ0Ffki0ZM/ywTO66JsxLC56gYVlutsM
BVtQ4vlLCYEutdbPVQfNW7jOXnJdBmuXMLQJAYcCX4XUuiqopSUWd4LVDS0j5RSjwr3LiW5y2Lo9
dMoMicDTlBdaC/9XnU5NheAMeIj3A4q5WIEOk9EQmQ4LIf+1/Qy2LP0FT0pHjMcUtTA02aRhspND
59TygQpF62ogZVeM/RTSRbhUzK96t+kREVht2FaDFXERZ2P8LAsGp1L0A455Fvj457gqKE5dZh86
QTpEUUaSo1DQLUXKKakGtzMwEoQcGdEimtFizYNhM/3uYyLsD5kPI7mtrMjVdC8bnXvFbQXGC/5l
1HTNcvpdvjqIat+urxx/33bBI8VoLhl98gr01mP8T9Tqe9NpP1usTyb6KV+Xz7bmHlcZTbFkS+oI
WzlYSqiMqej5IXOFCniN/ELigU4CyiRog4SHNr9d2W7lFjS/QZj8PUGvlaR3nVLJO1+lczDKFDU9
a4+G1S9rbA9bA4lI/ydKUPzYygJnTPMZRukqiZ6pVH7N24sk5qE+mzMpaTCnMWJdC+tFn4fC9/Lx
3GF4FflGJOxcZBL3q/zKbuihvHYEkQhZfi3D57CoLhftJ0y95svraBXF3z5JChYUHxoM8MQ2AvMz
zuKmLdWUp3muKHQe6gC9susIpp5ME4CTEb4e4Azzos3+BnL3TOl5H2bbAyxuHiQ0vhOqIjADMvzT
IG07aJ/Zo1xjV1BBKSUUuC+6Q5mi4CSmvVvRvB2l05eEOOou9z7VipGr795E+LfzkNEim0gVj6TZ
WY4hTQlPzNXOwq75rBl4lzD9zeoTmslKdaoIr41eoe1h7nI3FYzRzYEu+Z/Us/OgNUoglVbD6vhG
RRsMQyoAdRB6zBbp8a48hUYcM7WmccQ8KEln2ZbJ761fHYH1LOgUrc5vzg8T2oXUR/4xUFisYRCj
D93RNb+oNlU+sFK40CBhrB/PJ8sIwdCTZrFiGgrk3sR0sOEOS0fNprKwu/IcXdzjbIIx9y5QWQKy
A3dpvZXuolVJo2d1A5Lg68mso6fPE8y8SXHnLjxLYsUpdq6Jv0jTbStA+QUpVg2PX2q7MgN9vNBQ
XZTfzqFVFBEJb2YQkCFAAzZsOaRWNNkTuvpJsSCJlBPCNWqLtSdpCSYi5queOLp9odFFUIjKfmbI
pTzXiaCNmBMm1gSSw0yFmuc323+cbBMTy6HpU+bJhHtXRD36n0kbLM5/ZLQEhtJpmX+mh2/2DH16
Qp+USDAf3z35Tf8GFzvnREeoMItGxVIF+zIc0ovsPOgXtwAUcUacJl811Ga3wFLxS5gAjTggOEfM
Rg8yeGZzvBWPklPRsny9Ke443iNejmrsvqVcpwkM2Dv1eIdG3UaTDJ2+sLlCkoOBIBQ5yeYyooqt
1zpT2FIJWm3FGuvE4+52sehldoMlTTA118WrHITA9QudgB90qcX517Y5qF3o1rbQdZSPcnka3dUp
DJ4t1KWNwbq1hdnDn4z+jHhI8RoJuTqLGbSOKhYJLfTE+9/QmmvdiFZxwpdy9J3TayBQI/qXVrdk
R2IOcyQKsf3FZoVxSo7n/4+E55YTqySafdjSohYSeTIKl+TRdNonlBYR2veB8Q9n4wEnJt6tQlyh
o/F1BhKwiSCXMMCEobthD5L55VsGCesLJBaduV4SG3Po5AhncJCbC/kH/wCutp3Ss474AbWTCjov
XCPu6dRK6MKdM9dmkxfDXMRBpmRJDtNKFu1L/h9/YcNQcZUxlMwFyuBhxZyvUSAvS+g1SvvAmfx0
uJyBc+OC0QDJnj6pCV7/SFBuycdkoLJNFAuJRIFlPu+abOm/GFAy2BzyyGjqKZFUKGexCkdSNYxg
8Mnr+5k1M375mnL/mOG2RTawlqNcPmXbhl2p5UozjDqxe/mbamQkk0NNtVv35j8VNFnsBafykCtp
6IpyjcXwmLwdPrt9dqZgcJZLEUYQiGqeJnHv8WPYmP3x3OE2A+iE1O49jXmFb84plMootyjxyrcS
C2K49WGxyx+f5i6aJNUUp5zN3V6MomnRLVXN/4/BINlexGcttzU3KOodRh5Q1fhS3KvS6h1Yr7NG
xuQY5ftj7bQHNXVzziO/zcGmYL9GVcZ3Y1tdRLGCEPngZQwot+G2cPUOB8iAQXcofwFCeDJfkWLl
91mHasbw2FQVee1XBOVyR94w13GzvI4jMu9OiXoP3rpzANjxC+BB4aEDTF9zEXU89NjzSKQpS5+I
K5lZP5s8IhPCocAntPKK9zjKNeBci/VtMGL0yoF4hBQNLwvBBjUBhJ3BkGyID/mCAgJhBjsWhU99
fw7NYbK566unFCXAIWrjGcM14lNy0OmnBrWZLnHLYX2LgKS+8GmNV7RnriVp55Msm7C8UNpxlKXF
NERcLtCnVp/HioRg8NYkScu2+nAZadDaYryuSbddLcR7lmwc4d/04aKqnxlGgO9NwO0lUqKxUIhm
uoA44pLMKWA5bksaezAw/QdesVRpMiWh4t2M+mFlWK0LqCi0cFLPrBPY00vITzc11vmUkeL9Txh7
VoAesZ5p5PxNjay3T5+G8pc/CBRmsi2c7bqG5RkVMbeTNlZY/ILC+tBIw+rLLYaeBO9LyobaUiAq
rez3Ho5oZBPrwuRwXh0ePgBEK2Em8NmBjKgEjD1m2nKAoY9N8Rvj6FQLx0oKo1UaoxqrKaujAiDO
E+TanHxiluu6Vos9FcXkoMGAr6xNrBdp/fpg+EoTA9pKNn2uuyDsN6lkt4s0WGLdgiUBMPF+wBTO
mEYDhbJ/7o8zFQT6jGKRCOvkmL6NgSLsT9eDuq/3g+t7tM6a2TY0J8zvVViAenZqL0Lr8xy4Vqf1
YU5Nh+1wUq5ia93KsabyAswPStJvZrCJawv+GgER/l60TOJI4GhOvTs0C7Nqb5YCupIzhDb3HZoI
YhUMnxapsqGMdffYiKur0p/2cpf/b1uChG7gJ+TTq5Uas1B+SJjQhytz/OKL1XIVPMeJ+pZss7pa
+6fTV8MBAOctkyp0TG/P4YU+tYdpAn+BZDImUA0MaAzjCIPaazFuyxNPRU/Ea5fuw3EEsowJs9qO
9WT2hKyEjqqJqzyWDrYRxG3hJldaeVcPrESr2YmQJXo9YN+anPHW5SnzstDz6B7bG1LRaie0RR9P
l1445ZHTnNqqkjqz1j7U5KE7CDk4nOKxIPFO1clQ8H9bnc3XCQk7SXrsEFizVKVq/K0MVY9kUc3y
jv60VCXb9tdPVUzd+Z2RpjaUb4Ua4Dv6NRB7Op0Py7/oN957xSJAQ9WeBqhILk4fL2KdeA26E64p
IVTPwXoMCT3XBAPP8QKYnvS5Blg2rKLKahnLz872uSrv+EELv3/lwdnsd+BHBmfaYRfeML2POONX
3GpjEABZFFjmrR6Ek6lKVYGSXV7jQ/9Ti6kYxhuD+Fn4z6huTRNIuaCm2/hrX9ERHdrGl8VdwBkY
G5iqEbfQIJnXK5TqnkkQpqCmo2BEYG/VkMlEa+KDX853AcDcuUVfO7GD7sNH7/eyq/ZR6ou6z6ZF
tA/bnaGZNllNZSWgGSzpIRRmguX1nHAlRfq5CiFZNgDIdYNJ/+QD7x0gSfpcP7yuFtgv6COVh5Cq
8pFgBuR6triurdP5WO5SWA+Lu5m74mPi4rQ6bu9DB+9gSpbkMJKS7iU6Ua9BhD5kjNC/nl06e+8c
MWJZzNhrcwHgQu+tJXNt1rsJSBpAnnYwa3yN+R3RDVlLOxXd7YxHV0iw7cX62b3L/+DQ5mG5g9ap
5JoiIjDKzv6q2v3lW9zGsfQvdrakbliMtbrUYSMGwnQid2JZm5Weqvr6qfdNwL3TLQRF+MUx0coA
XNzjnOBzE+kp89nYWXh5dY4eeSJYinvylVCzPFhZnfnpGXyftHWEJdPD/LFk1z9d0nKJewzSFgsK
G3snbgTWxM5tixgjcwrYpqwXFq4zYsguuowQYtLa2uCCbXFdFevE9+lecL7jQd1RKV9CVA9AovF6
pp493XIjZn3zy9X9Tmg7i7yEayn5jH2XDmhn34YEVV5dc7zob0om7c39haxPQ6KzrEut59Hs+eUS
7RulrVPy7S36e1G+OgbthS3mhiVTTrBv16G0adsGknB68jHuq2YakmE9EUIzmYwd1ddP2kjwUNIq
Fdeh5MRZ7AnTBMba8duAhBTMsUrU8X5EK+UTnclimRjrIOj0wJEbLnh5/9UCiDoL3abHvNhycnRi
mw5qapPJ9WrBhiNyO0pcZuHJ7sAC4DT+zO50DgwhSxJuJd0hLV5OWPwjRQAeJVDzJ/Faz7pRlJMY
Q2q2VttxNZzHh6qHFy75uKqUJ4DHGrgmrupBCgVuYfMjGIojmvs6Zf1VB8vL8DVwLe/tc1hwGkMu
lIP60Yz65bH6Hu+3+gNaL1ZL8wCYLcgucXm7blMJw//AJ+VcHh6LJjjansrcP71DZ+s8/3FgV9Pr
l14wOpsVT6aITbf0jVd9LQCHxyHUpwi53vB2HMkohurlOMgmz2gDNfBJ96zF6Vw+NIFszS8xeEAU
wSA3zmX8D2pls84HTK68j7PdmNmGL2v/uqKXKKydBUOzSGZGWnNr5FkHQaSYiqFc1CIW9kn+XBCP
/VQVgipcRwTF8ujbCRQDzZSd4DSyAsJwozUoMr/fVjmy7EVzFkh8p5dQpcIKbI/yMBAZY49KlAOp
xPYukVM5TyzZVGi7OrGBJYdFv591qdjAXu76r0tVA5FWlC7Nm8mWoZf1HnBSTGIzyrFVm34yo6WH
zivf1u74zq2fLGMkfGMhUn2dnJ1TjNhyXCmN7OcNtMiZDVbfKbAdAE5dGn74rlIXaDRu/iJ6o1dv
9ev2Se6ZOc2X1JpPxbK9RL0itmIm/M9F2IfZyOohhxCRb9ItkXGigfm8eWqxEQRXvtRae26EyVBU
Y8RreeJUmwrzeLtoSH2sQQFcdiWGnNmeFlx/MHi42L1LFIUIjFOe/PUqFrpB7hpuPN8EN1I1S+B9
oSCWY3yVfdhvMzTZjd6gPzwZyjptf6d0Pae/j11WE3+P6lDtJHEOFgmHrpfIbRkyMwO6hkuEjMoh
F7y/AAY/PBuTQNYu2YZlUV0L0gtHFqpnp7KCOZIpPI7GmJOvnnpK76SVlzFGO9ra8BqzcMcNTM+V
Kg/QC5vXcQP+/oZkl6/sVjvp0BcB3deKcT0y0GJ2dGEsSljwCX87yzzVp999yjm8cvmj/Qg7/1z4
EBInyJjndU/YrAHejDeW5sf7iVOzDgoLWp4XK35w7boZmo6nYNIo5eLFUjwRHPyDGdhKN894xagq
wRkMZqOG4EPtG9reOEXMKWbPQef1uzaNap6fK1T9qBhfgmEKEOCSIL7dcqfGc2HL07TmGDfQKcMw
+mPbLyIGC5xvwyi8GEr8HD0L2hiU3bgtbReftfSZfV6ghdyZ7ZEYBJbVgykNU2gKdE2umSZOffDk
IbBOx5ANAGUv5+876BIVhdqPG+S7/1GN1W6zucIpqsHijYYLtra5M+u78uInjFfmeI63t7BU1rAB
AAlcq+smTBJE13kbtln1y8la082NzzwfKquTCWk7QUmrj6ARAESZjjPtzUvt/W7L8gl0APyea8Pj
v1giGDB6tEnR1fDMdJZDfGyspByfhVAeE2eX6V90nJbQYadM9dh8qtRPhjo7fwNCplwMPkLojdwC
VYPlq3+mJ3GM7qjUosW5vqfy1AMLttei0fDgMG+sUH5UbR37MWByNu3gQKryuDV4Yr+KSMN8qLIz
YzqKDHvDNFm6Pa3BH4K93ON5OqbyPg9+KXgOsg2VdDhkFw/3LbYLHFF9JHqfeOViu0KUJRR1xUxk
bm+zlaxK2ehvrmGMnon1gSv+Nnpt+grWprH3fAMcrK8N9H4BH4IA7J990mokZzpMCc1EtznyOdgg
/TnpuFCf0WutmJ5lPq1J1knfxvf+6pOkv2K/wENKT8WTeDVLcSjcEgwN9tAPsTMXUoTae05Br2Uj
mMpGoXh7h42Dus9fi7c9zOVGkLAM4cuH/+2nRxgGavGbNCC4fJ1KLciSzaHOHqpAOyFh9VRAUogn
Ay+HADMwyTVqm0freb7k0krZPVF9knWDj1Jraj3EClyn9xeo1ni3NteWbgZvAWPZOFL0Tp7aLa+m
FwiLXsAchoZ72MoPa3Mcsh7/TyJtgIVHnyyywXd/Ujdt868vfvrD3Zz5MjcLupLbbNc1JMin945z
kq9ZpLT1q+33VAR48I1UL8ePJKul59MxQ1LQkcJ2Jrm6Yi4XIv9rQGAtm4szD+zoCBjbFNBDOfWm
6krRVq9+ETKx1nPav3aNrCNqMZ0dTG/77Ov11KbwjvDOAZW8jnl9skhcdqu33ldOmOCmjOxs0PYy
82h//LwbwXeN2nWNzhMdVAsru+qGkpT+jOAFhfw0gSBC0cGNyWZaDDAoEEQETYRQkVjGGrZaVw57
O0Cuu0ntPo097N/IIiN/E1+g7Ye5Gpu+6HSpT3vj8SJMrNaaLjtdx9EHtsT7xBahh6Jl0cHPr1P6
Mnr3vJ8rZ7ooUGIPemB7u9HqhH8pZ6jW0TFeBd4tMxsS7EzjV8bM0h2NKkioBZnGxkPEuLSoOVSF
gOF4bzK6fszzDzzNgqghin5CZs/Uls76xeo7Eztv3Z8eZ6wbTONgOCkqel9fTtHj+xi4etHSEMIf
P10/bXhGBV6fS1+/uPIecn3+c5usYZC2RVuXMoH3GjTMgCty647cBjXsZfn1c17dlnEmbJoWLcJ9
YElE7Ywr+cJyXgUnwcAkEK/I/xN5m9SVcxcVnhLTrLzjHWpljt3v+LsQ8t3N4vXnMdzT8IW1eH1/
fli7b/eAC6kq8W9ymOOrIywukXeSa6iK8gxdXe2gI6WsoutdbNTjN2d8GIip6WiiLbEySbNk9bx1
eIhSushAHNgBzj+2cTvoKadfL4uIceoMcgSnwawOSfxlt2+2fkHYbgmFeiM4X2tof35bEj5YTaYc
LnkrTudHGkAL25JC2A+nP0KAa6xex5vDfqbEwxf8QhBMKaCgUZr/yQxH/59Dfh9makasvBz53cpq
xTNRUZxgBeNswMhFIfFE407dxwGyPm7U/jKu8ItetByrugbfKQUGsxhqdt5fgNg1rR3n7DA2CHht
rFpWcjneOR/+Kqc/wjZkaQk5kJRz4Hx3NyUD+0bEMPKyD3ca4JXFn7wt6v6vtYY1UrSZsZr/8g0g
9N8IS0/C+5iiZcLFPORaw4/GAcFodu4CWoB+ZmSnEriIFKigzNpofvi/TV+rRcPnIt93CLG/hRXO
TNVTM1GD3bVU+/GiTAYv+WNpG5EWmnE1nC4N4x56LuIY/3JCVxh+emqxQn27PBe+qw7mFZSFGByJ
XrdMOElnSnxEbsDUykY9SHK3mB9BUqGwlPFY86PXnawJV/NA8jn5/kL/spS4hU8WwPIwyy1T32qA
a+egy1EUZQxwZNLNZkog7298Fj5eJzBJ0vaDtlunQmyLJo2Zm26NiZTmbjw6gbL3iaUNY4Q7aen5
Fr1w2LSOatGU1Z677bFN2AQ9hPPvlfnZVHqjNpvkQuT0vyzbob0CjHk076Q3HntQ/FUd4IeWXZdZ
r2HkX92WLMA3ysMs+WrPS5vMx81XCdpObqx+3Hc0+1swkk8sCr+aSqM7onPaOTmRDlI69lWLtC26
PFILOFkTmwAJA+Vn7616zjaL/oEdmL4rC5UYmPPqdG69298eOSzr9A/cuSka9DvGf4FwxmEzbRH2
as/RnsDcw8tHIDpa0CjCLncqulvRB/kM1qRuE8ObnmVqnJ9Jmsd5wTNPiClzlbVwCyz18bLOL4Bj
bH90T3AGSAp43orhYMdTHVnevcZ/kBuP2cbJnZlU5oVvHqCR1pxU1k/pJPBB6FKjuxlxdLTG9T6m
fkK+zOOBj40IxodRG+/1Sz6ZDtF2SSN1tb/qx91rvwkZmij2YxqPJGT50adRnXzPjCrGJxD10I/A
Z94qlO8G6g7O/E4oLreTYnzhNKTt+ATYt7lwS57oHj9+EmkkcS5eDOIszi//Xq5EExMv33uwuUXj
askB3ClHeOayDZGnQKcyvgMVyl2x40QqbRMIVKnkYiADKYCAVVKtCdREYzu7Z+k5KXr7mgB5DMkb
09ey6FvII7bV6ZtSfVZJI/rkf/POnPF5mDB4wUFhWj06PbR+tugYnGXgddyJsnDX8BaEH3oQBjb2
NjEpkb2dqj/19BsPQOcUiysLQ8FOCfCl3v/B6dz+9k6lo+N94MSM3bOOpQNvK8U7qJUH+IoLcJPC
jH4FEzWm7DdDgyURFwrNq4MnL5qhs2JXNwDkepCM+7T1VVaI0c6reYTA+d66OYtDprZ5pzUlDL6d
4QuyUe0AoDJX6fSvl3Vrp/kDqzxOjlf8WZiNqJSsvSUE1yekNFPYGJWPb/kIgN2Pt4555sCeY77D
pa1ZHP7RMCPam6NuT72QY+HwtPkQPjJiNnl0qhAaxN9srAr3IwmKRLRFr4mYFva46+aH2nl6pJN+
RHmOzk11iaU4HcNwMzkUmItNc6CTdC/Y5XPek3OoHXwfVHfJWu84ZXgEMN1rRC0lJtVRh/ZKLYYs
Us8gaqHcvv9+aNVHMgtmI3mOq4oaQwW9qG5A33Ga/tC/iR6lyKAuF69wjKoA3NeE2hCq1af7POZu
I8vqySIO85KLxr3B3AZP9UN0nQKCZlCJtP+dhMuy2itUh1qUm28Aw30M+OGcBFFkr+JDmGVAlkNs
ATzvQ04OCxf2Xr9kpNnjZ8FFTMVuB+BjEPP8jp4ow5CKtZP2DY7YEsZ6rEUhmsq+utcXyyfPvkrM
8HjoB1+qOTfWboDVJAmc+g7mjO5ojnAtjn2/s/oae5VHZednBvuJAr2rdUBm89q8gUgt4BKHljCq
tdvy/oJE5nAk5zGEeCTVQfNUHSiqC73JdlX0VbmXU7mAOVAde1kWmtPOOyPXSNpSmJS3cNPMTFQn
ndlrnTZzjGq9U6l6RCBTDnjOAQrOamjjCjYvdcfp43Sg2IfovV0DHqoqJ1CmsgkFGAFyykHl8h0G
7gxJf9twQhWPOaBPq2gb4qMjL+okG75OD5UpraD9kCJko94Bniq2Ko5sxbfO6Y2I8CdP2rFkWmUQ
HehVUn6dPIp2/qqcrpK2we1kakvq3q3RRettCJWtEX8ls2DKt1fS36rEi6c5lEF/38+3heCMo8uZ
OSz9lSErjyUBPQ3OhKr1CszGt061qQ2XwiP8V/KJr2k46Eya5pc3gc22hGx2GJ2MkmoWRA7UjSFo
poVw4iDyTItvsfUQpzYjwqtLLsZ8yCLB6wEFruja0mAcUrPLvEwyEukdq/jCVWj+yONYrdyNgXC0
1jnFORavjxnnMw9/b4b8pk6njF9OQZgUpNIJjbdHyzLKqI5bOqdUMogYIptcSgHYJYe9p/RVtdqt
Oo9z1vd2JjhR3EGwAwkIEM95LQghVA3Isn+PWWzph1us9+LgBcvDM6LyRcnDnY49azYgqDBtCABA
TTZXjG5d259nPQTm4fRzOIaaUA8luJyz33lhl5V/xveNbQfj9PjKDK9U2gWnDkDqe3uXUnPt58aq
NXA0qGWqcQgmrKxKHgDS93gcCLjf1/OPkZve/OzTFUQEfu/TxRDLz5aBPR5Dz9Afp6LaLksh6T3s
8RYnnFVJSTVYIHJEKP0GczLN5mt3ggz9CLkzjZn+4EEohpjWGz+4s7Go+q15dbFUoNRypRIkCAO1
Ysl2oYY5oXLN5RPQPM5shV492UPJqWBWeuUmjDaZbiw+v677nMuYmj4b3pgCmBp1mI2Vgx4N1XmC
AlvKFOZH92NF2P1nWNhlAHvmiSVIGryCdrFovmcvV422suI6KkuIPd57PhU9jFrg7KdUQ8P6p1NL
g6v9bLTFgMiEAAwteRMJpE8mzJWs2NpbRtmqyjL1JqNXgXFGyAUXgmp1/J80wdbwtnsGnduBDTEm
a2Q5vz+SR0cMdKFa3JDphmqd5KOKOMwgpTpEkabVUg3e/Z/2SS35YTZ9tyw5Yew0c8TwrZD6s9h0
xIngYw4fLXCPW7jTMGkBl8CEayO3y066L8Tm3UNsSEj5jAi6hIL8Zi+T7ji6er5e5Ev20hy8cxYT
92DPfPD69kYaVia20ojWJyf59dIVs59KI+nIsyGtLEmcmD7GAJla1UUTjTmp5Wap2s96x4RpcW4q
O0Hb6AO6hVjZWS9bSmjSMKBWbX75M60coVZWh6AZmFa7yZ42CurRU+BUOwUyukykls5KVIjLzwad
iz5SubnEviXBALApTpSIuXmxDP2rGgf6/xWSQ7DhrxV6dZOnYMIr2H3puu2XlNjCexKeMEkO6K72
aRyWRvsrHBT9loKVHDEwyGy4X3CbZisN85HUFppe32a1rgOR7pBZQ2acFb9LixDUmkYd+atvNJWE
sahhquvTMF57gXHTFsCCcgdZSFD0kM/fBE0WjEwnV3t/eH6O0rgy5X2QYeB7yQfjXF4s9OVEQkQF
GGausTXB84Z4pCfWqJhFm5bB+ZRTomLvN7FkYxXxWctu+3qy9R05f7xFpdF5fd/W3yUY0SQ54SmM
QPllJbGe2Wo2ZtDBXkT+Pz8zDJIRp0kuGUZSMLqEX03RCS4mjoLS8J5Pw5M3FIEM9RiE2vyNhv65
hOozc96ol4R71WNXNn7xByeXmGiQWfekJn+xruatAjQdWh2U3UJVMlFcq+uMpgH+9tkGiWM5lcGy
tgBIZhu9RdmndOw+JTXLv+cG9umNyl5lbeEvQKRaxbL/VNQ8gA+FwQ9Hj5TQ7I0m8RLpVftQTQdB
q6YDw5hFXQqt+L5Xclp/WLSjsJ/h/BL1v1fbVSsuD4NVCNaeTsxQPEwg3VFX3bpNB9PXpZWCZsvU
M39hzBQoOo0SNssEie6DoHWKfLbYbBXhonVKLDua3l66Ca6Evj8/5RicUaKrjGwHQODwLa789+yi
Yd4kO5GDDYzA5+6lPRgghjZW2YtkBKer4RU+ibv5N2tzR4d6cpE5NRL1c4D8S1PosXoCkmo570fG
g0NxrKy86Hp4QS70ZeacN8SgDNAIo1ZWQA6LL7OOQHBBACgg1B/wivEHIPJmSDuRjZIZpusGzPf9
PsOcJRSEvREvJBOX6mGhwU7MhcBV5G+D5gNXXcwN1UgIeqfjCu36r2B6TLTyl3fdQDiUT9Gt98TF
vDC/YPpHl7rcVXEX6KwhrIvGup1gFWLDfejZmDtMgcLfiUs199JYL8RuCWmQGyIVNlLLxn/odhL+
107BwmIAUl6xvH7yiaeFffS8jXNBrjVE29fYAgkv9CAXrEo/tkM6Yh+2GY7l1RszfWp6ErCKhp/t
iKbyRwBt9IObK9FRv5HNJxcZrPPH/fXzN7Mka8VG9WaONFpXzC5i67tPMvwwRuSvmORTPxs1hOZf
QUZz7FGJkuKeSvwo9fyF9/lFb+2FzQF+HmOFzMfNrtdMWs+kitLR69LNb5pe/PWtyDWhYOHvJH30
xK9Dy3/sDkj5XwP3wYc8m5IsxJdrgmBHy6Hv7vuFFdqYrm8t281eTAJ4+p8970ov9NOBT0MUrmuk
dW0qbN8Lgw9R4HwBbr3yl8ma1wHZzK4MJHL0hs84KMNS9EGzDid1Tb4wTlpN0D1XWemj1xzJDkIp
uIGcT44OpWlC1WqvNplAe2ClHtR32WucvGjZfGM8CZel1aKtpREkxSHrtwTyEox7jzELfqRQxkB/
eSJqD4tKffgoyQlU/UsjfUwtrVU685JhB/uqzHc/c7ZA0Knb5nKdqUQ9t2mlY4k1AopgIQhHtYPf
fjsvpRRL5+rzMojz4Wsl6nhWyQFPRTT1Sb/dbmQzaROLPORYBWaX/Ix6JrEqoTx8lmsgKivkrLYY
/3n9cJFbYZ2E2UPffI8sk8ZALsy3njU+4SnfR9CQzysXWdwCo156hLSB2R236bMoGXpVu+9H6mmw
nBy5WVRE+Jzj7ViVLIdIFj0XlAThqGqluutnOiAipJpDqzP2mfwMBSDMEDHw1cVgd8+QnhP3aIHp
t0VIQo6/EdLp2xKkVHEqHtIY+nOhaWpIvDz8pRNhUheCiTMP+pBrmSzR1k51uK1Xk9btXGUWs6wt
K3L6I5GpGZoLblmofG+T53lneFwzzG0NyrgRzJHYRyp3hyomdQNf8COURMHY8yyc93YmTnaYUbDi
1ghGCqJK9yOpy7pmOv4dKVp+kProb7H92xb/x0nlS9TtUcDo4csvVE3OpE42Qg6Y7B1/gseq2k4b
v/Mtk4z7zaZI7qNmGyVfTYBncMyF5vdrlnbxOlEZjtHPsi0MZ7dkSpOrs/+sIJ4ho/QrV4t/KYy7
p7QT6MlT1lnuJ9IukJUBnjvd1OoRT1XFMgCPZXvT22pbgcczdOw5y6MG6MeBfR2SyO5CDX57Vz4M
SSBVzAwO8aJK9nGH62QKR5gnm+sCmzfndxKO+pQI7dxP0vkxilofMae/LgPNw/uVNLGFbXIOCeYa
RXmSYpM8FeysAXifQ/cfBFNmw57I5xpVXMoonttXeGVkFW+IBE6SDN6aahczuysQTn0ume1DukrA
BwfD4ckJTPCRTkWW4m8zZzGJe8k9Qa64qLsz8UfT5bdCNW1T8Ps63YIPSCQ07BIBDgzRVivClzmW
4+Wo1IriZ1qqmlbP1VLEfDXgHi/7Nz3L2p1+3kpXNKbEFu2lpKOeIyr+Gt59QKPwr6ORrq+TiEz8
btSn/I9x8SySl2LjHdcVu3JjLMUmxujTJNm9LlDI0ek8PdLR6lSabH4w+VvmlFYggQKJ0Fd6dJHp
S3sf3oIdETbEmfsZMjxFZ6cG1DLsUFxYfjphqWO0+0t0KAHCc2XHya4JbbgKwK6g0f8q6mryY6Fa
LwyeXWzrahfSP4tjIgrVP10Ee3v2GZ9a473QtWsDZWrlDpXLP9rZrgYlLt6obtetpbmD+nXTBYBP
SaP48uau4MKOuE+QXlTnUacPPZVNK9ULSBzJoQZhbmFBRjEh/zniLHX48A3qTt2+yEJPnts993Y/
D/r4bteAncjMCp/e+B0keNuj/Xx+xOIFMiYPwsSkISAMEOrD5RKCtiznQs+dO2LWrhXhrtIQfDbi
O/Reda16jRrYTtiChwU6AyVaomJS1Fw9lVhFfSj4XqHyD1sDuIZiDNdE/AaweoxyTMXmeP2Fg7KQ
lJUEyBAs6zMIEROMerrH5QrFM43S4gMDBxF/rQ5e0LajwIcX1Q0byeSf8IaIFnGThRo/U+RSlRLf
GR+fZU4wNT2prSDj5JYI4YLk1Gm3M9Mm0nSvbS9bQdAz6Ki8qcutJlei9KHDRNmsbiDqIpbE5x9R
vr2jpjKpjO0tut7FFSXbOwOCP40IWwsg0MxnJRJ2w02w2l+tG1QlMGiR0RS1VKFZj4b78NKOvTmG
22yLvEs4cfxoi9q46X0kiTN73m2DS19u/y2+25Ou6rVoJuXXTwXsxU9bIwQwRn0HJieB+EPt1hVL
3zACOQTMK9AJ5KP6+/7PH1ZhsGiXgF/JmsCNo8AjnmjewSEJ2UWk7/O4798H1INQdZ9oeOrdNph4
aCnoe97aoe9HNeJ2GypPEYH5OoPeGJ5yot+9kqpeeKBDNyd69+2va9i9Fo2VAsQssu+DH/QWZPbQ
T6gZ/rUvGq2Ulj1aDQQqI2nCVvulGZatm6Mxen/QEsxcMeQvGuC2RKrlg1IdhqUWtrFxeBl1BWpd
VWsTNAt1jtg6JeyjuavB/dm8IqoDGz1gDl6J15GskaA8JrogT5cm+H7U2txzfxIBbk04yzLpssv4
0svWPdV9ZykiYVP+zalsIokzeu2kly/ZcoMRX/mcFNUt7quzVjiczuZ7pyyK6ggba2Py6IbJ+mCR
9MYeoZER3zq9dnu5DMRjokkY8wy1VSK6xWyz32aFNPKMrZ//afDGFc+iQhjHmjpI26J2WnJuWODY
kG9AdXnUjdKKu+4+5MUKEejw85Qhortv0a6WfkNdjUmpqgMywNYTK7+Oj/6deRuDxHUoqYCDSx0C
2dXBeZ85ypt5ebgn6Ekk5K6n3Wrb9YbIS0YdIO9pnnMHzk9qmCROIWCFb//jWbFZ7lLXBEKKoQJk
4FiZPt2yf92IaBov4zZgqonT8qHpG92+3KX5SzXm5Njm4nPwWK0m3NoMzV2HFkFFbmJBlMYp324C
W3TAcZ3yxyg26ohVwrKst1UTrt8+DePb+6jOUrXiSJB9PvirJpLbu8FNRwhIv06l3TLX6zW31V7U
5FunhVynGSt146yTFXODYzm+8aXvaJ2WiYi+X9jG68gwFHhGe+/VhuKVZCmINZrycjax6OwTvkuN
3x4kNx0zcM/6JWi+iNZ+7KKgBYWaFarJ8gBogx9GiGJ5b2VFDHKYFRZQeIJIexQYRoai3vfbi+/p
9/JyAOoUUp3ykCWOUnPPAVihG9RYZMtA3XNydTsVVdvQhUOxu9aMLSJQdwwCQdw0B00Tqj1CiUzq
u09v2O5E6zRV7QEhCaN7VbL8UfvwHxb4hbm1UJYkYTyw8c2wIS7KXASpvgUqRHotU+1u3CgMh50p
4TrjPFCGrgCtNAYyShJ3DEsYaJaiPD8DVayyLkTYvlzHAhvWoQaIsZ5zdGDlONIbRrBeB0M8O+VC
+QN50a+gpTjaShCSnqfKciF1QlgUrH5Dmo0M2o8CNTtqmYELZDwGh7Km2g8ey6EtHTdV/SecdC5Q
Q1mMsy3T8KasPKJbhK8zXyxIChLp+P0VNmECW92C3XV9lijS4W/q7kLbSieNgBT3AT1FAPtQAfKt
7AW+pWC9q/o/xHxPuYhP3aBVS1a9kA/vWUanAYJzrtnlQsj9sB15NoBNeYqPjG2krjVoU2mpfsem
SUeA8hxqVLUVL8gTovJuACp1ECgu51Cs95FJnJ67cPa0s5Q7LeZcs123fu0tuFVA0AeoXnEcq/Vm
7yAZkCcrXG6KsDXsfht6WKT16J2AtPuymHjr+ezSJ/Rv7vRzAUh1xyNazOuamtVfyuZjcOnv0h2D
NVEuaA5rgWkW78qY30cce8sbjaWDdaLhX8sELslgIQHmfLDSOKW9JzgnrtFXoyoAGGEbWYauCxaY
7hacDd3EwJBXL7nn1udN+VxIS7sLRWh0gcQJ5O3fcBfi4wG1rcaUMEgXDZdgHRSzF6AkMImh52QQ
VRMbkhq9nJWaHvudcc8dxaDx4aAHJwmJggRIZJeAi/CLEV3OaxCN1aMNhaLEGpQI2GlpC5tHCvHJ
/zjw+P7+1hCZd+T5K1PUgmzAFNmcF1u3cQFAf77w1daxh5QMOOB1FEI9LgZhlV5Iq+esHw5b84FZ
6B1veXk2TQAZd8hDfZY3BCgO9k2ZR8ECKhYFV7m7BIbwi/OJ5camaOhgS8f3zTy0EtSv0fFgGD9I
P35Ylk+M9U0FjWbpm1MteQB1wCdYLKM2l1HpEr8ZtziQf2cUf2WFfdkZ27nk4pLFkEKKOEsxc8UL
MXo0bwXOoXT9QwnAqdKpU7Vbk7b0Hp0+kJhjjKGMMbcSCg6QWYC7vwfmzBf+j+4bk//nwY+NM7TL
y9VkjwJlleAt6/cjzGnwcRPqVlXo6mLVsGAsLWsxSSZjdD5bWYLdr0Lq3+6UD1otn7t7fv+QbGLh
z+H4obpqywfgCOpjT7FKi0FxOfVRCoi1Nz8fmBZyLuwhQfw0iImxxMtUGxOPUYUPKCCpENO8Tzi5
TniJWjKbozA4KpUIv79yQYKoCrCyz1iDX73U6PYZ7Npl1EaEzP8DQFlZCtwQOAW2R7NWWQTPOJhk
R2D4jmbEJ9m/a6R3mGNxxpfOFmtD/vxKMHHWUO1piZHNJUyOlbw0S0ZZa1nGTqj1zp/S+iKVzCJa
jGjUJzFimXbPNkNQ4TTFW8N3Cqyr489ASZzukTh0udtNFPLMZEKaoBDqvabgwbII8z3Ue2l/43qJ
QJx50wF8kTQW/4ayra9gdouE2Q3Zv440qCLgZkns1HO/km1IWxbhsqR9gbiJFQP/Eqr7rcY60AsR
MtmUh69ikSEjjZU2SvxEYVTjvZndzfn+Dl5wOiYTlkISKPins7k134jsJxzyJs5OV2H07J9SIRGl
rUZ66IBXgQksXUz2NBQF5u1EqIc93nDxVPt3Iumr2BDxMgpcIiQXobnHYopu9feSb483u2yJkmk1
DDaN/dG7mP0r4n0hasPHTk0holz7FLr8bK4J/ynP9BDr3tr9c+NUdEHVq7atzLYdp5txVaNB/YWg
iebAVKlN7i3K2Yx9TOzF4dUEPx80mOWNmElIlncJZBhpnvpiFY4A5Sr7qmhD/5ZWC134hjtf9OFL
tnG8hbe1uwoM6dsZ2sXzP2soQnIEeMX9qAxkYtIFn3qMvA6JRxERYt6SFiyTIa+vtsRiLEH0J418
ctGk/qfeVBc9fvW0dKhKODnRip8Bzl+xcWCZmsp8p7M4e+mgrvMX3y/eMSuOlUSovMAKKbkBGakb
BkpXcOGkCeInWyk86rCqwlIi7Tiu66XuE1+R7nN9+QbIN0w8aBa65fMH3oTm6JGR2wgYNYcmGMg/
f97uG9PQ4xGVOcHgExRF5LZ+7iuwekW8IVVBdPeP69Mb7GQ//8hFI4Y8ZKnvjIJxofDKSrJ9Gz/A
avpqxE98HmeYclU2o7G6KX3OuhxUPwSGLU/GqSwTN6oNN3+IUpkBpteaucHJ9q0GRTbtMGm+cMKv
Ng9E9awnkcx13IiN3h3MpL/cfkQP5eudYYz0Gy1AwsPTDbIz1Ux4B67o2pF8WUmilFCHCTm+Y9cW
0mCJz3/ReS0h+o+sAk1hbMzkBHYbe7lzSX3f9XPDQWgzh7rlo/8pL3I34kr3mQoqtSJTWVJDkTA3
5RzS8l0DVLKaiRl1NrNTSjWMTKbTW5ur/ElUM4LG0lQhf6Se8e57k5pSvC/tPmxcncjbvVKRdD+e
anjhRdfrjtlqWkPK/wJJWrsXMezxOwZdvOnl/gB6QBNsmTjY5W/Zdc4w/70LT2oW8mO2QjwRNdmG
knqxHheulpSFsG2J9NSFuY8pvpoq8R3xRFApCcSl1uSsv2oAVZx44Vh1+vFyJP0s+ONJLMlSZAFA
Dva8zIegYMKBuwSoGEnuQPr062Va4qxiUMrsxUGjQkyoIy4fl7Hk3urVBHcH/uUtDg4zPZqd9vae
usS4Fvr/TPrf5tFgN8lL9LT+0Xj45jtn58RgHEtsezzCNWaCkM7g/SFRcrqYTbTADHFqthYw4UT8
Jl/0tZlwl1Ra6fULfWFotwRrl6Hjn3MRAMCJKw1oL46BM3FG5sdXlKcUvAPMex4zjnBFl8Yosv3K
JRto8EVBXd1rfJwC4C7m6q20AUyEJmW9G0EZQbePESmlKtOx/W3jbULVbkuRCTviglNhIuRcCo0F
xi1+5LpfSmc4EwpaukLp5HLgvdJpNS2gvfsTWK5xNt+io2ovMEic2Fd9/Bhd9zC9pGQiRJGYyF37
lnna/9t4qBavUXJbdzq4okO8avI5T5ZQdrl3j0asveFamBgB1vdBeLs11///KWryDJqRc611hMx+
7PVhvgY0aR8bX8npEIYkXS/kJnpYrJQlFUlrcuVyBXZL+vbYX3qEZNl6HhGlIbrnlaMw+jQVe7oN
n4ba9UbaYqn5mOgW5xC1vDSgvUTZdq+wDTp4dL6EezXsJF/dkNtNdYSY6F1f39Y0Ix9dFqgoTHGA
BrrhOGDhvYlGB7a/94fqwCZvbGIhsGeL50tzKJHmPE7YQPt2eRMoPmt0gAQguyZx2slHsVTxqpI/
f4lEB02Ate70ZmPQEgB9dFk7CABC6+2rsKd9gHnLANYS93SKzGQfLnj6gTjqKaP1H4y+MrBcIs1+
KFN9Q5eecjwt1oaxx0CTQ60WEciDu1qV5OMXgHijrR2N5ripSU1sXUxG82TFtqQOozi33X7gIhMR
nmYPTBrRdF+gd+U1CovWgILjlwagnQgFOUZmWURMYbS+P5cEkUK4Tg/w9aLBPct7vfLvS1/uxGri
EV6hb3AtjK+xD/qS4EwpB6FCeBt75NyrRxyec15UWisxYHBkvYFumrgHZFj0lUHQSLIknbd8/YGj
jzSCltbDx4FUhu2NNg3OtsyFcWDqm5H//aUbU7CE3bJv3iE8qCkQGB+WxJnEkBOTUTWtqYAy5RDZ
pqjZl6ReUzEp6UMbUl+6AmIr49WDF98B9zNF4LnSqjTWPSZhKraJ7Bg25z66D8aQtwlbs684Wuy8
eEwNBPLtLyxx0CWdUl+nhFL4/w0wCtPBq+5q5Yof4n6f6mEZKNkgcu0rUbKeI8YxMXuHtNshcoXu
08uMEibXA8Y9A4+/LPCotj7O3kKh3+okZ9OpZNw+lm+o08JToqmC24I08/Ynb7RedtbBdXHjlJg0
PJNJ1IFzyDkx0I9xZXrXuyJtRd+qDrZ71Jc1ZAZzSPrtXGW4A4EM2AUge4tX7inP7exEe+q/CQ5W
h9e2SsvTqu4r/1tPVS/hVvb2cFe5ofSf2G4Tj0J9LdMoCOq7jp5mXpEjFvjbTkkSjKOzPj0CGXfv
2f0XA/jyWJVzfKRuwIG0toG/GTyzWy474ggs/7FkuSdhx6sPdIZSzwMZPyt+cC6lT/g0wV1gevCY
MrjRz8QLOQ6ZMtPZ+gLyiCXRoVTB24jqyuf+pR7uOq9EDbM9F1b6dH4gfbTZoDxk4vleSgO4Czvu
SBZy4CBYQhIgWUxi0Rr8A8meiv9qzHIjBsrZY/G5l6AK9D6VuINiDzcLrB0Hj4hcRXkXXn1DbiV9
iSpeI5pxwGdjWmIEReZS5bPLqdZNdk0L1EXhb5VXCacQ8tcC1IQPu7+6LW/7CkYRgeoHyyAKbhpB
QzrJYU5wVMUdybz8AM7oUcaUnY8D4hvuxxRqHng+C5hnBbbDHhRmT6lLdR+CdPz7yDCC8XxTCz9u
/pVeSqsvKR/RAcFtl7EZvpi2fIR0/rI/9+CmyMzFr6vg5vHnkJIbpNFXAL8qfnaoLBLmROFSu8tw
LUS6x/dV34JEBLAmgguIHL9T25B3fs82cLUT5Sv7Wd9eLmNqXi+HASE1XV9jXi8A3tgGR8nJO7Gl
eop+tANvck2n1lG+SrxLsUJqrp5RFI8KKOtYYQKCuJhVpJxulXNX2Mf5mAfS8jNELLMS+lzfMTor
szW8bRsYB06JkBkKIcGRahrK0z2yLx5UZ97sSkt9InlO9O5ftJLTM8NL/to/gYJraXMisRg3JhWm
/OjFphQpE3wo6Jxf/SXZK5V8irMfEo+c37hwYRypqmTmIT/rHnKNyA6dg0eXeWP+asTaePKz+6B0
KGDsZ352JXQPbmb90HREKONC8t2PhMgqaDQS8U8G/xHWkL2JYeX684W8TYSPQWOJW7JqwOvmedUv
XByKWVnIHVM6pH0mOrEeHGbQFJ53+5hiem+ZDc5M/rdFfWR3WzfCzwMpWCEyzw+0XNHR15LcPynU
ySv1K4pXjxdFJFyf2GGpnEfFBTjxn7RlNrsgVtpZMPonZhk2kKhBP7wlWDD1+R82dZfMMWSE6qJn
oyAAscPa42nasbZ4kD8r3BxpqqGegqHmA8zH2a1KenEd/P7COi1pjnlrKfzn2P/OuIqqEZiq++ck
iCsK+s7+eu8BKAJbaWJ3XhxfIqRNvssvABdRSLWm6pgT4h6jYoqu/kt2lfWNcHy9eoZigyNWBNd9
3hmJdWqdytWHIWUMpfKGaQ+/XUVA9+fQ3S7/+ftH0bR8PuE20XfvEB/9XMxFzlEk4rPTsG2Somvo
4dxy6jdqoL4YUxxTSVUs0Bs/OIBbXKsrLvuI231OQorwEL0rxwZfhpqJLW2opkod+ztEuCuFcKvW
ZLdevtGPmpskZDBeo/5A2ocdP0CMbw1T09572QWbW13vDLXHs6uuqfzmd+sNzMZH+IYP6i/uVJlk
v20+SfqIOFe4uJmJbXoR8+UaUqFOjCGD3a5mmNnbDqtT4lZQxjFJ23rmocSYiVPP8HzwXB+UC3uw
5zFuHEYp4Rhi3I1hzTHImFj2aRw0Vt8HTQgE6Pgeb3NAvQ5q2z6sGHqTgkw6BuzXxTJz56yRthEf
PpvKCXYtUrWSH1iHTBC9IEGLKON7K884z0AWk41PAB1vvEhvipYVTD84jEMbby7Y+JV8cr3UyvUQ
sQr9dmAMdlrqCL4dT8LibRwUQKljuP5DR8oEfnJSki8jJIE7MIwq4tbL1KHTMXIwfWTTCDG3fk+x
nLR5sYLHZyr8pDXg8mYFBkiExuD1buk0+GyP1NzGWnG0oIuKsizKGB+/UNoxX0Sz7GjFmdWxj0jo
fW+iQkvGC7MtppmKGmCB6MzpJ9dodUE1ESRKEJFcI2lMC170dO+Pms30ngvZj7mith7xnTJ+w+rb
zt8ee04Jvoi5qh5XTjIKW7HZvB8vxaWyF+XttDoz14LeS4BXcgY0qnRavnc/0YLEuoXREBGFW3Po
u0E/58RJIRUHYUsl9hz+57C7jxT3GgfuD9lK+N6va1QmYrcdGP01q+nxqVnCOquDJCmB7Vv0w4cI
pl2BBeZHCKSKRE4wA/LYLhNzzdO9/zXlbTRYrC4edfEKnKT2pv9vrS/+GaxmcPm6+gs3d4vk8iwm
qgIUWeurAtl0ZW4w/biOEFX6ZBPAaQjQgq5+Zz2ZqdPnqzjyNyZZg0vK93Hbhi1ePOTZ7/n0J6qB
HcZwWf6XQNanObAj/dy+XAIkyDRMuphmuJPuVGz34Ex8VvXyOFqjruJu1LfPdcQ+z4ZBgAdax/qr
9beP3k8050NGiTeneH6IIQK6DF4tcHEwnBbvGboV1JOYIH/tyxG9KL4zk+IdXnjE5iKaAARAJwMD
1y073NWNmu0j0u+sZc6v2LG5cLstyK5pBEvqMLpkfm8a90U3AsdMiY1OrfzffpsqRn37hysBVU1K
b+V9/bU+fcSDTHTIwhvy+lAiiIlvJFoxkWg2Erh9Q5bjtGuelrLaGgkA4tq0WE7LF1mcpD+vpoIE
GciJ69CQ91fwng6G8zPZpOck/SAQR0YlRLL6oGGQu3yLO8EZNbxfmPwT05YBHtsp3AWYLTDhVGIZ
QIbR4ons7z37zBEg5n584bvmbZLQhEK0jp0NGfiFQ8mpzbo3gsdqiGLImn17285CQs3YnTb3Ip0s
x/rUg3u+Q4KiP2Yni1bZxD1VqCBGev4CIB5V8twZDLJKr3SfTpdStjR7EWsCNeeu8gOlUwdkMNhM
54oi5FlY79y6hgTVr/0GVO6LZkaMosAeE38pZQnSj2inzTlxKrgSS0TV1FaJoiZXxUMXHVrH66B5
YRCwMpXHehEFf26MMUvy/eYXxVY8Vs7N59SMbjKWjhSV9o/bhYvJgZL46t5LRailbvBdGW/3EORm
xMqKQz9HEzsGHaNPT5P3p02gn55zMztdgyAZmx8JGtUGDD+BlM+5ph4T7meJF8YAD+VHvgvRV0A/
2yJSiC/xl3NSgZYq7rshoouW/9jiO3qXiOhGjsfxOD5Cijw1RRL32Q0D2QUjB2GvlPIdpgObq0mf
N5aTnQ/CMxUy6lMyfG0R6Jlb7QTacbBt5iwMYBL3WDSG+4m7Cb3eNZrlpFaTLbTe4xaqT4OO1fpl
58x/fAZYUeP5Oj7Lb0ll4LaVQ6qGUQx7wbDrDr6M3CNR+91ZqHNecd7HBrerwmY+CQwjJy1gzhGc
w27dBb7yubzoYIQ0pQ0E44N5Xn6HpTPuF1aaU3QcpyveAYDy0ZW5YbfwGv4Yj4QTnqLoL957gY0u
Vmt3HK6ov5svA1royXSUjrwWQYxNhuURutRTmf5b92PqO0yFaohBtXjGr4TdMDp3/L4p1yCcvj4q
4r5J407WEWCW4kD1EwqA+js6heeIHv8hPpI7BPK88tKLLhPMk+qmm+38uyI5xYGwt0+BJPPQPjX3
HyoWplNBErdMaRy+TsXyXu3+URJohojsYLpMR9hpskbuXNLAIqV7dZOW7zPRkdwwdgQFuT/JrTBX
OteDd92jziCXSnmX+YK/T+iMayQVWs4Qwj/6CTwparu6Z7aIBSPXX37Re0zdJNW1d3LStTy77cNo
lnLsYm66rJsquLsRkxjIobo3wG5p7xf+shnnQOuVYAocBvldoZe0EF3dUHsyoy9RZbfsv6LtCRqP
sMLXexY0vO4ZQ5KX0s4pZ77s9GKREUnxsV7Da4Ev9abFO0jfLjWxbUY1iGxa/hoOjysBnJrMCnF3
3zxHVrOi95RRN6FSYHcsI/dM8hD30/o1CDLokh15YU8RMCDnOoVWDeOM0fQ3CKaAoeLI8sSP63ju
NJa7Fs5v7U8G1xA9RPaLpntHvJvbNtxgflbEM0SgjQ2r68752RcgmG2wEJ5GrhrKY88XXdvx2f4L
0h/3FkqXWC8bYZ3mwoIhdnEXj2E3/5b5inQMN6lwyTuQdgIhAN0MZ9BW09Yj89uff6BsOOLgssoy
Nfi8B0pM5wd/DpzJ3vSmaP4hoguV8HNCx9omeMKr5G1zcJZ2JF22uCBQ0zfV4b+kDDTQ06cXOspV
9wi/ILTYlWXVbcRnfRnYCiI2JjY0DrHm9s5+uWI2WwGM3VSrZr+tzSc7eq9c5R/TACzqKurbhDpZ
m79O/ESaoe5ZRm6x7bxTVFifsONKtc7QOezZZt8lNlnmvSAX8t/Lh4JLqSfX1w62lb6H4lP8RHGG
bPLU3ZgSZDTZqORd49wE5tI7LFRXpdB4/LRajkqZm1IL/N2PWvVestkW/rRQXDguGytyVQjZ+gjz
Tp7y/mXWjiK7P9bYV4ZIbNOmqR2fp3EyiroYtJzPAfvDt7+fnf81xhIcvOTmJr97arXGps0mgUk5
Vi8Opp+ZFYPG5ufnAZ7RR18JNx+Uf4cYsezBsDqmQOi2bVkgGtMTCKwbAyCggAIF7wvOKa/KD4Nu
8vVGLAvM4R/JtPuhNOExlGAjqLAJdBgEjkPK3ZJXQMrCYa74GPMXaGr9jf0b19vR+57PzG4rFQix
W7V5p9KaW2TLOtNJD6Q3RvNbRMhvqU5VKnavxm3IeX8pwM3VrN0JsGuo/n2jplCUOPeeUYmrtUMG
d+uMeXedgyOJtyvbSBeLe2zWxCk2fso2oWuSlX/wf8YyrpiYA1OgXcjxu7MrrvlCCutGimQuSLiI
9fWS5ZE9LFsOO+EHwhTnAblhMYc9mwgP3AvxndaciRGTW/1nBtBI6iulpdrbQt4ntVksX353f1CM
3KpEx7X7xSaKqWD9LpKnA3Ako0BUv17b7JkbXuRvfQqE++i8zFqdYPilXHvnxoxgBZifg71uEkwC
KIX0J0uFXWnxyb0lTzflP2qVTFcg8huVs6JUMvTewWII5RqZIJ457EA3KDjDJBHYThywci85rifG
hGJSxw7+0LqOjdVC6+4BGg1/Wu9+jDsG/YecKkp7m67dHGjvr9/IFK6eKsMxK5wtVy4U/kjYzVUB
G13LGdBSBm7VnwCLBxCyZ6gKqv3CRZ0r27n+Y8r7U6hcX3D0fMtPSKT7iuX8xbh+aryZNmIUBto/
rBV49G81/Gh0lULh8z5TyjW05GAAj82J2s26IkvMiBu4fbxAYmzvhQD77IaXsmviiqu5dZefhnwV
Sbo0yBjZKvrxVhRGOdLbmMIcT2NliNwGfsAPvbTQQ964c/oX70x0ehKTe7A0gWWhmqLHFRkneOB7
oJwoncN2R8Z+8K1ZOSKChx0TSJriGis3lmTtSw10nhfxVPvF/vWMBbMrRKSug2ktsqtHc5L4f8+k
PE53J45Fv54vSF2GcB5zTlN3jUfSD29VSPVcctIJVmbHPkx1Sw+DwAoF+PykpE8swIoFh3/BytrZ
YC7NPkIpnoUlRdZ9j2c3BjBEejX1oRBnEnBM7b/nEf/6YpvfoOGyLb9boPmRkKFfdUJgDWUk3ok+
kjABrGeqbc7K3jgDuMA0zweESCv46wHvM3cbfZlThUKmDLgXl3JdmmNq8MtbylAHxs6udNJI5EXm
phj0GbdbtBpsv6vi5G9dRw4RTtrk0EtPRVkiVukoTrU2GLoXOOg/om/VSoh/h3CBQ6bCPTqHVSo7
t7P7blLV+yYyjfwMv3s9HlOvpm3UZ9L01nAYunKG6ick0P3d9CjKp3S/mSrejBUF4lfYktqzabc6
rcttATrgGJLMxIa2e+6MCKD6bVEXjjZDtD98fqnz8GmLRcNF1pmmJEw04JWzea+m1VPuLUQyVf9w
5pF5kEPTh1h7+NoRMHf17MD1mKUEMlSQ9g4DkqPWQfNllutfsa5LRKwc/qeodZttEnV4s00AlqM7
H1qQ21z85XGoYc1ZgHB785Ki0Xolx/16BinutX0Ky5C0krurT0YlA/r9QFCnbeHk/670p87a5ell
6deKPvM970HIAodO2JnEsutXH8458pRc4DxnXPIXn0kG/j5X5FDuRrsypqV2jgj5u7V9IYcQf0Ct
Btt8DfP8egwVT7t+MNbwZpHmtmlXDCcKj0xMsp3kHIzXgEgkwKrT+mWUAXHXKHU5wKrUXcIMmN19
oDhUI5Bx+a4M5pyN72YyDN7tayRehiFgMBYESmlkQ4DcxIR7vVx716lAUBc4hPRoBIZ5mspfug1P
/pDqCrIMkWMOihvOzclPsUsr/MtuLZSRe5itc7GqQja5JS3RC/691eM4WMsRAfDA3+dJTiLTL9xt
8B+T+5HzOx6zsD/JCoQ6JZQWk8DeogYeZaMHwBpSnZRg7L9D9Fc49KLgvP/yaO9PSBT7gG5eRHIO
0LqMlEkmMvJ8DPLNMNUmJ1ywLciXbExIUWbz+KSfetpbvzDEoPX80kSNWw6s8EPSShWrNz8u06B5
iVda3sZxt3D5GKOfZ1O/u44jNmYQ2SFb9JpFvUhlXNgRd6s5Bob2ehaBh3bR85j9J9yaLXdLsNMq
+5dmbITUwnq2eTdzwhMd8OSZmjJHUIh7BKPwhOSGsh1UBmbI/Hjpn7EO0eAnYjnJg8BzeLHCi1Ol
zBbfhubntTvfa6sa6pikFYy+e65OzmbjSQRA+vRkoJEYn2q9VQY8wBehqvL/F3QWdEwEqScLqhsF
60CiWb/ch6HoIIA/vOzy6tdseEFx1jC2IPrJf3LFPqK3SOajVYncmUMnq7GxwzpH4Zlm4c8k34xZ
CeU2bauBNdm/RA2ko49hb8gtj5avWrv+yLqyo1421cPtrMc96rtt17VpqzoalnRHSG9Iizp0XWa6
+3x6/dhugYu7blWI5xvWKOvKIHBdN64GAaqAmlCfIuA9aWZDPdCgR4v1hMEF3py34k401MHfRecc
aXPp/18OHtUCAY+t/xCcCDBk+8c0IgEAb/fFSrGdVVwjozpJT6XhdoO1RXd9KyAKGFtzl/4FI4Ly
6YsVPc+Gg6S5Qe7WwgazC7V3kUi2krD5aqvidTC0q61eHmRa7WT8dxL4oQYnyT7unUM4xqti45/L
DvPrl/HAXSDVqm2+Ghe2pplDyeLGUoKHClKD0JsfF0kdPnE3vhOLykkKdMy0dmYJ6p/+PDZPgWw/
hKf6MI2Z50uWbPhKXJ4ImQzNgzgWjbgbvcpgQfek90hcNHpovXbEzDOcgj08CpbjvgwoAJ0dlFAh
ZUrin+hG523iBPdfrpKSB/zX5xSl9SBvowUJdga8lNanELGGgwrCjnTMyQQ0hFWYbZTNIeOY1wON
uHObTyVsTQtZYta+QWuUSC54ChGHSgr8Za3Vg0Wv7vEL/xLPUvJekc0kkEAKs5zyJ07jrBadGclQ
7/e7xrmyPMX9pilngyVdgzBNodyd2JcW0qowXr135mm7r69+A59lXW3UaPK2bhZYdMrlDBjleYLz
hwg1++6PJv1LMoVrNjMl2C9QAy95yJLxS+4YHBtpTJRIC0yozMSC9RFw4R0QSLs/O2ZPwWB2su6U
3nDuiVEN8akeb6vW/NAfxpHH17xLbQZN8GdShHp1KPJIDaeIEh2Aw6ID3pXKAZsXzIm7Up1cmXAg
Tdc04MFsuXTSM1hu38N20vGU5emr/WCDU9Ouyt9HTtMJmOf3ffsOj73+q0Uh1LTHSCESku6ZgjV+
68r7ba2BsTGKpYh/HMa5LW1KcY+ie84L1ZEHv6BTLTyWq75sDVxqO7YtK1blkM2MJxUCKangltzJ
q/T5bMS42SKrXl5kZbj7pgI+nUNuoHcTOoZyGizk0D+ZdWh2+mJ3Dni6t4EBRUdkklXMqicKQcDa
7x752piMruxrCofIs5xkh2D2elnvkIr599d1sI43Z2dEbyWVPtwDOk2hfRTojHZ+nJTDwCqTr+Fg
pN3dK9QfuvmqW3ZW/Geag1UhsZ6QEIGVHt1emRHewSiDNbmxIxLVfDmVJnplOMG9R9eJVDBzoTTc
BboY6X+B/LYHMMCs6mVy1Sh87me8JfXI7YmcSvIab6DvZvMNURmpkvmAU8+inXu1k45JUAkLnGV5
LHgVlMmcjRL1bDKAJzfhzdOSdIgUyu5DZBieLJvkDX0nYP/AckQwJSubfXytZL2Oz09n8ExbXlMA
1iz+iDBG8YSz5sC4SlOKpz/RU8ZGfVCP6cZTTpvNTAWrEpk2hF6QOXyTZx9DpZ1pOomQkVZVzKGJ
2F4/Bff4DBDDWoi3dsnQN8saGkq/h1EQxhGMWpxcvtR9zbSFM6manVqTrBk62Zb783gPZuzSy3/l
L5dnl7f1jhUPwoqU3FeqwrbWWIebkmxFucjmbpTvG6z34ggMH3W5aPwvRFmWqoFvTbprf92R7txE
zA6k5YEJbMxrGbzfr/LtCiSTGJmil/2vyYkM4FGLptKDKFcKcVbLLPiXUtP57wHDEOfl7atRStu1
pCuoX4D+Cact47iFuGn7G4dB0pt54UogTlm63u+DbHXWhpjTngGhnZbr9McwLKRA67B4gkJWW2e0
e/ZMaDjKrVHfRAWtv/wIyGcK8zMBIW8PmfJN3oq7jzZBIX6fE8rCN3T0AMtc4GOy+306DRRqO3GN
pRTU5rSfseUpoRoBcSuP7Y136zzjNWkZTPrP1++Oq7uaJyrTNAfIMBDhDfx1ypA+dl3ATjfqndkc
skDcVT4NVCMnGQThYcbNxYWl+WsCyc4xI4NLQdYLEjZl74d+A/YCA8VEH2sKX29Wam8xZk3iiWFY
Ne0BLnTZNT8XPQ9+pgSpdsh0Bn1H7XeddQdaL3931bS6KPM0B28Y01s9gBqws57v7JIPW7jlyxnN
pQf1a1zifBOu92B9QQSnXeuybWlVtIhnXwsL9JxEOrxLVT70Jve17/AFyOzxgDCup5DOEZVgRtqW
k1RtczMWJkoI4PGIkK6nfi5fpqdRNsehqRSy63eSGErtVEC0bDB1NMVR4abzp0VgcSPlBN0piIkh
BNcdpgonJD6T5CNxXvZOBULqQXBF7Lm/PbQGi+28MXF0qCDkrUSLMrOq0hDm76qQxGWTMnW3B27g
9kdlXqT1yIXw38UY2FmDFeB5a2SGlBl+dgQ9/u+x4emFmCh27HNRfbF+4ya1P+ouxjD6Udjltyv6
i5ctdzyfCUgXhSko8BrAVY+KXaVzdckI7Lbmz+VZ9iPHX+Auq4BBi+Pln47Yn+pdrDgoTHdu3Nod
DUYn7cyT/6jE5VRCiH9H9BmzbWmqLdwCL1I30JlmdW0FlsecZWy6BsHYnOYjVnM134S7FnlQpy0m
rb4fWfNizGlb2ycO5m+/XwFlr0/pdod4ZxCGiseW/94g3KXVJYn69IU5taiXWvz0qFM+9REA/gPD
sGfEGIAoB4bD6/fVHd+fzqxPPDjW+Y6p1dmug3KxuZG4YDQ69CZjaTJtoIkTG7YqkINuCFRawk2G
i63w1cOYMUSAZFewKS+A6WNwlxS6hhWLPFTWbJGUpSV/AUtHuYmeWmOQqjL1YJQqLdamEoJnrlHO
gWEYCJ8K3l3TS09zB5ps44RpXGxCnI2NH3SQLBFwK+3FEad8/8Lh+lipC70nxorDUGJINwG6IF0E
A3QHN/vCfncTLVmmd8YkUzVvPHY189k19Bxg6xhdYQzT/aO6s2pCch/0A3vndWvZRaI8tjp+ONS4
azLXfpFj+7K1gGjFeMUBxmrRD/kXyiDqa5wA+4WQVDgFnZxbEnK41l4YnLli8Ys/cIZQ5lkd3Axe
ErccCqWsfv+u4dNwuC+tXmOi7Tr38FtK22rrxhIeNsba/t4FN5HZKknyj36u5aArVKAAIhhOCdgL
hdowNrZJ8aRfky144INv9g7eQ/d632FkrzWb/WjLkzby4KoQODyk1Tx7UNR/9YUWQ3IG36l8ZwLN
Q6d7kwvY/D07hrom1RtbCaF2lN5XQPY3tPbJTLcT6tR7nM7a0cBXjoU+CxoGLi0RBnSTgImqY9BI
gsoBsBvXjw06ZhSW0i5uLIRU2mWl2ai62quXgSvAkCX+LlPDKMIi+UuvGizQ5iEvIEpqVvc2YrOS
2tmXHBlBFtW7rxxY9CdkcSmcjY7N8ygczd9S7jPk/1iQdVSzFEpXf0aTxX7+XCJkOTLrjnr8h8x0
tD9TUT9BGiOFlgkvTYwbUUrbDdmJ1pJll6FJEhp9/u3idZj1Db7G1vGNTjoSd7G1ai6ejByqG+5m
Ar29wNPgQ0I1OLzqRREnY33bbLZGJvvVcj7OJ08uy4yo9/YZw0qhy9r9lvzOAbOVDkjS+PuZGVBl
OBCmh4zvhG2FI1Y6ZWGxjwgIIugUuU0SRxvM5S/OTPl6JypgpusBy3f6opZSFCO/3xUpQYbvmSOi
UZWeuC8NMGp+k+RmmzlbYW83wZewmfXHnCawUu1dXooXnwBttlPQaUtZpfrNhPghUgVB8fUe4npK
CLWt8BH7oJ17FyJeIYR8yg/rPw4KNPNHJF/2++Kld1frPH5zbMzvw6Ennsp4kWq3QrK1uj9a7J9X
KQefRvO99AUtZCGREbW1YmIKR5ecffq0THyX2WGWWWIBpNnbKLl9Mo8IuNPvQNNprr7uPKdQ5mDi
k9+brpBqw7fwM/4dPWZ9CTYj2eg9SRsIFQIJ24g8ytEixJiCwAsBYk9aY/RrNTpRRJCTiA+CbTai
STVcbDEwL4Gc+GvyYBUWCXQtRXNFURY1Ez52lLxx+6DY1MfCllhRVSKce5uOcO0IB+ZREdHHLkOV
7qlxlncUqo/3nNImiSr86dTT9jGoahfcdOtlhQhFJXdUbIPZY5sX6+idDBQKBKWXGn5Icgnq+eFv
/3XQSk3/ngtCDN50Ro3pHYOwPZhKBUmNZkO4/oNJQzakwbtn6Q2oKSMW0ZHVXeOvVR+Lmkt8feJg
CoFOvo14OsYlkOW7ggY1bJINnI8glltV7O/e/do5Jh3z58imsTMMxZ/g9Rma/2mxvKvFHexKSiU+
Vr8iyyDLHHcoTifTVprVxsIZB7Mx33ODE9ZkblYlcpjA1e8vnJIxt2ws9sLULcR4vIX3Jb1Eh4I5
L3kPtRKYaWDgAhJu/7ky5q+PnvEJpml8n6v2Zw/3RBLCeSgTJWhy+TvZsOU3FaD7C6MGTyzkIlXO
5VjwZCPIZGIsimx2O6YZ6PWORdAsFDjFne2A5SzFENwafpXxIi1evxoP4VBI5N8TLMWenSYhRaZS
kWhvGgdrmn/k1A+zgsiTP+rSyHFaiJxgdxQ/UW6yd+BptuyF1yEIwsrr18Dg0esksvtzfSNSebkN
ya79mdW7sMmufdm7LhmZG89YS2jR5NMd26+3bnIR7v5XeSZWceDzkC8TWI27wSF0QDC8M6EAkA9J
LasX+EqgP3PGqK8gA8uHTsFQ7ZfYpqdH7WQEvbEJ8rrKGvtrOBCml4g+IKLNCG6gyUIzcrA1Zkvg
UYzUImwAkUx4ZKdsQKeqQC4hgJpQ+KE7RGABhVq3JFKuseL8WtjiyV5WQNhCnwyvZTf0lypfa6Hh
y72dd0g/AQLI3xm+ZOzpU+xVjP+OBgAhVsC5MISPKwVJ4Pb8GEB9mu3ohrLnVCef9412ozfNw8N6
iFbYOJzxS+a0mLyJXBGLpT2J4+GbWXrp2KboioiJGxMgQbLK5EVgoY5KcWLCWuM/7oLQQ5IPbpRD
ld4W6A5pS6bR//gUdPnvX6oHA2vPFPaMn6QsjG89NKJl1M6l0tr3F5gc+WRTmUjJNsmY44pLGW5O
/H6tpAJvd6UgFg5I1PyPmsordXCAedDNhCCu/4XQjAa7Ad0UoefmHBbrPLFXi6Q9ya158g7v6SAE
VnqPfeQRS6qNo7DXNZJvJtd136f+5FjSN13FWZxqO4m1sKhMVtH5sfAImNx5dLyxMJo0g/k7oUJ0
43PQP+QPAn6WLECQjoK5KPvEOMKU+20CAUqN4ZdenGWtdQjT3l/U/16x7kivwabBLMMuE7/DCB+4
ogK2YozUV/RQW5bqrW3uUWDoR+V7mve+3SCTRKQMUNwiqyG/fAIHl7rnw8p2RjI1wWfoAuQDHcTt
F1zRZaG/NmaHio+VXRhTnP4EUbNtvUaiJ7RiIxQNHiQY12UcugidBDG1wGl9GuieH+nLJ3RjgyMv
Ve6pDbjjdQT5ZtATEdhIPGX9oOrf0GDkgEx5qdfd+oz55qT+5++zcHgZOv976jbm2aun7hvVb5K9
aXSQ+hqCADbSZCoHgAiEMvm1Aqg1UE5Pzz3L1Ub+cryyPmW1pRi0L+69n7LFOMiJVS3sLlSx3UeT
/QsLxR1mxLnyH/KDS1mHwxCqoMt4mxYlK3lH9E7uyxKhs0MXSaWw8h+vS+OwXcR74TBAOVmUatoQ
yd64UAf6k9w7H/vcMG6scQqJWVm1xqOrwmK0KpY6DkoZS1r3mEUpGLFMN0bMRF5ioGznjuyC7r05
Z/niygojHqmmtXwQS+UdAWjJZZA/L1HWxxstA+WyUmuWNvILLwk6ovu7AVJChOrTwUsxLtRSNiln
81+9xLomRVEs3zJppFlBhn/qFOLwgNfHPd3owxWrQKyB/IguSEAZOPPh9keKyFQ+8YzRMNDGhG9Q
EWv8I8q8PqsHPwjQQ+If0bpNRHGxfV4vxxybvTOaPoeuWfz+eE7FQFWu4pKpc9mmiKgENdLpRF7d
ar5438h5nTXulPa7Vjuz2Cum3eSYndLe3M6WqN1SHiCNrVQlOWnziut6kGzY4W8XMw1ZlwKxZego
u/WzlgrEB1KDYvRANJcszHh0TYD64EiT4EzAkswzr5+AxOuO2ZtlcXlMq3w/Ptn2LSJmdcGUVJss
ILPKWzjJ6f3+4Elqj1KBid0+JW2ta/CYQNUtyX66gGW+lzTIOSVRw/GN667oiG9tSaKp7aA4FAuH
2ClDiIpzuIKAoef3QaZcU5QhwxoDnYuqZB2tWhYFgJXdi1cydOZUM/Y/CD1ij76HjcvvAdYUs+NY
xaLWqkscikkJI54+GTLR3h+cNEblJ7ivOQYiZp3O2tNDp1ddEQF7XwP/zG5PCjf/NM0VAvbDzFpH
ErG97ZJNIw3udo/XlEWVwrPH13PSWwBjKJdibxT33Ry5OlYeexja8UmelGtjZ5SjnQAbC/HThQEw
rmy7BW0TELzEtRVfYaNXP+KRwzwx9WjZ3TggVCVIB9Yko66jIk65v1NbPtRBbM9U8OVVeZPFtm4Q
sFP1yybaM9DTXIHCwo+OHPCJ2VRJusLQS5NkFZX7oZe0jHoc08iVqu8piX0WbU9d0MsM1PRk+kdf
T9INsif1w/XuHoFiD3vyjVIi8eZvMY5EymmBaA1I0a4sOhizBi7rdKDJ3UTcFkWauort4W0OJzmi
6zNvL3eQTRHp7NwO1ym5wzoY4xbPio4TVjTgLdJGLNFsKgVKEREv1t14T7DxDEXX6FBjmrjIoqSi
ciBIT5zQOzNSGcUpUbLFCs4lQF7QlIhLBaSS7iIbuP/F5qoJXKrSwORXqaSP9YKZewlPdZ8HDHqS
tefSkVCF83KQKg/i2oUVextiG0+c5xhQPlHKZIUyj1TfDW+ugIhcCTJqU2N9jcDoHMcd2sZaNZiQ
9gqoTL0RQ9iypMr3t/kBVFDS3eCu31/tNaV9bg0jdviCRiEYHpZ/e1J+LqSza24svJWoIXDH24rn
UuT4ADYmy0TmX2Nrjgnmx7A0WQR+FlcOtXF7DQuKD8FR8J/2DaWCUlF+8aNMtDKyyoOAj/d+ymgd
SH2OAyPkU7q2X7dDS4T8DyCKmhuwKz8HDcn/baUkloUJ2OyheHUh7PDsOWI4Nv/3F9O7sN6Y2OOW
QcVsUo5ElYDO65ODHsxkxYbZTd5VpXCJMQ9rCLCO4hsJqwBJoXbbTnH6VDZBtpF6erKwBLFCMW0g
wDX/S8c/IfVXgdgmOoOod2q5KGeWGp5gg2/e5X61LyC7WGOJ6IaDfwnYGTVYKAfw6rYEbiQP//VI
6yj7NR2qczfQz1+uFYDTDIAgSgYs+9ZvH1P3csRACqpV1MC9jm6b/LibiyX5zGPeBOQDNCowZhbh
4CoE4hjRXD6AApguB1DsctdM5307pImBxbVF7S5rUTgmCLoy26ISFRhxxKh7b529ZT7kFrsZbiSN
arGLC9ShiWqKs32JrcP7rxoQdbypJpclrxExtmKgdRR42zG5KHkvNrGGJF5VBplZqN6+s1ANfW73
uDWj03/Q92LaHLGwKKYlpagE27xolQg4q59/imgRJ97xQXHITyApoekN8g9VUohxGakrGBcWuNGw
Gau3luTdRzKY1/zoRiSmEc+x0e23OWBOHI5gkSElLMFFaZqeWrGWa0TE9bzn7J/mPKNoEeBW0+BI
rWeYhkk0IfXABb6R43TSQAvOpw0eRr10sTC3VkrbPCObmpVJrKriTB6Ojx/48FmgdqnHc7N72N4+
1OM5qB3jhl+Nxo/dKO3m5EjgTDSqZQzJseScZk/0JOBdBmnpZIk65T8+pD1jqocMl8/1Lr2pDuHw
yO8OQLcd796mefJbhK00LIXnjIc4S75McjBVGMJiHhPXn+EPR0SdDJxNtyq8riZCFPmngvWTNdjN
g4kKZCvWGEoUp8PiAAhaiM2wGFHvsyVXeKyFAw3hYfAZeUAuHh0jijX9W/V6CWQJOza84XEPJ/uz
XMvtQeujDnaxEq9XFr8L335sii0GzYiwcMKgM0Sjfaiuq72YtfQUcAcQe0zxWQnxS6o8Q63rg0RX
/5ezLisyPrFctHgXHwtVFdmnTv67IwglpyEEVu74y2wvi5RLq/ijBEtV9IaoHTs7rsiTJzV5G7dT
irc6CQj0HPsaBGw9eW0PPkRBhL1B3K1ytdUa/QQFW8+wFAriygt1/wofx2v77+vSeHc0vIqeXAkR
txixtW+VDHgsuOodFzIyWQbIlLRTI8U330NoEqgDzRJMri5NkX+QWeQEjSPjb4YEVEGs7JiyS57w
7ChMeT0YDsy+zOTAn6KvTPUZhsaaB+aKLR7TaGzL+8amXsjZvKMpL2NR1wyltWilkF+HWNRvHg3s
7aTNz5Jm76pdXpT/PZp1QFA9VCEH0kDE+9DGYU0dX7YxpM+PgjkdlRNyB4ynBV8x5xH5/AfEjs2u
T2hdTuZqiXFAeh3jV/N3fQ1PGg7kW9So2JHoVJq4az28Ke1AmgedVU8PkZtM5a/cIEY3eB2n6r3N
7+Z3jybmsAXq14yx30cmixotE+1ww9+0hJk00i9el0wGxFa/lxoI07jM2mRp6MLwqnIuLO/kBb6a
PhQ+zcHVXIHJp+mYm4ODAWx6AoZkVWplDIbTBSyrOYZtAiTgwGVZFlSiMO/2WwCToYGSbYdhKjmX
S3KB9wO7mRlickRYaXTGkxwj+Wnt+LphTVj2E+ZbkEzXfAndj9tCsyo6+cahjD4Lv9ga2S36Mths
Wm1MFWatM0GaTig9LsJ6c610VCF2xABzK65YTHDv2JGZx8yFtiIg0I0AAuvLDeIAgI19euW7I5b5
FAmkrNJe46WujYkw+KHnTTCqF/TwMm3tquKnX0xq74GdCYCX1L/j58Z8QtdhJDjup9j0YUt47LvT
uyZwggHcr4InkQHhPYhQrXOZB0NqMdHC3P6Oi3LhGcYufNvu0GQGhN92en+ZbhpHuYqxt+QIS6YM
aGn9dBFa2zvAOO033jBx0LpnutR2KHQ2yOvAmUNDu6IZl0D+njJCYv3NSB01jclS1RN7zGxU/2SN
zdH45Mt3p52hug+wNQ5rixUrt1gWP7Pmfj7MSOxgk2n9/pugBHfHo9Rt1Sz2tKzI4MniEtcbBx3o
rdaJVe6+fgvcUznd7bsGm2uWI+N8MGazRivS2W1EWFiReKlzhxs2t197EaPwWSZ3jXTsV4gWawZG
0rV5ilmZHVaNBJUIhYgx3GzBHlZMdDvBVVfLmf/TRz+pS/JyUVbkjiMeHd5s9UgKnZ+Wxs3av7EN
uVAYvaBecuuaFi1V/JnmnC8Ad0HjHimS11MjvAY5SDAc3ffmFkVAIrIuZyHSUpFo4WJnpeM/bkx1
NgSRienHBOe8runvTmGZxy6x1hMn3wWgOe4+QGbESfvmOLpfeAfa+XQkYxDeh88cpoG1Ci5pAUZ+
YLSmCyvizDTeV88V6c0MpZAp9KspAnzoZZ2JVoffOLd+0yVRZAbb/e/qZC4XHBMbqfaCQ4oX7Ocr
m6kW5bHgfdgBfrDLLF6EZ3VLZ4lzSauqVfc9RFVLrgeaCUzDwhN4Z3YF7+0OYFh3yvOkmjtcOPvv
Vq6TMBXCkcIo0eC8R8oAthP2rRs1VoJ/8aY5SLz8CljB2eVafUKFnavo++yClfI1WhkYmUVbp0tg
N/leVjRLiXPgPOx6/g4kcyuPH0M4KLttz7Njdkuj1bN6cDmgxNDw8rillJhhMqoex6FF6pmwvpQ2
CDuVJNWtwSiDxmvVGQ4kfg5fBED97aM41hIwf0cMK+zYuJrsNGzNyX5q1byOaZ8yVghrheFe2uyI
1rRUnzAZa2t9XJIB4jqsm/RO44T9ZxGiy/4y411aDQU+E1IGNEL3FvVOsCzoLA4DZvt6Q2BAUpoQ
NgIe+1KWmaJQ9xn+q3F9J/BUdtgsGZW3EUgmMxwTDSHBuA5t1OQXfoK70cyziS1W1nRZolRH9yAo
coX9vAdVlswB2b5TVdt/8wGbVYgvW+9ls0SxUrnUSZC+LM9wVPa8ankdd2o1aDdwl+qWhse8mnTY
WOrFZJK40AYdBtPZd99VnHalEiDhsqzMLb89j35+r862T5IPhWLRYmKqy3g7QImyGZ9sESfTKHkX
Ed/TZlL2yi0e/MyXjMXTuXXiCTInyDxHs2y2KFdGsBF0RZxqMEyuXdIrDf/V3gDBAM+ISl9R1u7I
VVlcloeVj4OjmhZTPYzev6z0XoztifzLeBZoiGWM1EJtknvaaKIlK7mEfXagw8LJQI18WNRDycgG
TY2kvz97/qYX4EXnWy2oexA7VoTOiiWiDUBy4q++cwzfOlIesosKg9n3bpFxdh9JSxfQIU9EUoAg
o0fITRpvgKneM49ErYr2PJdsJeImPscORWdcyGaWgC/vgXhHMeOOmWuclpKbf8xgXVgmKAtCI1Uf
YacYuhyVk9Um96167oLouU0/C6DqG6sgEExQfYwjee6lFE3Hl3Xsvn4ZXo9LB43wb64elJcdAEpI
/dJuynfv9PZcKKoCS+mE9qQiyTxtjYlAX5dnRgeKKVMvT2NuGIOJ7eNgU5gS2oFmj2n1qPBzlhoj
adjNpj9wqWgsODeXkW2OVt73ZZuX4kG5q+e93wPASSQMdk6mH4/5ff8SxgFiidHWs/DpGvKp5lLP
pWIJEdYhBOJf/mxcu2slcyVJdtA6yL8m8+jK8402gKfjlLkrc5nhq133doxunIXXts7SWIIn75/9
txitwry/eO5F0jAOr3q/N30MzWxeLASyTaW4x0rbCrZ//3r0i7X1gvbCDnDZWXt547XncD2sHz8A
rm5+W/ecXO3uxtXtG/S2Iq1wC3gcCBlIXnEnNlBKyYimrrpWaRlmYNzOlXDV9DBl0ZRR+RbmLb60
EXaZqj0mb5cjTo0ZY9l2tfcodaMjJYlu8kApDHiHKn46Xw2Tcfyj7f2a/HWKj+Cq6gW86inax8vl
HDOfK4Nmy+aU5cS4dPOw337NOJYXY5+94pFiiQVywziQl5n07qH7i0vI0hY7xxFQB3J1KstsIzSD
8lUoUdzOHYTQFFYe+hHPS6m1+hGSnIaeNeLECYo6js2uO3tSzYtZHaubWImZVQO0vMEUYx3t3UG/
9mlGSQ1AJXowOpyurZVg81rzaAdJzTQ7aAfn0f1evKFGpdgAIioH8sVkVbeKcrhRrCIzkmfvWsJV
C9EuV/xinMHAJR0gf/DnP4y6l3GroyO6MEFBbPR/lay/vxtyF3BBKzr4UcicoDM+PJjAqF06FaW2
KyAKm1Sl6I+K6RTqlchdVvd71jvwiYxDdzo/mPVZFiZMsd6T9p/vDwLDIOy37e6NGYRfFU13jfk4
pcawEpoX5l3HUMNhmFaE2vGEsOef/CXQCnumTt505DfPN7JdQt90s/2wJ3sN6OQqOoCE4yPzvDFT
FjJYawxXoLQvAoYwSW7Q7QcNaBlzllHp3Gbw3HO59mz9PFta2XuFvtenxLxAR10N+rTfBzvv1kQh
/wI4+B20t1QAIb+LevxetnYSC2EnpgwY4hTI2bFx9T0FW5mNJcCEJURDA6HGcq5+ioiqXFCcPfPM
PS+mMsQcCEWqw3cj5w+Ub10u81I+vbXjVQKWdZzVmDFP+M0hiDKi8h0PoOyFZOEwooVxeNQfRBKl
tD1x5HJvhifSSgKPKSEAoHlDgckdWaYoqVw0uE0UTLwHjB0heKRdN37DKj5S+5ohoKXOPC5r2DRD
qvKq4J3uehI67jUGSRqr+5epaOOLFPLF3QGUCLoYlV/TFc3XY6nleRBFhDaSiP6/T8q59lWu22y8
qKBFyHZst7AnEmridPzEbrpJrXsy2PCsu08h1jesLc3OXYnaOYEqv2nFNu/OUFgCbRzAJPp4Qo7X
lB3M+E10yy6CGO6yN4wvYF2EBguRjt1W2E4zarxiv6C8yi8dL+XPvcNMrHfwDdrIl3BAMQQ/vksm
mKu7aCHSOPPpSW6wjGoHAWDGYFA8or8KHahYR+ZmIdId+IqULpdwHO/2/b9HeF+UoMe/2BqxutzB
reXKpMCg5IOU5nGQ8VXCD2bRG+p8SF5Q8S2D9QJsx5ANZpozaoDL/LGVt7EpvbA089V8osvSJqeW
ylN2sUQ+uxrTDLHoaSce/CYzHXp1Vsm9FDNvoKby/rHQZz2BBh4yO0ZPGL+1Bhk/v/0VtHyvVe2j
bS/bJ1DkJJT0PC54pPvsXjgoYbogKsnmDmmPO8tUh0MvNXM+kp/IXKCZXeTiPzAk+fOwNiyBAqYr
+u+q1Hok+rbMfn2v36BQn+RltC6KSTr8j4CySgYgHvhZHAsrxGOSnT9r60W3NZoIRx5JjycAYaWn
gVmDVZLJFsfNey3G66cik9Q4JRrl0cwPynoRTO7PI98F+gBDeh5EPb8bdTT4eMWj2KxPBBPhofTu
N8hruMKl10Tk6gyri2ljSEJ8QTbrWVsBN7IWVqsm0dg7MSggRxNOrOPNj4nF8UOLh8eUcaiZ5GZq
liQiw2oWNw5GKPpg7isW0k5eo9Q9TsSdXsQ60YFojQWZJn5EcCZd70WVyootV2iBY43RBIb8X9yz
LJpG0hSAletv/M7Vm/B8hq8NsrmlvRV0+xqYT6C5Ig4OtxFwCQEL9B1UCUg1Eeu+NmPmwZHxjMqT
GhYu7+O7LgwfGqv5fXKsv2kWxWvSTCwSdzUZ9ySS+XfsZpA0xyxvL7Iga7uxXnnQs5Tiim2hMhQ/
bdOt2SH/jg/Yks7XY4zUc/I6Kd067u9UNZtb08XBBUYlh9MAhJesWUyOVMSxNHHfdYI8Ueks5S3V
NHDlLA6KGMvqbuVIaIx7T02p0er+bgT8WiVyq9YsVXQlqkE1YJoOQFwaLZCM1QE1mSPGOHlXvFZH
OkRd/D1+L+RbV/23WB9WmVi8iPHizeJ1hiLjomg+bWxv6ECRkD+TCZIDc27+CblD0xH42Pvqgq3/
kmEuCi0jIUIUz1Xwd85dI8exw/5kSuwgTUAUB2Pz0hB1vh3hJlQbj84tlV+TdJracBta6QM+wtox
pGh7AwgPhkS2SHlhiL4BPjS9ZtaewefciwDlSbBJy3x1TL/TRuIIGTQMK25jAUUM/hLJDX/pS3Nz
x/ZYhGnZHZQoWNU1yRBOd9eYxUNUisg9NIGoqCc+pdRBF3nmtcZhwDXpLJ2EePJ+Fs8FAV52u252
3hbGLTGk/GDj2jS91izrZZ8/Jm9pJOK1WzYGQ1vm9di8myrkALzoZ7EH/FdK8wbRY1l53gGNvtps
hbl9G6wFoMokFcMu+31JKRQmhbXpE+rm31FmKOmdv9ScJfczoDLbZWYqbMfIFU802B4jTm/wy0Rp
PFtSn7ZGwgL3ZDgcFHQUvdPsKUBdlJdkB8q4byLYXSGQX1he8aj/J2wlm33r7ddLZzbiN9duEUrg
R8cLRJbq1goTqasBDOv4Uzes425AaSxDDhysvnGysJ/FazX3e+iu/EgvkRy1OxFc4+Ztsc1iwe3h
+ZeTzmxYChx2OX+igFTjhl5NXkQPK/hI+QMPcYLavDVUICnm3QlFgfSSaS6Nk3bNbSJI+iMyWhTg
mttmIWrgFnt7Y3/hVPFMqYJxNR+1/7HT3SxDPx9WVJMRMl7b/D7SkgDzDs0Y5sBgUNV7SJNQh35Q
a1WPnFmMQ0pAbQVvuHF64LbpADBppVY9eHuApTtPjBCTLcV5qlA05npPhMD+oR3Sm7cQ2uYzIAiz
L3GN8juZKMgl7Li12YyVVS2kCjnf6wKy5ImR85Dza1pNKvMIP2zswtc5b+ugCFNFM9QgaadeYkTk
1kza4HmU4C9TWWadSLN3HmnLFShRJNds/ZizODbX+MkYJTrH85P8iTcxyvb2bXxqQrHZQBYi45N9
Sy8ljGoZnSGDu4abkErjPHwV+lcBCFuv1wsF/7yWwjxevXLxIIGyYPRfRbIT+xx8Wl5izseqpy+6
wz0DGARA2QPcpSVJCoj3Ea86a6zsIddqBeZFGWGoCNBKubLuzoa9G78EaANp5lvXA0GPoWiN33cv
E57rTwBtnSkmuzq4MzUQno1GcsSGFN5gpJeXbb53Mvpp0yMmsWCbiGQAtg6EfrRCRwG+tVkWopIR
S3yw8yv7Mg+4svSihvT5Cdq13lVrXf5kMdfkClxdGuu4Q8C1kDt4Xhor/Py/sPHK82+skB8jUmY4
jLZfeNoj86hdie8ZgaPvwJBtfnOmMgiTlXjlH+0eOFBDew3w5cnXRSftvFrKkTVkjPMEu0R0rrxy
ohIWLHohB20Qnrq8h1qfqUXZ7OGAXMQkOykWBM9sAbqLrIvGWgJQf5nxaquoWV5FI4G3u+KtroCh
0JDmQRtBVbZKX7Wef5oKNiHA95bmijh3zhq5OMIQTmhw48XDptTNXTmxaPRA+EdlWGwldeDGHKj1
70P6hqa9qOiZreySMPWjAwJFlMSZUtyhMS1QUDFKExtIPQuq+/ha4VqSqzc8ZVcKu8r3uXMmVirO
CXNCNb5BwdGR1gSjOhf/QSfZLkOvIt9w+eYvmBNTKXAY2gJHQVwpOC5thY2Bt3mWZCplL9AOQgYt
aquqp+9vj7AVfuAwa4c+sn+Mcyz1Byu7XTqqlOEaTjmxY9qb9Ogm7uo5pMwophgtAeZMMgZx+fv4
ZR693ustK/piqds2i05vD+rbnphQMBVAe0FuFnduHuJ0vjov6PJBM4DEye4vI2EO2KttFJV71ZNk
V/J4hSpYT1Dfp3Zi20V92pB3BGKt+OXFcPNjaLqz5/3afcRiSNR8JgU40fH5w7RjiX04eLSGzODE
nwCEj03axvq9SyAbrKqyTtHtdmqlGy6Z476QlDz3NQwW8+TQA4gvKGJrqQeelCBezybYk+LobFFh
QwjIt6+Lm0U4PTIACLCaROsU0l5lyaXj6zSqG9hpZE8sy7yt3etYDli4FL//7BAk1VTT+c4obnl0
m+MtPajxGg6zf745bYx20J2eLLoJR+IScoXyEqRzd9s5uiJF1XeKQdgiWBrELT6eAQLE4nQvq1tG
7eLDLgHm+9+7uUy+eACMmCyOwz4kiHXjipGLhgSmpqLLCHnQddu1/Sn/j0EMGnasfazBylGWGyxu
I4u4hWTnL9ifDvvjEC0bzbrSLfZFhYNDKTIqSx5Sc6p+XSHH32LZ1TIrqK32VJ5ZNpdLhqDnIUgM
t3GB69AlGWNMHeonQFX7ch+kd6T1tht0YT9EWZezVHsqSVvc/iJp3rHka7RRLbo7rgcNPQkm51Ha
LIW/HOYUQlMHQnrrochVb487vN4OyBsmd8xLYY2XabnYTIjDsAuib0ruwv+kRxQLQPv0jjgwdiXV
smp/2kKWDT1AZLDJpqh3KoumQFzym6Tk1HCALeTXWRUijhJhBB281eEbwtLmUnOQWW7xWRoObVkO
p2Dgzgc9OAZdOASY7FSQzXWBZ4dV3z/tRXbh5dfIet/JlzISNeuy/uhtyPc4+1DJjydAgkITtQlK
06cSDL3KhlO0+plBGm/GjCDOjVWLAdoepwctTHxiw+3wlne3gme2ZaSwt9w69VOsmoN8OE9eAS6O
5ji6Unec4APJ3FTliu3ENEJQYoT7E53f9xLKFqik7NXLEb1x0s+g/7YbwLyzx3Ye2l6HAwe6OfKN
A/RGyzlOyozf0I+wbliLPKq+kp+0ngOrE7WJ9so95Frjrfu3MoNJK1DmGCbM9UAKxuxtEp6ikwLa
cbOcjj8E68uMM4SZvpqfALgVF25H2Q6EbHo/sPo8xUrdk04Dc2oXMkHeBvoSSrqj3+rmu0rCOqyO
9hQWB6MLw1XtB5PMdLna5Osp7H3LlPpeC6Lk7MrqLb4jx503+CInvOMepwTDIAYC7YdHFZA8rpG/
XC35HIfAs2ywGgNoVBlO5Bqs/tWaBEF7s/5sxY547rkmI4x1ukmiXFOsoDWFYgZ8NV9sXfVkEoe9
Q8XadWWXbX8TAONYxvZp2WE1LuVYxT5uCqDiX/Ilwj3hLfI2oa8PQaOFiXf1iM02Rn9OTSqrBmN7
HYZCwxwJP0oUlZUyBWlWKSBFFksFGrK8FOt+/bcteqJhwMcRj27vGFIDP+H91UbFRMBchDmSHbZV
6CqHXH0FGMuCE5qGWIAPQtdS/ALu2JQc8OgwE169cqm9cC1/0tmTTLp+NE+y0ycnjKakww/rGK3I
aJnH6MJ7ZLKUG57iXhmblJnzq+hW0pAfW0YPrmBdathinjUHSw7G95NEhBiWHaoMhn1xwNLblVNd
WK/GhXyEo6sqhosiGLwNpA2vY/+DCFkSebAF0h+UCifbWFRlGECQbwzrljfseybLhgOtrgtQ4vup
gQh4PTwsD509ch+ifXtNAnaABbCWipzboyhmJeMHXpU9wt+rOw9hrXdBK2kUe1MCDdFZ55sH0lpX
3Oj7wtLaxqiLYQt0D0QnB1XH5LhMQJ/PniOhiOOUKlOPxtyI2PPZqp7xRzI4PfkTVQMshXm4x3g9
njquUHDkXJY0xKKCUV/fOpvgaMepO1dd6qE5GnoyQmyMuTE1RctecqhUybL3UfQnXy+Fw1iXH7l0
SWjO0CcdnLvnRarwdUZ849Bdiz+bgPDnMo9lMf9vw8vHg7iSWrVkOOO3vjdKExFVp3MafAD/7s9e
w6VJUnBlVNwabUDakJJxEGQ6VmQg+Y6GiVp4bbx/b52f53wlMvf+1Eap0tR/Seeqpdoqf8FzTxto
rpnJtIVupbqG6UnflbhItLQnectV/6Gmsl8FUOu1IUZHzKeq8kaxczflCV4TQAeOPBZD5rzcZRxt
CEyc3IhcmUvCEgre++ZDhc//Qc8CggzJbOMeKZ92ARtBMl/2b75o8RE7WbztnNA/JycZughlKzLe
QGm/GEOOY/zOiJm0ZhFV3K87FDJbptBEb9qBr7t+IepYj11sViHcV1LumzsIJAbc0brMWYuAX8SH
hNWh59fEHGx2/SDhuLH5cKILaKZZ786bJl0dSm88aPWN1rZhaBKwMF/wbYqRo+xAzNdXad5OVl9d
FgmWLpcF+p//vBlXG8FEmpsTYXfB6f8i3fyRnGZ8Km1JafybxMkjMh/RiJc+ttml/DRdGuA5FlJ0
Ong+vesQJjvAX8KxpE4IHF9j3AlHtzPwDy/D0IGk7ro/gkfYDKZLF2swPQbI1imdQ53AQhlxW2iN
Cz9M8sVo1uMLUHoXaAvzv2hHk44RBA+86kZrPnRWZmYoFvv8rNA5AN5Ch9Zb613utEfxdgaAP1Rl
+mHygK8zNMSEn1cl2oNhgwyXkqgjkfVpiMTyw4vNarQ3C1S91Q0ICT8At3OMt23e89peHrHdc34O
KYJaas8fQdjOxkRICNj6NMHYZaes5RuX9NbzlozXpT0bpGvj2HvrOGEEai0I3XzXUKNfrCHnDUbK
LvQe/LuON5hKKlmd4oXj/o0amxn4c+LkkpoJiA81pJy1smNDQdhV+LLBPgYu6eZVERq8cfAIlIr2
3vXEfdLSLEZvtij22k7p72joByk1xX9VGjnQpxXK80IzmhS3vzhJ8+NPrbl2bZBqLsqvLYu5pYgJ
cT6tjBb4oruvSLUbvZu3xU6yzQxloSqtS1gteZGzy+BRgbGzPe2BOpwhUGj1Mf08Z4pSNlSjOlRp
yoi6vHXs7XcBt45HFaMhuo86chTtF6EpDH8TNuURsXb4GN4zLD9kqTgtdveBF5xoJ38jud31oKxz
F1VSYOgTngLgAeWzUG1Bfedaj4nemClLUK1y+VqgCDYLH4gxGiTsNPWdSdhjlSaN6nzzoZ8mCrnz
C6MmDpbeFzJ8sf2xtLE3Tg+hhZpa1e0O3GNmpn6H3ToXumqZQP+1itn+kwO1TsrfcY9bWeW4zgNw
XsxpHxTqeaAOA8j5ghgyOeKnIwZSfpYH2wa958P1Hzeyu3hAeDswkYirITDWHuioCB8lJ0iYPdkz
i6OA5pOhSTAXLBTFyi4jqPPokxdl+SwRc8naPpcrdV1EUQQ+fz33h5VGT77QkkE+u6qBor+lYGuE
fX8p0luHG9lLVkPKMm6BlJtKCrdZcYzkqEj4V294HCsov41/elRaczzbHXYmev3hnfA1hk3Gv0Jl
vk+HVuUtpMlWsBjXsUa+1Hfpwg+85629x50vPWmhtns4DeQaYTXD039u6bdWAOjvJIfFYJSPUFlH
lEVVMnM/7UmvPKd0lRANwjaLiag8mwos6nHZGd/2CZIvmrp3UgnRqCjt9mbEQUIVnSbJKbaEgvkP
rxszR+R4QNd0CvfCRAo9aSj76KOQEj2MJGaTV0h/AvcW+8M6C3AFeGwm2opbbNVZpkJ++f3dJ6pZ
tzR5sBGljp1QlZnj5fNjJ5TjL27IvINi6wzLEHr/YeAa4A4VXOGnSUtWXPJbAB4eZxmqWm2ZPmea
EFuE74VNJXuVwEogCKcTNZy9Ay7NjG19ifMps40k0hVeXoUk/17xt4b/uaD6pixahlunbnunBYvF
DKuF08RWW1v6OsVfCYsenrHTN4aZF6ZjSgFcYEKd+jofl///YFAbuDELI/4wN7W6dkprOoSydl1W
2uaf2x/OzB2t68q08+V7scn30nPGWLqtA2fRQ8sPHtGgrsqZcmjawR8aPRZscXdARNTALyZ8OXrv
dqmPQGIDKWPGERzXopbM1UdVapQe2meGxlrAF6r0A2wBGgbr0FIiA2BOX9dCdrNsAnckpMsFIG89
4ETJuih89PIMKi9sEElLclr0xUqc0PTz9h1ahB/Tyv2F5kNSH7Ln9Q52tDwf6dqCNnETt9SkQJK1
qqT7PXWnYSO3Xn+0aF/CJOJPmpMYhrKTPR4E5urR8b6GeP+dt3yi4iwTLmlQh1hN6RpRM4U1fGb7
FYEQaX5L6J1UZT8N836AfNw8t2nS7UVSPXOSJgjMfEzvDxngHHimaz/eWLo/OoXn4JeDL8HK7jXk
Sy0ydDH0GMCTiQuydJzwSrSJbssD7h8++m+XnB3NApu50Pia6jQNnnwV/lK8L1RT3GCnXYLv/phH
wMzyST675yUB82AnotdKGcUORWeD+EuuH2ExvcEcgO65xVBfleyXK0Cz+5rBMC8fqUpr81lvlxaA
jZpttB7QkGkT9CHpHnwHN6cnO4E1uNc2nCYi4iftfNL8MCXxeUkSVpyaymZX3P0yJf2YvzS2NQZQ
2V36UWFTIXvKfIqcnDQENJ8BLuJ9oS+dsqtmab2/wesWLCwfVqqWy4yjIpZfNgHCI2ZX+hRxI/oM
FOpqMreCsqu45JKkUc9Qu2bMuL8Y/Lgz02RIWPJWNLgh1OWV4a58owafhwIXI/v+6HkXL4+COI0C
9GMJMDRRbbTyoWqbUsRs5i9opBj6kw3HeUl2WtlTIWt2wUoyJm2daYgklJ0q0KIHW7RZBQR7qi1X
y2/ZwRoCih+jblIX9TjC8adiMtQ022M9M14zCYp5ZtRZKyfpDJGpIIWDfE8ozWvO/oSvTWjd21t7
xrR40R1DSFkak9YYr4kAK56r4OgYaPD/9HG8Z5xEmMrYn3+tigVv9Hh+zai8wiLxZ/4RB+H/LHHy
DqfueKUJCGaI8nkJYvk20nj5lhPxHZr5cOTD8camaLGhtf3qyG5ZdwKNGVK1IqgmKnqpW8LIVT0+
Zw+Rha6uwIXwS2aNjZtvhScJMqirhm8B6WiqQmrq7lv1adr8sEKvaiBs/6iG/cIj2F1hPYiMUsZZ
pUvQjclJWvVs0NU9gokXRcliRyA2wP2ljEty9WOFp6W7pgble6IwfOKDmueghInPE+5QOB8IoT35
D5osQxqKkbRsDEzQQB4j8FfwmI9Xe2/2fEZPjYsaJVtwzkFER4wIATfNT4oFWkNoEyQyb/7zWPXt
ioY3kb7Jr4mAn0sQ7TzKiZiYGj9pPuE6zQ/+WOdbgRvR5JUccgTmL3nyyvSzY4LobyR/DghHaALH
Mgq9FtN01OPC5Ph3cx6+qIkZkIsDk5kZ8W/igOUC56I0SszdG5OGNHT8Zb0841fpvC0FJvhsXTwR
OqgKefKvkFvJEbq1Whf6ameIziugwl4TCZzRqDslPNdDy4TC1kP2CvXLxMUsv7YobWX4S1pXztTp
8W+ayoB1x5FIiNL9lJWnveD66glNamlffuf3I+WtVXRlk75JPhRam6Q5aainHNE3JMrgPrtndswN
06ZEK50EbuQQEDe9rTSmmVLRpIY5CMiDpW+YCHd5Yy829oIt/+YR/t6Y+QHiARPT/gKmDv7H7CMy
KOBLWsx8qHjlg4fcpRQSJYAx872wn78TNHi1WK2ZgpTcyqCN/aPSOzE71tjiumbfxYNidglykPWV
rBWFcE+pSCkdjEB0HUCB8Gq0hR3X/sAvGGvDz3eBUqVdZm5F3dHWJgKGIm+jeqSxd9ic/i/QhlIv
8LMaJXPCM1X6iSnBawUDVpDtxcB3GLnvkvniNpkJ0wRM5ljOFrGAPIe55srYnvxwbddNfiOF1GYr
qTqRmhNOJ8Pi9wWFdWENBAVmm9hYRxR19Xn5dhsgfDGo681IYm+YTDZIagjrFp4tPPy1TsBvk5UP
TrdWqoPpPhQoXYaT8bB0f2Hq5WJTp5FoUNRPDMjX4z0D0YjlPaKX3eo9GQkAhS6T/MkEtu/T0K7C
Gfri+a7W4Ys/3SR1fYzhlApC7c31fHBES/47bfCtcivcYiv/k+KJ2DGP7dt4laJ68bGxzBphiusR
R2KhA1v1LUe5GSB0EvdK9aZt60zPGYgW4AxYyM13su1ejkweX+5E1nQTNyJAkIjCt/JQtzuGdHav
QtAExnredcd9yqauix7MrULeZgO+5dFXfC3Y/UETGF3A04RObWdcpYkcxLVCjLhxusHjFSGjwilj
Jt4T+t3usYgwOReMEutu3SeeLBCKpjwimyZUEH06Z+Q6ZLsEh78bxH3iCHL/X+IzLdn4TsOZZO1V
WGEC+zropVSSqUJEpZFnE5PZve2qYk0KZ/LfZ98x89Bprl0kchPkT+GKbW4wNXVx8kZJR3Q2+z0x
YJsfwcw3P7MAZhRV33TmOOW61HvxyG4u1GdH6GwlTNgDWl/vaINwF0SBaB4jAmXojfGzem5xGRcB
TGsM/Gz87KHNfhbRL6Kcr/djNq8AbUrbCZGoGRMQq6dfpZsVzx/R29QnsvtGthaPyh+MQsZFpU43
EWv+RTN9+6fQPI+lqfYcXXmu9EewuopNzDnFcCsFv65LX3IwkOz//9TSpZcndTISEFFC82SSBPYA
o6EvMR+3ZoxVZhqgJ+EYrQFBIQoWTKNSB7i2sDWpqXyIZKINsupILd4Z7R8UucAhh3Uxm4D4wFTe
K9N0Ly8C2iAGBWlOAch3cfgZJg0rY//cQ7zIECGx9Nannyat1Y3idX4i2MYtpvxL00GWZtadrP3d
CBAXTxIKPOX0QAI+m4p4622NJ5ElTrDw4lgJWiMVNm97VsbtUfVm2dG1JjDzm3+enC8dlrhE7TQ3
uepIOZqZXXGieb4MP8Q5GpI1DrlJRVbye/1bxv68bzF83r3JOoAZE6NbWA+GbsPnE2LhqbeUlhbu
OCeTVVzPI79iGhYTThNGq+/Fp6Bij98d5tmxYrKbSvOBx9NYQKxKLy5Iz1GjlTmnUE+Q/mhVugTG
iS6rU5Y1LW8ZtA4+qLqGMkHEK9eL87m1GbqonaPz4m/SjjmDwUUXzZp48bBsJQhPO1l0elGMBHn8
Xp4viXyyi9lNpcV9wKhn/0dM1DMeQ92vijXePQ2egHu3CNtiBj02fV3oefi8tWbGzBOekJhnnMQT
Lr9JmJWLf5PquEJ4++yr5BvILhTVFXwFPSiEVH+BaPBOjVJLXKjoz3ojzXlocG8duoe+r5TyenCL
+D2XW8kd3NGHoe4FKcEsekMBhE9jxFcguOQR0mOq6hdPJ3/IIHW7oBmu2tIteceLMIbFZvkJt1bD
hwBEZcfEBCiReJ/YoXYz57H3yMUSeulHeEjszazfKG1E3W1uwLgMQE2OwvJbibk40J7DSU3+HCGb
tF/zBk6J0LMXxjBVXDea2jGjxg9fohUPG15eA5SI21uX5P+BNshEtQmmXC7ufmpsHJ6gBlzvO9xb
l4/zVZY9CB0vCie+Hu9ZMIA+fGVRmDdedwl74hQJz+SVq7IsloKE4YgqG9F9FoASwU5x3e4TJrFv
daTCyyJuib3pvr/NhVtF2AKJOmTJkhXJ6I0NPYW6UqsKC5Lxqs5VdnWT2l3e4LgrdAz1JOmcspTM
BpBjdGtCMuZXWIy2GsL/kZ1tcn1tshP2y1ApIY6+IYXl+gm0rdf4617RwyOs/chdjkxZStwOA9Wf
2m2gRJXRFkE4EglOsODY8+JMLVxotDjQn+/R2ItM7Z/gtoMdHUIDwUUWjNYKe3+oDk6584YBmc5+
5rP4Nja3OpLndTnXSIPrB9ANSKZN7CbH8s6Ad7qcLrXxx4f/zm0yPt2s71x/baIFG0kLe7MaohXz
URgr86xsEai3hgTIP+YcTmiCqRUy1wpzWFzEn2ospLqQM/sLx3VqyGmjYN5EAueJ2XQiv0iZ1yoI
RsCsmrFdDmxbEjbuFdAuXGvIxZPOF2jTToxUoCu6SklX0RdGZEdXzF+4SSiFIle/kHFKGHYJqru+
cgEV1Ne0CmlOcZcJaiY27iRPpCBlY7/BUcjd424w5xTjcQxlkd+WypTgJu1GwwCiu/SgUU3sfHso
O4nachhukR/6kEVJ2CqYUI+KxL8Xz7JLzSTYjAc812uQODIY0GRtkBIBwluIlICdqo2skJjIgjKZ
FEqTUOqctlbV4WA000ocFacRZ7v4uCoLFZRuLYIQgqWoTWqPewMgZWBKmahjHiHBFWJpWeY4ctCx
FRZM+Kh1Po7dz4fbRzFfhZvjVwN0doqvXQnv2/jwlR3meK1O9aPte/26GChrDU+4zU7WLHtgqjpb
z0AFu3ldd42R+gtDgAnytPpV5OU2fOIj10JLVdT9t+mk6drC2SFrcC623fqmfAplUeaJPJH2pH1z
xlZuJJZwupiE/IabZf0oC81itaVHQrT6VsrszU0tma6WMkmH/RpYLpgSHQTtxIfyiXN8R1H7+FKL
NDVgqA7+FzpPISrj8ipBNW8heosP4eqWmbCZB+eRnLN/x+wNC+ok8GHZkHB2YUezzIBIiEGOTy6s
uekYRM6bXEU30ApIgf+kL1oO31pEbpeA2BQZFgIm1OetuMTxuk3E8v+89azb41ivPHiCf8F+9yqk
uW1qdnVZ/m/hURnCvDqFCnCYuN9G3iPRDF6/gjmnoYe3BBJM8vG08IwXVuz96LOHQJ1w7nB+bu/W
iOcXUa6aRiE6SobJW3wy6qeV+YtUfUmtHiVwG8NQyYGyq9hQ1ISabPHlXSBzjRNfWCZFaL/bk1fK
s6vWJpVZ2tXTrJu9VNjSeYHpIUpwhdMRU94B21AiiRucGZ3ZbxYrowlcVl5+5mI5Z4dC20RLKlIZ
uL6D2xcHsTRss10vT7cAIRz/7xEiGEm5z+GY2WuXOGmsgqecjCk5fXPeel10eIk8RauzIxfMHuuB
ZszBxmA+ieHYed45WpgWXhaC8+aVFzxY3tA5rdO1tlLcsAGf0gGqlWlTYfDZ/SZRWjnb2Fquuy1e
HkQGR3jqZZRrqRCw2A9sVjhzXtIjgLHJPxiY1jAUWrMwoIuJq+1OLRvTqYLZD5QsaW8/HRR9Qs7M
I182w1zXwKj+50BRLOOvlqAf/JohgrNIPP6PxcVldjwMuM0ySlTIXAOWJXGgoNj6QpI4h/97e0JB
r+fs55ICu/1OG//Dk563KbXMXRloTHsVRN+k1BVY0AUBEoeH6moxQSrdEjJZDQIO4MuNjSkk283r
FzdwpcSpuwtfFYlConA0fjQKcqUslugLczICPuBPrrERTbPHDO1JBqRLGeoeDq65eV21IS5dAvml
6V60yUo9Dm8NevMwOhgmRjEFIOkOGTAVbwBpQRgxCF1day6PpIxbqATLzYcpHa8RZld1pQWR25tP
ngvJ2vQOGYFBf0JX6CBcHJenxionKhPvZCDCxkiEJNIp8m7JNZEpiOikLunfCw37MOb51W6iTk2F
bZ/VOL53wo/Bb0u8Xb5ZixpLgs2Y+JUKG/38DPv8PZLtV1K20iHU+8+pTUgT+Qf0m4DiFNT0WSx3
DXS1HGBanCDG8IL23H3UKvIRTBsUiywJA2kO1lVPMhYGIU7nW+47mjjg8SLXkH1GtKO1cOFLAhTL
FkoEP157IZAbHFufO8YMeu2iQzzqaCUimBSU8qOJJivjWcthgMWu/DpHF3ldw7yoaohvJi55PNuE
azxO77up5ZnWdUg+KNM5hWng7J3Ul7SnB+t7f3qbZYJM52bH1hm4f9++o/+VzLxQ5BVhP96U7p/Z
EbAZXMiNVeKPY+AABSXUmCB1CNcqL5OqRRcAz5cKQ0Lv/BJw1BXJe2K7zpxF0O50zt+LaDAy2Ihw
a3aodYevgvbIX3EmKKTsH8c8r02cnwgpEZPJq7M0MegXIx3jowXAymFGSyypuGYanOul8xwVyGG7
sjbSkXMb5mg3vVmUIjFhlRRT6+BFryp8X0sj6tkMT7ME9/BLW3Vc4IDpaFFFdbHeDQRH6PLL8JFS
Zf48OcZtzSywNucFPm18vpRMXGO72EUGi2XnpXGXkTlatjcx043bTwmgfd7/UnaxYLhHmcZGvBGk
g75mozH7lZ7cNJAVhzRN6a6WM4yL7gyAXl6zaDvvO48xU8E86rDtNVle1Sq2JC4GRZPLjkm1ttWv
bKiOtAZ+WcxykuQJqVkVSmbE+vJUDdSPyh53dHGkVWQAYVK/7I7nIBWMN2/j56cFs9YKTFi5EJ/O
AWPikWQ+GrwqaSyV9wEvantK2gxx5gOiY76LYbEHt6VIh9Q2TAs4JMdJp44h5C5bprKtrcl9oSzw
9WCCPHyzzRD4/LkA22IFdnbl57IhOoz1hNtHpAHeIHRx0+U5vRQ5fcZXCXdLZB5/i5pe+D9c3Dj9
ICE+ukB5jDFCwNutsyClCbfu2Q4DUAzfjb4g90f82IiGs2sGomySPYzzANLdR49t5Ufd4qiqszQS
tCeGt0p5jwHTNXhNOBPwrByIeqWpTg6ZGML/sGz+cLwqhaOMwfpbqTCp/FfJRpwPwWnO8PPSnt1B
SPeNypv2j5Cu0VsWadF0Esy5oQZHgvd2A3vpSm7jmhlnEL8qjiosnTz6DGywYRPQaNQsKTm54pNe
l+L3uXdJZeR93hf72TXuVMURv5sPyy1AkZJ8yOaBDbwq9DctRRHlM4nnjRRMW58iLPF4tPMiRnGz
/tpP5uz/LE/GNsdbI40DkVAH+Mb7AeVPnBFoOQ753wxgSSQtaHhzsppdw5Bev0SW2JbneFibIT7I
4jlIYGtRjKoWCf/IfwzGt1nF9a0rmuwwZAUAt2HOIo32G45j1CAjhCVkKOWQvadfcweUJxYHGioO
+48M7Xz1p//BAKxgSrew20tFMVnH6qcKnmoo4HklWzmn8YsL4KEEvL1DHVxmB24lk7hsZUefZ6Zb
cCyjSgS8mwQgMBVl6BhrtcJWoJMMs2f2NL3dDsAOmzwUDQGEJhnnk20NdgZpQfrQUysNcYiaRNQ6
nAtkUVZo3xHIlbT02y0WEbkuqIrKZxJSA+pkUiXcy5/E1LhcbWIf4N3SAiTg7mqBpS71x2sVZq2i
UdFFcUzOf4mTd6CZ8VibdsGrfYr3ioXPSmmKSEpYCq9V01uwk0DhyamvlHNSoDzZuPPs7/nRxiBB
jMhD5Zvgcb7RjoMn3UWdKp4D5LBq+omp883qGY6eIUBZ6nYMUmAyTXHWsF208Mr7KLLLu4hsYPNi
zreyU5juOLlcIM0yMQdkD5pJCDyAzyWxDwdPOxpQu4l/k7znYymvw4+PtZb+7sSN+bRcTEBFJYMW
RwPulY9OoF2mi/V0WoOZFN2Um/RwKiY3zo5TbS8rZU7isP8yNTIvgNSnybTLcAjmCAEUZq3zX58r
7u7hT8vsY5vRt/gMNufIlHWgmxEVOv1JYror0yF8SumWPrDFXUmDp1tvXUMIlYUmYriqlhvzL94r
tly5KC5oqkSDQNJDwrw66cyjl4O6hMtKnuikcIONpHgBNf1+oZjFzgkY6VPJf1rB0u7FzqtjbVUJ
6KhIzeHVFj9KtGS7V4iRgxrowh/rSmjhu3om1EDQL1+G+HZz7JAmLSj/P8PaFLChuBE3LxvKLXpI
iS8xYdcJ6vNLkeStzUFJiGTi4s5V1TMuh2N7i99VSZpQNQq3LpnkX2qr4mq7xAkkD0+ws45woYNV
jb+7dKgZiWYwM8Xpgh+R8g0lqmYGwWTCfYZYbOnE2hRws4rXhLseRnW6LSJcydf/ss145MhyDmaZ
J5DPf37RcDXyAIat53Ij6qoy4Ok3Zq1mFCz8mT45mw1rJXXdPd9cWZeuLG3HwSmzWUENRU4fd/eN
0Gy7KjFyrkaahvxG4XLGwmnuo9x4/uDRzJKZuihYB3WRbrg6t0STChi0PoRek95ZapjxgqrXLwTF
90zmI5AfcB2DAHJFhPHE+6OsGplH2KvRwq1MtOyqQkAsq00hW9gGdbwJ1R6DypP+Yn9RAtupsy+w
Dy7PbpD5wMUuxuthlUKN7ZqICg7QWX5d9n5nG6jwO+XyfTKB2W7Of4AWSc7UiMSasaufSxQlu8u/
AtQLONVajZpFkXm5wLgt8mmtSdqkNbH+B7W1l+UuFJVnc4kCnmt6bU/aB02BHQki2zBTwZ//0pT0
UpTtNr3Siq36yLTQ2ttktMTBI44POh3kvC6hhSyzpL2yskvIgUcuJEQwO0QFEu4F6UB4CPmDTlC2
Bv18bLBdfux/TNYBAWkTzSrFTX27atZpyN7gyYr3GllnYxYXfuntbs8qkhufSCH5EVDzMNuLozQZ
IUw+uvKGk+BFev+BELC406T8zu+X05wEFy/DnQVHrtIZa/q4e/MU7tBa4so93OUpEEFLBLJdhBNW
zbGLF26SLZpx/gY8WbdkMEOHL6IBqSRm8rEXSHKla7rcocXKOoXf0AUROdzCieC5clva+/V5dm+W
RMrYLiuwYkPScekN0qzGo9B3FvNkeJKSrH72xy3pQRS57S4BaS+2thdXFed2dTIB9Mti2nTo4Ww/
N3cZjjmqEulQ6HDzcFPKrUBSHZX6NfXn0OdnhvPdN89Iqrq1qTVzCabqgoPgwCGhlqov2t6wk5kP
4nDz7o63Z1uWn4yQ1mwlR31oEyHHefn9vAGiDAWU0sBkSHMmTNNfo63YT26JPmyNsotjdNCowwCT
FjtDPvpwuE5hxB5W8gdSBS6spAgSdTp8VHgTaB2KxrJcjlo6h+7M2ILNJ2SVIh8txuxviX3bWuBz
YORO0+Ta+HNSvJyZy1R1/0844IKWQVQBfXzjC+iEsj8CPvJ5TpoEhMRQdlA7gqb4jHw+414oMj30
4lVAYTfPreorH3/c18PB+CvleeW8R1ol7A0eD29t2p3/RSg+FLfWHZ09YTp8uCTOadR6ZSriroaz
nt8F6/nCsw4veUSDmldQg23A+1Bn0D9pkQ11wr4RYzwbVlDXZVH1g+SPkq+hkwofn/Hz1llOYhMO
G/gmwRVorFD38gLVXRTHUhZfVMGkhO7saGxflf64eG4kNe3YstCOix6uzT8R9NcKCliix+95TEmB
sUjGdt+JE1UK2OLV9KxDGX/t3VhMLxAMOt79aO2SQcSC7UeT/HvGPe5jX9KF9j9KrI7ccgZv6Qv0
UTquTeYNO8jbBLi6USUsvNOhh6dgkkWMwiVMHqojhxu8M288e3EEyCuh+QXZGpH+9SGwlERyGVQR
VzUJpz67evyyu+4tIKwooPYRXtrLZxq1Dum/LPWFKtylK16rec52JQlRlzHSibGsT2jMevRquslD
per13dpwGFnu4irU2KweSaz9JR78oRT7BlD87U84/DOzVfasWesxgRvRERnCwSmguB4e9okJokDJ
Bkdbr1k9tGLgnhetNJmAqx9nzGOkQAZCUh0Peyonohfuk/QGalbehu3KgNOAPgmU+FE3Xf1W+vQb
gn8QYhfAv3F4wx8PoUKVB2u787/PTm+8SgCtXt14k75ABQIPDr/nIy1f/FeABqrH6As8L/iDoguY
gx+ie3AYap7Ef+dM0CLHzbRaaJ9UlB/QwxXl6QjV7C17PHc+UC/B7kH6Zz4Gvtzo6QFlVYTkH6TZ
kppy3Au+Ii0Usyfm99TIzTkvsb9MCpbI4A1tDDYbkr/3OMn4B+TN0EHqSu6mqzZByPel5o5D5dHF
L9w5Wcv8OP4M40k6epojModzXWxsxy1Asz/dnCDaZFklo7PuBMlLm1wt6UaAwtjIgpXmPeJ4E+LL
DUfh4vROvOBc9DXxNss700zh5lT4nPlpIfbhdQcIii1/iphpb62wr8Gca0OjwxYM3dzt7HORCuY4
fl7AaX6Su7QajSEmTzuXTq3GTBxObigcP3IAMANTm08gKF2auD5KcROOzfifkDF2GXJmS09u3mrK
WYqwb//NpGPcwrAKIhSca0+foyKfzFuRGqkJZUnXTG121l92KXoMDpdvq5YQHt5Y2Iw9zGAA3c46
Dxv+CER2MY1HcUS8k6MSTJk7h6npb8yjIMr0D9zDphrqHmvvDtXyns4aQr6SatlA4cKQwcxymMXh
zN+awL06JX3IHzTeQefiFUqLlhWwMjPhCMCKo2HGOuRwd8k2esHelRGCq+xG54dm26exrEtCdDn8
4TYdHlBHyN1U1D/uawejmptStwC7Z48WaGtdUqgxt+8E2luNbybsxPWf5WrVlhgWn2u4Ez10MXS2
a6J99rGkvqk+YbhZU9is+Jnv182vjdcoThwLTVG2jB4teKiO/Gv3UbgA9FQtWBp/OsgUt+W9lwpF
BnL3ZjqcTF226t0L3eO1GDEFhEK2FKsXWCvPTLBRKWX8qwHEKtp/7/pYxwgHx4X0GCCgHgBzm0B+
6hG2YtZp1fP7UQ4GJKOQJ7AGWEnLUbUJuJ1Og6IQqolmLz14HITtOWGzHm6ArhGs/iXc+/69e00/
fYHJLHST39zQ8Ldl0GbSBEK2iGP283PQS4LVLmPQZWGSZih5PX2R6wpkSKFUt3cwDActjqzFz95r
cxv3RY9HRl+zTqxpVkELChq+iEW26kwwNuOp/5iWkOGjkXorT4xJEM4os2fGidrskd9qO+TuaonC
sXl3Ua+dvuM3ZoRzq7ky4fCtzxc6X5WKlx8VNfgFQkHLMbdNf1uLkpE9swcckfHmRJ+js7b/SY2W
WwTryzUYiVoXLflr+YBQeKdafQQIxkmdhnGtxUu4KC9NHVoIDBWkTxGn67q/vdUCUG3SEtN1c6S1
sIZHA8F8zNh3CeMatN/OZojGeDvkvECRmQRy2IOKNiId0HxgVcQmgYrue289xuDxSr8yVQchlU1e
3Owg1uEu1FRVZV7UGggnst2NQ94mzjNCz05TqvaczeHoZjvUpl1ysP9r5RvIhsTetK2Wme3CSqgr
enqMDZxakVWLAs3Y+B4SUPUL2Xv+iTBPDv9b0OVfQb1JPuQXW980s0FX0fsPvxnOKb5jBn8e1kjx
1xkU6dDc0S1ftiJrgx4Nr+Rf9GiuhUaq4p9bsra9jAPIPrqV+AfschrGXyyMzEKXgweIDCxys6lx
YBAziHBgw0ouAM9reCmmRAcCau9Sz3FY8+RYqwrCc5NckYWqpe1qZqQ+3//wXqnS5WEkMm3Zml1R
34B1PmO0hJtFom8y+OkFRJAmOpM9sRw6ry9dOW7muC7UGO1UyaAVDv3mKe0DeSDIk3A0/EUTLx74
CckaR73dD0HYvrZeS4nQeRycmVO56XViIp2HvMFLEKp40k9dInAHjm//YEoBJPWodWHMgL87JJfT
ny0sYlyZqnPBDYJcyMynnObhvxC3YQshmwWlq3LM8fga2rRzgpezT/heKxnUvmjJgs4y5dhHMi36
7Q56fHN+qOtZN0+Ne0NMOQCxQAZak6cetSoxdpNrjHoejTmD5BE4crK+uyFbHSgb+tS+oORUTnWm
bZ0tuGKxGQtiGQ90/tLEnuzAE+TJr+yotRt1iErly+cGDfdri5j2nUGo8y1xL9sBmJ+S8p1lywQh
Xjg7Kvg667iRXf8QC7RXRRVjD+RP8IBgNe4f8P3cRLj8iLcsm1xTEv7A1Lxi4OCNlsPZtb3Rb9Sv
gAq+KcoRaNkjYQ6KCSC8TrzznsX5rjEN92KAWSj6knAv2iACqOyH8g56iyZxuwIPO2thV1eUMgu/
DD6VfUBn2u8bT12KBH0nVERWRMcOBwy8t+KNUGygvwQyB01SKBNt/3+0BckGFlNi8NjCIviP+gVq
kJhV7nLclhilCXR+6J1Sh4th0pbKHzjjtXZj8gEStELx/aPed1hL3lEMbpcv+OO0Fvot47TOuU/T
rKnHGSs4kv6JTi/Q5++15jVJLOFEkShojBHMlLWVDO2aMH8hUdM17sjN9yerTPgtyz/h315cpzei
ezWw7hLpVhx3XGrGh9Onvmlw6d7/GWa0CtsHvCyJ9WVpB7BdtR7pKXUrFWWSOahgWdz00b9USfBN
pXioR4qIBDlueFemGpSJvOyWuEWNFWDJo4FRD+0rvFWi6DaBkjTlRN5H7M6CiHCG1nua7zO2rGML
ofLs2BNBSACnB3EzroWGdVteOuSgtuESOIztvkbp99SuXBBWaNVvWbi2TMtsvJA8wp3IUjMDA1b8
5sQ251fuwd7qfHIHg89CU2r/wK/YE6LDDagu12UUSjKfumyfqFGBb4Tr5TgBwkZ5BL44+fRTMsI5
mero0QHgpEZAejTaoik4qwBb9aWCGGvCtC/sjLVvF0qgDeZpfb81pjxccU1IRyTJb/n+h9pq3eJG
hqzizQQSeKNbeFzj9SHiS5uC+eL0yDQfa8O5YeWv+3+oWy7HrkR9MC1+9PUe4q/jG8UCQ6Y5rq7G
hrkQhHmKUQeIumJTDKgT6IJUMx3FvapEBTrgEZc9J356pbF+XI0T+FvKgi4mQzRlNKxLVa8HJ61X
J8O4wpZ3fPtEdk+wWy7h2GuxnGujuYN9DEfPJ+pKfGAplVDN9sdVBY5OpFjLUwYAKF/h6QQ1kj/e
kWtsoTCKlSjstbodtHc2apRrF3in2w1jtpWm1JS6ZFP5blNoe6osFA8mWtKbTt/uzPrpGWCOxjuI
jElTdJ8SATgdE/xKC0Fy0O0/6Btxi6r4VkmM36Ed85Z6Fj5DnYEthIaBtHx7+3vQq+sL1HFsXzT+
aLDxOn3lNCVEnwUMRCulDOOmQDw14A9505ri+aEO1yQH+JWFv70ItqUjVfjX/H91blA7FsvD/sU0
FgB7WBCD6DJwPCSBYDMIrb05kFhQS2VVL5H78WX1zSmpAzo1K4S5ovD6Tm/8GccL1L7+fQ5PrNNa
fw9Hq8iIWW9KTYDOJ1ye+aRCS/0zCH3mpiFheOIiIMvwvLWd7o16+MfnzjioiQzXDQXVPoR9GcB0
qcZB9w+co7sDnQ1LL6hA0kQ/qpGcSth1Uj6yqi5Ye9MNvLXaenQSqX4XLgOBqCMabE+Oc59+mPGq
Hy6oNZ6538wea2NKUkL7bSJsbR5n2HENB/mEnzuZNwYySTMQe34UxqVox0QGBsagulXLL+Ec00D8
aND1rj3E/LxXxdwL/PH244+R3nBdFq2Vu0hjQeefBff2/Wj68B+99k9lVo71rm/cmfv3pYs4jUrY
bMtJvUd+54jRc50Lu0YGkc7qNJ7VktfQFTmze0T4yuYopEkK8Obvhkce5DGq5r0DIw9v9PDUi60R
tLKJNCSm5MPQReVzLimP32To9YbeQv6wNgXNqMlGdPdIzZSODzBoUkVgBpU8n7mE7Xh74Gm9xlYm
Od6aSvSD7ETWmInK3capdzEyLCaRMT2aueRF6uLQ5WjBnMraHv5mlk2Aoubcj02OaepSxdZewrE7
D6lgG4YH+DoIZLLki0YuaVXhyD3b8rBrufxToHbHqHDcQd9WvSHm6jASpuouhdHP31Ne/YylqiU0
OUMl/0bjAg/+UNCrXWqb+EOjbv9QPp+JA2b3+QGI7EQFNDV7x6/lfkT/NBd7vk2v3/Nz4uRzKN5K
T71Oop8zC6M9jA9mCtQIAjLYoIK5LttpeB3Z8+VKHagw46BIVjkTbrj11wnt240nHc42aZ8xsFj8
VZtx63q9p00/wzpw7POZNG13+7I056oicKd+ymxhXESBRtxVRvTBaqIwcvTzeFldPN7/9tbtQ+MO
uvTYe/KBCyEUJjeXhzs7ac4FJsjhqBMKdA7pcuWfB1mTyvAd/Zotru2JEK0EEIXe8IdCYInM66iv
osvTv4IIr/g40Lnk9Q++CBOGw/gbokeE7k+2WYMRcpS5R4WFEsbAdSoztf5lp6JwTVFlbC6Ki1m5
Hr8b047Gblgao9khc1FgMM5WMzONJJ9ENzNtBOSaLdSl/0LzbvTvDK5IP5ptMVb+yLTA2+9oY0VZ
mSI09I3j7EJHXkE4eHXSB4rduiheih3Q4/VdcB4/E88XAqt2tzr19jBTVbrvBJavCuUYiAKD0vZt
He6lJoDd/pzDU8G2lI6ws8GFDTXmOo+Js0vtPgWFnJPVUoLah0ZowUiwX1o9fG1bVh83m8J3OgnD
ENygH8HTfxnAWLxkNhcvbHN5uoWs1pPb3NQnl8Lq50Ga5bYexSaa8O3yPhk/szrAIIn/zIRioEcg
V4b8lhtgQzuwniDHv5sRmlWlIi5M/vs7zwukDp5v46sFiGCpQ/AwdOo2kqo8e5OA5skmsZFPCMlH
fPQ7yQ4PHzHO5RZvd9n/M+SIJ1jFB8X6J0E6yhGnuheEXyL7dngaD7vRbUGGjiVXp74YoK61S3l7
2zl0BdViN36bFYFNuUrvSRgoPkaielI9Q1/fFZUT7LZQQyATJS+r0TbO0rNscNThjFPCdurnlJBq
CkNr/w3uc8y0YL37sd5Iap77B/SqSDwQlx6W664IrZ02BDMdsSnx7HZwdxQcd1rLDvh2/Mjfrzmn
RE+X7x/SN+EZwjBVjBM4DvviVoGc81VHvcJix78xWaXXczd5CGVHCKLfab2P2v/l+KMkD3A6D8+r
Fn/r6815qSMnipmNBracJ6phohYgR+WOZIgPwu0kLlyTAhXN7uIHPXevRVwx2jlTikPH8i3+o/FJ
V/cEbIw9Ds297YVE0PEUKlSc7Vx01edqnq62dzBJxgCxzx7gWhth4v6hQDNi0UUzdMXxZzL3qdDw
RZ77U0CIYjLr0568PloOSXvej2GOQ+vOuv6ri6ZmtHgdeNOn5MLPzU69XBoa6b3cHwMwZU0AfNIV
y8DjXgSdrMC6zC4/zSk71HOE310Rm1EiI2b5crQHsdw4LqcoE1HSd0Y2uPva5lqYJflojb+EjhPs
M8XhiJF16weiY0qWKg/ZFYnDr20z4sDiGrLxN6sNiJvqrcDnNk8Kj32m7KVjDwMxWT4YMtmyDdUo
Inv5DGF4CC58OeVd+qXflQaCTGfpvz/aSEStnUewgDZYd1Ksb2Y38VGyWm7zHJfPJ4aJxxpMe87S
hDQxoAdEzCdzRlFHlB3hjczJ5DQ8XkotC6QKlIlGdDM3jna3wL4FIp13fpJgcQOrjUoZAXlwErFJ
R3YChFn9JxEQ3vLSUoIm8fG5e51+MA1P4SNkJLdEpOOpI+8LOF404wDSqAZuMXkBECTaUNhmugsj
UY77oEGkbYYhS7uDQLbrod798xU2SYw5+mkvMLGqSHsU927cEDtSox7KP12YuRTdBQ65fMX3UZDG
jQxeFnPw4LgVX1Uv8LxJGmwm830S2dTClqpa2naPyKozzGvQdIo3fjhC413NxBwaSURbvymipSwz
CRsYCUUHbjDEXAderAyVBs6I8UUGrWtLdZ3bSISgpMgoEt+3fZYdrtGKROc60WMQr/z89tVoNeRA
hV4g8tiYxIaTEWxT3NLm3lGemJ18xPkzjz2Uj0GtNnt6RWbLyUTnBd2ROhOd9IFLgU/SeRQa0EEW
UXiPxK1wQzgWtYFe9Y0aEly8rUqT6i7Tk7XVp4Z8fJ91xPpdCpkVte8WJJFKt6q/6DU0KS5RIaOP
9VG4ZZcCeoeYRhIpgls63gk38tgq0ERh09qwYH/3fitdIvdj0/PwqDpRr7E7uF+yx2onTQ6DIkOn
AshP2TN1a1yr9RpQSxErSHCYcZO54ZL411lnI3mPLmTGLrEgW7nfr4piwZnnQko5LBc26PdKqFSp
FDPEZk9CGUGYFLk3cj5gSrwEQ6NTqPX60lu1F0zkxSahRidFRt06fHx3ZjOXan2W6ZrttuQRc4tS
/T/Ek7v+1UlAkxaAMTftv31BYgy4SlNfpR7CUROcbNcsGDzOZZJE82t6jqClmenFiWhj/kyO+cvA
kcZ7agjh51Y5w9Pl66EMc7qxZI2sGJEUDZ4uUSuyAECsH1T04eAxsqXhMwnPBhlgw3jOnfw5bD6C
Fm7szF6f1PR9KgeYDYha0+17LeykwHmU2ENJXYNaX46SijtpCkUBK9RucT3VDHN0ybT3exdcmuFB
ZRkDZAeBIbP+OlHa+vhvnoUrUE6Pl/JbRjf4NjvsL1JLiRcHPPNo8U5nwCCEiil5ZsCQEFUJmeTA
Yjiba58JELDoff7eUJfsxZn3NrBO2fQVMK6TKyun0IV0QlvDYJdThSMRK6fJUG+EFOZoILwhGaVR
rzldSk0+u0hP4LXjnQv3YyELpcebVZhzpHaQSmOu18t+2xifjB68Z7j/UJx49AZyHT97jw+J0hNq
EBuEgUAl0YEepWj1YaqhNnx8/p9L3uRdy2tdI0YyE/YCIQ6zYNAcmTEvtyQvpZa76A9aWX+vhj4X
CpjN3Y6KEba0sMzS6F4lmc2VUtbdwC5CcrYseyxZPB0yDRxPvGmknJmqDSBWkhtjzrffHdJiUNGs
+Z32UQNI8IKm3T17cymBx15a3zdsQ5gQDv1xBBCO+EoHfSAvNmEjVXjaZ7EoKsEMKs66J+RTyiYO
BcL468SHqyRPGOHApj/q/qy/OS+3YrvO9cTTUdqy65fWQwTfZe+EXkbu3XX1f07g2tn17+kejy74
OduHQ+fQGbqQxxC/2k7pRhtkv1/M0jFeheAUC9+x7ScemzVQMXd5dV65fEa3v9mWNHFpDNzup49e
QLjGU6+jyLMvWtUAdcNSAFhWap//fUtWcdY8ra9obQdbU/UhqfVm0oKrqHdACVZt6m5Kv+Zgj0d1
Lmy/9mpLlgeuvpPEdPQ/ZNSnFfCUh53zJ8LCM91YhqaU9EOj85SuS9TkQdKeLblyugFz7oVAhU4h
eZID+3db0ilHlQs7s/1jqudBj5cqi1MwEJT9IBrfGuZWWKfXUl6oUB1cAi8U7HBH8SqGtGU3oC8f
Dgjj0nGkEjLDdnYUcM8W6LBXUU+GpNj3EVxJNYnVxRomSW2y4v2sYOQnK4xvY2uYfGiLO72syEiv
I3vJFjHfXwkozk5crTU6Ml3P9RZRgtCxkPfOvpL26oQ13gcrHGxV9zAfYyxWpeRcRiOWX2/SQCth
lrRvyDmsacp/T3nxkDqamVsP6/gaAzdylyBoeg6XnsUqXihwH2Ivm09BGHXZuUUEDXBkACEeHKIW
ixQQc5E9JZV54AuxTC1jG/DYk2BH78d9aHHh11FUKil5F5bpj1GUHn0wZYcyMlNM+x+P35GDGqaj
lRE2HIamY2AR1OqUZ9ceat9khmq6rTpgqBnvWjuHumMM/EtscSNCUN9rDjVAg8HovqKeJW5yiV7p
YtkgYVcjkROGCwJo1bIBDu7Dk28pJQDWCSm5uSF8v1JAOnnNJCruWr4IlYFR/Ea8Xemzw2/l7YkB
Dgbs/G8OxGF7eQCCI4NsMJYaSXUFX9nDqsAJN423CGWRGR3H8ADrZcAzvKJmIvQ7vOaiDMIquqHk
+mT1SfLlOJ9gNAnQRLPnBQZIiO1bwJSmb3+h3oBPfH4NcARdDTwFIY4bTvMr5KxBQDS4kbY4j8J3
WICZDtXBEXfMygMeYLwXaLsxbctNULIMZLU4wEcJEclrZLxgfQRDOFlDq1d4r1SbJ+OeW7aj1vs/
7o2gicl7j+vQQKJIctDQSfYFXQx4h9vfjBSTPAc2KOts+IidoX/1pzc9Xbdzd2v8wIAY1f4ioxHW
2kqT9uZc2ArRp0RwfqKsZZChzpx+u5V/xVvrmqPoZ79cmQJz77AP2ZZ/xCDYEwMGDago6NeRpsR+
Cch/Nm8Wkalxwrjdd40fxErDHeatZ5lHrlRn+zUWuRHZGtHeNoFHxEmiJG/IwtOVc9ky6CpvWSWJ
TeLmvAX84pRlEfoYUXS+jzElvX11sOXEpUlsNTv4P9lvDxF6SLkbp2Z4vGzEteynZXenxp2Pw511
z/ZzxgyGAPivs8jUZYjI8PMKbvX3N2JAsXs9DERCxO0nPbt0Oo9rYCNrq/G3QZFY5Bi8XfTMzjT/
zj+TdwIGk/SgT4uyIMQejXQ/25muOOl9+ABBwuWY38FqcnT2u7A94aWZPsGJ+RhwbuG4kZz+851f
F+3eSk/HFdkup+BB9CW4I7trzOxLBYvRYyKv5FB6KWIJ5olpfr8l8ZODF+yr5LKtcVyrCaJZ9OfF
aybwJy29GAaZDvA6u6xULokdGKkQlNRhbmADcVGCKZcGbIr3N8ojtX+xClcuAs8CKHbR3fVWdcWQ
z1GA+7q8Z5Ohqdp9VJ+tVAnAIpYFiJp3yerCPUSbsUhsutYeQ2Rul4Ao0dcnlWER5Ul2fingasj1
pTXKZOIIKF1rF/ki/HSu8QCG2c31BucGEdaUzRl497ZSk3H88POG6FvXWXmSIk1cwhndQxbDbGDG
j0FaHGr6+gI99gnIqvSUpqgVYHjvN6L2ocTmUWcuzqZfYwQZFOUJmEnhLMTndHhyQLP52mTGDH8A
aOftPRmrCtwL7WquGhP0xuk2hTqk1ZsTE90PSzzolSmaquW9C+7yQj4w4/btfVYRiWGPV7BoaSiN
P73cmwIBMne8AKv1a24K4lfmoH3+VtQ61jVpMHFOTaF4TQfrkF0aLBnUhgqpZGouwb4gbqd5x3zF
BuxNNBmQwnYmRK8Wl2ineRnsAcbfDrBt9IfMYc0hHexJvvY13BY55EDJueoFRVKjBk2FW5DvmmF3
N9unZayEZKL6+tOtfuBGOLboMytD+ZFO25XUL7bnkzST3g7YBNJj6Yo558D5eBvh4gECFAVMnvqJ
R/PZLSM7fcgSTafrKawU3ooTCZRzyj5FzMET26JplM3qPkf+KW5VAI/xEQYSw07Y/7X4EF5lFIhL
nBqe9KEOBIBDAflQt9+PEXf+LX4YIYWt17F7ie/+/h2e8JUqVlfgsfgquWtiID8FOaXOfp/S+nr/
uretAb1xkK0MOkIQHCpcvlWbJ12RyXUMyykBtmQDb+i2ghBtuo8bJp8w4gfN+ZRCrXGxZ9LpfdxM
U8bmldVly/F5jtEJDJopeDi9FAAWfcaJ1kxqyG4tcQO/weXqpVAyml+u4BlDm/j/GMO5At9l9eMd
ixNhylKKs8njgEkOMp1rr30UFC2KH76rKYJY0EBNbzTUICn+AWJis+hFazD4ARWAbpFzyXsnAdV+
5w5EIJcC7vlEnOkw0dV9vl7RByZFX/hpWoPmrGq5ObxwoyXXNtxB4S6y5b7mZIpDEIkX+68Hm53D
IP9Uf3PXBo92NmUzQjOSq9XbuDoGNpxOtWDLsTKfSwftm2seGik9YV+uTdBhQE6DDe7sLq4Ed2XI
/7/8FNIFj/b4nNGHD80AwrYbsYlvgjBZgKXsA22oEJk6p4AieJgWe/JUAhzTfmkVvHbJ84mU3ITp
2OdNj4EoQwCzTIVUw/rnsaJd9IYh3TudRKEibvoufdEl+AdjnLGON3xj0cePcvTI1gaiHJFgt7vn
U4e4LyCP8NtBSiWFleIQcX2LzCLw16wMGsbKIBww8RN8WrI0ZTPuqkv/vobAKrwxwpv/ffq1UW08
SjjyoAejq27j3K1jk3ErSdFFVfmEJxep6KA5Ja/FQy8o0V4QiGpeSSiJmIrhkfOJypx2KCoYsuGb
Ncj3BRIxaFYPScv8Mb9K1gncU/CdcapFnoud8S4RfMDs6vBUBpnuaTJ6m+2dAaKfcqjFMyLUm54P
8fIPVhxMe6wkb2gWpW0XJCJ4u6EWv0898jtpWjW++ACdNYofRiXbWj64lqg2hBkd1Z3xA+kw0RMU
oY8se6QRdVo6lQ0RQpAhz0XrFM3sQ6rmNADl9FyT/GPwV9Dq1usOxKEnYRhlp7yY78YWwH1omGEl
23cmJx2mLc05ffagE/hQg4pcTqW0HspftGFk3or6l8sHWk2HusmjJ7kv75MTlR5jwPyMxitmZzNb
JocZAmarfJfYR6J5LX5xG1YgXbqG96gpD3Xy0FfsZwH81DWX+kZ1zFrLpZXlMUaGO4xoYkvb0FAp
5voJimsiL3T64FhrXoTLq1C6iHRxTk/0fk8me1qo4IS8xIUTG9S2aAjvXMMVqnynoOGhcdqoz2YQ
jmQEVPo1Qp1SdeClQMNVCnUdzsDNsNXrm7DShdx3D/tQd189oJ7c5KQTREcPp/+tMe6wx81qhRnn
ne6dG5FoaeOpe+VB5OR6d1drmeO8QaXnxPGLdeiEnBWvxcJssQEAJL99R22e2XM/NjPEKkMdIOM2
+w5bF6S5e4Hy4yZzke6tudJBBXPGW5iDZ68ffkzoDaadvNuKkgg+vPDT04yU6vKjvXZNW8pEOT8m
2CjM9i7VFRP/DdKgWfcVwBs91x251yI34T+3T54GxlnKqz/VeJaeAAK4APnxwqgDnI2sVGzThh2V
knN6z7/ZXBVgAofayeUG+8p9VIuEHDRjME7VjPhFjYPtvbnzIFwmO9fFIm2fUXufejJDanGA7px+
88VY7l0Yf0bXH9E82l7urNo16kCB5/XR7bJG8OsCmiCJlX21osqcm5HpFzqZOyIlFpJDFuA1yj2j
2GgukhWFiETXWYm1LLeGf3L3jxJtKVqHyNmc5jnzmqDnU3Kc3i8iDbG/EOOC6aoJd0hf5VicPQPy
mCcUxYt9ILewVmN+D4iLXyu6AO9UGInQJLpZK1JT99k/+v4CUH6QjADDgN1cm17vv0Cy2N5wJIhe
yNDR+cryw6p3D3bYWmPkf1eBZoWKq0ZkWb5Mx561m2hSSAtrg1JjfwsTWI0CyZOJQ+WgefLAAl6N
VjCFzfS5k03GFmI7kp0NhBoNyVlFE5V4v1b7h++Drm0zNY1sRNWgsFnfedal+0wyTxWEJc5wHFa0
V/OQgGiNMjZQe4SeouCLJ+JviYKJ3D4QiLscU3R8eLHajpuERflTc+pjF4FXfYvYTJ3ejSm3IQm3
PLu7DOfJw09AQh82a0Zlg4npYP1uKhRyzPrFbPz4KADYOc4Z+XIyBfQ/EynhZwbZrLYWihn9S9lT
5Yj/bTNay1I02Bgv1fcRu7hY1/adkcaJzBAxt4Miv8ruP8jtjJZcZc8/NB5Lcz6Lgs3J3u6oTDgi
ti0mpchApWb/+4jbbEp6PBGP/GIx9wMmiYE4BeIqhJy9itFu5yxAG8DiCMrKzFk2dKIa0/WeGUgv
NuWmZYSBlt2xEJmY3ZioVh0scpy8uv2i1OD86NOfIVPMmm+sk+u6uQTLv5OstWx4MrKEy62R+FbP
HCdPzC6OT9w2ufE6EpIVb5iF1BHnAAF9/s+QX20ZXA2JsPKiNhemJ6nQljzJQmAf/i7YBiNwF1LD
jEYBOSSucX7zjuXEImPIE1gb4sqeo3ATfYB1fHkJ0gW+EcnnYYCa2hgeVAjWT75u8zibfqqBz+3b
20zKswdCsK0fag3f8J5SM1scmqSAOPGihdoGVnDTtyC4ofbOXR40UxzrlKfk7f8Uz0uDbwlmbmHM
K8rbgsq+/dskjYtORMUTenLL65QNrAK3+gZ2lZF9OQzyjP7vkHrnCScNG8CzNm7UagIpmH6KoGmc
CwUs+ZK/cTxxCKxH/N6R3dca8XwVZVoCkXojgAmv9d1N1B9+qZiFANcs+81Z9SISzZNTfhIPZOCg
z5HKGAYg5b1CDDCPQ2e8qJoJ4e1VTQgbzHeQqn0vwmeG0Ui3wfU5pyJobeJ+QsD4Jx9AP7cFe25G
n+Cc7ylSLFsLUMKNJVuE58xUHeoxK3JU1YUYy3XjgKzNzSGkXAgMBohS5uyLJXY0/l1UGjAMMwX/
jFwUaEw/D8WQo1C6UwNK8XL9HFsePiLvHoCifJBsvGXbypHDP/dveeOumqBPZiCUR7NwLHakVEeC
yaCx1uQaCcbtwatMgTMzPrhtX2q+rHgwacY/NltJ0tSkFOMPm/ILHdL+VDAHK3UmARweDAENB1rx
YCUZjdRaKjIZaZcIc2KmHCSGSZ8UMlbbntDhNWPsfmDrJ3RiK/6qa/5EO0jJ5jltB9tUG/TW9LiM
2Mz0QsCk7SRddUxv/rAeqLZ8830QoHEq/C6bwdyHE2m0eef43cDmLBfC41OAwC3W/1jnr70SGQqz
G0SJCZHUyS8D9dwKrYHs83erV28HRq/koFJXhAPLEYjh8kjdpOoTd1yQ+UXAK4qJZGGOXF/0AVOI
X/HqraMx7ucvqGjSdJiAxdiCUy2a/Y2bvQnRMO6a0a4TmEqRy+mRomtwgM4fDFzCAQE9vmSPMIuB
PW/y/omRbmi12rYFWA198uARd/1N9YYgpxsFd3uRBA4SfyrWj+Me4T+n7+pJ2CoHYOVheLGGjW50
GnsPGDlHpnfqdYYnqI67Z3UOXrNGiQKdacTFdSXAJdFrjG5SX4AW9lILSsJm7DK1rsTNnH2wZFDi
9FQ6vP+KBCYWR6IEVJZVt6nS38SA9oyjdTFwhIgJNk3e7Ka/G7LVzAfBKssd/IEwZz2fSxCf+Lem
shImzI4QABSRkXVu7CNblz0a+brxE0AZMj0m0mKBN5t4a9jXmOuHctEV4fT1Nttg2t0eLtMOuW6N
XIra7DeDcyzqBZUMXXC+Xyivsp5HA2wOPykS8kw8pRjHW0LUCH01HZ98mX325EbjiaK/vSBjFmai
KshWnG2Xfb3+DWROyrH9/nLb9LgE/uLD4jMjzrAC1PNqqILMWbykx6HSCqIFeKMAZOth1AsCN/rQ
3F5g+v4vZbLp7MhFK6IqtEeIPVwM3cvELdSFkAfWuSPU2GK9SQvfQlJrtFfUJwu33nLPdogck3of
oTP6iO2eIStbjpmM+bXwOYjF4asWO5Mp7DQCy/+1LWJvV/wOAY7SWIEwxQiZQWDQEAbkE9BQjnwz
0IqAvaFg79Zp3fOuNGt8sKmyJLDpSCnL5jPvA2oJmlkJnQ7dkpGRzXECD5T32dx0zPi/pXr5c0Gr
lSvJdvPwDm7fIrhfv1wIOACtiAbJN5HnDlr0NAcIgoIEyqb66aAalDtfOXCfnLQI+a4QmWzaDHw4
cbntPmfbVMMmMzQTqLEZyWfpO1ezipz5/r8Pusv+91nZdKTy9cmppw1en9oqhd9NyIv8d8vNA72X
XLEHIjX3bE3KlmttXw2CJI9V0YWdbrEHGLvRAMfBqI4OS8xVzxYP8yf/5wDPn+lqvxzsYDwPdET5
7ui87HX8O2uRLy/n3V+oANyw0GhXgarHHvPqNNASit54G6E+ePqLkBt4dy0liaDTpBov0+iOwHfk
XuRglVZoTMlep7wR8KDT7mY/7WtvSpqutp2gbdMhyI5yhuPKjXH7rjjo47u21cr4E4h9NbW2Frzb
PvCVY+lB8raaA4i1tFu7vHVQMC5wmLkUSLGTZgeu1Vt8AGrhlyyYJamEGv6dmRdj8U7tgeLp2bKj
cjVYJmiyzGE9ShP/vkHXb7v9ECCEnV2mm2C7sr6Yo6EMdbVdS2MBSnjfxFb9veSj93xGjWrv4HX6
1Eja9ea8tdbnfbjuRS2VZAnPgmnmKHWkVZraxdZzBDqLZKvKCL2EOzzAJ+D1IknEH4lfEJGQUTXk
9TYweuan/DJmtyZHeuaAnqtfMAXWgkl9BOLSqiTlA/NyQPEME/bjQonrAPXEvGzQseOfkEgDj/Ss
N33mG5YNWD6+V2BB4i/RaUZyKAT9/mQppOh4MX+fLensLe9jgsFYA33xoE3izAnrXqhGVE2ncjg8
CAe0XohEfUGN/epVp016otgiwwEHnjvyRo9Zw9Zsea5nhw7hfcb5dqHsdcfh5pGewpjIqR60z0qp
L+s32zr6tVatjWkjpXiixYvdgCGlZlRQ4Oc+aHAnPfu98IlBB0FW/s3PzgJLN8hiQLZaA0+eBtUi
3G7kZkuVUq0fCg74s1H+lBt4R1I+pZ6Fzf08NbtPWstDVbcmpmdo/EbOHydtQq7PSauJZoROK8J4
C+9B+w6sL2+55+N7LN0G6vDtLwDTLz7LmAecboKSU2U0JvahcBWKTA8tv+9MOS0uxlV2UfuN3V61
4HdDvSBhN3s2E6VyKwlSwiR+n5DR2GRIV89CiA2fQhSWwEkbP3PwFbLoE9wuzbfRrvAbGnKqRgyM
mpazo6ZQE3dHR4JINw4hdrn5FTvwzhfqWExBwzTSbD9gj5sxBvIobLclW8uFvxNZqqDxUH3Ew823
vvFrYdWHxK05qVWbIoYOV7ZHDi9MykDGzrfYAGHjUl7Vdg3+dJmAYknUEWZyl28xP+xD+S7Lopi7
bGeL/juFMrZhKSU35b/DA9SksS51Yljknefpg040tOaf33eZFRxY+3Vcftt/oFKRkPwKRB6C1kO4
ZD1Pxp3co55g2SvOqe0vSSKj7Nt4JP7OxKhK5KKIa//rn8NVgQw5Ddr83N2/ETrANouFQIwj/B5t
QSoVbe1T4JqDEzmIOi1Z+jNEaZvyYk+SMekXfDSDaq1z/9C9y+IrCSwxueAtMqMnas9ykzTJj0E/
TagsD1axlB/z95N0+JJ6+XV8t4PSSp2LUD3bxFYgxQK0LNMJDNs1fevfEVOvpu6h5O5SX4WALZYl
fC+3RgdMsFZs+KDhi4iA2CG4Z7CvD401qv16I5spST/EPTw3ff6ZNaQSnNAT/XUP0S1cBx5Dy0cx
OfcmgYd82dROQ6zmhzFuNBfIlgu5mUb5Vo+W/SdNmuqUYeZi1H8r23novbOKuEIFNvo60dwcEdAh
vowXBs5Qh2iMwn92WnAWwnwvOyhyD1FmDpj9IKmlgwzgfxv72+civ/iXGefFPLsE5KJDktte4AQa
JCcvYpcPmfEPwHwcO8T2t4UpbgS3vtVYoNGDmsnNVJ5s/m9Mb0QMf/RpSoveZbZKwUZUxHEaHYBr
STO3BxiHEvTBURCICFljjbE9wcfNjYooJhLYTH273bJrog2JTJo3aVjKA9DtRHy3M715zkdwfwna
7nyNGRz5upL4TT86ODK//UbYGFQq56H8mDiOV4BDWyHok9VtWzRS+gmCljpQszlSnzDvq2tDVEK9
t9vHW0/CmAV33kUn8i1OxF2mArJRIJuuFHC0zyklAmQYnP5BsgHHrdst9+5FnD8QpEV8dDS5FhEV
QqsxQuKvVTVQU1MntYq6JlD5G7NS0hlnXSQRXHN9nuG0RBtH8SdzpFaQ+mCzhg2Zpwn83YRU6sgK
gmhgjKUmVxLi5p/VtsencAzEeWuBzeLOJxcSw4lAoS+BkYdTPinsIBAgWTqCBC7x1mUW4Cq/xjS1
PqaYvPqZbbsSaNZPxUJohmKZW52l+doTaTEyh9zGZjK/lShqNhL5FCSkeMNymArX27MkaI5/fzJ4
YoI2rviAx3zPygMN2KypYoVOe7jNGkFllTFO1885b/GTKnUBNZKO6bU7H7dXVEk/3n2XmUQciSsd
EOVWhYCHp1K01J86W9AnZ88oDY6V10I3zDpM8lLffU3R/35e8moiwzVg4di1gjSTGDx8IdQw2Nbd
E4kfkWyz3ySh4/rKiLK5doW/1s9cOmrIEvha/8fZD6zVYGNe+rj6fq8ti8WXhmxu6ZUi+5Di7L7K
eaApnjOI1zA5GvxKfTV2px0Vmc4GXeoZYP3j8orUvNTiRX8Bvv6oi2pZd792GI9XrEFWyWGPKa7s
r7l3RNhAJD2GkeFjyoNDziFcoyKyEmC0R/rGpMZ7wLzrV6czkQOMfRVFjx0loHyfjZnQQRLg46ML
vHokuuuUK/6yxxV93mfSEn6TLEpcM4s/IlAwMxWP5f4vD0me5JMd8kKgbi2RSZKlKrmbkUX7SZLV
iwb78AGNvpydmjQAdIihsMANaARHxBKcKF2Xc/Qfdz21eJLgQA0dBoVMZdrOk7A4/2KkncJhaYP3
SEoqj4xip3U3zJgPWWCe2sxL4hkpjQhdNGEZCj+prcc5QaQPBDHIEUBQtif87MnqYWZCNPAkP/Oz
BacgCxVQcHmMQcpVle1li6itIOXc4dp34f4XKjxH8f2LIZo6sbZfYVHUzcmEHf0HBb34p7FOu/qu
5IDGOZvDDUI5m4dAztggHQs8X6VcAA3IwjVKdxVl8EB4YGPBxIO9ok7KMXqucrTP3f/UrmXOCsuK
6n6cagZaPjUEvmiIicnc0kHTnveCiAM7LtBB5t6D68z9vqBaSGNqqwN80CX6whmOGL4DAeqR2F8+
xIOOAzqc1GVPfhz/eZYUsGAfRMmVccmKhI8WJ18LvK52xT5I/UwNDNJVW5mrnyAipP4nmc7QqQ1x
BrKzOX5LpcXU4uAkErG4i8I6qvnQ4VHVJUTtqXE97wEnOqEp8SPtswOWMzI5zCkRnJqEx4xH4PgL
pnhsyfANZTOyRH1rYTFYggVhnmbP4C5zldf3RXDNGkG9x5UYe6499gAun+UyXBiiuegPL6V7kwSb
HcJIJuJvyV7lpRSGJBcw0BB2/NeMZbhXAWifFVGAkq6s1S0BSyuHHA56rq63e/FUcTLU3ptKDqRO
ZGZEkbciU+OLcU1BtZ31UPTemCFyGtM+pCobj8Edg4IWxfyqPoGVKKdR8Z7arbRxN/d6RnjyOWBE
MSWFVRDbZ3lUYLy+Rv7FOtWUV4bpxv4/sYh1EbITseD1ww0cKCaqTeNu6PDo/ZhumGBBEJURCcNj
k217yNoyNTIpU45jnfy8g4r8lRy+jXHmK3MeDc6+lqeKvp01mVIgSjfOWGgCxu4ANr/NN3eZinak
5BjYjLmDCmkQhcd/nVHeBXpslRR6W4D3W0E2Hinc4gpzsqINqEMdGehixjO1Zkkw3jgcNcS+smxA
hXn3CzcUOrA17LjgGviHC8rnG9l1FXlONP4flXlwvl+BUna8+r962WlNcsp9O9XHL+2wkLQVSfAQ
8gbqOdjILVdzZrNqQBchDJLbs/dVD4urJbvJohmFOuvxnZG0I64gT0ox+kQb7r1iGIz4sYSSUVe+
m+49qb1FHdMIWx57uBpCXf+gNZsicf25buMrXzXOBUGjDH9KdoVTxgcQDMZf4yGoy3Q1PWFvj+q7
gc5WGBVyZgVmEVDel/voC+THE/f/AQvlfVZrJuHiV90TFNDeRGxUfTr8XizOBh2fmRc9f3XdhSNy
JCz5pK0zsBw3S6tLFbbkCg5O2lMUq4/I1j+b7hOeoewoNQieNSUkict7MGt/wKx+9GWwp0YH4W1c
e1b9jO/gSUUn7GqkOo+6cnJ/No9zDhdXy5MGpiSBa57f2yqWYra4MNKq02cBcYtQaCMGlTEyKJpJ
m9lIWqElGk4/GCv7tMfmmwb7mH/P6/0SRVzCtNBYuHYJSjez9zW5DK3ZLl3hJxs1S/Et7LlH0+hQ
yJywA23thCY6C7897nSoDt0gLvSc/GbNaij5MXTaBOe5Zg5t7R+OnZwQfwONtjQuNjIMwEcw8Tkk
MB2cc68feSg+kLGsVaIWoyvpgs2ChRz4V0dPGFCBfQThSYTrEg9Evmrs2+9igddvPEg3A9AUpVok
I1BzOGCh+svvX3APHto28JkXr8+jDH4eoMgd+DeVei8Fa/SlhQ8blNAyN8IuVaUx0xGnV8Z3Q6e5
OiNKMjmYbqiawgGvg/ZlTd2RERC7V49ZWku3btEYL7aY6a6kyEEuw5NpcmzK0hD5m4RGszp7u/xG
CV0fiBdhIz0OKB0wSsY24eNB/ShS1Ny8faRLpP4IPYw2k99Kzd6zEAc/wr4ZQdoZ6U7EXC7WZZ42
RsUYnHs2nWSMsebVxV+HlilBTBCei872UdJaP+9FiIDzDSJe0DuwuU91j1Rj/MCD5itr/l7HJhEZ
xE5YIQlbxty9K7jNQq9/8z0KMVXkc7vuPDQ3VD4iXiPZRaxiY+Dr8Sm0GUe9dykKoUdnQPl5l2tK
MBhrIAQajZLNXZ+2O8Qj8zbA5uUSR1YQJJnwLg/5qjaj81Ya4IOg7auwBSnLBZaYAdzz4ycsDCtY
BmmReFOvyjRXLwVNOlwkbwSdjTazVPJhDCcCdhynbI2tWgxtqglA2cHXKSMnHdovF7QqqE7qW0/0
nlR4Zg4dw3beypHmvfsUZLjNGHT4+sKMP2b8+m7pljKhVop5cMGUhGSUTZqR0ttOQgSizjESroPB
CuEQmwgFWW9H4e705ShTjOvRMCMWm+3nxmLQDm5ykoY3JaPgLyfT86Fgg2zkzjzFtCJR6uwAAp1L
5DmjkrRjzBMOp7FqiIagGwMSvuWVafvv5ZkFG5Eq49GtSx2INFGIZ0xY0Zwuw+iJQMBdR4KGicwn
goGxiJjuF7nXMFWwRA9/8dzYqqyVnl2Zdo97/LmEwKK9tkjV9MtX4ICZCYqL7v4Pbh80MQnULPC1
c+trxCRYfMd0dWhUg74g0XufCV4dqzkJWN+7RIQ7Zmrh4zNFpm2yPmlt/JU9w5Y2nocydR+znAn7
OkttOSufHk+ILsQr+H0JkOAZENrbocmr1jQYmdsSifb/CeKrCCbjHLuyBe3d3bk98VBmlXg1IWlq
bIwr5YfIGEJBle6imhwON3l5q81U22oCu/0lrfb3M8UCWY76aiVJoJBkVpTWFyzMtvh90aRY94b5
6gicwB4E/iw4TLkwY+H3NsdxeT+8n/upwSLhgMOgwSuLtyTuVJPNfcL1oEbbgkcRLKNad4/7hLly
0VZKGvbIUyO/gA+AhWaeLQB5UXUrzbE0s8/x8N5fQO0xILKZoLp9S0nz5A1Y0M7nldZrc00nsueZ
ocvbVoTnSkRvaa0Hknxp5TNk5YsCqnSUKUtz5OJ5BPIu5+t1S0F42pB2kNESc1lSmlCbvVwTp4d1
h8uaIcx42/hVZEA1N/UwlT6Cgw5NjDzltAFOO9ApQnjlK5jC6Jril9KTt62ziBQJZHiNcrZBP1vj
vVK7HhA5pi7DgNiBrwLame0deZgHv9vsknawku8tzMKfkzLkOimj76QrRLQJ6jA1BYrNYp1AACyZ
U1GPWI7K1QNZnOdmb6bfy5maUNY95anVpIPENlqpeYgBpsu+BNxuF5el0bvSp7QXR1U3r/abxZhM
1xCEoPfKndbT9VESHiTIp6D/XcZRD4wUvwu8J6lVORSz92sqWfrdh0PtnsKB5yn8oZiXfVeLDGrh
F9+bjYu5BciQvZaOvEcXa1oWu6Z/Q0YsE+J1oV6TLxcUShIy3+h/jgaNbcLTa8jHE8/fKoKeOpGl
EL3FZ72cwSUWRRw8aDtxXO+ZMj6r9qwj5ryUvnITNUPnXN713H6UbzgxkXQ20LCMTlPEABO+WqPl
Xrmk2cqQUfAhGyIClHiIslU/V8diV1I4uV7lGZzAQ2di/JAbH9EG84WSRoqjTbrqzDtRzEE9NeXN
8uzpCOFtF6+Z7ZdKFApMSwjZ3rwUUSgR8IVae2zT7ACnYxpv0Dcg5MIewkx/IZe3BiWdLT6YM9Sl
90F8KQEADvVFA5qHMUQJkT2rfrYbYuBlZkXENXKzhxwQP4QnhoXAaPag8lgU37g5dwDvOjFBcq3Z
7aRHcMglYAFeGbfojnxLGC9dBbO8/zhzikq0oZ0oWwzlaei1+PXu32gFQ0e5Nh5h1NJiuLkTS/5W
9Oo3aY6zfD0ucEyTEsaoqWpwD+XcBk95kor0d1aSgJQcZYZw/KVCIoikFMA3Xo4E/GEc9z2AQ+6l
qe9bG01/bmADPr9o9KEIgqhsVG9aOOkmUclkMBkJ8JylMgSWWLp5L8XkvLz8BRcZ5A1mUqtcNkY5
fPGF9M0xItZFQ39+8FeKYUd2YarCDH8dPsf+S9l3fzjCAA0iWD1nLF6AiGlDKfo8sXyfonpj/+fD
PAn5Hw9MrmScM/2n6nq03ydNxr3Dc2Z0UbmQXsPbtyU17qwP0nDhIYhxr8/rgsC8VEBLYRrUEypt
zZVWcGKipXph32jDRi4Iyc8/WJFpNMZkCcjsNEoGVr4CrfXs9WBMJFq4WBN6A9deLlMTrPoMdaCU
gGgBdPjOl5Ili0lTZon5k16dPLwyAG5W6Ngu2xOfvXOC9Z926t1aucZUqk65ze//hwqwZibzEggF
YsAksV+TnRH0XU4cYRA4dU8jDv6yns9nRon37WSR7dTXG/G2VUwVRNkXTeoHBKhbFccnDOsQM77K
8x6i1fsGqGml06AxFarNATqbNKqQyd13CmUCApmDMnL3WEnEHVBeyg9adC+8FozTVtqcorlXpbxf
n3CJU3Y68QdYGgQyIewf3o5RbRORG4aqqDpo0Lk+oO35mcKvVzGP5WKwBqfvb5fNVYOaBzUSlPdS
4jwUskQuYMQV8OSoEFDL8uMQucanpucj3Pinzpt28+YZgy7VPspIQg64UKCsfbjdgoRiY8SlEuT3
oNwY2uQc8I9az1W/1FGa83WuAt5Ln6FGMD5MXHAQzJXKA+0cD3Spb401A/BIdDCxF+HSd98OVIfJ
jfrhhTgYcA+74t1SMbcMNhnlBr30AdFqLQUnwHIoOQisqgqZAAG9E5YNho/ZzzkyVhdoHX7nqxhU
4UiTMrJ0PYKEV1dBOtMfci9CRBPuDWrc9JNgwIrA7oIO2kbzmh5Sl+wo760R8KtMLeVD12z6kNYN
HxLYHv/cwoApUNIEznIUrgbhSE8TCmxU3V7FEB+5J+a2MGwXeNsHGGIfnflVggV+uJzJ2CpHjw9v
JZjoABms6kXw3LyxJlV6Hp4RXy/KW3Y8aoK7Pyd+ZNDihr5ubAYUPqsoNce9TrZwLQHiocBNz64w
viX1x39lpDvayF6uteMjv0sBUSwW902cDl4btcMyU6l7tQgqaMbIQrUFAZZGsUB0nY08GImDImaJ
4JTjIOdBJ0vEqem2WTdTRjL0uUtBpHzQ71tEvXMEyYs0m+kwS2mgA3EPWHX8okiR5UNJ1oZvaq78
5R0FN6cZQ0lSig8l0IIA5H1ggytV1YndLDPnUX7DvpvM/ZPoAHrglBGGuYEe6jttPvqn75wIGg5n
sGeBE1RrargSyhV/KWW/lXJTTzn1fEhVHQ7IDbE31x+hfSJQ03TvfsKdI2CA7ipxb/oB1GQRnmSM
YjaeKCs5YEZPc+bQ6q2fc3D8tSbuOv3Q8wguJgQC563UGwH7gI2k1ivOfnuihcCXdkUxFdWXB1K9
d87T6z+4aM2SWIX9dJ2mCLytDK2NSnfBJnUED19+ptnyTXBHCkwEInt9q0yau3jTaGPTj3ELc6HR
+aG+JgZeJtMyhicktNX/JRmZFLw6qCCUJ0fE3x7S5R4e7G3gSzm7zDNHJroKoVCv0t+W3K/kQVVg
DY/PwviivnOe7R8BWr1Qxsz830hzBL0wEJfM4lBc8JOylJY8B1tHHtG4ZiwWtjQDzY5gBqY4kRjP
OBmcyL3ir+wnxZMhGTronacA3dqTGUTaKLGjhfCfQhL4YSGUTj5okEXGPVsCLjHRBmcWygFGynjZ
YtRkDxaFan2CC5M/c4KpX3XLGYZd1iJHzTfL5Xk2upcAD8j6TJB7OHFIGis1PABBnjXf6Lk5+Yz8
L7I6D7eeCcabltIcLvsGrcnrAaS7dGVpSk/1a9uYe8zE+87T6cHajOcsq1QuEfnORsvUvrxnF/2E
dlQmzBzzyccoPAmRWPshKh9CEh6vC3vXkidRMTjAXaSvOX5x0BVqWzjNlZBvSmmamB1oyI40ohDS
CbowuMBFU8fUdGJKKrc9l6/vkEd2pBNpI9kmwdsVDkMk00FcI4aeZbGblzJcs+WJyxaDjMo4+CFK
pNUbBIj/Ytp1opTfmnru+4Ery1cCRBD6ktQZtUC+Tk8rgA1DdHQIy9257olzOKZSbHLl+G5Er3xI
1GF2RcPcxT6JB/h3Lz1bY3aNwHeuOmFNSMseqDMe3KD5AgAA/1pSmW4lM5IN+oDa9znzejFzvmUn
kecraR4fxBzfkU7GYZQGNm63tCQP7HYqiuueccd6WhLgm+Zv85My4Xai57k2uyDH3X1Qc8gkv5Yz
kqfMU+JaN1q1+ykJz0dTBpXnphm9I+GRH4IuhYKBa8fHa9I75PvS9iUmYUGPru6+BgiDUuOZXw0k
gI3fMCQZkQVPaMXsuZINFFuMtl5SiHDF5he4S9mBlgdlH+5U54Di+lgvGpemtCjEUyW5frmK6Zq1
BNsRqeBVfi5pPcGBsrDXlwGy+5NjEN80E39KP+cFvnnFadIHBBTnS59GBdvB+VvEQpOHagHRQ+iV
ne+86sjw6VDJVBiSMyrpQkzKB62q22VUtlYPAdeSgUdqX8X2C7J4F+xURV5qQZAGo7oj3n4Sx1+H
2H5APQIjcZJgLvVIxxcY2ljJv0rpJOsu/qxRo7sxtDIwvovGuh5yYZwkMQuUdIJYiPErGh0g4f7J
jrV3GL9Do2f/bhmsocVYG1ewQMszcNneBHhCFcdffvmtGLAzScIOisCGG6VoXVel0qSdj6qVLGlH
A1/Bv0VeVvq+L6X/k6RbJevLNHNrwpghwLZByu6hWCG6a1YztfXRaARW2b/IiBq2OPKfnBzYk+R/
Q4Ln2NwLqrJRHHEVT0tXrMFTQHYwDYya9jrFUReav50osHLGgOcrgEEJGW8DzdEPHVwcLKBJwXgC
A8vnG2hOVRNY27EcCHqFqPatCyUAQvegl8Mi9vyRy9oSnflMI6dtPxHw3JHSr3GurFPskmJhax/t
F6yfJB0nr/fq+FG55peOAR/ez3nlzDhQfr4+NqiIci3HCHMOgmyuQfpPcqXW7LYGPnSiljvtG3Kg
jsRqpucXNL07iAP7ji22BvfZ4Kk+LIOE6WEYbp4zlwhuZldoQWnqHx+6ytNFOnacJn6wrPyH2Iq0
kzCadIrkYUbYyVmHQRPT1tE15mZMts55rLyfa06tDUKnjyBtQFOyn3vsoVEMPFQBzbgdrQK5yA17
WTRautLzwlc+MEM4tIwNe/QsQIq9QQyjmQL2RcOSHEbUfyp0I3wnatuuWqtupLOqFeZ9jh/0cOxp
6FCeOG5I89fOJBZ7Hd4292fztOhHvtl3ec7kdgtd9pdn2UInEi/ELh170hvibPC914DI3055BoT5
Cy/sfkVJ2V49On5LxFYLYtD//RTuIHKazH+c3k+SobgU+kmQF9Vjf1M+TqY83ZJJOSr6T20ErQwa
3Wo2msK3h9jXFKYEmiH14OUGfeHcCTZ4DfzjNMnOetuLsbUBYOT+72h0iH2oDsw90HH20O8oj5QZ
mFlji10LGE3qRqTwGhjLJ8N1ntt9Q3yOiK2MrjRDwreLAMihDdOWeHCn7Yqx6xNIFixHK9M/u4YL
JhROjt+lb7KinvdIoPRC3elkvOzyDbkCWLQZIR3CXnbmXjeDPNuluylKy4v1e/F38k5gxVS43xVe
xLTQG37mNkdIeDymuw1ytHZ3qnFMqZkEqcNQhe+ilAArTaf2De4PztkAF8KlrL/Sm31ee+zMueyg
nS+QdOdEB5V/mCKFEgW+m4uSpb0l0vO5nkspWpuYuhpJ1IJCzzyxMpJo2uZbDmCy0ecu7BZ2X/If
75FMwU1a/GVzTCyDsGMBfGk8ffY53BtB9Zk7/aT0//YaqJFmlkqPEr/4ebErVDkvNbVFCDc2FdmC
1ksPx81IYd6ZI1F/ca2s5peyi8ASnhy2QYt8m9sVtGu5H3t55E4UlChSEas+6SMCz1AcAsUpmMcp
sYJPY6ewT6E17HeleFo7/UsyIVzc5frOelujjQMmAPMJAQNgxQy97mMFZP0w+vZL6GlGVzT4UYXP
WsHD/aBC+isYUfO5OM9ZFD91quP2go210MW2lfyQU07pPP3uqtrmqBkhDD0F9bH/v2fjoPzMSBDj
2qJxLPjxe6riB0hdibDOjN8evXp31lgScvOyr/ahowwuVExN3VcQRdVjKTETHVJrIT+qTxuFNRg9
jZla+UVMw/xkj1ceSpBCwxcL17yUpOoiV5IJ2S742avCSlVzJOaUoh7wF2PrPgWottYKk1rpVe5B
EPccazrT1OFC6f3oo/sLVycNJsc4OYZJJJqMnPZFI8tcqCPIvsGtb95T5jNUQ4bLTFV/LNoU76wZ
7JqchKmfu5F51UmsJvqXnbLX8k/bH/+3tUb1TJyRKGQ1PV9LPxyzXTRO/W3vrFHRaaqtp0FYOD3j
0D2d6dvbl9K84h0AT2BVwOwIHKw+TBnm+E7iOXkfNic1DJQ7EdvqU/R/+NSi/GZSJEp3iyajZBen
fCG5mzBsvzokIvH6/aqd+LCT3DJKPdclkjXFNJV+sbG+Oe1r8dOFQyClmK+Wa2hOYsd3kSNawF8G
Ruz8+3tDP77JALMI48zg+RJ3Bo66GesnwZlgZgk365hOLK//tvaFV8BQ5ZK39EVwMDpSOE3n3KOo
7gu793Uzplz+GYmtk9Eg+OFANnuutdasqUCDU9KMU9A7ql55QC71WuKaTA+JtHnCrJRSTtGk4uz7
SSro3evuvqTTSQXfj/edujvYYTRcoBGiMa/MZBkW1s+s3e+WUIqxR5R1eTzhsOEutwmGaBEvcuts
R7nhsFtEPt/SH6YCR4xknCE274kZPHR0Pg09IjwniPac8jHjilknTkbdxAJAMZVuZQQ+LYTDQkfW
SHIdvCJ7hUuVd+hRGzTPbue/KZgmSfSKKTOSKZEeMzI5K2XpvIJPPNYptZaQCkZvriiIrWjhog7j
YOmFUCFn63OEIwJRT7di4IPsZifYPwbf9hX3MwO/TaApNlKJ6SLZ1nwqZggVgaT6oXUQfEizdBfn
z+3gyFLBw9AcpdVpph2qYFcoYhbcoPsDtso48Wwr17PKZW5yd8e93LacnT3F5EeeBkMD5YwMvJ9c
tPW+82nryj5RhXrtQBmBj4Val1PDgAEyYMS7fc6jfhxu74MT1y0SIF0yJC2vszmONkfmaTH2ENho
QNMASX1gfHT1V0YClChtZM7atU+R/+ltHjTLT5pJs8jCANfKAbt1BsO2dH5o9OQrRqcV9RtEz5Bl
EQykXhY6dbPaNpyKygvchTk2llFn4sTVduz2gSG9Hi8Gso/Ir8phZrYZGldcj7JsBMjvWEwSy6H9
1YpF22wlEmUNGHZaSzA9M+E8XimgALRtRI2EnF2XQ2PcZrjUxp+HLKUvCMLTdFEkJ27KwFdnwuKP
wwOfXQAtHYNagRp7Dl9LR6gd4c6U3YDXqiv8bqROXWvNCcr3TPamHBYjkcb1qc6/9RqJdiyIUebc
Ge5JOenaV1+l7WJAT6jOue1sJt6cM5FQdsh1HqpcJMN0MAK8Okf6KNxZfvuh1P7pjn5NjbmCCE2Y
KbHJbUShphd5KlD8eO+t/1UOJ3m2/6IZPgL8k5SMTbJtlMxWAfqPsaz4adB+lVj0ZVeCoWjFEf6P
fWUrt3H9QpqI/BlvdUJ/Rh5oragcWToa6jJ26u6MUR+6VSRgkZQ9PQFztrisdh/52CC5wygHjf/3
u69Q08RKiJVG8BWeTi6oLuzWNt7h9FI4AMYxc+x8xwcI9ZLzDXQ6c+wDeEvTSKzOODc4McscZkKS
U21ZMnL+yaMVc7ZeK4YiBjWzHh56it5kT41kCbOYwYn52nGpCPk9FbA1LPYeXBcGR9nqyC1HWbUc
q3jC7nU17wkAVQbQFr3od76b2dp6NljLG+vbRV43BN139FLNBibKlpIC/Zwk2R+DZCBC13Jq06pV
CO5qKHg7oG5XipTyYU07iiRMvA9CSaSk5VhDZA2NgFoM3T+RDzIeQ3rdn40RbYuzR0wZHQhIT3Sj
an3TO9aekVFckmKT0LbHiMD+M1gyccp82TDUYatR4iQtgxo2PP2OPHb1a/MIoex29QjXNeA6SYE8
lgEJ7sOsFcWdQlYxfafYcLCa+VunbLZ/Z08jJo86ICZ9yl+3HuHZD/c8GEoW8q7QINAyEQIIMftf
isr4HXN53uQ1z1KgTXfxs55mlljkJvN5WOalPvKebq6zhQP8dKbya1Q0UJJvGxUq9lzoVrWeBpQF
E1jjZwO2dqrHAlZhXcG5BIdlcS1n2AWhBo/WLSi+Y19acdBoI3kUWeDPNHJHXe/jERNSqDVFtNYN
wK35aUVXzWKcZt+CJsa2Mk0VW79pTCUQ2fNfe3IJThcpvbSupqxeYponYJwYycdzA7WCh41HvbWY
8RC3TzxBcb3Y+5SF9MopKvRD6PBSWyLIi9N9ciT0BnHl5eHQTSiPEAl1fHTtoCFNACgnl+SEdKP/
T+PEuOsPBV1DNpQqqkUlplanV2LMjXVU5uFhBWGWRISBEg0xSiZ+ISMI/1bJxILlGKJbtD2LMBz2
5TBXtBds5Dand7uCdzZzzpFVi8wYkVqDAOYAmV7QUj+FOY9YOcRTTjCpYLtCD75Zy3kzlJGCGFsa
BQAXxaeYh+VvCIDIcQd4e6tzZb5iYaAdJqQTXPr1ZuSU0VCum0PALGWL5LjuWff3p29rTe3VnBOn
mtaDpIm7gpG2igUjC9GB1Vn1NdiGyf4VonscO85DJk6CJRhMLAevgKddJRi68vIxv3Jty75k3rpW
slRooOK3R0IPLk7W7+C4K3JBSgnTk+u1hLov7RBDxfi4dFfO9rfQfc+lf8CP2O13nYy89nrfX2bt
81AoeUEUuXHDXoNE0ua8M80xfh6OtV6CDKUcCqvxzOvYSzN+p6EjKzJdtkYTr8gtPindI7f+0Q9m
HE0HiUvsELZjUAlwIvLgYMizbR9bTkGiH1rvZOECRP5vtKg25++sTTfKq78KizrbbxKteRBnlVSo
7pL22BONb6fzLC2mJJ/2y5fu1APFwSE7h0h6E3Mgw89s/v09d0Hz7ZCVUo7O8EyHQ+4HML34/vHo
DU62dW+ZRe77fUTi+h9MIWwAyj7Qa2NjTNv2jVn3FxnmNxgXT9o2bu01ylp1D150q9Yz2uyFGlHK
7/5TqCFln4cxgRm7wkWfsXlxeq7wm29Hh9s/IWhJ9v4ZdruoZiDnusfOSNhBEJOYnMzXHGr6CzI3
qgjnr6fnkbUArO3W5qNyfwbrM11BB/clfra8J52VKiA6n3M+T39Toi4sSTc7jEHUyOF+QFnP4qVn
3R1NzaNDM7fWyAdb8gxsySHcSoPtNdEklEsaFlZgq89DZzxXl1SIedDFoTm29JCCGf/bR5y0Alba
syGmf7ZgnL5nNwS0cd/t97XXhtXLlhlL6yDT+0gmutDkjAHToJ7ck6yvCyMoDQ0gxpDaSxLta71Z
Vf6vYpPTPUws0hchQ99H7SucTOWB67/7DjK7i/v7cKY+x6Hswmaj38jtgjzcfMRJwwN0YlDjv3lZ
LVEPNHe/BkaxmVlrUOuwabwvc+nsHqG2tl7imqy6PWEanwaxbIGZ1uSeMmxZMWoOgBocY4rJhoQV
6daCi/agdaPPihJ6Bw5JkIaN8cdpK4lcirANCL91GU2wdd8Lnek9lJHmhSiRk2G0kTzw4Q4TgJNB
AkPVWbvRs2beMp8Sgo/FY3b4FxrJz9YAC2yFKMYqTG/npi7E1rx1Rq8jrN9iyjmRNzL385SnjG6Q
Z0Rat7pU/Etuj5yDuBz04yrDMEOZIAgnppFombVNLEbgbi7r+b5vIqcRD1ssKOhBWHfHRq4a6/rv
Gjm/tKscYzt/bwcbZpQ3xoZiydQd40g3jx1mC9xa62gqjUVDVMXOJ9ekt23Dnw3e7Q2FKG2VJ+tO
nRwTlrq0ANPneN+b65nYNFxAL1rZvTzYcLqRo80NC5Q7IC8HUm5HOiUaaMzY5Jzgww97+OEkz2gf
v4Z1XU9k2rSN5Chg0/HB2SKEYnmnMjUxR4NRdJH0FDoMVeBTbVbEVjxM9WzrMrxM5xyExIcf0ftj
5GUR8RCNwR0ClVMIA74wS99mlr/8UoBLLhjemEKl4wfGYSSusxTu041yKf6hUnHVkX3K8DIBIjo1
gAHlhdW5Rx2zvjwmOXD+SZ5j3zo4/AKo7/snzKH25VbmyDTZa9pZfO+9Xz8mrLNvsIXIz1E5f8mr
ats3Obql+zKz26vQ0IfU89e/DOhEq2yVprjXQX+yJXL5NshWOYz2v7h7IfTEtD2YmjZvZArIS623
cz+C7ji3/gS1aG2Hdxm6S59LA0d0V8xYqFK4QskvcqqrZF7J8Wry1ibY3+YhRcn5mzxgRwWLQtxi
qQs+ICU3kVm4Qdl/fo1MYE8ce9XeuqJgIHQQqPHJI6T9GyG8J0PVHmjqhuXm4XBLKlytfHm0uzEP
P4PUe/UVeeJPWqyo0fYYtOg1MTan9PetGQl1UU+yaacyyYWQk5ketuMq+i35sVQFJduQFJAIo/Q4
j87ms6NV5ip4jk9cjoEWTbv1kLdXObzQuIxO7hLERQpVLw836Qvzxo2s1ZLmKCVEwp38YGzAnTe7
u7NJsk1Mi7uNeeWZj3/AQx5cxcB9zsKlVlKVGgW/136mrVR+PubwTksUnpmGQUyO3msAGSzJgggJ
sXCcUqtwwEnY54emRn3J2VEYZAkiN6w6k2qwQpIKVgj/spkMGSMKATYLLAfZP4T1mt9yO+GMxH+3
QKBq+3LDAWPRS1+LrxszOB0EtkUlEkxo5c0VtD+TG7Jm3zVtfR/3WLE5nOn2MEP8QhA75NnhgCqu
IsVB02wecD9SmOnLwWkcUqMp5ilrOx/JM5gP+vYYqQY7o7ZtzskdBojRZPxOEZFl+75wT5pPiYCq
eb+7Sb73c2k9Dxh44Bqvn7ayRPl4RIMJUkRBttQPJYrE660D/4MXGkE2Bp9rmQmvDjaxpX+2rO59
3ZMNN/0uK8xbHDgJRfDHyNEfyeoKXcTGgY3BW1XOnJCDBI/nQB/V6Rc6Os3qwiDorkWvvcAdJf5z
clVoQjJhZdPfoFzyUfKeqboj17OmebjsTWUY6AK4/+hvOwqEKkL28DwNQvwrWW/t0PH+nTGdKFwN
hVuzkppUOBNun/6AKCfWVXLUdZPfy/FC93F+mHiOZK4Xfz1VRBcYgvpEZasYgJzUVaGL1tGYQREa
WlBjiU8l4SBT/GZFIi8A9yuFzhXYiuWS7dyAE/MM+Uf1QP46xGm5zD0dcfvRKob1wBvrJX/ugGH1
vgApm84yGp59XpBOw0HF+Mf0/28mvKTAGeTzrfpokhZNc52bbpb/XIvlaaxfiO9Yp3MAq4mJXfoi
f5E5VxO4VIYzUJaSQVs4/qeyaRPctqsxQDHlyR6VMKpV8h0caQPj3w+bpFB61ztIwW5Hza6trmzs
19MJr9XrnAlSRC88JUeawZ2nwItf8KkCJ17cEbyRfJVCQJDopt7EnOmVLOptRj/oYHih8e6Unqu+
aQzhi3AY5fqeQCEbXD04XD6IFU1nZx4pXh4h2YLr5eWSL/1f/VGRR5hycyIvTiMmSYh5UE0BkaE0
fthj4nXiCgMNz4EQkm3BmkLWkmA2dGEulMbgFqBFO4JASxIksLpzBohMw5LEktdu9nLlNakO3adv
LJZH14NuR8Xsn8vzcDat/LQ5e6VPk6J4FxmLZvQy7Mh7GtTuG2z/eQZZRmsg7BTWZfj7nCM5ngMk
MYnkTDkkS6W+n8vLw/mDdOdk/2wOmTeHxnbowGWffL0cFTs+MLXHEhq8vUG7gCMvl27wJWh9S6DC
wYZDVU1OWzFSuwINIeqz7dScuzhukGfzdSA32N0gDBv7QiQNZRhnQ+ohsA6QwgUzROnMVxngatzP
LhnMQFsZ2CQN1fA9x7lj0O+v4zySCJAtEqpY2b1hbk80rqmvDGt1h0BoGtsR4NgQ2474hpljPppG
L2hHWR3/kOQmTlTt0p3RRutlFgtc6J+C+jeGtPwVMAmmXw8IxEarSAIaKlIJOTx6qiJM2hOej5NT
84BHg0r8jjwiGMVanbJtMKtIh9/YJWBPnYtGjmQcMOGFaM3SnOWE7Xxmd76mFca+/zhi3hRa1TCq
3n/fxcKLUBx5mACaYPF44kjZIiYN58k/3pjv3QmfsAmFGRbrCzixXbncpmGMpC+4yOGUvV2FmvTi
cXHt5EAq6Yy4P974vYz4ZIpLmK2HDTRmdkc3lbkm40kkQ0nE1hPFHYhldA+gBKKjRYGssC8S9RUt
0phOPgJP9Ef80IFxbHGZ2fYV5eEHgMfDE8d4jjy8en9EakYTJTq5iq3kfMVTHCdHqWVkgy0DFQKQ
iQVZYUXsZlBUMeptTMMO1LVXb8pvFoqeGIslFIR6KceAlTp2bIDhsCxE1WjUwyuLK6Y7QUAQY5o8
fiTPRjxTNVdfKB9h+ypGqYeciIjmGGypstGkBZsAFfmXyXPqzUPHlbYJYD4+CDGriDGOWaVQsJzs
mhbV3rx/H6YWz/GYPYMPq41xEg8pk8HuJmV0DQ7HhA6eS97BnQpEt+Cqwg//eB8ssJBZJeDGWTCn
wBnx0Z4NP8Ah/cHXqzfZ7Z/tSmxQ9brKVBh/nvjYXL1XVae6REPiIViRTXeRNOn3CBdjWKNP2rhQ
paKISvJZERtYOPYAXdpWKjHTFMRhhiRrjuGLz1m0dcFz1H1zxdYT4lBkIFx84c3qrd+/IV7JTWAV
n4WVGApT73/ZxJsOjVinC50UEiMQMr7l4+GugQHJOgaIrBajec4tiCfC7OhWy9+j7fx7g2QySCQX
F6ZC0gz8pNP3butoTnEpVkWpL/PqTojmsVjYCRiUEHYiqw7XihxZcFGUKAVNtn74sMTJDnx/ZWtw
c2kJKVdoK238wwr9Xgzx8hPdFDCmF7QgAP7Xt4MkU7FLvh0fSkGpPSEs2ENnsXyRq4Lia4oIs9xC
JQ2FkH78bqL87VskJFIMpdKBbPk5X0ZG0FvciI/QXOxLApGr/eCg7k5uZ9p+bGYLoIlePwiCyqWE
i9YualBfdtb1W0gie6aNoZpDHOlia6zlsFCxgJCceY7pKnEyokC1crS3tPm/z6m+BVqjIaZClR6G
J8jVUBz2t1KRYh1twknHJozE9s77XyXDok3bY5dIltailZVkRseP+hpzZ3kwN/f5AvD8IGqy1hLV
wSaT/ocVdsK6eocaFWIgWATBJC96+kHNWT7g+hy95FHxA7lmNbP/Lo5YW8wSR+6TVSY2THSLNeCE
wrGKN8zPePyUXAT/s+6D6ll2eKjdQQtuUT2rfUmayja0JJBHoE7bibFKfXyvkX2UhPSj7djrYnH1
R5ySXbiPJLHe6DvCVYhRcYRa3PxkOT5f827+w4rr86U8cFgb0Ft/dxEnf+VyhzfB3HpoZ9Pw8v/P
u3ZB8v0RwVFYE87LJXeS1VLxpMSQJOTCd3l13r0HCxsmXu37J/zRrIfP1Fl+p3jYXAoFZZToribn
6S/KQWAtC+hqa2+I3WbYPTQ52uZYyLznYDWqtx6ybkn7MwcbkfDDk+tnS3w7dQ752cPC90pOYxF0
Dn2T6Gn71W8PVxWX3uYykHrczhxHrG+eUaEeAeaZkh8fJa5I4Mu5L/rXK763+cNJ8OPdIrk0S+lQ
NA35fcNyZLgcFUTJot19fDJJbBmv3iJ+uoQmGZKVWZW03Ler6jN6MDE8Z+h49kEqhdDnJQFARJm2
QJcAcyxXAC9y2bQDhCzm6yNUrIoqGi1iq9Hx6tOMFiJuFADVVkAvi3qqPX4RVxzxf54bM7oL6dmq
XG+cwvyECefDgIvJvPwR2fHq1I47vfXyeKy88i+he0eAENR74uayyCLjf9eubMWMOZ7I/lGHuX9l
YU3qr7aa+0TOpbcayAQ1eNLg2cIYRw0L4xXmQ2dtCe+kX/4TEvZSsyA9NMp833YD5Z3qMWDj3Moi
462wuQ6hu7OY8qGtY3McFEGIhWv4bpS/erSX2k0PQmq5jZdSEE3OiI6MibycfvygI6nikNGASqzL
ZZt7yLKGbTtP0FCuodkLKGUZaWC1xKAa45GLfWaNIGH/xJN4QRdwQeygmvGPIuWxR4TK35looaoS
9YBn+ZFZBZ97fKS/2VUJoG8//pCfxRP0XhPh1nU7vtXu+98OsdcOT7ytarwn0qW563lQRaNL/tzn
as+2YEN/ZjoBWzsMPoDuLK2sOMdUgRUlCGXvBST/mEQTBa+5iFyrxOVQJHriPFLOgFC+VJV5QSG3
PmH2E7xPvj5qi7QlYXfME6ApzkQBucYWzkpcBC5wfk1n3W88u7ClOz73Sui5Ebb61I9wXlL+7D40
00cg454rYIW0WNRIonZD5X2YoLzvlqeabFHpPgMefmclytODpch2BpBZKfbm0H+VGWZHMus6ujOe
lXTquQVTipdqlBOGvORDD8Am1OYZwUz3XO0g2m9EBlwtjdSuOIyLFUvHinV9uoBpmIymw97XV066
r5lrBTHfFXk+raE/NN4XtP4i8lsvzJVLBmgx2A0exbjKhr65pMSKWSq2F1qSLNOWNAmHeFcnJNhp
MX9WTuygk1icPpmTIlFALeAp9IoMMCQgWsgcHPU55FuzsMwohL/bRI3q9R8LMerodGqs8jbdSBRV
oqddbgS5IneuKOpjHxFtm+2F674qo0Hr1euewwhtMCRXfswjcIk63LUgfzfGm8XjbmkYi4NPyR9R
1qg9wOR9T4362aFE/q4rH0/r4t85iYTi6b4e/aGVDNe/ZVoyxKremVUiQjXck59tUBVLVox5MGWj
E68tQMP7lUSBa7Zop8/Z2+/ylHJlRHpw1elMNGClGjAB1egqHAAnirEHqH3ZedF7BipDC/sPxgvY
t3I7E3jPN3wAc4UwVYQIrfskXtrsPuVCEv+fy6PadgUm5aVkRvcc4NbYMSIyzzH8AQtk+7dfasz/
8MsHkPeyNIWaNIY1bc5/zGNjCIX5/HYWqKj2Ihq/nltkfnKjMOHxG0+eZ7Bg6h+lFFk4yhoIYPGx
g6fhMh4rPCitq+Fw00BiF2NDjcve90hMCdgN6O1CwB6nurEw61g2THtGMyXRJ7CA3QceBqpq9Xn7
SzEx9v2TWh0PZE4dPXBL77R4Xq3V//Po0NV1evclGdyhccYF1rIt+sBp7+aNQHSup9zApQB4/PLD
XZq12vZQy8eYVy6mVCU8EDiG3HAOfWEQDLCR/6ZIskU+a4KsrAqYMY84K+MccDQXu9yaBBJqx1Le
V5r1ymsnRZN8hi1US13BQDgTEheF1lrdZgyYu8yIt+SXP8xfIr6MSjqFh8tKuOTS28BAhO51FEkR
tDqembf0iRT6U89SBaBnLbcANiaO0JrsiBCNjRqy40rvow+FhIjTnubAonXQrE5rNm23wqF7U+Us
W0lC0p15V8TNI2E71zBz+CZqOH0S66UmW9Q031BWkAamGIFyafP3ZCPyAVBSafx5HWX2miUYGAV/
sNgVyetSyRzp6Jr5O/GgR+741jIQj3/IDfo7EP+WCymLQKPSUeAlzrQCwqg1ILVvf1AtR4acOqEs
Mf71JHN6CqSXmpFjzCvG8sqcHPfSo4dbgoNTpRr4Svdrk/QoP31fpnQv7o3hdiowCY0mAwRGxXo8
crEncL29fXunt10bfRaK63aUulVKPJ0gurAO9lgyH9tjKnSGzNEnzYcyDgLEWs8Vg7EHqS8wTfuJ
qfFPU9acBL2Fk7zox9UxKFLZJQ054TEhIdkKGb1t1q11kjTrDALWRpWKXGEInK+fP5yBwnHkePxi
tzz86HBshwOc1dQxySZNu2JEjxn9miIN34qIceay+S3DaPLuCzXTqsnIe4w2V8SHSKN48/aMwlRj
I6JwUOt9NERtnDP+IoLLRXmiHQRn0aFwBhFg4gsf5qePrAaYjd+CQfLMG5cUelhmK35WR/rn9KXc
VVkCD5uB42oejuA+jxq/md0xcGPT51gSW2xySEM+JnA7xgQSEy2vtzNCL7UDrNKBdoZcyUqXPE3Z
u6eKwKEG/hjO5lv4Jlr3nVqBWoInh7krjHJBAUh/9V1h4CE6ddeCQ2gTOUSMuULYkC3LNIMb+EtR
cAvGdXDDzl8TWHtlN6PssFzeXOOuBER9iA6nD7qE7eMC+Z/X04ncXKdE67orbFDO2qX1mST2ypRS
Dp3LLA8dd2uaqWa4TQiRySQSpuwUT1zHvnhZ9xlAstIborzLNN1LHBTJHXWY7J2tQmKtbwbm4MY4
wDTMBa23n5IietbhqKSWTT+AiPEduAwtGZJvTWO+n3+hKlyGZ+X8KpAmVAchaajYvnI7b7jnovPV
o0a+ztWnLbWwWWxqbo4qcd4AN7TdQQM4nDA5qiOW0jPsnriFcPDnDDF2LSmrWvNEC+ulw2wNZbMs
xcoYyBlmQICi/bbE5xZ+JdTwmSiKs2/I+Sns6mh0b8+P7DOgW4oPb8JQwWXOwqD0dSew6L7ZRsj3
vlY1POeXVJjoVN0NXIQ0j7JDsgT/pqh53OGBNRV7qU1tXQpqkSBpaT6fWUG4hbDvL+LQCZeCTtC7
i82wEb59EpgYWqflfVsfto288bDfa8RE5K+mdV5eldx53yovPnSHKCb+yuaWX+6ViASvVJD3eqYq
VIgBeBhw0Z3hYZ3b2Sxa8biOLgPs5cwupN7phJUdBwHk4YllFMcQmn0ycQeVXPjUN/Bs1D5fZ3Yx
JXkwRhw/NlEZ8acJFsqpt9ak71o7A2KnseyPJ/vbcWptXzzEOFXQvT56dNyuHnmJo+doAedMCn2m
B1YxiUzqs+sf/hdJrfyU5Hh+Py1mOBRWAAd3lM1UU/xGdXNghXcQG9U7uv9xK5ux8NO5v4qDHjoQ
f4Okzt/mmBxjfPjkV4h775v/u1Mb4NsgrEtufdWH20Z/irv2csZ3J7OVfIhYqvuIpsA2KNkZvyop
GSrYwu0/OBQ9TYYVwbHZGHg9au92XcSQgEG97rmU9VXTACbc5r/lpxan56nt2YZ2hz2KyMllROYW
zuTmUKcmRp2l/YZVhxYdHyxyjYGSBP3LWZj4yWaRaEDs3m1MsMYP6ob5gWZSL2k+aWxgUT/BZubZ
JYpMi+stCCJJATMajLUrgPW7OFaLbSlANTW/T6a73rTH2FvuJ2lpCE6JWMa6sBvWPE+qrqlDcNMK
N0wCIv2a/bEiBacpMAmS1Y9pC4Bs4Djh6o6JLihTlW8weOT+5nKbLljYWA+cv/eNufhCGiBp0184
EsV8BGAtUSUz+f5uJpemQD+jTwgkYGG3zb11ZH/sProkk/cGZQ5jxVKb9QhBj3j83YsY56M8dzTO
u6pvHbOygrnV+1tD3zsHzwRGbjObE/Sy9XdbbMtYnfBDd4yiC3qi7RzWMvJ85P4r2WoJA5dqdXli
rV0E/qS8fD7PlA+4kosPwklgjj/kTFLsSs3c8+cPlfsBUaRnTTDcvCbUXlGPu7Qw2Obt5KmEfzWt
tVCrye6AFM0yr+94/3uoiAohtireCvK9O5AQg52lN/H9ziISQMVFKow65PO5TWF8wJ9hNCXozHA+
/fxlZcFJ0pCyNH2A0+NAEOPotCkKjMlcr5VmKQjAQknEZ/Nog7wGSZRGgaFFevgOcS4ofI0wawoB
QdnC63d4pKbgB8lO2AoqSmpEkHWM6f9sjylAQnCPVlghdhMeeoI+kAUeWyE8THa+smDgyyEriKg2
A/cBlE9pjpCwV8MsowGFFlLRtRxYwTZS9a4CVfq8o7LGqoss6rZP1LEb54L4aeNJeNvdPHkvoDUQ
kxs4YOF4nI1sGDMWPHtRDFFKzMzthK+V1cAiPhi8dv0/ZMZzJhmviHdMZufEMhXCril8Fgu+ZlS+
UCyHvYFUCMXmqwum+v5pyqdsVkVrjoJgc4+pOu+5nA8WqP263zXvwIfA41IzRNvtP5HsapOC2R6d
5RSCHG5X/Skk8Kk66sn5Ujz6jIBa0OmiS09NYNVY0o+rWI2oaMrQMEKdIHssSSfPIJX2UM1zDHsz
q+chYax9BkEYrqSeOhUTaxjPeUTT7w9bdyKRQLrJOD5elJtVfXLKXeNIZaTLctv1lhBFfakx1azl
4nRscRa1WofIt4t0Ex/1YNLrIQ4eKi1LReXcX2kpgBpkX/XJAKvClcHlUH6zNF8gkKmGu3bgfoAl
UUiL8Rm3mr7HnCeP2yYRAh+1tWfaYsLYyAQYQjamV3WEHIYgH7KWwWMn9zNs+WBEr7pPl1CCbp2T
FZDgQnnvgf7xfAeTkXtmL8bTxJpow+txSTONUymPKAr3DK6p6DcygQFwfU3jG8bfUXwlKoroGWlJ
2z68O4FKjccnJVxCPn1soGxO0I4NAqYhtHANEZM2hT0XPw+pQCvfFMsyKFFjYvIUOMnKgGuVj3K/
Bv7g4tkEVZ+29xWx6Bomq40vt7tBezvtG6epJi1lE1jZv+GGheBm2PbrZRZc4Clg7/Jcb+PmdMFz
UwLsukDsVi12/oG7dBOVzLUF+g1eUxavOJnWDgAsZAbS29nR3AbUVJ7F3eDwceuuW69tZz1VhoQz
xO+6NylwgeeZRzk93zTSRhGo9RD739cluvmSWbA5gMLMOThJLx+1J7b1Iopw/pvfNYo6ynTQW4fo
qw+O5BSU3h+HuZxZBwpwbt+A1ED44NGDbZkJQEkOrXo2z+hpoqcIdZbu8NfAq5LYcV7ksSG+rZGD
6v9lTjaK+XWLcjlSVNlOexMUcgfnibwKPEwhcoaV2dy7g7gdTwJ0qW+XkuQy5nBxXCK+EulrmQ3v
s6jPm5MSseJA//JAQS6rWMpiKDAVdv/ovrZU0/XY6InJeUOqBjwH2aS9uW+atWVunq4W59QrxDR1
rGg4PnK28rYTVhPo6okFL5AUhnu8EbOwlE1HYQrHJVK5ZVLnKfDMBEndYUTWIaKVSB4DKXAXy03C
wqivQO3jPy2eAGNClRlGJvDi1DvqX4mS+RWDt4loQrC/0gNhVvHH8uJRC3ecNDOV0Ee4aHiBKVEM
6TaHiwSco3mEOKnAw/sIMcpgaezLAH5U/AD2lylTHJlL4Z/M6HRMlD6cEMT7HRLWu91c+4ZL8M4H
7LC+wp1M+8wxuC6WmsIZBAwDabJ3qqCgHGeJY5EU4S0wPBPlFk24vN1lBOZff3hnXGipu7MxwAFj
bZDkJyKX/WT45Ifl2qB6csd3HebK0Dcwx2+Jf0atONNYFIxIMuKC+m59PolROmuZ7mvBYW5bJcRZ
QIZBzio4vXOjXUur7WpCjvERKaQzMZpeKnMcQ7Lhrt6twexkZ+jN6moiHGHbueZAzCHVADxoJoGP
koikjrVqfgjPNdFl1UHB3E5lS1l4Rdiya2HblsUNvKWJjLXoti+unrDccgSWhh41HAee1L1pwrpj
iRSvXEKIHg49lwxjgAA6kn6gLs4ThPzjVF4yXvTLHIYYZGVc7VGkV/0VhTNZw6unFsaMcM3n7HOO
d6F2Uu73Vs1k/c9+u0CqMLCrum5SnzbdXGURhzp4mbdc/VFvEo4T0e6K6GUEaX8h2QG1Hk+DhrvJ
vli56rGcLyiGbwmrrX1YSlGvEFzR0+W6G6Am2OPJg0IgmFRme6xakoMCqU+IoVvgb55zn23Qz6kr
smtMBDxoPkNjAx1hdNVFCLwtSLMJDRD7J1rX7hJr6gw5zHZpzSBsUzWKb4HTIGLBpzJOdkydU3v0
coHHW2ytmzse8eL943XGyC1lRP8VI9Mu9chAQ/S2KCIapuUCekuLlPquGKASvKVkLKk3jkpTCyDu
oZFyZlPeAcT8L5E9Ay4pdc7QNvcOvxhi9r5CK8mezSXMFtBaJ2SiZYlVSrMXjtDxLHJXYX8D11je
xvAkNOpI0UO9KFQgw+u9HoHHteZZsZkXHSlelDsVt6BOFowxN5cz/vxEPf+7mU/EiV8eclqxqTey
prVPpbWTO31/YwiL8pX7/v2yd/26vyjdDNlMXsQYyR1HAD9T8Ux0E2lfIsRsEoQmbzmX4RpzbEpV
qwPYodP2aAVCNDYqKApExcOgfQIVRxqFneyebq34NhEDwkt07tZIELZG0vIbZu5U/WDwRu/s3USJ
TGxtgyT2oKyH93ehTjukdZE3OIQf4mN/+eJdX2aMGDogVum1Dlx4e0bdxhwOcsRNhZzvEln+YNmv
BnhoaZOgDJl+4n6HW8hqltbiyigaYtkl+L60f757RkMDX8Ky968VEnTGasXvvCKkA8Xpxe2EycD9
xWFxifm8a/jA8jtQul6R6Te1d1MeliLr6ycDKiGhRan8LsUQPahirg8+FnSntAjhy+HPngYp5t7I
l2aHJKy3x8W8L11HXxq8xdxjmMrKB7xg6bB285r1m7RXD+OMYf2OjZwuqvjFqjakFEG6nDASB8gP
svGtMSumg7NfbrtMh84d50jYvBDqln9VDso+5FX/iCSqIgclsqpW7NU3cms3I/LtjiDU16+JDRki
AGDMZf8BK4snWHg+XbEVt7TScTbh5bJl/gvxTzCeLBDgc8HzntAe47VbbdVMOa9wSyNvqP4WSc3+
tvmYPVZBbHgxVt3RMrZG7dSxI9x2DWYMfHm1qDRW+0WkO39DxhNdVlXdFfD607/QgHEv/wplbRIl
S+En+Rts3HnyCi60maMBezb9mS5BjNLdcPyDb3ApSiN1/FMEwRAz4BPNoqtq6XY0C0scy10Gg/zQ
0Y+XoYdn6dATvVzlpdijW1N+RQb0B799MQ2vE2EsqqUwk8ci3Z5eXrLg9e1SegIWRb/UQXm0k0bf
iDv9M1JyI949Wl+0yABtptCD4jf8Knw+cpHlAU6CPEBgRlK+Y+mdLN2gRgx68jU9zW/a0BJh1jLC
wAT3wGdcVuL35UD97OFwlhIKa5XYMJAnhm3CLPJOfUmVXn2YvvemMB/+m92ifL3AVA2GG4FFIpUf
pf3Res8AbmhQSmbUH/kbUuQE0++QQEgFRr8CY/riy/VD9gSmW8tkNLR++WGAqiwrbJd59h1GdTDK
0WQR4ejK0pit5/xl8fFq0WZKfkaMflSTIcVoI+PMrGAMo3Fc//piA6/p66/2om4o0JMNKFZ0mejl
5oOn6HeHQrOntMoTY3hNXxyxHMheDDkxX2b0JlnRGkAJ0Mp7Qz7jrwY0/x5/Vfs1DzF5MCh/sYI6
1WhPULZdtvp+Gv/320P+mFtZcIcX08CmGAetbb1Db4GVKKhsVpGafKBxUNG+Olwn/Nbr3jAJmj37
411rlOO0H6NNrnfJISRToLTl8BIT30sX42Aa7jdCHF+rLPuI1tZmXN/nh0Us8ueZOIhDVOlKSuf6
XYl4Xl+41hiEsrLr3Wa+F2zBYNDISHfdgHSigOmSNsxWeBd0b6gHDX+yq08u3adcXbmf+urHUoqw
aCi5m1wuH6ZNA2dD/ob+EsVCxBXKBuuqYrWdfIg4NFHbiACMj6Zurtg4lnLrJng72LoiPbx/vcKM
WnfkLFa+aR8inhmULMFRVkq/oXLuHi3eDCSsboU94XB3eX29GNFU02aUJC08dpr6pbbr8d79g1AM
ksRwthCz/Sbe3iihuNJgBA08bChBbU5U2e16A0S8qK/P8thk9BfOX6WDVaZW4N0IWQIOOLWltm7C
OPnXeN0v5IqKlJzqd2uxrbiJB+OOUAcM0IYgC9wrfreDHvL5K9XgmdDH8VGuIC5IpgrfJvPh/xBu
CXnITkk5PbvtK4zAZk5+Xp0pDeUOq9QsA2MQz9hXuVTk5NCDDyo9e+YWDQWCecG5OttC5voN5hry
oQjWA4hMvItlHSSb85FDNuA8wLyRYbLPYnAdc/e59bNxUSFASnB3viR1746GN7w61CUVhqPgGNJn
F/ZHYF+HybH9Wtfwf3Doq522LHrnQaaNm9a9u3vb3e9hR4A9Z+q+mo8ZaGpoQyRY0Elr0PPMZRSl
Iacm5NRfUTjRh8qht+6+Mck88vkIMBbuRlMAXPaydhHyZu8COncUaxWFVqyQVwvcAw4TVmjH8IaT
CA6jZCgHaBIoFRi8s3ZSlVrqdEmldU+KoeaRBy9IQI19LFXN7TJIiwrcIqvNh4WwSLTC9BqtMycQ
LJEFMOkdi+ZVuM6yGNYRHmNr0WrDIlciTrKCDrOyVQ2kPgQYrufnDtwIou6l2IC054dqiw3sBh5t
xLrXG44TPILDHLkVkYsC9CR2Uf9rIVeX7zxWj7NmoK4KHs797ovKu20Ts6bM/OMsn8RGL+T068EU
JyI1s2l49mdKvXzYqQUAZ7WbBlcyaykuyr0d+oNnyraFP9lJOnwDRIShh2Wk0UD98H9yH8Erqc3P
xUlf9kyc/w8xjjaOsKK6e/e+T+an0VP8ipeza8h7DZO3aoHz9Gq9ZgaiTVu3dgnr7btY6RBxmQth
97Id+cQ16Rsv7BGe+CffObP589k4RfcIN/lNBYBG+qsTQfxW5dC4dQngoaqWugcP0EWb/Z8XbDKm
fpi+3H2wN45+4B7pRo7ipl85dbpsd+FNAmKeJcSMbIPM2VBcLcqRLeZdzC4J/nAvnm/f8e7IM/cN
tRpZ6zHizGf0rPx4suuBWKISxH7czxj6e6UkxyYyWggRRR3sPvH5Byh2M4XCvRoTZsJi0u/QqGng
ljnphYhSUQrbqIqGm60GoRR3jBmOc+NPfbm+7/MTm67dMbdyoCkeo/twyZ4h7vWsLguPFu0MM6NG
N1NetYQeDSipvy8xhb5bfzYZNBNQDmZoweGAf4nvB0yP8BQqXYeuZyi5flehh1EjnsK4wMilIy1N
brtILrymKGAcdY9HHkf82IqbvjPUCYhG3gLNgvYfvVgIP5urJzgO4Xd6K11tSPpUzldWQwymRl6y
/UftU+hKBYm0o7PUUn4/5xfQy8+/Cw8sqoto5x4asOsrBX8yAdnvlRx33IRgPFwdjxZ16pmwUb35
/H9HmB7feT9gvnnFYBKWxNLqKUiFBfcCN1F4SIBgTzjjmZmy0/z6DbKxBFTLp/zYzi0W8E5l95c9
F6gboME8IaUHwf0b3NzizyiEWhNkZEDcEaUTswePmb6S6S/IJx4ja06s1xC9Tp1qwPnj5DlAI23B
6W5XdQHWjs59B+O/gyzbJgXkOJlvzGhC+1zzEu2o4lEW50GOeNj4iFrkaGwb9//tTQ7Du8/l6srv
oMDWhPCZO2K7S/qfem4hBW7YxlmzlWkRcZE7L9GN24FEHBehRNe/eSuHPGRSK4uqfpXAj0+BEWXq
Jf0H/+sa7OL1MawF68NCDnanP/o55NsRFBRIz0lMED4W8KM9gFd3KKS3jT+WZbiO9gapaElRE804
It5gLgIdrhimUdX24WNHfe5zwy2mJEpEuYVclkn7rJle+ph80f6pTLcRi8BV35i7h/fDr9W0O9VT
I1ubvcmqKhTeczV5fvIu79eNAwozbc/2fnBX3zsvyyYNeKt778MZi4wq7Zh7ZkbKCPu34p7WijOh
djecNn/I6q81MwVD6odVK+lGJF4YNd+e/i9QsI3XPg09elEOHRzHJtvd9jqwkx3TbyOI5R30B9+A
tyhaqie6VWNUMTbIDWqsQpw9TCKjV0aXf3caEZWSgdbVH2Uq5TaBPDTdVJfYEIJA6OKkShRvYzPz
3uxAyXM8JKJUEe3KehJu19/MUsSEDOqqI5034dlGcOUDM813LJKokuhzj8N6u4ZBVif6pywE80lK
tRUxIvlIx5FLJsmsK/Ng5x8IN0V4I0om80Mw8emG5M090xhSfKr8jLca4zC+ZAb1mO1Qqkq23cT1
8QYj2x8hQ+rFKgpqSLQDW40PebCnZvtfMxhVdOQ7k3loLH/gI/3x4p2stMyW6NvBv5ZZMvuB0ckm
xC5OvpUsOvrCd2WdzMzQXzg+pqlXRSp4u1FfHmnOmQxyy/TyAOgQsl+eK7z7bD5/EHSwzGyz7r32
hLi6uyMW5/ERMO99WMBreCA/LFSt7vP1wGdsRQsmYnZCITIcbiRsAwSfBvNHbDMD11b1p1apmfSD
XBCUS7VrUFRMCKBoUVh3oCNg7+VVu0Oq5F5KfysvHwaXhgaBWa3vnva0AiSMz3MpXeZjtueZ39cq
RikwoTp5R8SSdhVFChvGozq9Rf1iG7ZQWIxU/h7h2z1AOsSGXfCCAYRHqRLkJZXzuncaSYMPDl5r
YFyYpIjlY0rR/8dQWFvNZLZ3Wj1fyvztcebf72TMXRPZb+z+aD2DLWJSYAiIMZnGDeYQfsLJkfDn
kD4RVe0PtMqLO5k8OADCcDGu2fXJHPqnEVSB50XxUy6aKLOkJF3MZ4goJo2ONy2VZ5gWYelv7kIN
BW2FU3gqocU+2jV9DEn0vQqLuOjqykI0hgCs6v14g2OarBlResVeB08EIuIe1b2SuqzObKcA4zH+
/fZpCVap8IyoqsrATW102oTFfuA1xlzGuLnFfEszCKc8rXNUmc3Wuy7p2mH8Mfml5yF5TzgQOHEr
VvW3XlzppgFTPF5bmVDs5LmENH/j5SBweOYCs7KZ1rv71UXnnlviiMbv7ZC6w4dZlYbU9DOqtJ1g
pjfqp7VotsYgQOnRkWI+t1d7swZBiQfHsprgZje6v9RSp4qbXFEcwCcDM09CVpCy4hzl1wvXmHJ7
6TkrIB9SOsL742zAFnKqu1qNEWFnwJkjNgfH55jBUgKv2DPFE7DTr7Q6kMkHpJNS29rZ/v9PAomg
kQumLg3ceGzjB0ZO64xRG40Bwqg6MFDD/8kgdU9ekkIgRs700QI5Jtb4PKDxrTPmeoQTnUkbffyI
+02CO5bH9InT1cUaR2qkVNF9h9g+W5zfc6/PjE+HCFGXbJRBQMzPc1TDIhLs4H8c19uFIQu3E6px
BnGlVUE+A3A5qjLzKoQlJCAjsX8DY+FKM+b/TAmzhPflTpcl+Yii6eS6a7my8OzKbpBi3UFNx8cg
nK9XsLSzL9jS7aZMkfoJ2ZUAykyRvrrJWm18PadRWdU+8leY6hAd1U5zVYLkgY5goDKgMLrFWqMZ
n1hsWEZwdS3F8nPXeYzxtiynxZvx3SJUxTN7lyngPSfifWTki/plMQQbPyQa2RYNugZ/DEQjRTWN
zqAgkHptpxMxrib7LWUjLbm8Y2r0aEpBDFJOEfSgNSTnGYgimM4aucQRj3Y8SduOG3ddWbDy2Y7X
owaVvqRbNr2QXgM60OHAUPtnCgLmmhar+EeRtUW8W0qoKdLyLTsxvN7G0SKPzStNFWOnTuGIYBd/
KQJ/yD62dQHcUTaMVVQmsduetaPj2ASbrQx+VD4Png/eRCzDWEjAV3dcz3TIqpsTW4fkhPb7Bfqr
NL6RHamxsSH+2CstSvBfOL26RsvRgjDDZR+8Czg1TiCXvlwv4O435DRb71p4XCnYWxUF5YPDAkt5
5UsHOUPPIjjJaxWFHbP0rBtkerUTJW6/wsx9tVR1qkMnIfj9od+KcXscyrbmcfB3b1WkruZvdh7r
XvtQsFWXF1kR4rz+BeZ6C44+3bUTSFv5HJXvfNCPRHXpLJfNOhiU0rdEV8tw8536nTtPWbz/gnhM
5mK13CB/aIFZ1LrjZs0cyiC3/YmJ0kK81/YW/TjrZWjxXtdybB0BLjiAYTIxynaPigunh1vH9IWl
oIwT4lc17ZyzzHAkISlPgLcfaxPaD+cu9uQjLmBF25ZcnawxYIjC2JxJmPm+B1sYp5AN9d5ewFkM
7pfv0x8X77fbbRo7lyENltSbxpaA9/C1hJkDpU+lgKkMD3pXUG1WitbbW9FvmZYyY7aqHavuSARZ
vkKgVsUal2FsYFN+4CoZG78TSB/b32LEM5QfyOtZeYxBccHyfd4jyU35QwdJZvRNufFiNRI0S0w/
87VwCtTy0mbtjy9uXqtcYl0U3RV7ResbiDdNiWqZEn0RQogMHgmWJGrjiBciuLjlHU+eEyy6wfXV
5Zwz96YQlx3RWz4Nz5wxGM64XhUtYJm9Mp6KE4zI5xhWg/udl1xGwwdOWePaaxbXEf2+fCUMeVkV
SFN/0B63Nv1vqBdiS+ntvX8iCTpj40brho/Pjvr739mo6v8qFwr9C+F3UL3ToqqILXQBpD/c/Ee+
+ixBuH7qZRHLtQvvETGQqP850eSj5fDktCqIfRwSQKSqsOkrzf8+bcpY0YrXiSQp0t7OUL+cDVsQ
u6KCW1TWowjqUVmiXZnfEQ/zDUF1N/gyihq1ONnuVGgjblIM9CDP1TJrFZ268mVvW4J6PKOxzF5W
twYUoxZ/uMqD9aHDx6tY1zH2w13kf9lLy9CARHMxUUgoqriy1SnsnnVR3z4d56bhJ8umXnAMhpuJ
uetplDC8pidCrrLuHPLkoXUNFai3MBzqyORzrct8UIoB0PORkWsa0QlanFZQvxNrow11RNKogAN6
JbnortgNjCg7RV3TK8SLepH60/3w7Xb9mmG3Jy/CQgqvCEJXtxqXSd7I31Aom8Zk7qq37hOwif7q
jKVNKC9qhvVcLSfg2wwvjNqkdcv8a0r8e/+vycZmlpeEtec0iMo1m52Jn+69VUUlAGirejC2gdX4
P1TSQ9YSVJlLfl+6eYQp6NJ9H8Nd2jp6Wmo0t7xm4julOwOGr16Z2+skQdgoq2krQBz/j8BtWjPA
7oZa4AgCFXIrVcdl0qoCiiRlsLxHWsJRN0EETytLg+N5TeiM6tCBvt1dk7cFtkEduEb81BB4rNuJ
lkDsUp32iEK2sGAtlnOKBiJKvvfZCmFGbdGfa4l8a74q+LEFADdWIfH1NMOF/iQ8lUFI4ItMeW5k
gKpi6WNxL15GQ04jhsz7hjBapvaAHraIUpQYWNzsS7WgpvIPi802uCMbXsdpRBggQTc8K7vk6Ni2
AzD5y60w365e6DcHCxk0g6vkaHldTPju7p3QZKdWzCCcfv14R5wogRxW+BnFMZvepBCtPajgvlXu
8oQdEoulGNgPDD6CGUJivaVJs6OCLcOwR2OY2rxnmEve/6XmxeR8rQPla76fkKpM7KPphpxhtolt
uHTg2VcjIfj+YSwqpCUjKBU4A6xm0r9+qvSwnxB/R8cp8MueTj/9x2PZGc9JVUsW6GvBQo74xXt3
s51btnWwGEdv0GpNJaTtMgwIn3N7lWMCSKT7nfwhyqyCh3xmMqOPF17wwrbznMfsSJXosHuqW3tn
H68BoSiF7pQVUL5Ze/A31d/RMZOx+PvEQs3Pu7O6V+HdBysSdzXToqDfjMHC82LWB0qcpviV0i3T
RLum6MPrhLkus/T6o3ZgWMXSmIHqESKLearHb79JVEwLspL3XiOtrvvtPU7Q88vDA5yzTaRkKMpf
Ap/GwDThactUe+z/G7qtF6XoB4Uc7XKyQVhHZ23gXcsZEdMaBb6lQKDuN1lvJpTnQv8XDYYwxbs0
VI8wSO7Y38obdFg1RJO8MGlRPu9jVmIXRxbQbjmsXyBJBbsHi+JPUEaBQvJ95BgEzH/0GlHxZFwy
b3jzMkx54oNCoAg6moHe95JhC+OtbUYXgpYjpvWMhLQoryrhEHohIW01f4cVzAs6f8UH3iuvUkay
L1TOfYHR+ZDV0PRgNr18VVU8Mh/johikwCqJ89p2bMpr0+U27o50lOQqGIiOMCPeI46CL+mM3+kG
xGa8VvVg+JDEewDOat1x96ytBfSncyNiFbTb007q2kUjdy0LxxKylUcDw6Jj4RkAlES4aUiJPaPy
LZWI+Hg3OWylr5UsjFNp/w0/4LbJ1I1SenJrCuQ/IDSJXRB0eWzeTCOf0P/76CFQ++5YWbHFexgN
v47AteotoTOV5EUW+XStpbS33rz3M2at4KOgeb1IHVddD7MVVBQhIoPdjt7v51bwH9rBhM9sotsu
POgADUhNmPI/S+QhxpCVbCo8ZKsiLCSLIJJ5t+2886Qc2SwUQxmb+EcoQRPrOq5OctocHmxLrGSB
vIzACOBTOOAwNHvrd0DjOML0gN2BACkwyR8B9OV/UKyzzI7zuthxaKOS4jwpJjLkji2N+hC/ub4l
nXkim9MCN+hCYTORNjC5uasQdRTgBcY6hfYJi/wx8dtMYINPp+3wv44rYWpfAp3vsnzgEGQPWdPO
Sfs5f8mjO0vjhtp6Vr7NqPr7oAljz2Cv/4Q2uN8OkcsTHUWWJGmC8eZw5Hewwoo9NH7AUdBU5pB9
4+h2uX9dPMuvZBRP4IYc3ZYF1K1QVrPKH6ugHf1xwY/hpGJ8p6PT2CKqOGdrMAXFwmviaftBuNRP
WSD3BtOmr1b5lWmXPNW2Bk2ueOhdfrcYL5E4zRXhpRnSrzvmnd8RXjttHlYIn+CtAWDw5UTfj6FC
hDMcIYhte3GWFT+4kzrkDYfLiOpqMnN22/MgFqJy5bmf8ABANVscfSUwqoOS/WLEM+em1Ppl+5rw
dpP5yTTil6VKlxbADWFXnTVFVDFQFQt5Y0OmDfgzeGvKteO4tmPAUa9rtW6R4fG07SoqJ9dP33vj
2s5HeaP4I12gxnyj2bXWmBrtpyqyqEUNle9HEmYm8HCjvzDG/Ve/7JgD+6q9wlTCAaVWcbs/uq4W
pNlgGsmAmU0LfyZMlJRRhSRZ/omnjaLik/F5EIiCnrLgc/bKHpb7xKoM++LwHbbE19NNhwHuVhMd
G3eMIBv9neAZ9vQ4VbgzlYZJmH9qIrWBvosXhHbRN95XcxQFLXH2NphmUsmLZQaH3LbaJ2wf1Eal
5sh7chd/+MkIneGgknH8UjMO8RZMeCl1PLkYFrq/RfDaTU+BmkGjHymJE1HxsuqR13AMEbPBlsB8
2Lhix5q8RpLgiRXV2N83NTWqoVzlhNoGDCQ7lsdpw2MZW9H+0peqVTe8ZRIxsWJc5/ZjIg8EMYCN
+nOEITwY9t6Kfgi5DCwmmUZqpAXsdmN2Y4Dc99fhfmoDTwgTU9q9HrbcIbWe1pkvb6mLd7njYkAP
Co3BEkZoz/nT7TXMqe2IVox6TLwmlyfDLHiadxheWbGgCJLSCizuPlhxr3TpVXypDhnLH7AzWE9H
70il0FHuQbwckXO1TVgSL1ecGsRHMKANngxr6VSZ6PWGmvYDB5LyPz3iinZwLvkKHf3isq3YqAdo
06Obx/FeWSgJLpRkxmvfAXColOCNEgcJIiZSP12FxNqA3l/2d6DLvipE9UqHweyAKtjou7YYHlpz
AK2TC8ClH2U8rhZQiwU87fxpcjhl60ZkAogRUgBSPRpIxFmUBRRhOF5fiLYfXkiuF5zW+caDtsWh
f7mxmqBXAbJbNIMtrXYZesb499241uTSP0xzrKsZkeSTsQS89YWyL1gUjdllXKQ285Oe0M5sroWZ
tB4A3oX1CC1OMukxY2nn1ROn1LUr77DRwIrx/lP2lzSxyPV4mdzRnhTkI3kDRTSefiNRnkG3EYwP
ww1uprtocwoouMDFUnvDdk+EkJy/F+Ij0UMh3ctnW5MmaSdfJyKtXWjSLkdHWmJNVnEgTEUvlirM
p+rZVdSjYfRb7Op+7Uv9iU/lqhpT7OhQMmwKiMnmny+Vn0NTh3rBhOFnxJ0mtO0mXpm+giJ6nXtE
4nx94C0uRs37UxJryzJTjFo6dI1Eldly7Q0RUrm7/lES9Pz+9XA63OCIOf4a0IJ0lBjwI4SADPUS
46OsU5po7fHlsHEKUMo/CCJ0Ag6HG6uaAgjxCbRCTvSwLLbTFJtFkN8Bc5rTOkKWYX8pX4Iu2US7
q4px8I6a6LXfj3X4CIcCXwgC9SVDs4XGHcvN/YDZLCXqGhXOd4oxIcBldlHxUYZuSYMDDjhAY1pR
6qgwAxb2jNT0HcDEW/873RP0WVZGh5LeSAw53r3eY8ZzoW4Usxp0pKEI26QFgj1KjhRnVTbZdCBI
1anu2Ijr48UtsDONzK5K0NQpF7FgpVcthZAnKHx1sCbIi6r5Oh7N1jsNkNS4GSHO92fj4WwyNba9
bjunYI0J02rrwAJVNJNBTR/ivDOgGX2DEYXmROCL38ckmded400rsQ7Kt6BOuSVGkuJ5yEoQU1SR
A0OnD7ktFa1yVpsCCn9F+bc6Six0EOMh1eDwi5eB+kxXgLG0DWJ8gQgZDW4G69a/WtZ2znplbPJA
p24mFTQ1kluXUtWXQd21aXFZqBLMiNmkRC+aUKY2T9KxVj+yENzCXNPeyN7WRDRNmSNAuOjAVl+t
yZ//PGlwrzLMf4F2f0yGa1mSoOfGQlOMR4Vw7zjk1qQHglNHHlNP4kld6JhV5bB4Qk9WfZbarRGw
+h3wzkQd++2LSv1ChbY3xjBP+a/o4K+ErjJsYuKgCBzZc3FV2qT8NtgRwLfO+qfRCAeX0JwEsd2D
HQyoU+EncGK1mAL9f9OmtrDFdz0vh14pR5mpXbz3EKzS4br7yhzs8dRWjbWrV6jAbh8iKvL+s8zd
599YOVvDuv0LYqR3X1KmpvLacrVPCQRENTfIAM58fxrTn3Kq4oY2/DlvU0FnHHZF4Y9PpRI9Ddwv
7elPdJNBOQRKWfwLYr+qe3BZGIafGfK5YSITx1ClVgxrk8LJDVtN294o0M8jD+8IYyf96u/5Y+gi
Ks/G/LqjUZrZFQKV+PbUI4KyVjxSSvkVAua7o18rwiof1dZ3PvYJjy3xdVAO7cX7gpZDBdPS3wuG
pvqZrPEYWssjSVn35f52rc5t/h/XX9FNaRPcrbR4gEo/HnkiBKGNhihFg3/1XpEhPWcSZBZm2TGc
FuPnAu2lyIDzsefEPec0fz/mMe6zQSdZIVPe4XnWCHJjlrj+khc+mlydKL/lnmeoOxnnzPcDZr3v
C9ibCz2FtGJGN+RmioRCFnaBjWzWSsmMbmRNOygg1t5Z3yJElSqqocZFxNQxcrjMYbi/sxDKk3wj
u5p0H/SK80Y7FZzqO1kQTqRKaMp4oqQocUPkIBW5g2qnvEBM2QKlES198YfJI15DnWqPhJKRbgRt
wGW1h42EJwrljk0DK3aG3C0nNZiKKXuOcXIBXcDt4TgzofbJyuVlVG7BYuSpYbFqp/QsNqJ9EfbR
XXg/HdAzdvAedQmnh6+zUZbqny2jFhdE/tw8wgVNOelspgqzaHWZXHoU+ukA/HJJj773DdNhY8m8
/xOeOfaR1ust0g3Td2OsLGxcDWASL8ljYbUb6nOGTDWTjEQea3L6FYCuj4XPQ9aI2MnoAf5UkrKe
tXpnsxgN/wBIn1P0g3NubaYz0RDOvXGO9hheyRV0EiNjoAmr7h5X+MQPiGgABuoaC+xgW3/p8uVW
S72z902PaQdGjdhrIzH6Hm24icfCiCdSMm7rUNSgtOSCvnskgbWdsQRA7ITG6S3PsvVkBeuNFlI4
UDPeyaS0z1BuIGWEImobNxhNK6iSZN8COaCSdfwQxkVmqnkwj6v3poU58j7jupbn55z09KocY9eh
LeET45TW9ZwWv8a2CgDezB2RzmnLydnGtBiMQN6APh8JhYMqbhwneleE6ED+dtWtuYDNs2mREI5w
WAIdGC7KDPC1O+iMLeuo7hewbJYTZAtBfNUq3ghiL4ayqOEteez+snarJqt47Nq+b7vw4PSTi5Mc
qJCn+9H/NDG3ZZjY4X+l//wOihgxI/Ub1N4z5FYM9CyiCbGgm9uM2PlFOzt2x5xGDqwGjJcOHfHw
CVcMNBLk8G1Kjj/E6xGcpW4z88ObJh6WhJ+H3dUqRhz5gMnhPI9Q+aSUnv1nGGYWU5p+bLj0NBWH
yKWmTIrSxkQC7dKV9hrKyAbqbdFfBzfU4QWePqwVI3Ee3e4VweuU7oJyjcgjaL/3yQt4vxKJcSWj
W+e8sFwh8DL87FhEtzWehxEnKyfosPULuAM91px0WDC8GBGlxSAZTGi9Zb5jjkygzxBn2Z//6ELr
J32//YB2ezGUXdLjTkExoAHdMOarvF8J6aAqkr6M+EJwNQJrJ5udNcibS6Ke1uSpgIIDmt+TXv+d
zLsqXQHc3OqFBqVLM/fj6M64zh/YUJfo/ouFHWa2zenFfGXiZF47RzNhj1juxQvXV4t4fYYI7lbX
14zx1nvfnz0EucNhihPXyvhic82nOlJlwA6Aw1y8cZWCYMcWY0TnOvqvsE/D0nL3Bv81XDLGdRCC
FW4lJtGKDb/yAT/C3JzAojSAVPfKpqkt/s2KDSFYygJHR+iTP9/ZnQmoY9efIHtc4knCnm6JFxUz
LFjqUWzc/5bu+A2orzVFa1AMRwzUrZslLcH7QgO1i+OfWKx7dEbbQ3cIClk97KC1rFlo/+G4qNbo
wUzcFAs04AlF+kAp+NMOGGd5WGaJrffjlBGMzT9C/p0wNeysShgtGL/OtbgSuAQ27o4Yoz99GYmz
4vT6Vc0yMfBa4toaCLDb1tK9p4o8jBXzYVskM6cFoL2R78Qjxxo+dimGV4/ADcuEOa7cgnxRBiXB
Fa3Yea7bKRV6uZZcC3naaQ0HWQxi+/OeAvQhxjlzlxDKrqu7bj81BCgBis7XI3KgIV2o1BomMWAT
eNLuPu5anIFAaovjmLJA+Epr51oYkXztH9m+tFsIFEv0lyFThoke/5QErcWvDCdg+YZOB2KObM1J
IcdW3ddcGitkqj9ZnWVr5y5pViWb8mR5cxD9Ax1LYsa+gZfamMkJSG/3HLOKsVr+jsLWwgJEog0b
WOrh4y1tX+c80zoZaP7gmGeouPr1b5T8JrvPb1H94GnPpjCBXZz1CTf+/A8jTmwhlI+oS4fa6yYp
FgDkdPcWKrMqbCuV93mova2fSnGySMrvO6SHr+IWmORdbv6tsd6QlArHknEZJLldY5m8NSq+VNs2
NiE84wDgFxDB0nB+nHykugENYO439YEvSSdGiFpiYl44ooqYcTopAsBJ7d6PP8s0+XAPlYbGyfui
N6+LKMWo8zQV0rdOmdCHj8yg0kaAUq0NZI1plLUfFZMH+GP0w839msBebIVaNimk2MDovMTbiEDV
DEnA5fB0IqcnuCMIwj2Dg5ocdojFuC8LMP8b4qq+sYfQcNzZ0ZfLxxZ6W9jKwOmArLxNawboO4hM
byLPVk3Rx2qvpO2490Q7b3VVsIIaERXBwE81GpJUh+HF/JqAJ/N4JFkUhpKGSYpGG12Crw1ET9DW
DtUHX+lSwM6bxkOr+BtSCopyama9kNI3A2Z7k37mkqbngkMxyvDL8kxJ4CL1Lgu/cUYQHYt1dvms
+7/ycCuzsRfBfJ9WXTbNWteu3IQGQb2l79lzoK8pVuZ5OUaW7ir6/+o0V8RAG4w9/U4DK2ld972Q
qWWt3R8Uics/fkqivXRNd8Vise0p0NSDTwCL4d6QgSkKQcWdZdoA79XxK3EWqRcfEK63DZ0OjLcd
6OJgaw3QtIWpl2x3oE9YNw/7kzsDsuo2UAXLOK5U/CBQ2DXvn24hcTxIUR8f+6ujGQYLei/C6dS/
pJ4bYwzJphd8NphnLyh7W1xEbGnaxwZmlvg4Ni7Ts+C9SAsz/rDgQqxfYt3Z7BMGAKgjdgowk1Hi
gR8/UbH2DkuhqM5kmtIkqvcIyuCtOryV4lyefjSgd2VNbFGmeOSsCefFbxaQ2EblklAQ5JZbigXi
0OiCT+bKD4RTXXW8Id/sr8CMM+4x5crUA4JZdROPAZeJ5ZvKib8IUjA499/iHej7+JSAGb7sfzql
vRxfucCNzIbJEEZVu8x3ptoPG59Zcp9Tp+i15CgYOTTh0rkMwMTrOvfPFu/XUxd/bvB7uD4WUYUB
uWM29l4SnLxv65/Q5tpGLtfOdJQSP3+NVaqn3OUGEhBr4QUsTykF9zCD0x1uBhvPeziquwRAI6G3
OjSKCJlCtLaTayumdwp0bkf1wL2ZPoEJYi4OQIkF2ePsitVax1zOFX9hTKZ+5oMqUWb1jJRn2n+Z
7f9lHKG/q1/z3p5PgoGRF0qBMp7TDJdLBf6uJKbvLu/U00ZmXGdMcXe3Ngg0vFvEnwF+g3h2sbet
6R5PkfGa7DCmDkAWjnxkOyOpQFIq6PBYpwXPgQQmAfxX0O7lUuFhKqs4IA+FhhI0qFq6JNiInQf5
zYKdCmMYNN4Y/UxWyKdVR380Flyp+eOPFkwmKfYj06zG76TEbc720Jm3V6+QAT9H9ewim1eNZoSE
NFkbP2Luzu7tR/JqiHxBTufrjGW/NOnFMRYPnNl+zdjboPg2OXE2iaXQSfaEgUnj6Q7ZDLiRoTqi
QLh0JJA1iXxWDAiHqejGBxDfKBHUiR/+KyC1Gp5hy3fLl8cTzYPhstgfJ9WEbWll6q+eBSEHoOfg
WB2l+5SgNh40lrSscsUIs2ALqbRKosgrGHeOr+7L3UTZSBblpxMFIIptmp8Lqmj46ZftLyMRPKhS
dpEhKLca0MxMOpjftCZwsM5bvpB2BURXqMncxsoRSVVz00zNloZAeTq5wNjlMMWlICzZAQU8H2U5
muL/a7falIy0mnOfeb9gDuc4fzUaeX7keSoWIut0jdt31rGf8/yTP6lue7ZHFcVsfuc8ROlUuDJ1
rITJrjWahsy14bY4nqXxo1PYLr91dirSXAP//xqLGz5Zq8N96cWYQ06if0a9NN5/gtoM3hCKx2cJ
WzGnGUmw92h7mjQiZqpu08kcQWydh6ZTfiQQqsrJ1Iv2vT+JnmaQt9bOUPJoMOUnnBch6nY+PyBQ
77z6NASUtvNYNVs4oA1YvyBEugRms0hefrKtHKMQN6KijJnROSPhefUnuxWYMcT4hfcacVxxxRTO
XPpuTncQLsUtIgUdq6/9UEyMnoHnFoJzWpUGWRtk9Da9QmGbWxrOmuYBIXyNmoK1fxy+Vn+dbcNH
6lVmeM0J2mV25uhzlIjBYpeMzeoKshIt/a5/xEOOHi5D/Q+qb2845QWMhYZT6hIinCPd/h3MnouS
7TEfCH5HJH3/xw0JG98/JqLbhiVLN9UMQcVkz7qOjLfMh0mF0eN1Ge+14VUOMYfNPgLXSei+idTa
oMd06shBnC+IikQYrgUnObMx/H3Dtwj8fkB9Oo4McWmC/+59dIM1Wr6ii/NX3WQVjxRCXoWXPP9e
qdrO9vZCp5+eeVOpTZaWNrDuN+ovhEgZ+5QY106msHvO7IXA2jkfdxCNhprnEb7JaTPoCPcb/z1U
00IMN8a/T7uXsxwPoeXZ9faW7fSEJ6oyN5nR2EFVU7O9q7Y1WRam1JLqtR3inQRA8DRpLNFtMwHK
iNx1f3vWq6W7dDwHOnsUSdcn7OjdWLPhSO+8IVu3G4VCbr8M0CYgToDURtfOuzP5ej5TDrfLgSck
LKmBHRRQ+f3nbt+96TGv7BagzCkFc8LPdRdrXd4UR8H1j2YxwBiPtl9d5kD0czKBpkrGf7BZmFqs
a0y0lQoZd0dNhPbq0EoPnK3vadRyzsuc0MMg+s0GzVc8T+Oo0jJyvtkxGQHsZE3VsYwzzvYzyTi+
K0MrbKMXF//I1wpvbP26OyxwD2rV1AFUcraFmSK6JinGgMckja/G30tjJkZcim40ugTrXjy+l5CL
mThvBZE4vUhaGR2Nq8eSwDldhzFk8HD/fMoSPsMwukXHBocTFOC2+dH8ywqgtOQWBz5sdq0HXBUd
HYxWc2pl0D1B2uX8+/JNw0WahPYQmc1HMSYrCNRrqpLWRzh7/3Fe8bkh0XuCdbnAPf1yU1vzhkvQ
r9ECcLXjDqvYQB8vW37yRH9GDC/YL1QSt0EyLc+Y+KLOmSBDV6atwadKumQnHHvZ5i96+pYvztR9
I+j+tqVEoHBn0ZjFV+2VwjCz/HpJsP2at8K3ngnky7/kYztXZpa8EdKmrtzlYZa7EdKqBK+B06l7
sTdHgMi84c9g9jJoV83EqZz9as4z5GzVdcbCfeh521vvEucgGL4NN35YZKTzWPMPhOO5pa1jT8KO
ZjKke+G71GO1ZI13XDi8MtbW8cRFhbY8KgS3lOh/5R+F5+5hpnNJNnn4Bi7FLQVKJb1dE+yNC5QB
EfLTwc4RHVCwKAu3vsKI88N63gZA7N+9PG57jz3OQbOAjGuNcASBI84Bl9KJ1+i9PxRq0roj+iSB
1GywySMKo52S9ce2Z6DqklUv9WIZtgoha42asoVJkGbsY166hKXV/xBwsDLEoQ8DZddRTjDWJyRo
x3COGgk4A5lSoRgKxsiOFBJMRaN1B6nWMmaZ6eYSQXn9dQ2h6G817WjRgoea765jy2UGsUY21AL1
ukWFquzaHuFZ3MoOKZ6fMr2YJ5+CuU9MjCGdZ4upJVQ6WGMg2eqiGpx4JvnaO24UNktipEieDd3o
0jJCVYmhixhoVoblvSg6ii5rdPM5tJedWS3tS/n4BBf/2wfCn4JCSNaWVdG+KMYLi/08lHtQenKt
f0/RLAhlO5cmG8HneCq10VtW7IUlqvdafnwlmtaiULPpg5Wk5dgYV3FmWiSr3jO/luOGQQ/Lhnlc
3JxC9nZARs7h8ot31o68ke6VzCBuV1IBcd91MTvoNotGJ2N+Gwq7fL0ZFAiE/uDHxf4YPadoKfxv
NooQeIzInQZsRScnQ21oJehuQnjMyDEqqcSvDDx4Llhq7xcxQS+eK1RWk8TY7pkicMEEHArEKM4D
TOrcaQlWyC+IbYwIA7BL3YnarcGV0zSnKuDgQVDMaeV7VgM4MUNM6TT2SUQtofCEk2g1Vwt/PBKl
QHTw2gp84fkSblwxSkwErhA8JmFu7IBN9KgwZRP2QU/QoHbDBs+67JV0F2YqfkvqlXWbKn6KdR8b
eO0ry96gnzhrsFX31YHjnqaRvVaT42R8ZPu16POuuihdQA+hAAAMIMAVtO0B9Agm3c7duEMMmxU1
VKzLTc72wUOX8FnD6nPUIc/fkUdddaLFZwvhcMVcfYeUziNB2YJx4JXV8gsz6Ku3ErarSJml1fuk
LkpFKm2c+mh9LJUsewB45C59nZvCIlwlgrJL9p41XBQATg7avva/cv+8s2TJqASicnMZCVxGSk/d
DufpJMkaglPtPMCLjAgvFcbg3OHkSdaQLSJP84GxgIDkSZzwO4Gpsp9vb7ZH7yc9DmiDr4K8Y9yu
yOHzEyFLhiyJNWWc4bL1uMqc8WPtNd1oO7ev5n9zL8C6MxW0j83AvHgFsShKIGLV+DJjUFu0Nv1I
hPhi9PaG9L+DQE0xYBMGvJteECfiqzh1rFWDxhvj0Sn34CN4YmjDxJsNO5pHXmf7ifxstViCWms8
sOyU0Dz9J1CEEOq74Mle3i4hT0vOSeZW2TdkqDHGdLFJodVG5za0eniHJmAljNr/KKFtYGwcJof4
wMrbpCbkek+dFKhegBB71xU/1Uw+lpuXUOq3HdqrFXjny4LdVzNL1H2N2KiUuvYwXGdYfqp4OT/P
BEt1BJ/xOmGRL0Ywn6X84EESMNsot/6Z2pmatqNvkcOV9Eer06uads767xN29orfesoqF5GlpcSH
Y8kfijPuani6o8o9Ouizh1OW0szYRMsareHWq6yMdQp+EfR+z4BN38E4Cey2ujvbSiLKb6wrITuP
4/45RN9+LOZCoCTlNbbWa23bGgO/udmH8EZ8i1nzUepkBZmx0+UHO5/oo5a7Sd39w0i2VLPDVFhI
WwGYrrrroX3lSoJnxQSMe99jx3W3ZuqSr0VQcgycpB5Cczrbi9ytqSU+2MBxk6REfFMNh2rRXTbs
9GgNnM+WYNsMf++7VBOueMWyNXIiV9RopAhpzHNkVxJyTvU1SVWCfjrzttbQFubFpsbLrupWcE4V
Stho4nlpjcNAtHFF+LhBPx/P0TpWF5SYybxjGdC4E4P7Z7cOuDSh98BzUpQZfagIgPi2owujDRaV
6LzXhtHmxGFkcGlUhZSR57e0WvAVwjBJT01svs5iLh8IQMrkJFYLwXLCUBoEYDIpy5+RDr6R3LWF
s47jAqi7glROoZFxlf9lSvjIkjZwzFLqKGWVJuLRgTphc+DrOEyEvFVt6SvnNYM3AxZ5ayzx473I
LPi6PzDkSJTCJ9S8JgIhzRJzoUrii3mpNiSKLbH2uOvKanXPafgZrzDG3rt2R092Oi/8fr/V9dqo
gYSVEcBF9zVwpHB/3EZHG3hqlsp3GiES1NSCMQbAkxpGgFeoTTHNEQoxiGfncQAraGkDz5odN1j4
o2WMXmP22OKTiMFuQWtma0AHHstW85jOM6Ufog2fOEMFdFZobrmaR35QG4xQKwLByXV0S5RyonTp
lKjM7su/0daYsPyHZTr+nQ8UsDaHxNlU/7OxmsNbMrywcqoFZbWP6Ur+PADoPL65XVqAOQwYDpeP
AtIvsdwKPWZtcz+syBMhzWCOT3xQ3gNBj/htpZ6ZT2i9mlOPIhfoaJ5y3cwlyw9QuBW9DIbI79Oq
NAdKhKGfkhm8P53u+GhI1IBwXwkWbLG4/R7o5mQEzKk8dm4WF5IUzACYO9ERD7fGYvuwc/dagBxi
D3GOxagSiN2F0zacJejThG2whT3oxfb3rE/39vXXPkVHAYrH9FPwatsc99vmqAUhUSgQBGD5uZEJ
XPnpay/Nvq6vYCMtai4MevSeAK3DIdS8JNAzMAFkLheK9+N+jazYoTcZ/02D7vchENI0tCwQWgIF
v8IFfh141vV+PgqFBtaBVkLn05X7ataYBc5MWKI4ZlqO9BGr40Gu4p6jby60QwPYgYAy6039kPNl
iJRTfcSSs/pivvnbtGMJmXKNdYEfg0y0JjJSboH85LBDdgycaVD3QW20X5Kl7G0MxeW/YUBD2spb
uPfYWgqK/fbAc1dbg9TXfJEObu5LFRaOBQcLhAkvW4Us9t4ZgSsztLnldFRqOiFzhFISZAO5D/DM
2VUF6/tT9bXQQDp52zgLwR8H1d7p6AnPLNl5iLP4zjQIfRs75uxiqdIPTKe9O6lyQW6sntXVn+GD
5jdpIHvI55g7MBXJ8SqynvTzreE8Xp2CA1SLVBv6WXTGvjFpE26Mk4LNsU9XNAjVKCSAeo/gnuGi
jGRV046eWjatZlHqlAol4o7dO4ipndLDr2sFeumh7/gSq7X04B6SqR8nNPO+1HhULlfKJwHVvTni
ReB6XMxRTI6PkDk0RJf2BV5GY4Xl5tlZFVW93QZXjNKFqy8Ttz1Y3xEL7Cr7Z0ibshcNmM1Cj4R6
E//ot2GJ2Rj07rqXyrDA2iQ7oCNQrFw1EGrdXH/eAHlwoYb1O5w/3SpHzn1tzuDqACC4ujaoG/tq
VT+wkWAz8jn+US0GVI6z/CGdkLlknbBy6EI2dRI9O5mY6Gt+0xhggvz45mKcSs3nF6V0v3ogtEbF
AkD5F61wVLN8psX9FMj5aqFa237HeNNgPHTmcEQzhnx4BPer5jUQrOO5lmdRwEp+FkZRcg6w0ls6
CDHDvsvMDk618pRXgzfG+x2z1EctYN4JL4FQjYOkG+Uzn869yCdY7ZypmVoQZ9dJ1duOXX2KAlLC
lPorhsl+r+EXj/VWAO/EHxubkHm03yAONZ8+MkXVtc/ivGU9pC4hdqWUgHzp3BaN5YKEWLBEQJ1S
3rzEwLWSBXpwl3/oJZwIL7Y0Oqn2CsMTQRzOe9L5edxO9p9zQjcGS/xxHxFDVVzQOQl9P5QmWlcG
aa1Xj7EPJG1/5owicbN5jQ9V31ScjzmCMWb7KUIXv2AwvSQWJLilVVpfus3hka0T80HO/E5jRbhR
b/1NzZ/Pzgsm/JYFTYnzlDKycfj9xxaTd1/EXI2LWyd/vHKIBkNqxILUCPES9KBMnQGTF1u5AE0G
806bwJCLbUJc5HX8e5MzQOwQ5IGlzjayentgdZ6PusX24V454ynq04ceiiG9cIkOJE/BqPLC61ew
FGviJPFC/HfMJF9uhMmJLpNk5xFAcLI+njbKezxOI5IUQ30+03W4HvJWbkqROfXEFHFZyc9nfyZm
fbdaQ0vueUST4B3MViXQPiQr85xg5ELiGRkFzXDcWUxTQkVQpnY/Kvfb3MOgENi2aCSozgnNjG0h
AZHhFkDkE5efFzBKdSdjbYgHfeh2fKqqQoXQznMxtLXjLFhwp/tsZGj1yyh2ed1Zy8A45V8oEQQI
ZApghzq6UYEO+X3K+zn2s3AwelKkCkRpMr4fNxdIqvOdLQZtfu771SCtm8ki3aeSerm+zhr5et4y
BmiriRo0JqH122FE/rCWpSIArwj5Evuv7XT0Ypp/QMp/P6/QSqisxc2HGNmWqSh+5fjik0ExFrAM
m3LGl09VTAI1OXBUBBaA1W4xO2IhVSNw7zkbmGz8EoXI5Qwiy38SXS15zjg0TZYdKzFfvEn82tOM
sjV8CppLBMMy+Xwos6D9zEpzVZENhLnk3XqbddqDhsEB5MzUhbgJkDamudxMRB3dQnVKyJDripaO
PDKV6FaX95YX1L4sifhjGCixWwgpDCxlQ1QfkBtsQib0O5/BkeJnQMW/C8oIRsSc/cCtnbACOq48
fAj6YOEtwFjPUREUcaE2VVJEv/VjajgCjubkdK2KbJEhn4Y9eqa71/rMCcBDvNium0G6b4mPBBnF
qb2aZJf46QMGW5zd9j3LGPpErKNhQmyrdqfdgBGRQYKonJs5cPQXQ6uTjINRJBGe4NPDQLUNHEJ9
7cPYnuOTZZGEVJdvRxNo7/oh0aXGJpTnOKm+E7x3NxZEexbs3R86rLfNhgMcJNFY0B6lYFqj4qs6
D9BJDh7JdsdZ/p8Yhcnx8KBfRGKjvo+S0fnOetrDb4ieB5PBgXNoyuFty+ciBm2rGb7XWSTlMEQN
6jkCViobcfibX9EOyYE2B1REc18Hu1nbrbIDz0Grzz018hNDLR9VgxZ9DN68Nq5Y1VWGDHs38UML
fRGwPP2keGzyg8VSB8tN++4RfO4uxq9/utBJeNjJJG65FLp2Zui3IpenKqbcmxZbU/JbfE+uqnRh
N8qljKEgRr/e4wnr7mYfXcB9hqwNNb4stGYaYL9xWbnefHrK5aooqFKRE3iYjDhKVd8+2Htjl2Fl
sl+3ZRhGKtNj481R9XsHMrgS3V8TUYjZAl7bTJW+XDacpDEe7Jetb+D4nVtkftitXVybcOjSlFgO
RMOAZYeDWVAudBUXqeqyzpa3pbI5mrr/uSgg+ubkDL6dXv/tbQBk0Mg22HP1dDkqNhP6F0sI4qSC
D/WgyQAa5RuziJURdr7mzhUNepHZ6BoeQb0ma7UKm1TlBv+6RT0rGosG+JVN1YNGYFM0XsMb6/l2
wboVP9skvVWjTlYVUjK54ai2zLtrQ3F1wEz4/F0JrKHQizVLzD9nxjmScs7q4xP0rjszDBEBwxFL
osYVt+tVirUmJPght64MBoC9dwGZ7EuzBBeprljn/A+J3U2L1Gs3Gzmpb70PfKIB1mHEiF3+SwOS
4gOu083r0vG7il7JbaHIEethlmjuT3NF2gQHOAfMjFvSC2cTnsDXd7muhUK/jysH+3Lpi+m9OGIL
MY8ceg6r6Ul3ErHbQ1r85QXyItH+n2eCfeTqMm71PIAcGHeaMbHdE0qd6YWOdYGbGNz8AyaxbcyU
31lolP96M5k6pTdmh5PwVjT9v7H/7xmeCGuKrppDOLaQkHdOL8/pj6iKhosSKB/Pot6qS5MReu7y
ONRtK2dnWzgL/S66R3cm4Qn2WbQIl7wgn1h5tfYlNJs7wdadI2LVFrhWxIBxsFWKNckUzycopsXS
BuyDs09H3vJTR597bhHSqh0R9fi0bbqYwpwrbXONk3/rnFLKYtKR5i+WSJqXK3ZPyzm6HMz+5yck
1215SFvrlDQgXNp5JAzGx+Z3U2L1YReIPtJX0PkVuEXi/GodmN4IF+Cg7CCxtqhq2oVldWjfhp8v
73E8vbXefKN+JQuVINy+D9qvrTkda438o93lQYSv4RUHwsQCRLJyVdHAlGqzJlsjVOqVjyRmYoit
QWZy/+vvnfzP12U/IajyTtaMTDx3e17kJC9OCafgvgx07ycpIMap7qZty9zUc9u/reeWxuYhuocs
dIRpSBpbFfOhH1uqicf+ylwnHvr7nAY7Zus6f4BsQmZIWnJzTAUuLip0jlpkxXhaiyLsrBXuc+uM
aBpW7Xr10CQCf154GiMoFr6a/G5Aj8EYdJg4Qu54qy2x2wbmUbeDrbXESP1O0EMSOiM5UGtBiPAS
I82lpCdU3OEizxhLxGVkuQkPajOnogDpivm98GxUG9crLCW4O4iFL662mOA5L2cPaouNOxk890Mn
Yf0bV86C25lJpE+QYCedxzeeqdgbtsAvjco7MWUibCBBbl8a2LbO6fB+VyF67PmDl4u2e+LpsyF8
kPfwjgWhhuftHwmT/q/p/gDxmQGY7rn3Fzmw+yvvUL1XMlf/ZyaWwI+/6IHZbfuCRqarZj2bua27
NyTqiT86vQTLGEhKy7UBKyId9+9qQKVqjimHwEoyJzswiGsr3GAi2NF07FcayCiI4RDoNsJnX9li
1ruYY3BbwpjB9NvFQC/KPs8nav/q0BZDGF5dHYuX/p0I4siX9uoqUqMY05wfkSIRGfVl37dlGGBR
Ax26oCCF+Ek192HHAURg4RxKb0fnu5OGWsebkgLnX5NbwGj1WKZQ2ASp+YFJf+BdFFiV1GL5GLj6
bEk/qtgW9Vua6UCLHpvzZMUY2eKRCl1Uprii9oDL3bm7vGFBaAH7QF+VYwI9D7A2WJn84/vdttwk
lCppzwkB1fy2ju5R1W0//qk9BUV9lmRMvWB9R3Vyhu1gPrsfPkrR04L9L5b9T5zwjdogLlsQcwJ4
zRwjwzEzUj6Ln4NapLyDOQoHZss3bod+EzyVe+LvVVFYKWLaYNSOVTMgEzICV9EfJOKhA7TncxhL
emgPBoYPVG3fc/1MtDh7IRFzl7nZKnGTJp0TKcVnk4+zyzaJKGaJhxGL0X6hVeV1+1vMYk8PFkVR
WAQ5pN/njC/5a/58cJ7cddpT+LvOJXWgJO7vJCuvLfkA/vN96D8r1UWuOAJX2mtt9jCO/aXRgLQL
25r3Kq/wdliMQOZE1OyfbrMqxz6H99NzXYTGaSuQU5UwozubCvaADUIsmROZtwzX8BniEBt9TkR3
wdfK3cYsPkZx9V2FIBHr0mNMVg/VSLQfdVN1cKMmJO6twWiDDq6ChKah3ZbJElVrgm0iVq9tY6TI
GHCFYE0PB8EZH0fKJr7mBjLeDqDt2g2A9nCoVn+uikq6eYjZ7h7dunITYZE1DNamI6PBzzoq4brO
08tzAAA+ANxuYI2imPEX98OxZEvTU0C14YwYQDQDYNUq/yMBQmk/WKiPQ3iCFIbZelT0nrDydEdQ
Fx/FVzhtS1ewFFTduK8yUy7g4ZSKp+teyRG3AjJHyUANXdLjOT2c8Hfhadld2cRU0gfVD6trgfZ5
Y/2ZO14LTGOgSgFGwxSqBDHvwcA6WeVkbi6KbloDsoS+z7ziufgXkW8WvjNnE2Cwh9RGyiI5ddRm
4FPaTH3xE9oA3LZUAUccWam96gpXetV7c185h/l6Hx4iY676ZHqAEu9DLqkG4HYVl4jFrzhINLWR
3sZ1IAOqJ+H1h1VcEYTTJWB198Xgj53LAnaf9oNEl7c0CnvO9LXshP3yqOcI9M095DhHwYZTxFvq
vAeM6dDWAesbqU6o35/T3GdEUGSwsdt7ZTSK1QnVXMU+3LsHz6SnaT+2IyhNF6PAilUTvUtWuKVr
gglD372cicIhCqASN3Z+41Xe34CNyLZjdUBgQ7ZovvUw8x3jEV57bLZJDTtoURq8yHiDsFYpLPYr
G0ZPjEOiISuB9Se+sgfAlxoiHCpbIxSLsg2REcbp0u4XYwG4Jcm6S9N2bLqGPJyr5gu4kuyas0++
24lHSnxqjDOQs+B6OT7K+tH9gRoyDhHuuVlldE7dotHGxy0SKe+mbbx5qug0GE+kEvQgrKtvx02l
6UNM8W+JRTYxDMSh8Uw+E7z2upmJpBMyokeg7/m3Tvv1YYXr5cI5K4HnjL4OlEnRosM/FA6uy0Br
GmgGt17edDrM4W3rlc7yUib62YAb/0vzHr906Ub4ptFMisNkCyKJ7ks11i9bq50QatEZkTU8oSnL
8FqlS5OOo0Nj3Lt0c9JMwduLJ1O/bmiEFvvXp0pf8WXrJwqAH/8yI3m1+D4uoxsV3FOgB+KrZd2A
3eZVk/nbPA/Hf1FJBsDYG4AG7G1LzrfSfOg5cdAeqU9RF9bzVF2Ft5r+TA1dT9LXMqcfySDxudM+
LPNZzpko+LVukSznUgOoq1QfV7FsmGysisoyo4pqM9dZnxtQWP5o+s2BvwZNvJBx6yVBA7ylI6be
rUbrslma4756kwod24J5ptGRwz9rgvwLKNU/YjHxhSGOoW4K+WSy38hFo5Ln8d3zupyqWGSPsYNQ
JVI4lCLuMIN0jJW35NcQ+ZzZptgsg8Vw6zuStn47mnDpE71/FeXLkauFKFNNtmoMOLJy0CIlWhFG
k6aCHQ2MAf3xK1OD5SZxaFTURQhOsNKG3HoNl3p5ZzpQRT1Rz1bJFfRpk5/zV8aQvey175sUXXHg
5Yf28aL9e6Unpl1v+6WeKalpWe6DED3ckDfzc2ZRQDdcQwz3xkdJWnCSck47hinyX8lWfJlAflgi
8KMWPL82VNPWc3BMoRlmpq6fH2AeWmw4CcWJ+4MiJb7Y0axP3PjeW6y+kQDQ/RFbVfdXjRSFBJrz
lSVyhujxBsMMCW8zK5x6v3PktERyonK5hi7LueUx6VzaPJHqy3D5ClwOO9vcHZCIjN4oZ9QeclGB
ygii7ibcPnpY/7Hq++CI35jMZzfwNaKzHYRgfxGQSnUm4U2SLrPfIGhxKoi6eaoRHIbS9l7IIbwU
vC8BEj1uG1nmcZwxDvv9NVwq9JTwXGFChamcZU2eGcyrg0sTaVljkfY/GkgAnzApuVBhfAlyNP3F
iNMmWkUsJJWLA1aYh1rbB0VEwJcKIo96c26x+E0gTA3y3SKq7eYaFMRy0LcaiaCvV62EUe7c3ai3
vPSTOk7KvDY8XZNfC7jRuxh6+fOdVJVCeu1c4ib3QmqFYrLsoZ6AzisoTLZF7W+Lh8SUtTkh5zIf
keoBCocWnmS4tNzMBQwWXljebQBxWVqhOfzikSWXCU7vGIJgKKnHf54v7PbIaIWYIlfkEirOQ5Pg
+gvqOTHEq4xm2QHDyVRNN2W4u8eTMLGMsXjZUwnPJLpBGCyHW3hY+HZNdQ1IMWsvjjcvWXmvXTbN
Xm/neji/5fS1fZKm1qMPGkvbCSOymlH9aLzP74JaDYOspo0vpaqcLzWZWZaKQqtQmkR7ezqE1a09
riJ3XnOj8B8UW/+AiObvU/dbJtOxxinLxb5c3MEgCR4cYBZQRuezGVHANDb0Wtw5SwWYQYspzkFN
mbAWtgOpQ+Zx0WcquqbUvDo+EABI0MJyVtymkaE+MlG0EBM+1mKTy13lBp3qKuOxjdKBcnKmzK3f
k9bc+5hcVa1xQpNi9gXWy6LqhAlwHYus8DpEDsSwMTpk/2bn/EngcUDHDRIMbhy92vu8jjRtuHao
FHEaLzTAbZbDdK4dNT9t1x97cIicqYzLbciAdNFfeCi1gN03cNhED6cmdlbgIvj1BcCmPKedTA4n
M/nA8ALVOoFnodFFlCBFpTkCQK5HUtSFIexO/V1/AkVOTVSUKw9ZsLfIFZ9xLQN78a+EdZmbAWzD
1u1gqq/NmGb+S+4+sNKkx+RlZ7yaC48Pv5XyhacVKzdMOlO2FPgI9TEVVo/3Uuxl3AQ/Igjm2XVt
i+exw7xkRR/zQmTccYQsDlGhs/tfh7o+oIDSvgquObfGry80MUQvc8dqru8ai5cSLXyRY/8T1EmN
J6eV5FzrIR6pxUEAz2PIqa2EpewL4HxsSk/roP30gk1Oy362GBboh5tSL7qdDvJgqzWHAjOgaebS
x/j6IDoTYVfbEGsSHJsSQIQ5NyxwpD0SRE46IA4+08oFa0qJsR/qJFLW9FyLq+hqnitCfbxb83vU
5NeWpVqqmtuXXLsWXavy/k+I+eQiWMMN/pROwyuTzWEFJycpeHNStNIQZcgKbUDsm8NVwhgtcGCj
LWsN71RR/pvIeZok/QuM7jsTfRGUgfJVjWKjw5DsNwDZncPUaOQa4hmg+iu7Yt/d3bXqpm0PBFuu
jFeo7bqASSc8ayjEp9231TgYqIf51q3Vh9TznqqP5VaqD1c9CAMKHMpOc8muQF5NdjONY1GeYW/N
rOgRCGz75+ORIS+EhewIx2aNM4XRTyGItS2uNy+IOG3KEqdqjX2qWhPdxPRUQuifs6652RNWxo3S
mT34F/pvyBt1a27oravy48QBnRhDc/8DyiRgIVa7w5Czw4oGxRsydn6Ws005ogeWI9XAyqxKe/cn
Vj1+WTz2/t6fBqcHgSZhTiYa7EAMSFNvyWVE2KPdnx3CAglwp3BcnbQnH3pLitNoe0K9GLgxD1m4
smQlKU1ULYhkL4sycr8wFw63fYAjWJ1hSTXoFID4GIsUTPC1bWcV1dPGYDlYVancUxhOo7sSL16c
S1BVhQ5w7hBi37OFmYCh2tWj/m6c07f0QQaE+vmu4AvKkHHbl0GTlu6iDiFdKY1gSp+HjkpkAreO
FlySTqpmC4wQkiF74iuyrcZNFbw9H4+/9sYUiomONKNBIhtbwapX8gZryglML8yBe+nokLSlkGB4
q3M5QwIs2rhgH7yppYNs1MP1Q7WdkKFZ4bzr4hkrzlpHxYqv4NG2csy0kNZv5VMT80TsD5fbXZqW
kYml5C1KL2rbIs9N9i1rTiKPsXhzvL7YyjiFtXvMjBuVCQg5DnKNBOGdofTe6C2U112yYmSA4bVv
ezw05wiaGbh+FeSuoLGzHYTe4crDnfxNHktAaDRbHQV/mLaccdNupIUHu2x//sXB/NMRH24lQ0Az
D/rN9iHTzSiX/Iiv/nlfndvqzfAtUKuW1wos4lETYmj8zaNVs88HOr7GxhFZyP29W7rk+yp2AQRu
HLre7K0WvAejs3acVBfKSPTeq5FOJVgcLC99sraFVGAYA9XhRX1Z0nDgqyTuVt0oKwp118kr1avO
LpXkdgX589WXsCRO8ogQj3C6iQRaBWZG9Xi4SNcDcW51+F39693kyb5hyv9KioBk5173QLZZcx/M
faXzoNNrcyC5O8t6PjXBrrRovFzdLWqco/FFQwSEdvZuwsSXxxZTx+3XMyndKePacqDUDFqlaiFG
ntjucG5tZATYxRbFIy9TwoYjzYnBhhKHExuGkxpaeNBEmX/ROOqAU5Tolx9BnY7euWTJBSv+dkm3
hwj7Z8oLga81LROZI6PQy9y991qQJOKc4rPIvDuk2yUK7myaZYu87WzlxAhiBMAyxqGth5TSq6j7
6eWhZEiusB+MsEfOiCmgTaD9NdBgye8YkpdbxXjUC77ADHwjULniw5ntwKEPD7YLZzpQnM+Hnv7F
7yiDAyc5u3iYog+1+bjp/16iplJxhgMqtWawWpYezvYlc50/z4mTRoVIm/PL9u11KOqZcR/Hb+M+
XBQW00856cHGDRA7GBgVnnoMe7DDhktU64cczjbO5KvrLjn+zuPVrH9MRc8iYKfkX64wnkrWscJI
70m6MCdIceYhCQEcFIGxOMIUKluogGi9b5Ez21l8b6qkwCYutmsoPnqLRUlGNmMiiosbtbj5AYmf
hN/pOXohsWZkeFead3venrbwIBp8789HZ9jvDuuWDc+dUsiqlpYqaWbmknEsBNayp5ivL2wC7gjH
RoPPqleWDLUbKO+nBNrMr5nLHpxS/7yp5rvJhm4Bmfx5bUe7vh28hY92j8ODOLc76yRIszbqwYCy
mV9X8oZU6mWsQ/hUb0toqMXzRUCfq0jWNPMVMqg9eFQdc55oqqw6sE6qnfE/4ZWMYCNZtYEmXn80
UxNL0lhOtPB8PuNZ15vv7a0Yzpek+Gic1yepjbfqsqG7/x7m1H6D9lUW5kGebJQfhpNTU5xtPNO2
hdnIAbJ+GpmpDXjadshP/BydWQKMpj5jK4QfCUqxQ2BT78o7mzev0y3wMCS+nEjxnCDcClAEEytr
Wki7uiIL0lbg9C2NPBtugHZcLPHocBPYWGAR0y+fUqRe/8FWxTcb9yaxDZCvdBV6Czul7GaKOlfA
jFTKGF+4DlXhh5+FkI0SZV9v2ubA5c9ghjrPpCP5HbvVdFJ1W5KwGP9K4Iu+J28ZR/+S+ga0rUOQ
ch2x7twmhsJM6r/RNug8DEKg1JL5c2jS/qtVibCemzpLB6EpQ03fEQjYmVhDkZhy87xC/FSDETY5
vANJrWhDavm8gIGbUVnRWzgayhFBFuv9rIjEM8RtpOtHG4AjG+EcqiUf/+4qlTALBV16gA3DQ1pY
1MJQGJ7p5XrLT8YRjOHsYkThA72CwAupvwBisRrHj5syIoixo6phH/Zy45SBxRAHcBTDB501xw1/
VKMhuNcw61QGMTacsLMWsPMMtFN0weWO5Ss6EkmR+rpUrjs1GrAxMwjA9TSMzgGOuIU0gs+WH4JT
Av3RCaZ/lxMs4QraGUisExqsL6gIPsD3WHRtsYVI+4WCVtT8mlmiZD1MaZ2vRnIY27YpeF6EH2ce
2sp1BRI3L94QTSRsa1g74ZILSUUaCVTdATz8kVAo/lqxv0Pko0J5RX2uylrim3FOnI87ZC21CJ+I
lUk3tF484mSunK25ICpUTNH5VFvuaY3ETUR5v0UvP15XqGjXCqiFRbxxTyPO7+LDU8CaDpzuueKq
ahvrwXfQCBZFHakxrz+NJAoxUn6N1fq3el4pOiJ98fjqa1HvNVGjoOm9JMBd4zhysSqDCS8dFvhH
mHIv0oMExj3hq6BCf0m0S0Si+X2rxIYBLMW0hTWQq+zGVuNFz3aBxWNFX2rbCNQHK8nj4/0Uvi73
AMTVy5lX+n3mYVdfBp47NA2xfHaH4sQGJhVSUnyuY/g+rbAqG8mTqSyk6k7/RB6u+cJ+rsE1xd9R
eNU9kwiU7RmOHH5AeU9AVF4sPss3rXBmNU9MneEk1RKMGB9fMoKkeOITuAX5VM2AzT+AOl8ryJ8x
kXjwoNJ/yGONWpVgGClbVY40tnTuMc5dHtCFWrPazD/+cyYuymZKtMyZeOgPP8J80P7js9oG27qs
AR+Kc92Hwe3BbGq1LOIEj7vPgiYd2ObAbfYncs1hYbBVNHKXvh7ouTaxvBLFDW6NSfI0khprBLqR
+Vwn72kWphEsen3nB3kOyMrZ7lN4Zuza9kXq6TmSWGez8BBlzLOgZFC303uvmBZUStAcdVs9UhAd
qaTA0ABks2uNoSesPspqfgjGeaHCRpt96+ew5laVQOmM4SNswh/FlwPKhL/GskdstM6t0DN6ABBe
v8iiX7RjDcHNISaP2htEx0+F8vefo4RO29GozW0RiNv5vZlWeLiQlu9fBhT3FGEPo3GG4qIKzn28
ydDaemHJQMzLFtBcdc9xmyyOxeK9EkoyJ1aGAUsLPnNjdSkES8dKcEdsUizmuZAXk7+Nd9S3MWGM
KNpBMXUz9nH5M3tf+a3NqCNv0Gb/MkXdYctkswHtOQOau1KVAXjJe9y4R37bYS3i3/zJqDl+CV/V
ZzGpU1AdVBx0MVdTjwgliJwkhT/ow20qyDFl9qgbGwaIMDXbH4YJtb7wW54btSOj3Ag2sIv4wtLQ
zGTeIUR35F1i7frZLsTZ5hBDZ6CzAu8yZbSePp37iiU1pY7l01AE3z+f4Dyvnqj3S/Q+9TbYdFfQ
tb+Ppd1R8OYvo/nPVHyr35fYxK49fQUcgyxentR2ctyNPkrBwpFf0xO4Fh54HkkcL/CFff427DoQ
JaCWqYC90hQEAyOIKo22I8wopvoocefh5KTEgOHesUGzcMkutYJs8w0bNsOl8vO8XnN0ULqlwHSx
m046qPqORVRlQhB/N0WK+ckoUEWG+2ZFfYfqulQBezIczNo/W9P22svOeQ9wBHEwl1GKbGhGBRju
OEmXnw4Cw0OIpN6PaG4KtIkqrH7ZlEgXDFkJIcYQe/ahsUh/w3P/cMq/q/hCBnr61lvbNHmEc2z9
IJwDOQuokWfT6HrzRTymzQ3dpocWnc1PoXJ60k8MCABwEoMts49j0F/0ciijl7+2YKk3Amhn7SqR
+b6Av2jnVwimxqk1OBxXnlzAr+9883xSholhHuWJ/kZfKR8gIhYvoU33O8Iwp9eFpJiafGvaum3X
wix7CUK+3pi0hUOcPuiAEr1NYMDWfbwc3ZZmvs5OSYZRfv5cJeIvTkPFadml6zCuBnkLBWZnFYrX
PKNgTDdodS9xo8aXGgfGPOLP8z7sUfx8gnWI43CRfoxd/V8KdnjQbm0pzQRPWiXv5ycrH/5EZkYV
A7t0TE4GDCNMUq+7TVGTC41ChwthBQQ0iy5PJtJ30OmFDh2T81y7Q3zhpCUYWPufY0pMhDytp8tG
yaA5lOOoqvDlamZ8Sbim5HBsAolpdEd19cjVyo1/ZAz+Te9JoDDt9R+GrT3qnN4+3O6FL8PcO1Dp
fjx7FOHJWeZiOQRikcOLPldVR0wFvFyzW7fP7m6F/+VxGpgNH5ne5RYz8gdzu5MOFNzjDsk7GHJ+
oygWsQkfWDMDSCo5siMLpzh7f8JnncckpN8sb6iFdrRm4/4RMVEf7Vn88KRejDNqR8Wd6FpDpfcN
3H6VxWNRbPFX5rviWE5fQmU6t+LusCyB81GQEeV8dfc8hLcpGLd7sUU3UDC77fH6VV6fRc/Ipp8I
/7uAXC8TBH/RqiPIE4MklLih3Zhz5d5NekNH93SR6wX7yvrvw49hc/4jfijeEc8C3KHR9RY4Xr0+
2l4EEbZAVbRBbXhOyiVf0sB28Afey9/Cz6lpN2b833A9NfTg0zHWbAkbDQQO4wbjZ0/jnmUorSd7
qZzdL52xZ4wb7Ii4xZ+7LT8xA8TM6AEsQsNBJnZ5vzV/g7q/hj0fEKkybMbVtCVEsqo6qGiFhS/t
JwzUc23SgQzsLyK2rLxWoTsFCMY/7mWrmWr9fsFhWdDSt32U7raUaSQFA6p8uWb0lumFLJkN05ex
adBV/Ugr9Bp7174PKQLn6uGReeewOxSJPaTo8VT2fr3XelIo6Wzu48q7Brrymu6jW2irhQ/SrfmA
VtztdiLv3de4y8g+mSToU4MTCGwzdUzjMrgacbXeS3i/XEpk0H+bvfPVhAeZ5SD5lPxAr8fxcDA7
SEDx9QkYHQ+glSppYoqbresVbHmXzvj4jYkn9Amny54yJnovUAr1bNOE4oVr77S7/tftPnds+AnU
kbgXHQeIngGVuedeEqD3c8ZU23TkIulpJrrYi+RO34cETl9ws1p14H0eXtDvXOQ49UuW0GuHkf+x
Ss12nSLym3jgGAsTj/P8mwb0iGWGaPpJBOkX5NMzVICqm/FW1RDcI+V2DdcVs0qspxMN831kO7NG
LnOm9mz79/zBWcDpikostzAdF690PELcSFqcNA2nkEX+FAjdxcf2u+BkY0NNBBw6N2Zx0FzM+33C
NxIEGzNp++RUbWKLzXRI2pKyet/ehUxmdABM69WNstgwH/qDvJwOXPT61ED2aGYAekupNDQCnp+Y
IIgwzEWBWVFemkEzqOqkWlVgc/T34gfi9EjflUGCWSIImV36hlbH+pDLv9vPCSKF6SdgzaCsS8QS
RVINTXWSojYrQcN9huyVsUcNQ0HKQT2Ei+3EJM0Icr69y12qc15EEOzMcxhtccovqg3fKVogdpaD
gyfbNLb5ogMoJTlSrfn2XE9X9nm0Vqb8XIvu0NnTXT7T5miavFsaDkewDLrBq+ENenshhQErSKXT
OB78GtnVkL+bS85AdFk/j8pLKOUuGdkiPLjfvHIpkcH1CQ6QLUZzXezbL1x49UtCtz0BGSXxyvxf
iZPjmo/blCm+Qn2Fvof3wAJccVeFx/REFHzbmCnGvsXy1x2OtxNHPHV1bRtHbmcWVeNRwqRXDTS4
c2mlUnV+5j5RF032H4f5N4sB6Gf1TV1yEsc0Bwi4iqKoZ3Q4N/2C7udGYx7WaxrsFQKndaZOokNL
ersrH2q9Rmwyo3+KCIhp7XJI8ULg/EFI4bW6S0bhEb3uOhawlkNV50Y7/9n3QgE48GEqQhhOT2Q3
LrUs/SoD521qyKOpJThK8deqeqX+R3R9uYoi6m2BmEGQ65r3YuZ6fWXuOuImc2t7kbRa5a+8VEyu
vG2bC2DYIGbH6ZRodGGfSdrRTdwPuFtt2MLXMh6GuLPrwOKKH6bQ72N2qFWbeZ0ofTbYoPZ7qWll
XxlrjvoGCHXUC0BI9DSPT5CH4i2tla9tsoFkMK3hzoQaMLATv3lRqlJF6cbc7TOWvdmnOpAX6nLr
yRZluvksA/ZnwpU5A7xc92/23GDlJpKZ5xW+URF97YS9UQ1+uaCH9Qw32NDnPUzTEtuwSfwwyqbf
WhtGY1lvZHb64CLwyT68dw77kR3qa3W+GC2xfi/ZROoNALEj9/Se4C/R2Vyby3JeWynZ5Gt8F1AX
p4gp3sv+V96AmhbJDempfgksLzmwpH8hxzyXBoSpSWjbDHNLUPQshEiD1OCp3VJZh+YNgOaG+QHK
6BLmNQ56/3MBEUWF+BB0KPnlVTlYIpGruDAM3a6etEieS+UuEANcf13NrWBQacPeh/Y8wDvTav4G
9qQA9P54Ziqd+CZDx9XzpRYfSESy7lniaTzZiMVXEkltH4l9PGkDdD/ylTpr+2kqgzdz5AwZtCPu
DebleoUBP3/1UUoC0O4HQ09nSwejVrkkfa9cD8iWs6QcKsZ24GSkPMmNS3avrB+dmL/LS8tHeLiH
Th6ZYLLqSLavHzcS2+ZF+46rt+ulRBPC1wvHdq3xgaX6H2cMQ0/WFS21mA7bMVi+2NRpfqUycMgg
x2Oox30gTx4CCzP0f8hQQ6JJFlKQGna5XYIXY98EXCMAqjtNdutotqM+xNZI1iA9LG7qM0QS/5yF
qIoWDMtifae2moVpii8qoEpjjj++tMKu6k7vvhULmcmUbwyB2LJU1M4WkkCcLYVf8Bikax/a2H+2
xq/plHSDR2b61Mu+wOApoLHNL15mUWgLUi4NZ2W38afyquXIuxatUKomM8WqGQPTqZuNi9Dr3+Pz
ZQKoxkiLCaTdld9TWWClFLCPgGGQmhZ3/pwJiE2QDxwiQhJ5MoJ312CmJdivpdwaLuyKZYDy1I3T
6FST+hxJxPj7qSlqf7EAVA/6eB9JoMlNXbhuRn/KUmfI59q21YUohXM8GbIb/O4LKWaIndlip8la
rv2EyNympXeIBExhsCEuM2DgXHwh/VJ8LpTOF1tGJNHRHUWyqdQmYUZXEUOYSa1FEqYRjIegqM5X
Iw2lJVp0mnmnjPrbPs+V8FCJXtHrC7hCXpqVZW5iHS0RG7eAVbolbpDd8bHpPKOhOudTPvI3asvK
puLpWLGbT8tCZZIVbDjDBeZVKUPxDm03P6IcHoGVMa+ofqa/Z4QvFg7KAKKhQcc3miqnQCJiugSc
QwoX+M0OmtkpJxwnvz8NJhs7ybejlZtGBPNKc61N9LW4fW1HJJ8aVsg8YV05uiSkfBw4OloguPSH
fWX/iFyiswnbb7kd7g4FRJVL2ZEL4HZxp0BNOpFYAd76hQdtE/SzHEFaf2PnYogK2WgwvO7IFQCK
1NTI0ZGGsrd0toytjc6LlnHGkfncaOKz+Ar5G1EXoDVjt/5C3uhHiqrf2yvFtiKsEAi0kZNpRk7E
Kxjbp5vuRqv3XIEV27t1xjY6F7SUwN8tG7dxCsVYvAl6YyQInIxVEophdLPQTJUFakGUwQHjOhXC
FjQ8RnRd21ec5i7KW/BTw/6ag+3MuLsABMRWb5RSCRzp4V6BL2dHkYyzdXTEiP5rMVTpsjq5oeYJ
NN5BOpRs8T0tyY9L8a9qWLrtG2ypBx/0CR6nWdjt8MUYD3r3Y3RyYUusStKV4j00LN3WMXseyyzC
7Z2TmWsWKMWGD1Y4sQewvt+D7u78yazAWmt50u4X1A0a0q8V7vrc8tHsv60zl5J7+9uobxMmjOU1
MCSrsxueT0hoPKI/FHwSuSLATiECHEz44pAJhunBvHX9+tZxC6Yb+aQHwji5/8S0GH5pQ9Q6dR/z
R5Jusb9eCoyQqCDmLPLjiN8Pg9lmKswHc5gUH7GHFkrqGKW4yKixCsEG0Q8WM7ydvHZpSHBvmo8h
a6bS7JBb8iiW3zb5nU16Lg5Drrkgjfv92vE29azVSyX6gYN73/RJrYXkqa4TwBwpSEz3JhfDft+C
cq6a7nnALVaSd5SD+VWveacTXAB001fjz7fjs/cfCdU2WkLcol5v8512zE+axLSeIh/b+WnMYJ4e
3M1BSHwGxaWpE6hqG95GAwG5TwVXVr26TF0vIVOaMwBMEzZzEUvpfunaa2Op7l3yBmLIs2lKzDrF
FV+o/w0DR9UERuwUjDIxOj2d+Bv+s/3Mf/mlWj62VkelPRUBzuYDxD9ACZVXWOj9kbLbJFvv9a7J
9R1Zn6valkstfkI4sMTlnctHwqElmwMsrK+4YayWRsJmwrpba2JcSbnZ77JX36hDKSAHJB0rv/5p
92FeDIUXmdEpv7pvl6t03VMjKK+I38za3YvZTe6vivcjBW3iEBO3ARGN1zvm4AtYUUiW13udQ5+0
HFUZvz6tNjFzgcCp6d+Vej+CRa2rLsZv7EtZaYGdBaNSYRVsh0Z/W1lJU9/khCCkmBi44ZicBqq7
SklKlQAW6r9L8YArh9e5J++TZndqFBbzUsFAJn7SZTUQo7ckiAFuFJIiJ9U70y5UVvuTwRh8K5Ks
DREtELrD17PLHmTS6G6z2lmF2ka8LXr+Mt5iG9Ml8bY+MaxFW4+ggW0KlMe4GSfUW4vfjuJxrSh5
EZySQCSIeOOJaxx87ohD20I7KLqndHTDRanekJFjAaEWePyGVZlbUQMBexNq0b848yBObErUf7wn
BrEKp9C+Lt88+NLyD1bJ6kFRnba6tWoK0nHk4s0Y/LSPrj4rrDd3tiYL4PzpzB6Lru9mbf4RDGIB
JC8kpZTyAxUgZ0fiGhG+UF/oyucn/MdbBTor+NBWy/SYpv9n0vaJLWyMd0dGo3bZBNrPvIzEnwGj
st4PdWsSUMZh3rLXPyxI0jo+FPWxBw3MTl+DZJAGS53g90QrrdgqKAz2PqwRKHK584g3niGj9tIx
YyWsxOVpd7B1c6d39HSQRktWnOharg1L769QIwRmxdvYkpet8zRM9duuY9yRIc/wwGrTWPi0Vhxl
9fwoWhHgK8SVEbrcAe1SiZaMuMNW8EmPjBdYXKqdgSSNWyiWs7L+6DRuriZFI/oop66rlBANKxtX
HQG6JNC9ZI3kRMjJkzP5dPfbgx12NAIIYcaGMDMNX1aksomDRu/RuzjK86tNC6tBXhDgJsVlWZHk
xLjJLMaxBOTsCf/8PBw59LPU0luCnolPvyvzaA0Eb+9eAa0f11012AAaxFWHqRNBGjw9JB6Z1lrv
q5yDCMegfErT2mQzJLdswub8fpMhFcP4b/22KYvoZQzoboOvz6F6+8OZBTXgVIZIx2nhPeBADuMu
pS2O/MKjygEK+yS0F6DVgrxvBrAWj7PQJ9bibYnOlyjLfkjCYuhdOaKwWu2LFucbOGMtidUp9zLj
yWqsv2HmS7JddN2nKg/rwQO+sTwGznnMRR5I2NO2TWTbRTMnhCDc/zUls+mH59GEuw7xsW73DI/9
P7zzF2x/3Vj4PFsLOHMoYiGhEkhVOaiP6KTi0LWgU+oVgDDxFGa5TzXYYFLpnC6pgP91lovNBrID
2ka0sv+eyxqdUAmGdHyCXkz97iGjTUkEDGuF7jL1Y3oVmo+IDnv46E63PWVskv5ucyITZH2AzcH9
UzIC4dMREqSkS3lYtskfJ44w7rog0SQRpXfs8WzUtMUJGcaM8uJXKjQM7Bt2L2w78jq28xz6XNYH
FB+wiBRBk/GwSWniN6ukn5qw47dn90qBvfZrHAYZ0Jq0BdFQ4Y49o0luGL56hY7R8qTSUG6mgCAm
dF5iutx0w19kXL3+1eEKBL59S7V3RPN+cR3QpQLwdWMlHLGOwgmnk+RsXG13eWBE4WmhfAJDQ3mq
PUGkImpLBpHOAUImc26W6YThxqBqXtZ7Wj9NmQAAhF5+phRo2Hrk9mwWTDuekTCVKZnNfXSTmsqR
NGg+f2141Xcy3BX6KGrQQe/eds5ML3I2W7ZSQAinkJWRClDeCx92IieICs+xTGVGEC+9LiZlK/tQ
U39TFHy/pA2iYW/7s6T9VYv1rb2Vo/nzfn6909/DBo+zeIVvzN2Wtybqj1EAq8hwWr7IPauuJBvj
oxescKsVCvIgrO30sRllQQsJJtNzMHg16Pn4lDtBzu7mKeO65zUTdVNQESLMThNZh60J063RkvFv
V30bIub+0hwtAozhTj+lkW4+cuvpqjoHSpiTFPYLn4+YtYGSUwPGoTHMu9LdW4fffi31ixvraZjZ
YMjFjrCo4/yXxqSWJconMCo1BPE/tdcQyZJ25AluvB8AIBSj2m1UxqiMo+WehpU5VJkR+bNQ0tJy
jtig/4TEWEq7UrduTC+vnxyG1fBfVneLQlfXHCeqBV89HDIWoAkS1V4gLvdDJAMBbD+q80Z9EHF0
Y8aUxU8DFsNt9wYo1O0YiBFWYQ8JOxV0wE/H9cgGOdyfR6qvITfWZesCIO6YaRr9a8lh7iDJEbLf
a4/isjvmRN8sS0SjiHUWAJawXe1hbbA8H49aB4r7nU4DTQZAZtPzw9yMPnm6gRrgNjw6YgVmi1QF
wb8dzXP5iW0OJrIYZRPeNqxrBnC/JCYxRNDKJi6LueN/tOCl3S5C/3MMYo5k86Hb8r3IzyV7kzHH
TVZjwTQcqTwep0aZrSoDqUNPFIereiSXTEenJfBU+uqNnTdMXi1VMuaV6D3AxV4O60F54K4UEYYa
93+eWKUh1rYsa8z560ccTKmBBmGIUueWdwI7OoDwcG9CmGTw9zqrYxek3ocVqOfGEvnFG1aib82a
eMgdpoT5FvgivllgyHNo27hlU8d+TSddd0CrDUP6obR3FLKmshoO4KnRVa4VEbPQ2VFa3fzu9lRn
Kq3rUDRBtrF4p4pBkUagVE0bSGj7BETchvviHlze+V1kLaA58A3l+4RCWoQmEHhZcBM7YdIZqcCs
2vpFzCvMnpbt4LtkNKCP76XSWUwGi2xFqU50LsV/ZxOPmnRsw+VVecmu5VEFjWMzRKyiR/KtKow0
Ds5+Wu0RKobEf3sa78nhi4ogQ0YCZGxIXWFzFXN2lxE0q370N+k3hvnNNUJcNri2O5D4H9AWwLgS
WCIOyi0Yq2QPGk8egbNY7x8fTI4h27Xtl67MlIQpyBZZvFFmS6zsI4uVOD77b5n4A3CCBNbiiUfl
EJSExZpNDDCN3YbPGhgWaaXJ9VJgoYXUhKNLNSUVRmf1eLoU84VClPbbfGwYkSJETM7VfglHnteP
6WX0NbP8xoxizWnonAenRr4QCaog+7BfW2h/NzCxR29vFjSWTPTAOzQgnCKDp9dyN+WSEvX3jOwD
gkNAOTdi4/t7vOyX0no0T73skIroD3jQFLbFJ/CaHtKRGuVt44iRBE9jSZOl9ZFP0BblDZqC5v3P
2ApX+5Z943m5V7j7+EaOmu5MI1tjY5yVtKWf+iaDAcgrkTZrUnRsmRACOSlIRs6GGfQD2o3afy40
Yv3bnDblf0s3JlDvVT1nb8Lua2zzNi+1zrOAKml8vZi3tqoOVFYw30AtN+co/AaN4rDjJAgvCGxG
1ZktXYDtf2fAt8yhtcXdmyCUa0STt82APHj22JylvRDUWx19PD7Qipsxv7a/qyU4hJ6Ub/fC7vlf
5iT2osdAGxmt0UGXE15eZj6BA6YBIzckFy9fNC3E7mvbvSL5fXoFGoF5G6ZUSBM5s4NajvHuVomn
aJVM7lFvtKSSWA1VcCbh90zoA3iHoxSjqJqcZhqGWIHcUiUBsBgrc8rfGr7K5H1QX+vGlmKquGcY
L0R94pt1wmVTtjZthta4iO/OAMhCNaKJnkrFgBX6qOo7m0UMYlG5+MCl97/A3VyMq3KIAVMUQrla
YVkAbF5zOKV5tWe9+yoaD3WUxTMVgZWTW2XLQ3v9NbHXroeZ4W/IsQwW2Fx6ADt0T7iYHM5UqGLX
h9V8HkaoE06AJHnqFHRcAPguIAM9UvYFxZAvAb38N+7jqhMgt9WY70R+zvIjOXPYUDS0EKtHzdY1
CO3tISkebJ7C333H0kRMHH3bRYhtCKnXPh/Xch3+jQGnH0uXFClOcNAFrk+EIUxPIWGoaxA9FBp9
X0C3q8IbEvbE5blzLV7MSnTAUZI+BftE+G6rpx713FFovcZ6J3pyk4ln5FvX9wjzu9BsBEDiWBAo
x3nv10BAvpLDZct85KwbBR2tf77Zrl/lCmpRdnJUt4DKoXv11y/JR6FQDecQT9PcO8+vxBzOGBCd
7tsdn7U7YCBifqv3bnLYz87SaEAnSytCG5Y2a1z1sH+QHAf53Wo59YDoVJQ9ijmgiUmoyS0uKgj8
9Wy7ahhxWhGVk1EKxZscIW9TTDiONHjla+G8z4VzrJZc4jsvB9TInjUAGEmXF+35cw00u5dMaupR
zHtBs1eqfLy2XHMbQZOTfBrPCZ59gZRaQ354KIMRNIg7tA/X5IwCR73WZlOzXc7YnZp6WUb9XE7J
1jnFrQE4dVngS9rvEEe5EvI4Qs3AlvRR8/p5bcTHEDc6VUkE+6y2acp6sdf42WSwRgmaTC9Vmi+9
nX5w1j/s/XyBG01thq6NxpCET5nV9sk+MA7OntRq5EYbWNqa+6ujQMFxEx4coFNGCyI8Jzf3zRC+
beipqse8YgT2L93Y+jrjTvURogICCWt+VzDtNAzO8ZWQjK8/fqUvoN9MvhRhWcFZvuTKMO+klmJx
dUyMw6ibYPEzY4JHFyvJElgLF9wTQAohRj2yEROfyfesN9RzDRu0w/MErgjDOk8boLFSi31uCJiU
SEUGhoagojw1kkzRvmQqgYFM0MJkw26ENfp+QhA6Bowjb37YOWQBg04ReT4tFSe3dnhgUemf01VN
hvSfKT+W/ju0okN1yU34aLYAJHvvdPGKxM9AU8te0JkPb1oMhV8+3ZhGKzyqcziGhrVdJ2L7T1Lp
5QbvD6EFooltE9OYQLUKqpzleRFVueq7Y4DvB1SlX88ORoaL2ifZHK+9SxGgrA2DScR9xmd1Ec4s
tnGe+H+4QbqjVAN05hZhVHixs21d91BeVk/tDu5+K/HWPKjHFAJCvXC3x4rTmPlev+M6FBy99YXZ
UhP2RXhoS3LDKDpJJ9gw3T8JJ0vgWRvVnGsMXZmawit7Njn1nlT62bC8FHxqcFIvWozkUN/7f2QX
fTKD3gwdAU1Fg/+h6pcDENIiCNMXTDmaHaFTuHzBqpN77MwZVzSp2xMSLQHa7ipJ909cMGK4MJtn
I0BA8pDJo3i5n9h6bpAzM0nSp0fW8a5KWmUC945cid8XaODqK8NcZ9AOsaGBGWnUB3w+b6JA7M8g
HRQsu4Gl5TcOLYkXeJM3LasuJjBwN5oplrMmkUMSnOcdUXFzq8m5WX7Vt1irNWl6M5HvJcj5ZtKT
ekdskIN3w6qJTjsk3/4iVV5KOiEcF/rIn/6PPWq8j2iXUfweyWoUwDdcs+MRknvTRm7RRUAhGC6R
EeYMbYXgxGb1wsxWeUHzw9K8qRPXQxkrzjvliyZx7lQ2q0+eJybaYIo3z0keHMIAZMIHCHZX8aHU
5PdFYZUMcdQhyoTej/+kjTI12ccBi9JRQh9mA2F++bPxjeIybCZh9TYFZyBLkxWdKj6f3QV1aMnG
RkpG70QFPV8kbf3Gab8X3Ed9asCShQPzWUDjhH6B6lBwnVnZo48VWIHPA1zFEuwKG1AXeqoMc+Yj
mOyxvlvgJE6ay6d5f9K2pDoj8lHh8gtOGqyFIgnjGTZvaZCTjQ9qvIB16ZkaxRJ17RIy1dEx6Hbe
q6OCUrnhXfUmpBOe0fXQm6zsmyEZI7gGX+Rejwdwb5Z9DXcwnCvtU+Wlq2t9Ho+8gQ1d8BmAM/Bt
6OnSEAgBTHJymidwvLNx7QUoHvN7hQ1Sacs88PEz2BuhbxJYcJQoQ1ITs25x1G0dTS6VV0w2Q0oG
EUoQux96OIH78W5pzs+rrJr7Peeqk9ydunMe0daUQVMnSOd38opb+ZSxNRIs+4gKaDK4Stc7sbrD
/7uUG2mP7leMQx8qCVn2ItUzNl7u7kF3f7IYwJ9aI5K+6hIq5qVddmVzI8IpbuEz49bbKA/aVZlL
ymL3vCNsh5XhTQxlpw6b+P46LEDaHncBHJPMCtS1Re+FpQgRwoT/da8pF2QYawn4a61kxas9RI8o
9r3SHYro9jk/o2WnGBo6YAQ6aCGUuInl0TDLcN5nCys/az2vWWY521ngSqtUAtKSjOvYZWrm3Mqu
fJPub3vCh/QOWYcVXN3bpOgUwENZZkOdE9pIJlHmv+gLOQQKN7dm9+EQCL1Y5CPidhq9BrtEPl81
yfdC8ak/2TEwIKIWAaOmo11WFLme6icNtntFdqUN/5qp2qJkjKsFbBtp3YBa8EchX684/qty506P
2LwjfN9Sgy3BsAm8tUbefGP9qdc2bcErED9W+Qy2S1QQvddiuXmD0JZaLGQE4FZsLxK/uJqmv5e6
tXzHz8VJP4Mx/3jXc8dgzupL9kqI6fAaXSUQUm62JDX4F5YNZBfxjHIn8lCZfqcFmaqo43ZMzMO+
k4WhnXA3+5VuXJbXeRw/lghG+u4F01GM+Y9x8IxQhGP2+B3zrvKUk66a2N2kM50xL9SjMXcG/vV1
SUzuVOS3IBGX+CIpkGjoAEp0DC4kkm1f24Z0ste0sl/4f72dY3je646AmDwO/EQyGa2DcweoxFXs
A7eQjuGFjQzvd9/9L3Z+exxiV5HqafadXFxvjaIHUl52kWgS1Fs5m3ME60HGcwDTEmJP1K2WY9GK
iVGdWRMPByrCbxsc2w6USNVRCQVuFsjog0vmGTPe7NFSTrCotIp63oumo8ZP9OjbORJRltTG/GXV
8JUcLDZYC/K1HHS+CsMdc+kx1BxaLUCLkjyCJ1nWQp35EpXF5mxXHJAjbFGBFWvyL+ezvSIsSAhO
rdui7oszm5OCCyvH6TgA1+wu+WFW/HZ43lSBV6+HLXENmBBBW/wmgvn/6omBy2DRmvskDVaYWP2V
DqW8/Mjx3/BjatF6pcfGZFgOWDqTEKJoikeZCDjkL5agokbwxYQXE3EU5d/nwVKBbtLekhOx/bMq
rpJooA40q3efGFPD6FMUziRIdSRS6LQosDQvpYoxDTydhmiWqcTuyF49OHmA/LIqh7fVL7323PfN
ooKKe7DunilKZHo2TkGIuFKDH3oIU5DRl3JQ/l4/n5yeDOU40VZ2wRbzEUEiB/MOu29dgblW47kM
xjE14QZ4BnTA3YeBTy87S9xGMaVVRg9cGYoW6aaWgDo+WvoVehs5hiTHrzfi9Vp0LXcOObb76Pew
CA0TZxgSWeVhA/2+tGf/jN1n0wV/Ir+kKbWwou9DkNHN4cTP1VDXzzFwmU2DJ/4uTl9mLn9iP/St
s2/X8YNrSCUzLZkfemDTwyFrKjwpqVHtJI8V8tzhZ/Y1lo4Grtx+B/w3uNt7u1HnLGMJf5a+PQUO
KE9Q1Wsbf7PDgwXkfVJ1FJgnBdxDPgOavdv2JMrz9HkDeuyr4/fT69Hc/psHaNgBhQ7BZNlLfzoU
QT6JhLwoiCGTx6zCoqsjuEhy8kBXv7enNdARYNdPIUATmdIXlDC9rJQcsHxm0+6ozUG9fc665zxE
6Fjs64Z7I5mKsWffTKo2VM+3tAapJIOwYeRMEEua7T+fhCANPHotL4cu3jyJ4ykVZHDk4SR3jNuT
ZYxy4FzoUNpjafbyNz/FuySK6VB2+oeBoxYcLpsv3jTeDb3w8hpvrcHl1YDYERSlpjw3HUDzK/e1
dvka+Mvt7dtFYlfGSh/NP+FcUBVmEiVs4F0e9Hm1cKX2hHLVavp1J1as+Gk4nHyS9pt8PxGxJyP2
+NOzBR0ett0flAzIkquKNI/CgSEKk7VovQVHj5hHhwr1I2SCKcHw7YQXzbFNO/AwoRktZnvrz5wM
QaSUvHRAgurav3GxSgZUxhM/s6VWzH+looQaTiIzXfpL/t5ier2FUTT0JMOheH4uWsstD7hUMWxy
bjZMywrqUi9TIO4VTIC8AFYFZcb8scvKT2+DCYMhngJKfmUhVXy2xuO2QcfHedJxq5ibtRfJ0bic
jgeUb5wJPuaKZTpAumeQHLNQttOw2DO7cn68pFHkVcApMAtyoGJGnj6QJ576kvqR8SgdnauprvIY
2RczIZT3NLy59+0Wj6JQWt/noz95F0woyHWyUFrQWx5w8f8Qh7VafJWnOU4rZJnwkAsQDIE3Y1Nv
oTEelsp3Snk+i1Qs7zvNOiKgGzBNzB2r5vIjWgP72K5ACiB0x2Uk5bktbREvCLFceWEwTVvqr2uX
0ljIk6K0ENx7s6J+8s6aoSpIC+YL6eidk/0Q8I7OII8Qt5a5lXcVe0PnaL1YaW2XRmIS4MVyd9Hk
wfaYVAfLECSoEHZ0A1CIBxLIxqkhplvIU5WFrC2W9dQcybbadXp7LoeFWehhzdj40AiSVuuHoK1+
vj+VQ+M37itXRHooqQXUUo0ls/jK31WwREBk5G6f0zMWnMmmo38bUSmkDEe3T/Kz+R5c5HM36loO
c9bD/UbsZrsdqS5yxYdQHfzJhUrZedshrUPl8cCflCvnpCSD1xJZh3jEBw30H49BNJh9bb8sGTbM
YmAsnuKv2KeLQNqfo/uVcvrYh9w7ghDd6mfv9BkrCkgYm5PUQkq9z0E6DSx6nJgTQGg5po+HTjw2
1AoWCdFfWOek07goPTPJ2NvVu66xAS6/n3VpC8okkxdRvG0sCczv0+gBKLSn8bUL6jyKO3JE+JSP
OdfWC5TpHzDYzf6jlfksiDlJWoo6BbohdGCWn0oQCcEhfp/mNbz4nA7QBWfKPvMJlPRew6msdJoF
Xd7j1EKvsX2PIz/7EuW8AF/z2HirgmbsmBv5zWlYdHfj29ojOR5vX+6iZn/1HG9z0EOO92n2EK3t
YsFE1QDA5kC8Bi5xV92f2mHq62IYRMTmYWI5tiFt/P3xoKUceeEWg8T6ZQ7LG5n0ijTscfAcVTWb
rYdicTGwWpaP0Z3I/vZ4+A6WeM3DZEdA4pO5pZR9s4nK74oUxZ6d1Z0Dvsqfdup13mWOHExGOO4m
bTevy9BTNS1umG8oyA957yORUsyAMu6jhWnBqHjK97xGh2uJI2MxZiYsnlMCiQqmE2zHMC5nmaCE
I1iU4GeLi/QYZDtMMt68/gPLvolp88QfCuHzDb2qKBVg0AwOZyKrJncIX2Qhvag15sUd653lSDBU
mkQcNQzu18SwGsoXmOIOQqmvKbTcgQShJ5GQCRRfpukoq/DP7USsr0S2tLL8PcgCL6IFQz5zkiLm
+9lvedKZQ6OC4vqkkjmi/LHQtH5AdAYEpV802Rcp/7Fx9ofZJcX8yrFlGouACnyD9YjrMItEEHk1
uk5LZMjfR9kP9A1rie+SZxTry0rzOgzZF9xIy6csWXJdB6OqMoJpRTcqttIvHnIrJDD1tewTSMSr
/LCHZyznO0qaLbOHsYrv6vcXOlynqFvRuEB557ZUlmYBRjvElLNShmfjEoomIP5jwqdUROpfEs7Y
kzVdvgK8rj1/0R9V4JLDRRQx0hPIeObXq/bsg7fP8M4Aa8iJ0nF+RV337P3oYPgErQPbmJjgvGZN
7lMtyiWCFs6FLawZQ9d80xieEnPIC/dSHyN/sjnkSEYafNoxLNVMFS1TkCBiEkj9VpB+o/YomJoi
L5vXJUNQkP1GkoL6IPeW2E6R9lTHbG7Q6RQk37TQGgSPEPAjzhdzN67cEF/7g3XMXFwYbQ9pQ3Uj
gJeC2EKKFv3+zI6XZIBVRZmyk+L5W0zjADHeHyaBANs+mlkBHOi0l80nX4ah5tXt9NzOc3yl3G2o
+S0hh4cHJL9mWAipD6ZlUmZ63WBxxTsm2FvaCyGkbXde5MXmz6jBJF11Ay6v4yOmudyKca55//yG
ZqfVF+Q90zEUPD2nwiW/Yuq5R0gmrxQqdBJUnbz61o7+B7ksXokgZtJKddPA+6jPhf7BTi7x91su
1b+O3+zslo8QSJpjz438hgfsgl39Ee2PAlF9lqLy4C1NOegDEnyF1Thx2IeK5cQfZls/fm0VlThH
bDZM/9O0DCNSSrS5kck5YqVz8WHSrlBSTtJ0CNvahGm07YdoF6tcdkyCJam5htesiq92tLMqQxto
Cs3HVT6P8sdw83xWFZSp7mldmCZv9zvkbw9m/vDO2myZOv2dpoWN4S4SDjZt6tFLPMhh/ATFUqz1
6K4sztSec2RZM13Qt9LbpjPhKWPofdET6ZbvaPDTnyDe19cammUngwNZf5DyUytnZsKNQJt+ycok
w1aswTd86df+eIN233ToMM1CNXQt32O78u9Gn98GWGrwpAGjvSu9QqaWk2vQq7xIwgdHklxyhJg0
4/HfdG9Syz9Nc27FjOA0VmTW1IL+hm090qgwRWcH16/zTzUkoaWrJSaAeSz4Vy0lXAXBldavpDM9
WoKbt1D2yPBFCXq+nACK3jX1q60Ia+9VBwc0iUTBptuAguRGYb33nFCuyPUQujofCraC6GpwvrCu
q/gF7y2n71HGi/2W25bzwQjoxtZKKq3fkBvs/3pleVvr7v+i5Yf/1BtoT/35zYvYe/JzwYjUfEeG
Oc8LapvLKEbQmkBTfNa4CWzclkWA2mMyOPuI+7FWo5qlhnaMDIX8jAxxrck2jqdjpWFniH3sVwz4
n2ED0aYS72I/k0s/g0UX3vRZ8P4Q3mm9DCA2KjWooIM3TbAdvuHA7H3zc6viSRT3ppJbRnbrCYQ/
tgUQ5y/70JKno6YSNV0sQ6hDlW0pQ7n37dHo2eoaxKh9X/43fHlrGQq2usL7Yg36Rgai3PPZYq5k
dlxUf6ZkpljD/K1iaZ+ZG3rBzsrcdOeJpYEd3RPeDlK9S/xXge+PHNbAO3mSAmLmRJOFPt80c1xT
Rg1FZk1Xeu4WXwVogyULIMBuvGiXl00geKdoInpptt748SppOgjuewvrqAnEenuADAmQP5jLPWUX
/WZQ7PyrCU66zSIk/J2Q8X0YTTF+qbzlh6+RaR5WdLT6dw/RtVtSSGBzt0wU4qZQltvlZuqBkYtR
bNDOJ2G0iFcxTBCBpr3Gip1MAgb49Zc48u3LDbj8KBdi3hlnV/CXoS/OC1yj1+UJcyBqFOCwk+ka
G6nuIJG32XVN2atAwPVeLPw+eRHyqRqan5DxdufCN2R7ca49OEvuMITSwOGe4iTtqaWQv6PAsZbF
+49iax/DyoU0oOqCCSR5t4/QkNPG2NMBSdYPfvc6Z0OTrEwLm3k8QLklhtS2t/NdnEec8UoXd2E8
m762bGbWMDjZEHa0am2qRwe9PNc+K07x8YY7yccH59yOrtRxnwO1JRbjjCxw7ozgU9W1Q7DBU32m
21Pka2sEN83l1w815PoqxyiQ8+wVbljwTROEQoT854A7hbFRD2H79A1EzrUQErk1MiFf8G/K9tFT
nCE2S27hxQfrbjBrlHMyereh7/PDPx7aCAI0C2Fo2CGVKyRNv0MeekVRb0YdHfsFDITN+UqsS2cR
kTgZN/cO5kuOt8iCwQa94az+SOv2mkjtP66xl0lzzz52sO8xiOhwtrWsENlXOQMIxy7clkLD4JcW
R2BnbQC1AzIlpMwHrZzTf+w1vi0jB33p7M91Pm1XNkNgOQ9QW4NPp6gBgL4H85evVYBUQ0uML+FT
7E+4p0tpRfxPxzgPtNDw+QtBgOaurMX+/TQr6SwyZq20dmd7Du+OFiuEDz1IcBC9PFuzn/ES/df2
PPDqLTTLbMEu0Tz9H5DdaeB+KLT8yrr9W9CWcCSrDRq0rqRYyCdzdCxk/hgASqfDvU7GguQdEmQF
WRdb0jh+++G1ubmYvJwmDTXxTBOlhcIW/8uwDP1Yy+XZdmW2VNXbNkPb8pATBqpBLV5wADvsBW6t
Mot7I+xKGj1YRvtrrYxcC93Az5hPcPkLV5cjlMGbBF76npl1mHxKHTPjo096PGSRxqfX45EgNc8e
n0vX7bsTuRwrDtN9a1vAC64Gm3fsoUDN3d7exgzF7ZRSd29wrbQeMvt/eHmvVxBTd7dgo8476N0e
g9RzV4jPjFlq9ouyv69hcuVlmO3O20x9omBui/eyUmE4gPY4wn4M7Ryv8eJGpbe9mXaNmfK4ADpf
qBttCMLuHO5rlPOYJZ7//taA/1Ai8hPXQnCdPx1oGiD/i/FGEHhRq6vJPX/v6GynPy+CJuGnSQot
MxOHzYHQ50l6aPOBi8iv2F3I1v160qqq6VXBxXoTLPwOgCHX3lP/manHIc7Jyd3Hj5rEoMfXN2uJ
wEmBA2nqxaH39tdDNSEcpW+MrJydris+ysDSofjpY3JR8lbi3Gsu7RqZQogDdF8G7ls4cxm8Gdru
cW/fNeC3t9QkFcfEm3HKkUjSOhk+S8r+vxBKRR6NCRvQ/uVBEK4tgmPXQYbJvfgMmVRNbDNld2Cz
CdJSEAfpJVJQCw/clgfmxJ3ke75gAu6cZ33/cl9w7ookdSn3ijS1VXt6cKu7sBImCCh9T4L4mU4s
FpttPUbZZzzoxNG9Zp0g6wiaNXWn6xYayeP/NDYAtj4xLkFAoOO5iOqYEGh6zm3WayXii6ywLeug
dibylMOY7jge2NU3Y3fiviickcSUOAh6EQmbn1K25N2DGpbpdGf5LmAbR8t0idf5HvaXXRrSbPQ5
MLIfCdGfWbI50hHba6l12gHbpHB37vaOKPN8ejAiplmuRyoGRmVr5kdXYpul0wqdWOfQtlEcgbtO
tq/ID4K1Dan64ZvK0p8SzbWsGYYFl7+4KA+8rp7CZYGWfyXjsbMhUI12Gt9YYw0uYWUJEeUBm/9F
ADOI/BNecTAL0Es8tRGSANEMBVyH36KtQEQ8X1KTtzq72ZopDiIRvMh51glZ0zDIezcbMpr7TpEO
zCopEGUq9XpauJ36fqOH2+lcSWeFGIGYBPKAZggV0076rrDPR9V48AbTOIU9KAiCI4GkyAp5HVtQ
G5iD4+nQc3nSkjopRlshgzikhs6XToSjMn98nBPLk3We7B9UU7O4fEDEbvJu9qvfuf9uoXLqLwDE
3w4Z4CbACNLlHeB11+dP7ZOMcdhw5sMf9GJSClm4z9friQNYNqYahUR8Q7pGoESGvFgrA3gfr8h7
LgOi/EFtHvtveULyE/GdTLX5MvOd3nsUUjrY7drI6jjOslTTznsDy/JLRD8IlrlBV0vw3W1ZY5Jm
epKyqYH5hmAZ5I82BXwjsExnWSNpStUbFKs0kQgomK2AWT2GJaU+luOo84H/klFpSaDiEvt520UO
nwsODCNpZmdJcx6KAZmpsabCeYC4dVdQd5MLvyePUlmGEEHoB5Tu3ImyZ6XvXngT53r1jxMG0GT1
t/7HvHJP0gGsnJxSmUIy/zP5DFGr/QJTMlIUn9Zzp6IFbKyyEa3Evt7y/g/9troO0gLYVG2lREhb
JxjRZP1SdJYTRSz90dntu9vbyYzOgtyzf9EPsnr3LY9UPM5CtiPeifufeFVk2vFh1kG4GvVTgVMD
RWHnnIz6FWhM9jFNs6cSOLO/csq5vhSQYtRtGt53pGmgNpbqyvX77ibYx3gY+MGSnYhohA6K+xGj
ivEB+GeXgJBSB7UO+ZEnhbc/6VibJuEQ+hJdAAtGq+uarc3S282k2IsDdvO8qiwQuJ+ew/D/D/NO
OEdoEn8hrSv3fYH7smWxJONALWcvp0+EwcusyKtpiAegmI+QLKnVksyj+oMDnJjMPT9H+eF2DCJ3
SuuvdWjgaqVnWKggeLCdDFyDWL0rNQn4ECrHe7E+QCFeHCWfcWqBTguvMnGjKMvBgwn9+fJcbaoR
RfQn68b1qglYVfMNGqwsx3ws4LLy4i9s5689gbtMMJ/qHyG+xudwYXRCfeK4+GWWWNj5SeqRy87T
ZLT6D/Rs5ga8Afp/EDUJ3v+P5LELkMfxspxBxMb75sTuGbvDA+n3cXtgwZ4+z8yMwkDKvEkwQk+4
L/MekGSVOWn2xtukwOkMjeuy+LvukxOyhetUcgdVxUanfFqS8TfPP+m+p1UfcMM1wXhGnJXAxPlq
z2MNcMYLG8wcPKH+hhnyKNtEW6nQYw+lKQoeeoDi5kDBtOe6M70UyOrmi0TLkVN3Ud+6UkK9tcdW
OLTfn5S28132yUFuwiQW20bGK/YVT19IMQ9jpHl9N3ac8d6AGqKElQloM7ky5xbCD3NrXp/VTdNm
6lfAkkUeaTctt8A2lUGKDDmvwWdfNOO99oWFZTGuTkdSsFZVvxxQdLRRcn2o+mSNZ3U5U72DOHEF
Zr98Q47iE1K+wJ+n9UgFh/XamDpmM1lo/GOdv0EOvT+eFI9wlWxbXhVaqrwH/0p0SObDZ77weDVo
SB4k41zrFqyd8KhxnOHnh2cZCbtimj4d7Y/TUZn+nx5Vnw7smTZjofNhmBJQCBK5p65xcoZjJIHL
4U3/j2g0EjnhEjqNZ7WNKwM/RV6qHqGl1fyBJlUrdRwGLyoWX450kSmUIpb6dZbKb5WtL3mnOEHc
1iVXvExeK1B6Mb8wbeHrfOeMxM7Hk4tcm9vHj0+ABiGFez5QlPguInpDgXjhXZNM1eD9KZb8lqEQ
kuPRhaJlWK/cPh8U3WhF4JmqwE2AYBvRYgKZPeHDu7sBKD7E+fb8uZqx3ruZBU/heAOhvwyw9rAD
f2Lmvn5tMYzoPkJIWpEg13RbsSK4HjE1rlzF6Nu0/0yeJ2dk9M97wTC1lqQ/BTZMJ4W96pAb1RL2
+PTm0HFhI/vhPLbEtLxArb+re3C/bejzKJw5jDHybqriW8kJtFZonXUf84DeWZfey6M/bGAy+huO
jdlavitgenfqrwSC2hZPHzzPMU2ac5pDSQEyQB+L3VX7Sh0w3deH008mRJYMd9VZtDqVB1GK9EdX
JS6jU2m3yzwFj9q+MogzSKZ+mobgBx0waT6zbSbsjL6Xg/+pUCQ5Y1+TZqz9FexxAukur8ViypJU
a+aon0F+jlOi2BdjklV4p9kh5KWw7wlvQiiPuKOFsTYGk75J/FWk/WJgHywLxHzfwXGUo4wBGOZB
yYygRA5DU2Pot21CAczmFqr4g7pJ+InijL/Brl1WHHg/eSWEehoW+J9LP084qwKh3i5dDi9AnEuI
m/QUq/lrQt+FWNl5tI0G4zPna3cKXI9CGB78zhVMVmk+/2cM9eBMJol5FpAxA6Xa/6bqhS24XGeF
aaMkuaqChnE3bSUjI+jW/CAoAbpV1ou6iIqvgtlJxSzRZ9VWto9PweDCWA8u3IRM+clG/L306xwY
vjwptd6Wann1LrrK2oUbusu2k5ZuGc9bF34lKUhtUxuou4ybCB6EePuDAzPbB8gwdw/azaIBLlQJ
3gLp/yb/eca/J7a8S1CyBydSXM+JW23d81q8Jm5c6wIHFWHgJOcqE08X2cZrvLWc1bqLGGKYlqqR
1nZUb12DFxxcMtu/WfJfRDzowOHFu/3tYeEzx7NpDceqfPl8pe6ESpvUjz0Kt6wM3oXHKXzo9j2C
e3KmCrzC+HWUNGJZ7PtEAtw86uCHTrd0UVRLQH3E3AaVVYes0Gqbp2Jh3YgBc5a9OGTCnnA4V5Ig
aecFoPUAxPGbmiVGdZDB7GGcjSy9Ma4Y2SuHaArp1Xv+ozeErY1wCUShys9qYH2blxeDESVHxLfm
XL17gdE2BOaT1KS2ZFedLZbmtbzcwFvrNpXo5FYfwf+pgg+yxze834w8r3QEsVosfESQ2lrU7Uqn
3xyD8ugtPwhgKQVv3Xa6kfna1tDgGrSKbYZoeJsen8Pydll60k3llwmIQXmybWj6Lgrynw3v8Uym
e2UmBI6dqEqJfKksJmEbH/Zb0FoMc34RUPTHZ155ut+cEAkRyupbZMNlm2UYRucFxOWzI5Q+1Pmf
TFU7Bg5Ggb7lQCTRtFfIBvZsMyYp+dK24KBdMogCQivt5vQyJ4YzI6B6rAMdKZ0yeGsjnZSZL6h1
rpwbGAKlzJo9zvF9YLHRjhTIe9VmULiljJl7bjoae/6I1sZv34u0q/82E+SdTNbz9Ov985scgbmp
6Tp2+N5ftvWeZEA6ASqEAhxXeFSg2bQ9AP8dlFDqQFZJuWJPTfia76ik1Mns9grGSB5gPnhxPAjj
kKHBwtvTzatlTiHXc3bWDLxcFVws13kPfuxzvQCXUxpM/5ODfmFXb/RKZ6fiwEB7ninp8FybQRZF
GphR+XXdkuZ2UrKKRpgXpZwP6PT7TSWsZSAYc8u2pl2AAaHsWeKlINLcWG8mq9Gix+qFG7px9Vxs
ZtunYv7Ociom9doU9gcejuARMtj2rbpwIkjE5ZVb3g8cpcUF+ebZNMDt2DB1bDL8lyeVx0y0QtMC
TMOa7U3TRLc/4aZMDFL6M70jNbLph/LzggR8PC/Nfe8mLsKHs7TlSRdR3BabgjEwtlOgEe7Nn3lJ
0InCCSoAdD+5a5XZPqdCDO8tdRrvH4Tk46NaSQKdV5n+HFQ6oFWnW7L6mb+w8WIj/i47LyY16Dom
xiJcwSxIcVAfxgiSZJ8PWu7zudjaPm6eq0cUvfUEwmOw3gH8cKJ6+2nlVs3JdlqHJflpdSUDnos8
jJeEOcx8KGLf05n/qL87GH6LKB25Xi9JZO6sEG1OoUpbdLD7DvuTTt5tzHWEhV+gc5sujhush3We
0z2V15Q+8o05Gg0TMQNJrZzb/flgU65ZUrnWV6uoKVrUYjww2/UanzcfaFZOxM9XrrZNr0dZ6Ghj
wmrt2SPgl6I19IEpm9SoCHIYv3gK5jWp131NF7i1qGpgtKI6PUNzz2wPzwu4oDNXHatMEeNRx+Fu
F4wW2QwHMmzZHKLJq4n7bUp2wOyvplI2P64SDNfpov1FtqQtt3o64t7LzfOWcuJjHTt9DsHkGTCh
ZlwOcwBqvvZetUJz93KMgCCLG/tOaYhMxtcUK74GNMGvDc8D+NuCWOXzQS2oAlfxc/1/NlwpQBfo
GNNMVC/wPID8EcTV/iQhJPoVd4wEeHChfW8JJYKd8Jicfn9QQJxy6yvxydD8gcytH9Tle9XycQwJ
rOHY9I+hNIsUTEWW9sc6J6yV0AOc2ggDH6KLvKFf6iIcOADJm/AgnEKm7lRUOSShhZh1Z+OYlpIH
q3NeReM5d8XSaUxc0mU5T1evPyhTSFCFN7SXD3shrzfvLvxn/Nuczn05HuS/kBtYyZsBeKHB2uLA
1E89tbK/LBf/IQWCl850suN9QIILiaKtcj8qjbJa7vHpU4CuLo9T4JD7Jr3i1wzIkWUo4T+E9+ml
LhS+p/2lxgnQcMN68P9hsjZde0NiPMTakIyE4Gg4YltoRM/pjlNL0Cu7DQptK6WPcg/lCl+hhiYI
hEoFszMb6sVhjY9jjajpoiamTopdKCSkmGRevmZHajl52c9q5mIo7BMxwRsSz0MxKf8KY4R7iSt3
sucUK6ztEgUdryJn/uKJmVDmgGguV9zQ91SOJe/7x6WqzHBpoZp1t2twFIuS82PGEcoo4RLx2ddW
yEqPbni202OvQT3LTFk/TToZxkDScQNQ2LufC3vzraYYri4Ci0jCf94ITOnc4W1pF4xRi8BXURC+
AZwKg1EBDT4NWQaZm3681FhZ0e2VALIG/F2qm35iR+itiKaDsvcnnNTLWNS/7DmeAjPwcci8A+ck
bga4xPCnYs9cm60IL1p4CBlApxagDr1SdejbF/ObUHOok+QIltKO8GOknZDupozgQBiHkT9uBWhp
1qD7iI0dMGWWJK0rkO63y7TuCr3w68i8EHhvf3ac+5Plpr5vuj5QVgwNtFnaC/2SKy81iPZQ0x2n
vWIR1Pgr+gdvjkvd88yQkBvZQ6/uJCQtKfE+fDXjbZODWB0+Jt7GKCHTFPRxtaoE9mFffnfKXPCG
K0Nx0370cusPjYFPPVdElRLwBAVx2ZXYMdfU/tWhYn2JRa6SOD/hDghLb//GKelccpiB0/t/7/T9
aJ/DQav6t6flyrLM88pZYCMNoPdzix8itZUpoCDpkWDGM/x5vQBiIjO9+Dtse7FlMxsyBjrnv7v5
hqJzzq/KRxwt/jwFmZYrwi+WoKkIRF61TAEHfdtPIGiGWgvDPvCvJU2TpExhbec+foHvw6CvIhQH
YOdrXRCnAxDeQyfE+qvPyBknMHdeZ4zV+BHg8p8dDwDvvQ67Rr7JYsxTMjNpJw6fXkVIOrTww9SE
WtT4CZTAnacYm/FMluSpZZa1eVQtmHsF8AJ8/XmK5hOe/wFcbEETSr7MdyzZRR/DCoDDbaEnuXvR
j+FbBDVXn9XZduiJwFmy9/lZvOyqCXqguTza5gCEpDJWJPtRSQuOg4QbwLrqNhURZTKXLFjWmy5X
hkWDbFId1KQXK5nW0pkizKH94aarBBog+yQpVWynblfxxwdcOylvQTqTFg55nx7cZs9UaU4EgxM6
F9oXOrFSrLXIhTX1rGzuwtyQ9WCnoA9uWC4UBTFvz1hOv7SBu9lhk9bqzgNEmNot1dplRqH2tHPW
PJZI7BSM+9PPiDgIutQ++1Fxfru1LUZxR83tvFSlmu/Cy/4pSgsK8KKVuvAikJzCfdC90WpgR5+J
hMHF7DLGylH8ma9Kdw8oBEYehXHQ1b/XBboYfRX719Aes3A/JaEBscJqOzrdsfeFD/L0DSenvIMS
F3fZ1vEUtgEmKxJtc0zJF6rj8WsYh9rSk+titQVEnsHaORPtJKSLZC337CXZnpFQbQTA0fzb8b9f
LbA9UMGeGdr2brdlp1SMeu9KbjCaRWscDBDUlIx+OqxS1/Qu0E2aboxMy4QGEsyPGfLsMEgfmhX6
1gSX0UB4FoO1/X0C9WlsyKadj6fzWiG+AG12k5yvtSz8ZkwpHMuk7kcqg81ItSbbypvufavr5m4o
4dG8Pek3CkGLwhDAK7iTqAq82TtUPBUhGyzODlMQnGj+/BZQ2l7AUNsmaLzIZCvXg3GRyglh502Y
ktWZydC5DhgTSpdiYe7xKnwNqKCqsUongZPxKL53Nm4S8OPImEvVKFyoOTdaTUeXkXN4/Y6PtgdQ
blYQJ5hTVQPblolVJLllU9hU9Nu9LznRFDV/pLA/XOLFb1gOknNd2YpE6XZIMhMcaNGFSsWldkDp
mZ3neZqcE6WDNFSzJdHXdXypPsgfDZgpuSLzqoJbPfvzWrBDtLKe9idEl7hPAZgaswauJ2f3s5Zj
b9B1Vvwjdph/Ggq+usogWq9svOmX0XvHVtm3nv0YBdMp3pLp++CVXaFylYFe6n9RacHEYqQ78zVJ
TivpOTc24Iv5/FeudnAenQExT5JnjLLdLRdUIMDrrdZmyRhQ/nDbohr4Roi2kkbXtr4Q9al91swC
8XamUxt55XIIHpdjOvIxjWXkeBw4BLu20Xvg4Yhvow1N+goIuq+NvDjuoXHPKepdN4uu7D9WfpLr
RJqDtedB//yIxvKckHdYl+Lv9YBTl/dTgTqle0amkZTBeZ9oyYv3cbcU81MVplAUV3M9KCHQFVFV
Ux76e8zrHabf58bFEi7Mm7MgX7wC4V+AY088OBhgsjKfCILch6NzydwBTtiUnYvRVgq+x6HisEVd
6LRP/n/6/lxAycHfQ+Be0g7u2xn9IPVKXnqwQVKHI3Pr3s9fSWzrnaQuoTys+KkjIL3hK8E0jel3
SXHAZO6f+nX5O7Fw0iYa1ppE0IvDm0GrCrO/hK3O2nK/RmJuhSIM0zQN3xH5fZckYrsl0BuJITO9
bqsdV2W7jW9kZcx/slqtlIh3fa0tyO6AZLxtTrf2PkOAhlAIdJuz4T0mXdpAYt0zKmgM0Xag1UpD
FSWOYK8EZ1nb+WWgOSFXE6HP+zb8K0w5P+qsq/sQH6Y3U77gFlPEN1wg8Wqh4uCCohmD7ibKFt00
vhOnklafTGy5rPauymT7hi+cWyv7bvRWqkjGXG6wgDDttpsnZbyiuKza+Gz9VfaFeY+eyt3tcNCE
4h2dUR7d0XPvWb+shAG9tzcMX/YWAQRXWorfd7BYriGKYp558Yf2ZIkpt9JwDbHDZ49zLnahISzb
TcLVOKaG/G/oFCOwDwOqAN5yYzvl2BAzQ5zZXzfU2j2TgPwkuHfEquZeATITOz36tBVtFMYdIDdO
DUoUC0s3Dc+qpmGhSOvlU+aq4fd6PY/qhIc6y/Vjnif1CTPOiKlgGMwQL7E3VRZPfiU658XQ5gpT
Fu3Ffrw1gsqnUrxVe0ohfIg0FE6to53TL9JyA4eMZbx6XduaqIdejd4ZQH8WrnN+6nSc6vBQ/mba
L4EmOHePmuPQW/UlA9TMldMxI1WRtCaMEpqhct6FIasnyxl/OaEXclumVlco7kQbUV0dn6J4b6RP
96dZd4wMGuLqVHhkpJl6j8uKsqA7fKLuGtjcicy8IKuC+Ip3JvbPXXwC15oLMdr5qSJJNmhTnYKK
b+rznhpBKMCJcL+TPHzfCuEwk/Ts1oVtHK5O8si7LwKXTYFTZtNL4YuWDmPnbwqg2l1QprbSrrjg
HwUYqqhf2yYzBLwj4UlMWrJRzhNlfgL3u6VFr/z0h3RvZTyHiSCqXl/b4L1DzEXxAGeNCrCsj4Jj
X24EmnGVVkccaoYWVQafLAWkqibf0nKPhf+D0267JnbfeHUcXpUVD/pjnQWNLZkurKbbXaSY86Nq
mOx3pXVvDDO5O67V0C2DwumI4TevZUkiqCey1G+TIdUZELiMPwVmHhxzGaF6vZNN49EceT0uRuZ9
l3Ja7+TzqBK4hkUDE3FdM6vsKKttLqDm7FC70ikouHS5+PgUsiqpU1qe2xOOg9vUeALUd65Bh/oW
otzNSI4t9De0jTnkL8PkzxzjalUJksUzndq7mssWpM0NZo6zFGHdgLKLXS83sA17Hh9X53Vyj52n
NUKtVoDnOkVwGJsTvUoCXo2tP4ymb5fJLNpQAcPlfav7QFEtm8euMuRfggne3New3uayhjSY9QWY
aPTYQVUhZBQheuWa3O7H3j+1EZmTM2mZB4Q+xQS/JF3SQQMK7uihqxpVT9e2YgdJIhvzJzboTXPl
7C68iPdaC58WNbT6CInNIOxIZm3NGis904ZfZuBd51BLGmchEOD2hi/wsw7jX4ivSxWUQ98WFls2
nzMsKeHDX3ti4RsMPoQEVtNCoaqZqHr2FwiqvbrK2OMNM+46Ou3W4dStD5CFWBzxIxyjWebdhrgt
MaAsQ1BdchkCcL2q/JdFHaTWnegNnCMBs6hFrpWvwOIb0dnDzdkOdh0qQJweSwLRInb/1QJFB85n
8EmyHTqPw8elfmj2qW1pLrQ3pTQO3tuq3G6OkEu/n9yWDCGkndwKl5dgROB6uGcHC00lM4uTc2c/
26rHMl0KrDDCSDvJS0l8qGt7T0aR1mUtHjy+JLGK9D5sCLB8e+yUoJr8nckDbItQcmtYy4rBYfnG
pPSqdHZWktsKGCSAfHHhV2V1tEAHWK1QA1JLWEHSA2QZvGFOxVWn95aJtiLc2mk1sVA64XCKoJQq
+zAXglZN7X8UEGvUvWpy3kErTZ44gSVSxYcyFQn+kzVXp8MfvwFDHNgOtL1xXjk36mnEDcJcKw7v
zAqBmUK6vFGpNohztl4NFCkOmqfZCFaxyfBQOOfQo7kKgspYqrZqSohCvWPUKqxq7r/UfvMzrR6F
YApxCsmDOjJFeb5s7XFg0XQyeWMxOHcBsvIGajUvOvT8uBN7p+ZFDC+806uI+fHiClMhMruT8kwI
MzkBO1CuSBwm+Bv3c1qGWTb/LU4XBG07LhvIxcyvlSThCWOor2/10ZJe0yd9YZzBhBMPyOSQ5Eel
doTJ65lzsIh0Yyt7BeznTfXCgtYFjvnBf0isnLxDHKeeseo3Rp1muQO4CiKK+VK25HMYpUlAACp7
f657Psp91PpqvgS2vxLiLNBjZtchJh2irh/6Z2CrR8De1ojo3mEjBSkOxPOyhzRH9vNKfxsoLdOL
jU5Bzrd/ItZer72LQhNpyDH0hGA8qpP/cKBVGL3sQ63M6cQ0lUswuuaoOwLkZ7UZKe6yjxzDGz73
Hdmh1VcVTmawE5eqddJPzzrwUT1ds9mado7KaOsZabCFVZeiHx85sfj1APWoCEgV5HEMZRmx+sWb
mmWmgadzCNYu+hKNlsh/PbH7W/CDTYxH1mfwBU680KYH6lLq/XvPgEDnmSk1bY8ZurKfMGmSFnJu
tVerc2y+TXKXcqP6mVuRhQJmN/GuBPsMYX/KrQRESpsCxyt+3rrUPX9VsFApnTGy9Pv8fozQDMTC
jdrvP5+yAkW6rPcr4Ps+aelro7gFrSK63b3UU32JFXkBlfd23DnC3B2o1y57rTzd6gsj0MgcfE3g
Z07BiPv4RLlNdVmaggDAwb2VYL7kVZFadX2WF26ONT48G16u5onrI7/8KgNSEpXDHOebIcgCKOPS
wbu+pXkcCC2cN36zH3q/ZoydrfrMcrreyO/3CmoSK1sriwLvOJB5kNP9/vM5aP2miySJ3rgK6L9o
lvNZ0EoPvmq/4RuXH6ZE74kaTyEJjkjyiNwzP8EmFH0Xx3wDSHade4EKA1KS1mF7KwZ5hm2tmpwk
DPcepZ+6Ow0aozbDGqxuJSLRvcGm2ck1DLfO+t7sxhfXf6UEoVOZTwxTNPkxAPU6Zu6Aod+nBCmQ
EHTwTa/YjgOTsxqOilsErOzdXCnQ0XjG3kdjw8+X0KsVg8vPb2y4QF/5WbEcnj3H3f1lxSflILeU
dbtTfU9Rs1vrt1TeIpaBRNc/NjRNrp+cnXafoM4bv55du/FQNKpKf1SmthLXVCE4Tq2QjHk16zhr
5HzWgmCSUVkpUcrCt7i6kX1yjnus29pU/Dd1oh+ZrjuawXvcJTJUerpDHrFJKtyszyO3Ny5wb799
P1Wr+OHFqGiSHvzCwW4zI7hzC5+ItkkIJfmfnpA6XU/QVX3ujqslhYXtirOiN9+UHwaGydV0Epzi
B7MO8wbOC7fP6aXAuovJHIoobKS/lDoUeZxbTs8J2q3FOTq+YObvYX42Z7MeWbV+VXB+cqsE2/b3
L3d/HxcU+ZkxeU2KV7rjmiBLqVTsPjKYXYrdrHpsgcTQfmLfDMtBRK8utFPFRWxDmu+wv8RsFYEE
D6yhXE0yrLtDatfpe118xZr9qoB3KxAPS2XW13gxme28WOFne2YWlF1zbx51yukkAB54Cj9TDI8p
cRe1NybgTO+l79GOysdl5VjxWfx3X60BTTv/A5y0plC58n2Yi4o7l4vn+/xw0Wg0WMI3DjTycJA1
1wPP1A7yxeJm1ka8VziuBYB/MT9mOn3tZEij8g5ys+YB3bqA/ruF4MUgt4oZt5xZm+Bs/Iil/idB
N3EK9ZASkGUNS4XN18M8nM3sfE1xrdceLPFFtyBrVFRM0xLOuPAP8G3ZzBg5Tg0JSqr5KBktieIA
bMelO4Jtu4yYj9+6E+usPr+i3JwcQ1tRTfOEikRTWu1/1wkRdiqGwbeJJEqXY+qm/5f8J9/JMtzO
x+ZqwoYc5iAC0S5efyuJ/VYQbgocCMiWVpqg2Y/ISWpYBiF6RW1W4D7I33DXDT06YbgpBN+OWRFh
8M6/6yOox54sc+m8DtVFboFN+qmzBw4g6OWV2dLRNYUqerAxwmQHA9cCl9tANb+O6xo+RrSyVcUb
33+lpv51ikEdmTJu4skN06l9h1ynLnIi90gOrUFDC9vHh64wStydDdlqfQzREQfc3QYefRfKe8Ri
06ChBFf+pN2tsGDcbNacp5bRPk0jR8/TlOAySJivB96l1yDTPl1vxEsBRv905/i2Ew9crS3diPVQ
IzvAgEeEfqjQPTqRlUVrWpGTAQh/MJs2/ZJGWk5Yzt/uImMyvRkhnikM0GxVSwDjJr9i21AdEDm9
1dG6a/DRe/LgEvtJs6yIVdKfV6rjtsApN9qx9OmdaOEhUYtdR0zie4NKl2Z1uZC/8Mqhi6dOLbgH
i1YgwxRAAMExCNnFXfFOxodsEJx52Q5sTInsj2FmBNkU6S9pWN+VgtQfno4Bdjcw+QKXC/PVeO6Y
uxjYwRycSN0VLsYWmVDX5if/7XgYj6sHrv6b0L+y7th9iC1WxWWWaaS7bm0FvedotawIHONykbyQ
CZJClCuhKyzfOf5ZqpU5qTvALW9TjNnvABD26xA/mFli+0dV4X6EenkE2S//oLMymU37YE1QGbcw
s4pa2J07OKmwiK7YFmN3qnB8Bpw0+nZ07BqfFxmbPzTgGVe1FU0zvDKkkk2IWMR91Xg61J0tC+ph
TNU3F4TcwOSbZTIv4zmGZYHzrvIeDItDxD8Y8wCLKc0vhveeebK7BjS4Ofwq7ug2IltN9SV+YUAm
p6SfiMCfZtbw6IsNhxxxlNty1Mqmj1Yft+eS+YeOF7NuI/5KBPsh3naa9AVEG13jf8KLmFpojRsW
mA/6wnW4wjHK2cmxxdHjMlPKNZhzw6yuBDWY7Sw6ZCTjnH8Ee5zxeIqvX9tSIv4mLZS/wgU1GsYr
TLtPVU6NE90qyIgUAVBEtXGAcZOWl+/w5MUCyph9J/3SmHcMlzqhZRYTvSOM5+cUPZdejS+ycXQA
cKd0JZHd2UXzM+7E/fJ8WBHYi1EzU3J9bMYfYllzIH510CH5EnLSKauikVsNcFG+iLTAK9q81jfr
yWiZFesJo2N3MKk2bC6M2zCPm9uDYq4Ph4SnJkwJbXbG27GT2LYaPdS/lYwxjTFhaTkLa7jxOfko
7Fzbiren9qweJi9syUq8klxuBZCARr4VNrmIorrDqPcfY8drLtJjf5goKGEz6ZxjOBwLxqig7c2p
zHHb4+1gueY46EAPxg7TwXiI3mwNr2QZ2De3fDO72FSWZzE3Ts7dO2J/yZz5RTjoSp1wHy9ZM/Xm
bdjzMcUseE3lZ7l5DrIeABcw6oaM3I3NCdmGc1ohY1er21J5MbWp3l4xEj3ss4n9N1HplZSqtpIe
wk7lTiHTbLFkV8m3Ut+f8FQqTTOoVxe9DpLusvegiY7qIgRg8YMQhJH0E68m3GAluEyoJ/OC+dtV
z6DfCPBKKZ8ahghE1lW/pCEIDmzHSkEqvdGX1OGMfXrIGXGEJq2exfq0/xfjMiVUPUvgRzW6ahcT
30Ri8YcUoHjOiqCVUs2/orfyVDiY0RMvnOQ/OTQwNc4B4almhDMeftr9xr/pXsgwNu3QBrr6fM7l
GwY14A5dyiIdWqYlr+zRpLWXcv/nqjRzXMo3ep8tU9R+k4F8EtrZk6pPhebuolBZxKgRGxF/1/OM
3GOJ9yEAr/QbX4b7FfNVzGOFzKEoNEPil+K/lds1eJKiqgj4OS3hYKkNeKw9a03z3YedxLbtHzAS
BjV0/UtusZe88QeJ6/ivGBArJN/vE7A0JbRB3F6odvZgcL2Z87vjTFyLIJcbQ7WqoSsndrYrGpUz
n80KIqahtdYsYKcLqjBvci7lVMpsKYqQzIhnxqt5BYtHh/j6iXkKL1QUDJS8Ci5tRTCLKCbZUF9w
X5KuGexmf3wcg6KaDOrvbjR1YobFqufBbRRKjdxUVyWk2Xua2WZEZ5FB/f/t/ZtTKOQ+mb0yAXBL
0d2lygX3Z+Dc9oqrgAYsB625DE6QLN/SKata5V9bqhHvpb7fuhxTwEujkdY40xq+QOMpDtzosCMl
qadE3nNwO+Cg8j7iCKqA+NqH/TTkP4fGmT1LECd3im28yTQLl0AhyCNiIP1Z7qao4UOxBeCl+ttD
+VM/nIvEHUVWyEXJo2lPjcKd/t3AsYQibu/L75horxM2ChNO1NZMn4z/2TU1rrktW6wOOa6TsHMB
mBcNcNkEoU2YLhs7SbVcJB8rEMFU3d9hn1D1RnG/GpbfuX59yDD63lI0DP+b+L/gbssQZPG3D2B4
Y1KmkNJ7F4N6wIxg6Sqw+XwGfw1jKafG2bBeZLNOsvkbub6y0R/FNbBrHoDgp2Nmdn/1QMCT//VK
UkAigSqNBgKgbG9Zy+MwEGE9ZYn6BK6COKBZUdZJUYmr4vGM9q7Yruojbj1fFotiO515/pr5MkBA
EJEly1PwI3/ziiPUv3w+m5Hko3dyrWVCLKyWIR8q/sgvD/BnpKEovmXWi7+EUU8d83nzsGyOnj0L
A+/kspWFw8OftlxSPFoXYJl+otSLq7Mo1ygXUoehQxeqW7KN4qJEU6tUNvDOZlFn0mRzD9KHazz+
wKKvoEitTznepO5+MgqAKm2XKZQ0UpdXHmKjO7IADpn0RzMcCdArdtgmwRL0ggLvWLl43KzQBfHl
DpOG+Co6lAMDUgFXgIFl2lwIaMQyk2SrihFZNroKxqjDs5GveFmuZPFVMwPRxaJ7xbB4YrQTMCOK
bBAAecMSek+l22aAH8T4q+rA6jAp5jfWZRf+I+LkxevzIqvI18rBfVpcsjfpXcmMnVCsxKcdybtm
Srf3NZp6E76vb7CHjc+ZKnlvkhQVEJGvgLNEvINkW/gPzaJnQDNPWczgvOwkX+W+b4YuNeeftONk
v9gJnTWVJWprRYedIKxTAN4l2RfGcAKOEJTMRVz9XMRWJxibSHBTyOXbfDpod0zy/+qvHqBdHHti
v9C49c81DxgVEVhbVebSReEutY/AZTD6TAa6JmRNsrm4oiE+6G0jyNHrNkwvFazrjtuwTclc1vaw
JN8sib3a1oDknKrUWYxVcOnXDMeKfvePtuEoSMyEpohMXJOpOcbe2K1aDVz6nPamqVmLJ6LUGyGh
6MO8pIbOux+VRMIYVbCtEKF37IQaKTc2YD0y4JIQsVYFifoGVxQXUUOi0lw1yVdndZ3nA/YJjoS9
dtL5B71a8wthBZquAE3vGznyUSHvizsCRwez/7Y0wPCflMSVgyuv2PDrGkdSoRaxl28kUXoo105+
IsRSbuH5kq0cO8KWYSwVOcw0Y5sSEBGspPX8mNQfFR8VV1OKbxDooCnb2LelS09UbsTy0nwTpuh/
Gxowv5Zq+n87zRqmeWqLU3pNoK9EdwiLsbn5w+SRb2Y61korfwUr0l9nCld1f+ab82W2zFj9OmNi
oggvkErmHGlu2KjEHOg9XydIcopFNbPJ5dNxXMELWV0/VSX1wjFPdeZxzJFa66Pogw3um8usrKqf
7G6zNP3GjsT44WdLg46etLGxL6MEFPaNM4zSGIpij4XNpFccpGgZJTbDleaopWINwd90pqCf+L/G
D+FMEZH7SuYi+wxflJZZGb05VNRkC4Cki4ydEAwc0Kd8/G1g39/FQNM/2RVFMyXeJFJCoTaIMrz0
C+q4VY8Iz/eyvJKJFDzZjfSXKFmJATFqXp/CT4KgsHTbBH9D8I+NEftAR+osfRYrP4n3+QrkUQei
OiGl7bqTo25HXxK5HfJHArs1V2Ox/iaADB63X6CTViIUm06Qz4L/PsLyZ1fVm8CeYwQkfnsTwlBl
RpHtgwltol8TWwJABXvTVovECgT2RJbwuRtD79JDD4HM+P8wyKq6RGPX0ghgVXQ1czP0JPOQ3DuO
hdnc8+GqWYsKPKZi5iO1OzmEXHJCb1RYzFFTBClxUBv1g+KGGN5xDkN8oC/wV5sOSqaDSnTK7GeC
k5LCMC4uyBk7ZbHqOx01fWYzEX/ktAlFJCNeJ6WUeUFy0Hj1KJNRli6JoeOquTY4dBeZYfINld0L
QfoLrxbp0nu5dOTPFxbaWE6J6Uq2CgNp045zr8164hrQBqEUmIurB24AuVnQzSxJerzhM1LCsU6G
De060aXRLtrmM/cYJJluib8jejRRrRu91OXkKXrBxeWLokBWkf+1EmWgtXH9tw/9ue6MahaCoBYS
pFhk+kuiGFfjHSRFhCpMww7MBpuIb7cYzdr4PzRG7BVruOxQ/qLnAsEEEIQgb5HenpU0cPyFGHp9
lX4n12GdA5QkK7WpDYJt1isVIYZZuEF2ElXnOXfWQ7WZ/pmyWiGPqHZIJ60f3d/v3DbkTe7FoFpc
rG4NN8j+c+lM0an8RSGOVJC+l8X9pNU3YjtSANQaw6CqXT/2tAi7d8o/vSPKUcQcEbL5X5G/upiW
d5UljVvWKXm9eWviioj9pH6tvp5CXdJTY+mXfaVZC16RZiIeute0RiTotjpYHbgsACU97APlqLeB
+5lc7v2vYcCk3cjoqPC8S/Bu5b7VccASU4c30GnpAvLVUF/jC+YgNeJzkp6cebi2PPHXmZA4vL1O
gSvRF7w19WnBcoVt+w9RnpAXOjaKvjPpgH2Bvy0oYdYRswTQ6AYmEHRqvYu3RIJZKH2+/3P9UNE1
vh0U9sEFzCgCWO9tHm+jn0PA9GxpKKgFXGuFAMDBw+js13CnIUbFiK24Qj8VYgL/4FLGbM6M9R+O
ATWOc5Iu49uSHxDzc/uN4R1tBLiOqW8uprGXl5HKpr2U/gc9PwHrZaMQYJMr0SmJxaElEjE8Gjdr
OQAKGMAa5xz7a2dWDCibWrs/WV7d+vcJKG1GqfiSJ8zfDELP6xOGUtOFhdSDfboy7guESM8jozA2
BKzuTVUT9V9dayMaYgdGQ0BVze0llNsilQnvcAyl2BWUQ2iznOSx58n2AjtIYVSKgM0CYemrGB0g
9j4NgJjqbw/VXNLopo/7AhZczjGTYtTs6BhUqT9bbC9+9FqRfO8a/bFv9GVaoWPmordxQAHCNxzf
1QJTGJQGxCeABy3dg8pZOtnkgqN9LPCkvhcT2JptVQ/T/b9k7f2eF5WxAyusBXvyFBqbU7++AGnA
3OsTgUEgQWRYpCcbNIS5KFckGG/6iadyibx/4oUU2xdHP0F0pIruZqBG9DuhMmyaseqcXPyqjwEu
YeqBjLB4NA9dH7OZBWxw1J1wrmimP3ND/d6Edw+aWjf4ZBiWXAx7axBArtgzYpr/RxelR+lItSJQ
4AwlKP6BW+savoxbtc5PuSIJniW+DjvyME/4sA1CzRXryHtw6bZF/yW9vq6XmNqrjMtL6jQo/35e
kngYk8sGNVv4efyglwqDfecsT9t0uU08vLobgfU9n6tRTOttHnbwJCOtYEhZmmv0pBMnG3QxSjAF
9a8kJH8pr/wXI5pbvU8cEQ6zQw165SEEylc5OiMH7n3qln3VdLu73Pe5AkXfyQqSWS2qpjP/++nU
5McsB+oYCO5uBcwXRHsoG9RV3dVQ9+AHk3EmhrK8ROuWILt2LpCK7jSdWSDi6V9LTlAL0H5Zbfzg
5IMmZ+7ketxUACzHIlpXfnUqvR71yaAjUn2vG25LuIC6h18rjC3tk+isBnf/iLYSc1IUQ7t9Skv7
3gdR3ObKrzhcqZnqtV7Nn9Y8Wig+Ms8JSa1abiATTKP1fNr//R7gYjXo6L6kppjSvWJcEH69YA+N
uGVmchCk0dSVncdEoZ1SW57klhPiDgCPcPC0NFYqsVGJ8t43z9frgeGJafaD+z48O+d15ESQnLU8
k5HHP7R8VP0IAPtGUYMgqTcKKL+qN2p6dBgM25cWyNw3YuYETdF6kWihoTJ4gaob05Hg4Wa9IEJu
x0fIC2tJZHixRvNTFZK27y8JRUa70r8zMquDpO+a0jmTqBclIhoH+jSDVjLsS4v+U++T9EZQMLGk
lVXNSKH14bsN1C28IXW9rwn/sYrEikOsurrOwTLK+GeXN0JiYfB+b3NZKtQrlHa8SqIa0G4x2xiS
WBPibGSKrmJFecmZywMuR8HS7Yyj7TKk2+6hWmv6YkAXqLUkOtoBEnoQ8xJo9cxPMWnoLM7LBSgE
xj2s1Bfjy8Dhsd1sRqnzW9Kfw+rO8ovL2baE1cbCiCtAcaymBRU2qggQSeFS5wC7mbfsU88csySP
dXwzPqMnxfCRt2GXAqJf7Naw5x08NTuMt6vKAaCxorANlu+gHg0cjLWKeg3aR0pIiYj4fBuh5BdW
19Z/4OqgFseK8xdhaEapPiyi5lKpv3N9P/DTTdSvewq43ETJ/W3hX1+g35o/fQ+u7aVuSJlyLRTD
K9Us5mp80XQOd47AU+h+kuegZe3qjRpag8eCLVZnKTJAOZnlvo7PhvoghrxtESY5yKbXujsYP2xY
lt+/qfIq171C1lbVAe/xq1/j6P8UrYtMnw2XDdFlQ0ayMW3UqdmtodPYMnnRv/jp1ZUPArx8fqKj
DuTI5PqhxxHk6Rei2MUGajNd/AAdi1MxvB95y+5YrN+vmtHEiQgcLFgVkXMMxQNy7efhrqmFIvzu
CCAThkedY2Pod5tsCZS1egO6LeoDQf4zjmSwokN27UxFpbxKswLBOnEbnU1Ai4fv9otKoasUoLG9
GrAhbVOdXBUEOoXs3m4SWG/8OwifHqCly+P8K4YPPrrVENkQT46PBMlAhr64fy6odFt0MwdX6l0G
zzmjmm7qNde14PHyc5TpOb3tzkAF06mM7yEfQbynwDWOrlg1wJdt35mSleQQCB9XVmxxTVFiAuSc
pFHRAwBn/Uhg8iQpHjHdv3sP4D94gt5PfBSffLBxQlu5ome/CQPlnadeGoCtL/kdA77Qx01gbUIs
Z9ovFe80EtoFhWn9vv1YmqtO2G40zfmmo3g9w9+NGb6d6vubuaYYUmRHpKzhY/RAwhJ+knJAouFf
Ox31VMAARFLsmmLFOXVqMLUQUU7P8SwsJh36MyYO6/blFKgp2c3lrfBcAJo1/1tTf5DtalEUACUq
UqBXX+hGnzFjyyskwTShHNDEGYh43iQknQcFK9YaXYcRol0RYjAKbQXwsbhTBFbIFeAnF6MpZXu1
Z4mTYP//8q2vlOMtMSs1dDgXJ94Qi5M76Wn3PuRiadaxqfckkGEheREqwzQkyKhPCjUh+2CJ97y0
vMOF+DkuPcgfF1ZSZpMbeP8AxzEThhlr3lxO90vqhaUY7VfJODxDs3xHPolY8fJ3vpH5RE0ssLv8
TilA2qk7ameUQGMZqhxni/LHIpPKjhMD5b8XKnl5WPz4Kelx9+Ar14spEGRBv4Sc5iV2U6JwhSaw
x33Z21nVpMIPpcNDm4CKJ6iQPZTpTPoyxfBDCuv7hqLKF6r9m26lkS0oa7V7HXlUTlem7Vi5CRd5
x/vucc381APBMxJUtaHwc7oioMg0jlIDn1EAni6lYidlVR3q7oUj0D+FNF4a7Cr6mVMZBFFKl+oa
3l3NN/SRTly0GciWovISxZDycCLGodVovvt9JL98HfFppDi+yvkGQuHtBuWJXMOJ133TCM8zv4Gt
+w/eDEq9YEaMMQLT3pDitDgcPoMFQqmsfonlbXfTDPReP4vl57z7O67zE4gsnDGt9iyZ5nKQ0uCq
RTFLt+/M2fYQVtaKBFaczY7iLhoGIYFQEgTZXmRw+5nug1mYPaHcm44CrlgsqW8gkOErG1UK/Xzz
Cn1O45m1EJT0I3r8qdlOfFavqAOczitty74B4F4G6qlTB7SlqFTJlridGettbn7cZUweVzqFJP5m
g/Elc2tHFc1PrFPMcXTKIbu6clMfjjQPmXFzYnuigKDjBS/5CwMIf/K4xR/CCD1rGaDNxq3DT8M4
TAVtU9xOc0wS15RVk52tP1rGf1f8UualV74/q3YmulBzXK/3YtKY2KyzgwJxUJDLmo3emPhRtJKZ
ND7MO7OW9yC0RwZDwnU5pTt5a1OA5N+8yETg1qc1ilJpxQqM6FCIgoiu+j8sc1l59QpvKlwSI26T
aQY0fflgqQT+Zo9DB8oSGg6DGzkevH7+1u7OP8VcCTXtAunWUFbnDpCOEcY8xRqWDpTKH1Jc2Nzp
cbXsJyIrqn2O4gTIG5GpPbvzlJJI9uRMZYGwvYFR+2ZBId///XYQqKVGLpAc10GKoggXcMWZTJmt
XG4ggZqF2gfyxDldKgIxWggRL4BX7IEY6Bu7PP7CE2xvmPSwX9U85VUAzJhDxL/KA4J1a7w7RHFh
kBs6yO9TMSqvABZYqKE+xshClWALBo0OZctCNiPO9dGuZiLpGcwvq+S/H+fMov64Hikwlt9EGPOI
7lEbU6pt4DQphwA6EvnbS0rfCKlFLD/aO2DIUEoma1ui/s7yGGICNCLb/dKtxRGFi8Q1kPrWs4NJ
//wPCMeRqiaJaGfPR0YWVQxhNy3Hf6bLWSJ4cj36WrOb2HTXmG+vTfa7ei8KXmDdIx4m/f6c87KH
vagNB138wNMAs2mlRI4UEmhx8nkksZFeIjt2IcUzxs/4OpUYEMJMjj2/wNMGuLmKm+/NaHKRr0e+
AQq8iGS5fB0otDd3Y0e7Cdl526VxV6ovicPqsjGwhXSBxkP6Aj83+nHrF6l489LxqKFjXKe3pHKK
w/5Y3o5ayoUaUwXYqGVsKsbTVqzZG0LpbWnqiJcrOBF7PNysd5dHR+YfI+UywrlMjLJ4dRSZIVyQ
EwVt5i9d6FUvZBS52BBjV20mGI45uLDpAwdoDh+b7UfFXNoO6Tn7qjx8y9HliM+LDUILtrA8f3hQ
+AbA1oxKfE4JBjApTTzwakwuDFTDze+DNQJ/N4sUUe/rQBgAosYCA1gdPj0Bp/bDgfivVL8TzIoH
PFoeFP4u0IzF3AhhPPgn8HNpa0s59Pb/G0qwoHJc4gE86T0hysLoYiz5L1HqK/7QfXxlAzQHmWdx
b610+3DOcNRlLA3M/m1qmjuFXlDNKqEcLDMcv9t+DjwV3/aFxjsY7NJsD/Nqiz0he698ojFmUwAf
K2T2PxKtTp/3dGdEY4/IK7pzWerAAh5OOWs6w+bZl/rAHXinuYoYADubosKkAgca+dL9hFpqz68Q
QD2y7G1VL6WWUoFCEeq69ZT9t3ROIoAsUBgCAokt5MfZCXtOAaF7b0sYHomz4GGPOEnd/NMEfu0S
IE2hQRbFj6o0euFXSKZP6A836N5OUrjh1NDhwnrJyGncstT98UV5B+V+rRc2HJw6K5uqeNs28njt
4UZHXruqa6u0vA3dwxekDY4KWP3wJ7fKg70hbwEYb07zonLlVjoS3shYgHA7ghywNT2idcCZ0WT9
79s/ByiSIcVq1YYmpQ48VxHoiqvXcL6S8BqBacKyFV4li2F5yZgJtPeduyQk4vRHJ8B+8g/4tYp2
Cq/qawwZU6HAs3ky4F6QjPc/jkpgZ5dQ3+2ErLrhWcPyMGEBDo6+9Gz71fsDIkKqtrzvS6opKOYU
12/qd0nQcdTVCzf3Uk3565eMNzFcEVx/BQ6mUmSYIgX1R8DRWbT1VmJTR6Y7wYrwGUy+uSIU1HfI
RT0HGMyj9/E48NLLDLuQR4pfWrmyZQG/B5t8vialMCoUyWGJkmEGlxOMlcqu2h7sC4sW+dESqPrh
9sq6TTOefawZw0dEcmc8D+2G+nIGNScg/61KeRq+k6EesUDDAEvgQ5czKm7JkNLZpXsd9zN8kau3
hLefInIfQGt/dYttsKuuqyOVuoAIkq8FyGBTDVkEQ+LtljTtBR1Ex7Db070+v15htjD5r4++waR8
C0TWb2XhLqA/LI46l0Y64sKYER+A0CMwl0B27cJ5s3aZ82If3AZEbKRdWVzxhqRih4libDe3vQIc
depq6SMxAdZmBR9RKzw8hieiZq9/rdBcCTKm2P1ouFyKfYX6SHt7uMQY0Yxy7vAKPi57f3Oa+OOp
bVzMJoLvTPqR60PD7QqZx3zw02QLEAbvueLN35MsxCtFubGc5jnUg/3UHxUOuVZT5p7WELMKDKmA
w7yhz7IWkHWNvnwUwL/7lC5q2jbltn2Esee7ulXkRE4zfBQMvtdSMeUNq/UtMjfdD4MWXZJve+VW
+tYsYB9Ltn6qqcyD5J+Aww8Se5JOP7M3AUgRJO45mKcrQM1FBGLbrAm7euJWPpEjb7Cp2gzoePq/
hIbwwH644Gje351xPoSShmMosCdNlAXIqux1OFd8TE/R7sjSSKWuKN6jNgjrk+EjLeLvBhL3IxtA
a1lbdz3pH2SaBSaF6EmwpZKEJSOk5xuG3vj5CVdao9m3X4zwSdFfMjqlCdATlSi0c1bZhPAMQZ6O
3F/uy0UgLoC+LiSe/KVdpOXnX4Q/RpygqVOewmE6PqHkZwSsYJpY7X1IaGVAtlh467G6+4YkQ3WM
2b1CKE5YSMDqVmODjZ5RDvw0oeZNYjrnsb0USX+F/3cZRFXyT124rzuQyFfki6qNruqWupXyWwbr
kdlduK5pmWX4pqL7+3PqnQW6KbKS6Y2Pda12Zk9qTOA1sM2Sbn6KXnnRHGClDZY7Y3apTbAh8ZFD
tv8w6bhMcZkdUtM/IxH3rDRo5ACCmxMbwqiYkNf9CtHfNeNfG+ZPornP4lZhzqLbJV/v2nUVKtor
naS0W1dMD24O1scjbZUiH0+aDh36cIJH/l4WNqOE1LVbrzQEoGh4gyaXmKctDf727Qv1HjkI0BPz
w3dqfeACN7LzvVCtc+EqUOYvgD/JJfCNJGG8rfLo6CdZK2kN68usBsQk3aWreenyJ2CUcBSfGlqD
tmea88NiQC8V09VbUeWypruVJ4gp9AtNVcg37uATOzHgbj7F08JXt5I/tYSJueRdKvuQvpYUEhZq
clPj8YJByo/h3zlV531yfBdxGZtr5uMAVwrieqtE1l4i1x+TwWQ4U+nOvP/RnhBHrlt7eBWxHqr4
3KqJ2HEdkXDeun6de20IcoAvmdcfjUobvU2q1peZcqQd5LdDijfk++kk+8X45GEYmhEajucL+s0g
0y16/yAMXV56e1+1NpEBqf5U8nHXIJDcsA3VifSrDODcmagWeFMjVVCpB8XPWJMrIuVJSBd22UlS
agXbILon5Aq5EmHFZ90Gt0Lz9XNmPRvZbM5dH4ix587u4CH4rCSmgcWDYCZZNaBo2i//lYjKhsFc
cKJN+9CTCo21EO3ydvXkrrU1lH34JGb6eBXE7uGcjpsKevwEZndlODJbaVpRGk3V3Q/LJk8h9i0J
KJS7pZJvhatC1BbjjIedtJtJ1h/c/yQQAf42RCq/dVs0L6EV1/JSdL5SQdUWfnjqCYTqGw4VdY53
7y4WMSf3bJufTfKF5Akj9UZHZu5tBJtR1JRa/WN4ZV9itjRMKj0q3japft9B9I74ANCD9dg+kca+
etlsBRRS08njXU9qf9bSKchjVl5fdvWsYHH/SjypN9gXvBvNymle0vS2XIuh1j1JP+bIQT7upsY7
J1KPm8i81dzo1fdERP+vaHA2OxZxi6Cc734nT6ieMDyA507oHvMpUIG9KYc7JrWz43waQ86e0k4n
G1Pq/DGXDAhlP9DKb1HM+3WAe8mvJNeyzXnUQuAvwGki60Y8zq70PLtql5haIFV4A7ao7kbpTh9d
H93wPY42SE7YHV7rMalRkjb2duibn9SCVEqM2yBSPdqQM+G7i3sZ1hao+R5oaaw6DRldA45+xyhN
vlTjITPMuQd49GFf5D2uMXyAVXvBXyq93sUDeHcOok/cQHxzmM5ybk0m6a+EO3LobC1Pq++az89D
wZ18cQ6wmsvijCcOVq160e0qCRFpJ9hEp1bMaeloyDuKXu7fcKws5wEo+azcM6e/exQdZ35i8rO1
6IAgoEjfiGm/8tLXDC+rjnNbVOoqfX3l5OXVPlh3LB/ThJenMtIMvu507cNbn1pC6oxZYvLElxbY
D4z6gWkgR2jsJzUwj2hXz9HEmQpuGvX/A0kBHSUvaus/Ijdhf7VLOKUD4LPLZ34zSrTUqw3+jxip
bHuuMteFjfAm1UdSBwfNpVMONLc1QK3MBwjV+kAaqu3DEqU3+XRXppAvx79Zpuy8KyLMcGnzvvI/
JexDDwGWSOB2PmKxnsf+8SD0lJtD1OPSiVjVlKxrRVhQs9ZiERfJko4v9OcSVBbUtjpOsEEU37UT
Pyu0WUPIkN9cpfidI77vL1FQDVO2djnIqDCirF5MU3ET6V+dksDtlfqex13CqQXqaHTNkPdN8J8U
Z4T79UCoMeDktWr+hC/ovcZda14bsrHLpcghUrXfgG4PAlVzByEFBUAA9jo6k2tRuk5S0xzzQFVQ
s/xj8/o3nozUzsP1pDkJkeuImGpb9xSToyI4jKonm2zKwxrhXgUViWMO0nfqO5TvBs67rdG/sIZ7
SNB4uXfDyRdWoSaPfYrcLuLS9RDUzUoU9VD91/8MyuT5WAm9lNSg4uELitDlIs5tev3vMAngr0tX
wbQz3lt0tumVMYTW53Ws7yhaM//3M5CW0pbDMUcpg6YS/oRzUyTdJ+V7NpkXQHdo7nMcezaWUCAP
I6jE7UJ0URTbKoyvNgTAmggnZCX/6jGgsYoIP16HKWCTRvbQHh3SEjOnF9mcbtjUYQbiDtVaPNuF
/ofVLJ7Gc5sV6MQ5ARTO3viWYEjNRPc3k8r7J5boG+SJ4PuWCJsiJBarEyIWZnuHWs8ufDQKRzcJ
FaORx/ZqVJDV3TuhFxgTYBqp0+hRpO1DlQ7fVi/V/pXcuFSl0nfiy6CIxCGxqr3Hy54GIxCUSxdV
pcA1nrIdtJBWWS+zhv0k1fgkH79O+/7XO8P9cNc3o/s0bL0mx1KztSHU8YlNt/uLfQU/TdN1izqX
gOGebny5nbG9oTVbid+QgJuCG7rjTF9kTtu7PtSyzIzTTeNx0Ra5007eUhSTtGwTwOnVEcPp/EXL
4JfxN2E934E7ALkNQ0eKHdZkwdMZN4i2Md9BePS5Sbj+3S2HBfrUy788u0Y5ruVTGTGTgi/znbpf
fFjK+kwDkAKJ256J8Mv254W6Iv2UTEs2fcQCkSGI8eEI2IDOnLNddKrE5umQrwkZlYDhYH/U3ToN
upoGoEJyZx5DzhdWBnyALon6Q8b/vvBcsu++RIt1OV2DrHq26nmj0s1Wngjzn0SkEUJLvDAZNET0
9RvHnW5rWbyUfUly8g090aX2naezoHjCbvxDm41p8zoKoMDRdt3UaUxPlDxYnGg5npaKqGej5F3p
k5GKxoGjSvAdfV8Lf8RRB7FH+CYEFMAD/JMB4knSrTYW++tuRco+jdNjIRuCGB79sJ0AqHj11AKd
cNBMxAPGkC1XMF9UPVqeK6rKXI2eL9Qts8UWMeIgSeglA8KBa0P5ii7Ugo32nUX09MIWh+YcmPwx
HEdUXRz01ohVzvgf/+vmSjUvYS7pIFST7WZ55/vsfoy48m9ZXPORiFoH+MvcG21eG1HbsoQCCLrq
FSx0OU4riLbEYuG5CjCZyo2+ipzpAEZ0xWL7FTOHXCcADL/qs26bkO8h/46P6rCb0y6qHzRnsLBI
IxWcgCWV0POX1sYc0wmDyFCEKpbwljtzZZ0CnvpKwIa7fWw0c9ECzefDNLKz8sR52E6+WraImaFm
EnYkwtmSPQpkyc6buPjGwJjNfnIP8gVOjcY59mH++NxWJIr9/2/WuuXdcQNn+ygA48cHn/3d7h2t
KzUdLj9LuBEO3xPJ6kl7/E3hHVTMvmeo3CBUi7BIHxz7FEdqC01jH4Zc4PpIcfNhu8JbrGWm70wN
Ac8fShYyYb+20htNUptE/8cAUFr/Gchh2qdmoPT1aGS9WPL6sLmd/z5+YnY9i7OFaScx/dfX6eqf
bG9ZC0yy8+TGOWlV5e7d3US3Hgib8Gh2OCyT4qpMflEnfz9TO0MuQ+PGUEBD13tVk9EcrA1HQNWN
J1NPNHcn4zpfaT1XSWdFFsf8nMqVOMnBOqcyF3fJNxMInkt+/qghy8zRIw1nbQfkh9CC6uQqIAXb
ZZzTSwIsL4Ms3nwPMnjeraVkxNH9j8fzsLO3duBEvsDDluYcnI1l/jo5+2hdTfKOULw1yLeoVup+
EcSL8NoE2PxJ0Bay188kU7fgoCPn2bHtYNwxk1zWnRL84PElehYcoDqvj9yMefCGimlQugVUrI5d
WEuauJc+TIVdN4DB/qVteT7hHS63QKy+74qJKQhIrqeCAJqOZZoP+xIKl6xd/smuxg09MmKaFfW2
TkyTdgVdVAtJ4NpLg8yDwYx5noyAgLZ9J83tOR+iPag9ZuhrUTqeA9sh/llb/PceCNwZF3Vjvu0a
Swug4qM5xo6Jb4xNeasggUvQQNBKfy+JWztP438by2BJImxjyRbkX47eX9huR2wknfk3Y0960+IL
J8cKHfozMrjeBlX74tIf3czviUjdFv/JiSdjkkRKhT+SF+mpc6HUiqcm5adCaFFRPA9LgRSM3Z19
tQ3D/XiHBAg5zBZHHaZq6Vdn7xSu3LjFq1s/cXFfY0EtN/K5ZEEjQ3GMUU5oRJIerQfRvPSywCE/
lCW3yRZhgEwX8gwfps6Po+TUbodp365zr7UkTW13LjG4oHJYOnUqdfNGoKPNvsQcolIJPj2c3Bg2
ddtZ86k12POzBUXG6W5mAG0dOpwCh35abJED5JTKDM/r0wWP7VH6DXVDC0/A8s9IW+EnpfGpEnfh
zcyxEjsxP08WNJesnem37fzJ1yK7AiB800zO5B5EYr7PC1xFxeN/1/fHUDtJFQrffRJ9yZ4PXHF+
HdH0ZcwyOGZtwiqvD8tuTzplnqzmMcK0iRC8kAeBOibQ+8QXorMDlfPZfztn/9javBVORnMBCJDR
1YhBnZ9rsrWjrWy01Pbsc+Zz+CLvbOIJcFnKsOtDzAZk0jVrGhYcFynoRr5iNB1y+aaQFomyOCLs
30mmfZklkrnA9Dg0YendGhLGur6HPGU3MrHSNkUnmiZ91LfX8NBCtxKrGPaPb5gFDsrpPtFKDegX
TseTS88bCyXjFpvD2lhWeFPdalp1AQCQO+Wo+1ZwFh1fxs/W7p+ELGHpDzyfHXlZMGkusPv56ElC
7VQgILMKC/lsbPF1UVlsSWn2q2a1luAeb6DJABqVjtnlYS+6sCoStPbWab9lRb3Mh4sKwrIY6rx8
8zfLYNUNwmSNZDdNN/MX9GXidlEAoN3jYC0bJOxHZe0SeBkbEIJhDJbjVVHZ5Y84JzuX4ksIv5pB
Bm++wMkbhufA/R9m/KIrEjKtcverzWHOz2zKCtEtVWquXH7Hc0V0WLYMDLyCsKOl9ttMJ81LZI3O
nSbfsjmfcLc6boMI34myU7Yo+kjsMguXK3ov+RSABs6VGJskD/IyjdGRb+A2De6kGDjfOpWZeCMZ
26rIjq90JSmiAOXxd0/PY0HAy9J1R1G/+YgRN6sOfEoSBfdtrzsXSI/I2iwmKQEdqHsylRZBmX3q
9yBOZ+aVKKK94qG9edEBiE3g3wqv0FR9Wm1lEqKXNHHNwZM36DrVn9hs/mUdLS9/jqYwkuZvOPDB
qJ0b7sIxUASjMpXj2kuIi0FIiL2eGE5x0pZG6QVDX1uxIVLCAQArij34EjgY6U1qzRQJXLFCGl1m
3XKwYrR102L3UtQD9CQ6AF1srIGv4LPjQdQmeI4E1DDmmWS1gpqFb3YqwjVkmX+C4rkg7h5OEmcu
+HFYW/s6OKDrf6NWGKv422EY36OK4TAUhCNR51gZtANzSIZE9UtqCCYw6EemUhhi1RHaqVEefAT/
doH+OrQPeR1bW5lRAdlf/92SH51il0ry1Ia4DmAEfVU5Qyi53z842C8dbZvgia2qik08Z+UKxh8t
yvmYmjDc7aYuuwpYw/ncjWzroKHX5WgzuFM4h8HWpUCLZ7CKORRl2RrMJFOLtahFoYzalSHofShm
poEII1igvs0Fm/PHGtCF5UAUkpWroidbv5GCbaNCHqr8d2zQ9OmDNog5aFY+LkWxjSGhydPKSwtt
GkHu/9oSGig9zRqXsbo9JgVe3FHD7SEm2SiESfGvs6fDsNpnjx0TRh2Tw4YGMjrfhzs6iZBQ8mjm
h4Ii+z2GUYM+Os8yQ+vQ3KDHvg5jsiE6H3+fHtHYmu7IB2db6KAPwCgtEfxjcPzzlMAnpbzFtHmc
+AAzStpS8kpEB7BJfI43XbWLWhPFV9PN70bUJQVLjCN2Zrjs+3by2Uv71ca4yCi3uRdLrnrxCeHf
AGMI/t+0BUPDh78rbqvbeuSH0xbLav0JvnN8gyLiQVudIAuIi6WHWEOesk8ggHXhyPpXP9gcjXQP
9ujL/wWDu5DS+cV7yi6uk70bpRE8UX81iqnv2ZDEWld9vlBAzQwmSgKW0NvEgQD/M3U29XkwSZ3q
ubsj+yocZbSU8TEUXJGUQhYf42Wfk7q5iVgfnJxHXrFe1Dac+RzZnPtxckgyXv74MKGwepsNfub7
ceu+aFV8Ic00/2WIhvraOFqI6mF3UJniBRz7FhG26ZsRb67+uxqYJKaWKtPnBGaD+usihOcx/w79
f2IsViK/X8UIfDxEfj8qnhMvXieJfto24SIkuMYGtbPmJahrr3rklue7/tc7Bh/VNTckNHlfwtzx
BzswU8FcINrrWH1FIAV9YE/iGsqOg60gnDcS2PvirzI8SRFk4AHoh8sC59MtbiVyib/EpqVCwo5F
yP3iJsY3PrHQxhawRjVTCsiztD0QwUuEBo5e1z8JETJnMM5UOxPhoDKiDp8o/kGdm54b9XjO0GYT
QQGEjveecYs6HFZ2FYpGtxTCfBtQ/iTiiXjN9d1vAM7pJA9+NjxiPKQcp8Ocnq3tt4QfsXtdF6s7
8qQkSz362VOk9wNT20VALAFH3B5vqt59OpkDLYrCDD/pB+APomn1rigrdPjXAlAVZIy7eTj0pkLw
/C0Ol9PT4f3Vfb/0jiUPBC8KvZA+vhxaNBH4qsmyP9X76ogsK4zZh5OorR5sQ09lO/f6NCAE9D1p
qlvm08ljh/xtMuBYj8dcj3ZUbtW1xuHWDtOC4T5bkyRYwPQUqRiiTYoPQl0u2tf6gAkRbPZoUSdZ
wnMI+gggnct2MQwhDKJUXXJOWaGgS9LRfsqsfshlF7vFfRthMiQoWCALGWVNiJ9FDIgsJXMWHUao
vBjk0xKf9iq2MqiL/hVeLpwQYa/nXnp3nFxuIVPwAHT0DdwvL3NaXqmil6t16nNfg9dzuOJgJG6F
XFLgwBrrfwPgVxLcJAU54e5nR3kT+gMgZdl+g5siB11OmizZkphCN0yEpNLsQmzWC4kQselk5Fty
jQ9hNDrhDO1BrGhIPrHl9Ks2txlv0coEprcPD2ZE/0ktbD5tljr8hOfyWzO4B1Y0pUy7x0rE2lK0
Qm3VLLgn+ebPkVhqRaw4LF3Rx2/vGShrjo8J1Rjo6BjJSPA/shWnRV9KVfemwCZM6X4qbteOK1P+
LcFfNwHj7mbZ3eVzHtdHfYpasTFYmcyhtc+MVWu5Vz5P8Er8w9T7PvxAOI+13x4TQJ36o+5dt8+v
Cee0OVWZaSLqmFcXOwwkV+dSGvNutp6IAxVqvQjr/In737wkq7wdYIsgIovb5HOz4Zgi66sbkvUW
rB+1CIsFqf9VnL+PerLdbhhQwjuii4u0nI2Ozze8wbRsMdNOP2y+XaKK8d5IsyTxwUHgK/gRbHBP
37cLZYIs7QKc0TCwEsH+A7gptbHMEwKmwckZc3ESxGluuauUq/aCaqObxf4ra5qyr/V7a8s5hRdf
4XpOYvNIXHHLuRscULkybBN2JuHosae3teZzOg9fbxGf0XN449AGT2aFBl6B8TAbdT+6TdnqKtho
pmxysKYI3H6Q7aaeW9mQnbPJ7VFG+zKIIhcnNX9LhKRfEsL1jpUxXLXQJ5NyJtvJYJj2a/zwun1L
yvthPMi+GbAqnR/ry447aQ7LyAJfm9ErqxqMtnfD1mR96GYUQcJA//9+iuHXJxW+C9wp7XD4Fi+6
TUuTEcLuRP5P2PpqDUP1b1y/UWx+L9a7FWmwH4mdJvMuHus+C/o5C/Vxv2CAqo7lfeaTV0A9LIir
nn3X8za04K0+SG1EPaI2IofL2Oa/kT2vWLpQo45HlMYP+uE5MVlJic1O7JgYpeQYVfs5eCAQXrFT
0XTNFZAA/4nIbW+jYh/tOtY6Z1980CVBWsu/2MpRcLYRb4zsw9niglYcSnc77AhDfqVglVXn4akR
pCNXhOEUDxMpVOu6Z1nmTy7/BVsEQk60aK6bts65SqBlzzhkVgLAy/3EPjkH6pt2YyEb6fscYf+a
tzU7oFarwkR7zYkPK4gRADcFRMpC8pnd4r7oQObNZYN6PHv4g6LAJ3ZG1UsptH9nvOrTWpprsX6X
aU7QrcvIIfeQOviJ1RxbzhcVD5NbKV066MxerS5HMPyS7cGjMid3vf5+LdrOaN6d0d+X8NbZGovM
p/qc5BwnhNaH5UdE7x/7S0zANlNCmqM9hJqrMFgv8vEBEGD+oC4TWhKddQRASczQCQONse73tVNs
sg7JlhTY013JNMoZBz9SJziaWZTWDiis/VOzW2+vRGMvBCOMN0Tg+NEWXPb9g4RW1nwxUQvUeJXC
6zWglLKYCmCu+p6rRUeJtrRvbSdc2Y4K4L9SZD5NQ2URVPg5kagM0o2hFPrINxWpm2YYKhsgHvKN
+PkeRUc+2JvgRXH94k5LbtMXQdisr71O4I1KfHl81DCBcahwtgbnASwvR73GzFu/7o7i4Jbth6rj
7XwJsS4cY3gpeJYcPbcl9Nw8eleoBsOj1teWjd0vkG/oRi2GX3vnw3yNm+uWv3/9z++If/zwlsmx
2yrqA7ig0ZeYx1HxNXIoZqEuRyxR8xs5TEyJX2UTbdDh1SVtxgab+8+M46i4JxJPvyJRGWa+kvpL
P6aSVgDZzfVMEYqRGunGz8cXEKk+namCq5aNgRQTBUchiHbTCVrOcfI6JwKcFc7epkWL3z8lV9A8
ssKXEfr+0ElO0paF+KLQo6OXdLD0hFrJKD622hazzFLlOovZVlUYA/rtWODfu0OoT+BFVUwUsZNO
rsrL89+x9u2ZO8OGclmFpoBYwWAsb6cmcbfTGYa4FQk0rc9r56oAjecu6Rkd1kh524d38DDVMSEa
fD++UrjQyGvGwnjp1kjg2VrvcbIBja5m9dTlQaH+fGw2sXZxrVXC0qgUxnGYQDl3F410jTLBYY6c
gyiJCusd7q68j3+yz5PO8wKo/F8PQCU0zNL7jD+hvhrRh1ibYBo7TzCoqf4tvg8rrtS7FoZ6j3TO
Ly3f+X/XtXJnJCgYF2VHQKax1eCvpmBaAK6U/1Y3IfCGiyO+6NbRqCztCVETNZtkL6LNkuWYjELW
6Nt0qRf5JsPirlOzn6PN7Q6NCtrO00OP6sG8vRO8YQZy6lIXfIbkSsg7CokoHs64878dRv0EjEf9
YPNg6hlhXZwqf+b3l/3Yo2Xf++UkE1ou5rrG3een35lOoRfBHXAezLcjeLFtDMtolcLyWHMaXNcz
FDYb7phZeyCs6wfsJosNM4Y18JN6vxY/w6cnF1+dpo4RA0Eij1BvrQd96hDldWHLST0WMpD+ehBN
FHrfbSbCxATp3cge551TMCsWKPEx0qHV+67Tb8A2hTUDWYxHO9YbSR6/PW2ALbvP/kusKoAzw5e0
COd2UL8tGyVWGzXtryU+0fQitLaX+CPww0UY7uHdFgui6dywWgVOUFBzG3NssTjfU2V/iGCpe++N
cxBj32Wc6ieIYg1hcVCmu4eET6OYw13QcmI106Jn+kfSJshSBFbc1oD7QYze6nCi0/4W9GkNceKa
1UGr1yEtEGxIWpwFxHCbBSzEN2k2zG2KeuBgPqP0LFjZ7wcUvxeN1NkzgRCxwvUDinS7ZmF4LC/7
9YuXmAmSvc+xBQXuCeOinNnQ6k7mWma9nPD9/fJD5fsBTVNcbuH9rQRyXs6heKtk9qc2aSfCg+L8
/JZ1Zb8rc6xzTeRbIHP/76+4KsWktABuDYt29Ef3+G+MOt4BwcOwpBaq3uuqSiWMNP34cP872tUf
aU1IuOxTxqh9DK8DJY3NLIxNfet5sneURIOfF5OEwmvs/zVo4mLm0+ET0jbfIt/pvqhV8ydhBLWG
HPHcFgi+4k1vHzBQx532x4R+y580sgC1dJ5H4KuCaIxXBlHOpQc3hqv8LSRV3vmWk7iQYQGDiLYJ
Thd7IZhxHtYATVs1TJmIhdDM1iEteaedWI44fiaRGw2wnCRmg5YornzjEzAc8GT8ERog5dr9ezfp
BPd8BdPdJSjwCnSCTAAPZDYknHB6jMUa/7bnnT8QmcxkJ/WdtY3VqpOH7vRqQhN4pR9E9ys+fwpp
E7EPg/XDovN5bp32vbYyNJLSOkAV0orNjGYC/xttfMq/w9eJousUX2t7AzXHtIF6ygzKdIwCpter
8/JDwqk0HcGeeo/PDZ+9PcUHaunVUPERRa7XiBHkUWdBhl3P9D3AKzSKNobUUkmudUKJTjM0CXBu
qqU4bsDMxvIuXbfKnZ7TYlZUecNXx75PycypD5QXcbPYAr+n67BVldbaVsorcbGcb+xLVMSp+bmX
B5qSaa7Q2r9vycH8jPaGUQBAiu/DDOEMUAJdYrBge/G4/qsI7IOr1+X/NeDc+g5/fFTfYOt0dZlp
KogrmCUqAWcelIhtaPqiMYvGE8Cd8Whhwi4Jiu9NGdX5KIMe81cld2X+3uvdt1m0Ei2gZXCGXLLj
PTtoBFXHwCvnGaxd/mmDShGApdd/yk/9MqGGE1Wuwi2rEe0P+TwDyAMmilLzVS+IkGLHybGS2N5z
XOTpJQvo6F3e8fEdI+ja1u5ld+ftoXGAnTMfuzMAgHoYkhwKAsIZTP8k2m1lk/+6AdEUi0nPiJ5D
XP9vx/+Ul+V7kXfPvAxABRkx4cr0bnK2XkprTc93Y1UOTFjpBmpholz1z4O1dnvYFaIG9S7ohvS5
C/Oge2o8jMwRs9vRsSwe/pIwyLJiS2fipd0p8hjf8vcbwiN86i+pB+kclRzMoi6+g1iFlCuZ0t+L
Ju5VRGOBmpWwf9j6Fz0nnmChyihuigr1s44k+zFdkulGAZobWP5qHyCBvlEG8BtJmKLl1Y2yz5nj
4bBn2MHbN6UD88OXDwpQ2ILCXUlgKu/Y1oRGVH3M9p0XHKYhUgjpXeL1BCzNm6f+e523jxTlB8Ru
2YLI+djzsCSpJkunysodIMBWO8JKlHANc3ls4K4295CtD3JGZl8zWwesGxTGFbYhPU6UurB9U3Wv
O4BhAPAMILRZ3bJhebp86kO5zi0Yo+n8DrtUyLnYBULlhff9/LFXETZ8WBJbnZcV+x5iopYNn+tu
gvCWX3JqqLNjld5X3OitbxtIocX4763jzlwPrIl5qKTc1NhiUsYI0t65/0MyQ5q6u8D5e4ckFhOd
Xck6yNlWV1+SnI1r3LQN/7ZzPX36KVjx1qq+a/nC1fblTpt8QNLYWjgTtaoUdoglXgbzFziXxV/8
FC+1brCSAAtj/DR2UvutnPXduTt0XoofUye6JM0C1xqujWpbomIt27HoFGSTDhUgohvCDdHpV4ZY
zrZlTBmGU1+h5CWXZuyPOGskBHQhUwl4mcQ/WNrlTlSnheHLXzhU0Et9KaFq5kXJLVl9+BqkLEnR
as0YRJ9SAUSp9caCUxaGpTJhZDnQ8ldhsZJ3moJbQkR1EbccZhfpk75gJk93UxyzKDZvNGS79B9J
TA/lFYN36M4qaYv+FMdETgGXxFHs2EwALfK9X70WDNvpJuqQ727L7ZJ+tzIwqanYcQEUtKI22LW5
OS5xE3sPlDMkvaplbBvOxN/FnPJM7zdLKEQ9PE/Nbhc6Y3ZrF5TZjUZpnhlHPW2ChZCtOSRaavhX
GsQRLrBDh03Q+d2ZOZ6jxNpdU/DyOxtaSLAnfeNiAtX41CGJfzCOsTNeUXcEAsqHn67JSIe3KCe/
oi3+OPBjTJST59D4l72o8x5iBBE24+btzm4pN6/+Lr0QPKkAFMN1ksKiw0TbuNVy5JfPpva0ut71
DminZ/r3g2SPbkSyYHR7g9a81Pcdw7tmhnn7nPKK+Oy2HNasegjoijRiJI0rANkp9EUSd9+MQf40
bc0bD9AdW8UWFwYICwoWgoBGbkUj4TmV+Bsi9jQOtHuz9qjpZl1meOJoI9e8eJIhkVqsJFUtd5mZ
W2unz0hzyoW/YXDDQ3D1qze3BeXRfh+jWwvQ3Gi3aCyhXIOl0c2o0w+mKJ5kv1AkzzOAA4Hm3QeQ
ElNoBz873Ep92Y08BxRGuXepW1y2ZnyW2v66qd8aVTXV7vzNJyZKAbWgclcIoMsIeLs3fAl4RhnE
gp72HmBwMOfyL80BCMvfzr+q32huqJ1u+7Bs+59gxnnBESps6GwO7MZjgyP+v83vcwZFbSr6h+cF
xSE0mXDNcwh5vEdDaHhw3E78HZYz0FNldh3uPHMJWR5P4d8935nssZG3PzUpYV+MEPa3HRc97wvW
3ly9wdg183Uta27OIYTdil3vr0ycw68d46Oyc3p45it7d4i6u9KWzUAG37OfM1GAYvqX4cMFiCm4
x+q3e7CdxGQouAlMYa48nUHU6piBEX6XaTysrA5qXbhBCBw1bwi88b/8bb+JRC3IsbEvtvLcsp+x
8GTL8vSyrgW/LBAVg3ODDB7JCudvcj40LjuPqvJzPRl3g/AytvrqFmhUhZZBkkdqrQGcWln581pY
WHTUqxW0T58pUHdu5PX7iQd1k6O7Xr2/NYuqguKs3kdYbjrrEXgMcd2tBe4MJ/HYFS0GzFjAudr9
Fz2wE9+iylNYREfxz0s5v0AABuxUH+t6pcDlj00MnDWE1hFPBcVwmT2xNmvKxXFFaLtOhsBSEu9T
nTHJCZoOV1llbE4iLKKRb+B4hNDHR/0p+esf1FAAJYkw1QRdVK+z0khfXRa1Bj89ZMea5pBjJDcO
K/nM9eNcwZbAqT6QnR2ZBxaRNgrAC2leuuTbp3T1ogtSEqlDRY9I+KPx1YQYKcDUnudLz+mgTgHj
ErIkJGVOaWVh9BFmjAxpoznEQ4fWB1sSDH7kQGmfDjv0WmALgU7yQqgAnNfDVyytgHKPyHRzbMzC
i/D/jgmDGpIWRlSG/a8sAFIcJ3bCd5yi0PsmJFRtKS0Hy8WIXC95+kiBxPDNB4F4xIsN499OgzR1
8819UzoVZGAePgQbvE1GVIW7VYbzQzrOi+QaqCxYORwa1jSK+XzW8tdMKEniQJyzXv2nYHKp75yN
d/WRdbr08dQOZqZGTX0aHaj/jG5iWI8XYMBrHMxZqE0oiDi+TanOyrzMBe9ghSauOvPlwOA8TED8
sncwI+YpbGhD+rEk4A3z2fxr0qA6pz5jvnz8kvEb6QruDE2wsG6Yw46IyrAYsMfibgq/n0GEvnPm
n6pMjx6eAMMJerykLmotpaWrf0tWxNoeMlBqUivqWb88OECtUbHRLxuSk2lq4OxQClXK2oyDyq9x
QG6J1JrpdJ7AA1D5GcxtZ6miezqTmquGb1f0PYUfLQqnxcJqTcX4krEDH6RSPhmCqsQ5qzxyuena
so+XvTAk/bmgxYa9thEJE+jUjgHUInTc1a3LCka9E+Ey3+8vqhUSdxt2qjkZ28kKAuxfbU3r+0tF
ga4lywSx/1qDsA3ETq4YTFvZ5ED/UlpNmdMPOg0St6Ek+V5g8v/8QnEkpgEeJXJI/Hyc9NvBKU+y
BQrTG2wZ2pGKUv4GrxIxgE2ocI2LIGOlq0FXveRrnL3zisUJVAZ8lbVORBOAihzwszer4TvbZKPS
4WRJuk1z0ZLTGIYoojLINgh3dMeKJCGftwMwqcYKQF3qn/vEkQdgCv6JmbbXPcQQcISMVfB2Os2E
5sEbNS/ldhG2h9reOD5zPj/tBt9rF2//Nzmr8sXtILa6WmxbmSJe00tpXkPZ2QX416nZYIPEx/aY
b5Lapr3PmlUt+Rv9YipArVbxzAH7ziyjo4osEhD7xSUHP+rDaaZkqn/JOU4hIVH7W5/C3baMFFEX
SXOT3QUJ2e0AhikRjvQKy3erwdPiB8ZovxmlonexvX1qXfSViC5A64ozTTObH1xUPeu4DnOkKe1w
gtfbtK765QF4URd5tgyWx1PlaVQs6N/62bNZRPTUWwupPEzyJmv2paltu6v4IFzHXGoIW90bFK/S
5l3SVWyrGE/qBc7mGhZgJWGiN/OjdrRTKdcuNNm4HV8MkFcAKxRBqxPQKnAIOi4BBhZeAygSqXoi
N8LxpiAiOdlgVGsIUdC4iC0szE09Nzuxh5SePXpbFv/ehKHkbRXl2ZWd6Xh4lyk8yes4cxte2uJP
b/68HNk2PATHhXM7LnwdPmExHcsB+uVCCYyMDzfhDCydLhwekLV0dlw5QiuheF09Z6phbT8KxAxs
OXaTnRxWK6a/sB4mxdUVGJjcB+XaBo2uFhgXzKTzHgSkU5xEDRTf64z5oRBM/eNe3tFUT7OzA1HM
oo5xpZx/AJ+26kSBkBnEGGCHBQ14omdA6FuUDV81moHcu5KepxgpNjLDet3W2Ntbtao5l410Ibh8
eLTg/8wxNG8ff/H+MOAAvHzwKSv2CoycPWvhupwSuy0ng8jp6OCAl3U2aI5FqOKpoi8H7WDQ9Dvp
WiGXL+MOhCs1BoY+BY9C/aXJScuV8BcBtwxCstl7NZ5PoFfBD/JzN8S6oFjkJn50eQ3/NjKYAqIX
5R8Sg/GqYP6nQH8YsbO/zPXU+ale/NVcH5qMvLwcD1ZELVGyAOvIBTN0Q0AxaPABue3QGxd+DHSQ
UFoNhgGOw6pUUSlu0CYcT6L+3RnPb8YUeGCSYfD4GqBe1bwFzno8FONLE3jLU/6rNJ29ZwqY1eSw
9fw4C5aN2FGdtHvDhdQnM6MSV2ppEH/sxK3q7pa2ckZSeXzQqPworiCT/cl9XK2dvPvn035eNsgR
7vSvGjsiclYTfryba6yss7ggQGh1Hp4gAAuMIRVuhvUX+A1BqegMeOfLxUFMhc8M43GH8++eY9Kv
6wWYJNZc0jitpLLiZKc+PLDLZ1GeYGL0TzSFzKGZdM4jldLnICDZD2UZ9v2q93OfjU8ffmawQTUT
sfHRmQlsrmihQ978efj2OHvBbbdLUsXV6tpUF43HkHcUOCGmq3tx5qH/lgoCuGhX4aggCFUo+k2Z
0k4RMk0x8AnI5WNw0p7iPyLXJi6dSZv2sv4UXsdUemuIfQL0dINgra/xaMYAaj1aCX32tYYYtDzb
7ST9ls2kQAu6rWURCSfn+li2YPst7oVQNcOEbsL1+IKH24OKX4uz1A1dzTIroml+O6qcl18MsOUX
hklTonMQ/c0ggFKU7mPvpohqTlme3YxYKXfw//7oZnFFS2h35ggpkKn2/APyWP9XRURD/eRl0tvl
4rrrYrZ/4N4V/8aXsZAIbNzVGf4XkNZDGjuPHyLabFZVL71Tz7SZiCYf4SQXYTsdVDtbFLvjqT9y
DWiw99oooXo7iHaBRt+CHGMOW9NEdIvVKjyaux9fUaMd6Q41s3HeQETNti2Zvje1IOMvXLfYAkHa
3h20lv2G2YgxvMJWKSOvRpM+qqMmTfsuodSPmf7N6FMk4sDcuKLAcK4kfVsxWrc3IMVfKu/MfcKC
ZphL9tlvWKdB2ctLU9QcMsOJfLQv8D5x7sOAVd0JYJhikqeEG0PNes/FXWk4AOYNXT4BYkMy2y0Q
Pj3RxdkHf9VJ6yz2nrF/SQQcvTgdMdrFaOm+iyfeANRgfAi/BtiycqOy+at4/1JJ2+CjjY09QEqK
BkcMLl9NXWIBZWoalkTQgr29yzavZGRxW2G7mNY0HKw5hPSCzB+ogRCzsRGJPCKRzexQ+nJl3gQl
gEJo81KByx5cNXW1IqFOwE/aVEhMxfPued9iHltAd76LSU2pvV1MgX52f6YXF4RdcxvqoyQytdae
H+wzTD5JevmfB7ZUvQy2jO82eVNTDcpNpxVT+5Ap3PLTfBARi7TOJVO0qX14N9ZINiP1o50uAh4L
87DSZ7zHcaz/HpO9HrjSACQOsxi4giE+uVdi76qpwCTFLDRgrdbYO1eIk0j1xgZ5A0GryieTMgkT
XDWMN4oTn4+4YO6YZyZpr4dv1WAZiMjfY90hUTjbL1o2XhldOUZHa/nswGX0o2iy+kaIvZNbkdYF
NYwGK58Fi4IablC+84snjkhoNvr40U+FfeFJO+lx3BDG3sddsTGdCKJlSAvQbGUf1wXgsoXIQ4U4
OQm3Ky/AEfGY2jHX8IPX6TSzCXVLR8beWipCu+3b0ztpJHuaVZz27MC4EfLve/M7UhrhsnowyPm9
MU4Qxd2wTf+zdvX2uaEPVyDYM45eo1DQUFPHwLhUMujdu5LOZomdOP82wBcpqVZnqB3NxL2BTI5N
LqcbzzlESK0jxN0z2P+ejnf6ZVQXpV+cF1yVPiCbtoG4Rq7nGEbD4tDsFffbZxMj1uRX8+GVztMs
aIUP4seIuves+12aaegTKp2hDp+vVbWurGIwpw4gsv2qEujDxS9FOUNPHC0YdyLc99m9RL0yQew2
sh4qhUxVf5aLWttbo6GlC+Gsfp/H5leRSxA5yx3x5dy3lO5eIPvL9ghreUtp4P0g7AGMxcnKORuM
5Ka8j8OfPuzcKp1fbq9glvNGYTxfsIq0aDjVYD7erkB+cvcaTYGaEu9hCvq7xmHVeQMtq42z4nur
IRZe0gYCLMJJFCDbg767PlX4tAh4kw0PBP1/Hd5DJPQUdWGPJ9nEo16DsQ1uJceoAPu0gpjMujjj
Phvr+DBr+nrfDD6TevszshUyKG4jOpLvmMBLq1KRwHk95g++XatxNAm/7Iqq3njhTSSPfNqwcx+y
anwRFN/UZ9cO+3MtEOKIWfnVBGUBNRYXcoIsHrjMsmYUehlqwIMcRa0mzJsF0XVO/ofzuua+z13j
uryMqqeJ017LR/V9BtMDjjI8AQSsYyCckQ0osZTRHzEkRvwIN7xO1Bhk/zl4gk3Z/jXpE6xzVBlb
lYNrwSWe3j1VpBzBBulEhGjeiHOFw3OydA2G7GW/Pz6d55CjrShMxDY5G4OPTkNViXrLOITXNoaS
BH3RRz/zd5F587p2keUtKMx21p3bszYwweEEghq01lsrsoaOcIBtok30k7B9TBPZY0Pt1VSb82d3
G5QY3lz/isllHj0omFj9UsfU9csSH7lqpXzhR8XBb2BlD1VF4fZPuxqL5WIdKecT+sBETjfXW/NM
iyJ4YOBMPH5VWBFOPrGzuZCwyTbHpR11OzNv2lRV4OgY5gtMmNwyKk23G3JTf91X4Z2FGnL48CzL
fOh9OJi0e/FSWzTr5wwjn+JB8LayITF7RFcVNML1jA9LSL/SGrfU9XV721Q7g9+q7Kx8b3Fl3epl
EaFNm0yhJhHAEW73d7K492DUNR4aq+qeyS91PAgmJiX6zqNUjxFuxg5OQ5jt815lde18FVI9ryun
28B07p1aagQkLL+D41iqMHcsjiNQx86gJ6t/KEj33xpPfmTT8H7yxtqB5NILl8UscjFPLPhzVQca
HZf4a8Zq/1nrTt57Z19Uoe4+JaPuJcpFty9ivvvM0hCfkkG3KjyHTgn0daNTvo3Q9F4uWwyrQ9kc
VGPUJcTlaX0vGIrNsWLkC3uLzX2AJbT3ZibeO/jXKqUjdAYyH2QvUxWpR2hibf/Q0JkqNNsCc5aJ
51/V7APRtu3VkhNTru8UXrAriubHVb9Xgo60ilR6cTVu8HPpovobjfCVeLtfs6ExKuxgsK56yfHT
salwcChe2HN+XYdeI+bS9Hl9nhfSxYQx3kr6Iot+vzNn0msxFGVgpzKkZD4dupaRNvssqo4gkNHo
GnsoT8hiaahQOW8hFdQ8Mn60nC4lO4H8prightFnjD9CJiXw4kbI2W+dKNmybm03Rfb1s+cG0qHf
kSICSPHg+fo8k5THdSul9WX9WOAKCDIRWO8I4bpsZnkGqabKKG9UVkv+3VEc5hUWs7WrPJjgRZNE
qmda7YNZBZufcCH7S7s19lNFIn2BIT6prbERfMsvN/mewwwMGGl/PAJvLXiGvziPvl87yatUo/S/
O8wFG7kewBKr+4N6g99ZIp9FGkFhCztGrGeO7qlrsCnUoJxcxoe+5RKWHUhq8Rs1B0RgvhGyH1TK
qTkg/nvMVj4DJKedcTU1RYHI93j30j2Sq6lFaqngH1tiD348YRkrU2svwoXaaAkxb2T6zw3c7PuH
wwWurqhSmw7Wtg+uM632vGJfUyQK0BlxIap1T23BEOONwVwKRuXFaxNHXcWiqMgLxcrIdMTWtZkT
wyTkqFNKVbgKmpdY5Z/Bpo5u9SQpxGpJmMM6kO/8Zf4myDDZd1R9na6SaI5rOi9pxeMd4bARmgE1
bECTwuVSIuCmS/1L80HHYzqai7aNBfUikfeZ4YCh95IKscgbkI/6PcVxt9ynOc/6aEHZCJzEyhBe
UQMvXY5bT9YwUvQqeGBeTvNSgB/HuQCXMZ1fi9UaZT6/5FrfL2+Ve8N5ghR1X/al7QQkn8FUEt/p
2v3STaNMAyCpFm7fd54KYq8Y9vli9uU76Lei4Wy27Q6MheEQQajxQk575CiF8rkg3BcmpJ+fPgyN
sOtKY1/nmJL7FB/O+nI0DGAS+QQK2UrD+VpzoJnMjzW4THW6T2QWtWofeMKUL+eVdtHCl/XzDQz+
X3Iwu2rQLVi1bgs9jV18xnn34lYMxy22ziqtZ0V0JYCG0oX3kAyMs4faFaZ8bgDrBWH2kpY4yvMz
BaKq2xZQ1GN9wWDVnUIq8yiyK9HrnPwNT40TjMWX51D8uaMYYyZ+8JT+WiCSQGBleK7frGCiRUA8
u9fPbaiF99Ed96UbCoAhWSFMYERIbBWhDNpfH/kMxYvnilCIjIqyMa6eeT4tUJszZQc8KIMiGh1B
7vHOcKpAcGlM8prZN8zE9sgEok764yqJft1ZQr6EevLVlCf0Dv2pP7qWUpQVLw7O7xIpLU6fbri2
nrc4rDGoqi2QmRtJXRC5VRVUMvnD8l+AZ5etOGQUBeG7Ivop2t9iEW7km970Xk25hUy6oJZnY/0U
QfsTm+Ke13EMbtyWz992PhjYfz6a7KnuCkA0KHHCc/2CTux3lyvsg5BuVJzxH7KmonnhkcQx9tKo
uZABJmrxUxHR0p0n+RF8pgvjPWQmSCqybPNtJbOnv02SZOVqU2LehsnDfCeNGPmtQbF2qtQbTMzR
kkmCJbEcZ+fV6edEsuLVREslj86/UCYzFET9yqrVQBmG6aHVgNz2hZ4hGYPefSVBAH1KjvzNkAo/
odRxX7Hlhe7ltH3zhofk1Hc7QIKphXVIzS4Bs3YJ1R7vp6ebRpTSxQQK9mD0XtYwkUuPWjLPMQer
R4BvFsWmj+UOkF2MZU2hEKM13fnRgTHPsKJGxPzD3srVcFHj5gXd9vfqVYRIeK8xd59OsW75E1r7
lRNJF4KJ94oqVgWaJiufj3uvyKzDLwpsWnOZZrExaaF5vV1i/M+cpTAkv4JvuBrqMKqNa3cTwozQ
+uVwq1RufExpewU/G+30y5+0Oz5b63sJSmMLTUrcGX6578iyktn19F3wq/dUUGCnVQtg1AJeEdZf
eK+CLNI5NSMehkerGRkHhJzBbXvruKGkOuB4lBN/NuY8WBfuG186W4RKCULPGCTZhlA48xpn/6uZ
ZGJYEa4Ux8HrYLvF5YfQMhQSJbpqHiHCTbWdflFLiudXAmKBnNgh2G8TSICdO7Nra/fC3C8D+Kln
IP80uYiQ5W/bD2xqrLDQ7tTtlkPCkNPoNyzrmdRDDMGT9g1EFbJ1OPVYYmc7UhSACGRjs/YBL2N8
PpiHt/24G6z9lwlifS3iOo3Abh30g6Tsc1uTTGqur33reVVtewInU1thSztKIWT2qiLk8b+WNUIQ
grSpy5DOtTz8cdYFq+IoOyM61Gglia4CuUBmep0M57vNYyh1qfGFx4/o/XYgco4uYbpS0To0NR0D
/jNs6IHzpEJciPvTOSqs44w1kW9CXbaqS2fykBR3/fkVPla4UW/XFzmBKNfw4KtXhWqTSKOy5PHZ
V7nk93nChSdXYmEPIVRm8qCFinf5h5ej/FZMinjNVbw39GcN1xK98IoeFQVd29senTk7sVE0iJRF
nbakN4vwXzjf4NLcglhNWqAq0hnFfQKPkw8g4VmC0gbaza1P9Qj+6RSTa0wEKh4LmiCZ8c1LHhmt
7OX4JU4YKd2lCIkp/LdlnoQXMIpDgir0yGOAbV8EYJo2WJ/7X4GiFcMV4VsMkSyDd4AttHkOTEVA
M3QfZ8bwbBQyEAZCiPanArAKZ6PMg+g0U3jiihXLsDB0S0si5ZZwSTqAqSGqN6TNeEC/fGvBjqrK
Hap6CLuTvDt8EGdpKhpw5DpJMvX0w6K2at0IHJWk1TXDgs0uuL2ES5d/AYNKaDF5CNv81Hq00iaP
/aQnMHVvIs+EyJXQuzOsFmvGBDc69DOi79+ikVl8+67K7U8srRwGXw3TlZ0Dv2Z4vZabyOUDRGge
t2R81RDQ64xFCEeeRazfYM7WRF7nyqV7DNClI/ugloB+1CK38IL8RgGcJNms3jNGOC+muqRIv8DG
B5DXOnfI2b1Lb7ASbopFdMqdOCRMIMda4mSKMQsb9pYYagRwwSoTiOTxBNX2Ll70HwxkfsyaYZ5A
FKXXb11FjaaC7iL6RGt4/VF1fYeKDWL/fz2lZ7Le54cX8mdnGuXCxbwjKqsSNnPnvAlKd2/t/F1D
W0pTqJfIhCnczUjmeMlL2ocylQ4NUcZt225wuoJOxBut4o+bC8KQ43cShiMXU0HkE84vjGwyNtuG
Z8P8Am4ojKkWHGyGbyta674eWz0r8LybjJmvBEktItzu4K/KmZMQcotUWYZgeD2Jg+bzSqh9VD9d
PrjH4kkXF/VUCRA04aKUChs873WTG3XsJrtVfAYhLsHNWJ+sXUW4tmu77+AqBm7a6Ml76J1NEldn
+1CIObSF8mbccMXqFBvCH18N1WkOBQbKZHAXc8tfM/fsr2kWzb/bzcZS8DmggnlviJM4T1ljv99P
EuO5i7n5n/4k/iW2QLL1epeawFEe0C0HoE89cynuuCNHPlMEP2jY1RIna1vFPh7zVU64vg9bpEkn
SPfObACQA5sO9cLHOsYtFS0E76Rqkt3LDpSjvUabYW5QmI/+9GXoiy5lbuhypcEKGsF2xkZPk/an
/Lfxjh+HbpSZ9eS2HP6+lxqt6GJ2x66kvMKGaLAkpQJob/KfbGz+aqVp1tSRuTkXKiIqYNFH4JC0
/0pG4fULuSVe7Rj2UCGjvgNTgAnY8E5bU3BemXoImq7PzxnpZZe+PCyW/Qa4bEl0zVX9u6KRlRrW
taZtGQ5k7jYBPXBd7NeE1MgBHa+WChDEzO9eeiCecbBrRUmj0ccsUR5XJfF5l8d3J//fXzyza7IJ
jn1koZ9cqM948TF27rThKk9FFYknUyQGVbsiBYsXhJbIerIxjM94djeX8YC/XfxhOfKCvTuj3vBO
6UqqU3Y9qnJzvNj/SO44eaJ6xaWEs9AOlLuWplMs/XKmL77Ucdy+RDYBMyL+yYMbHtO65wwFhgrO
Gf40P8dT+afmid7lnQQyBgGPJmYkYTlANG0NvN1OZzNYQWGKctGQV1jQDeJ8qOqCpe1fkZIfjuwL
GQnAZyy+T+k1fWxNOsBkObUJ9gX5bJcAO0YwdPFOhcCiOUYVce5FaK/gkUT2brUzPFAFr/M96CLA
SL7et5h0A6bYsW5KAO1u2eGRmBQHnEcfO63PuEjicDo3X7p2QtFj95itG4qy4qZOBYFkPsFISBn+
dSABdho4RRORZzJWTiuIC7QbLEguDWtwfX7EtZ2Pp3oyI8+DXFJ9DIXuvoR5siRI+09iBG/facT5
ma9Srjb57rxHaRUqwUfF1Mcn46hRfc5OG9ADDQQklViSliU2fVBOo0BHKrdOSZVSAxUXRSdqU2kB
MAXuHt6JjKUprszHkL1lImO0to67VtfLwmV46n7hH0oQpj+KH2yU7elvY3syKhC2vWJLv1EKwPfx
fTNFDqT1WBrEOXYw0RtD7T3TmU5Z1L2jmtwelBWa8zYl7waoruo0GSCKtNftxCPcSltpilVUyDti
pDOYi8mDDM7IuB710TPJd00ItifbBcHtHxIn2VYasrO4JdMkCo8WDFsQUu9sHjNdNhkDfuf/uRaS
rrVnk20NSAd6MyOyv8uaJzRHYe0SSnAUeUS97Vlgt4nSs1eeYJETzReeaVXIejZUbJuEWyZoj2J/
jlfwcuJ3UGnboQ1oKLR4VxKgP853/jZVaqWYrmBF08l06S1bX2FuHvSuxKad6w9taROC+BAADxzI
DK/ngylFAMFbMGerf0Le9RdbLB4fn19QYKqP9wsw6zvCnxUVusQtpBW0ZX6bnkJ0eke54RXatSsj
LLMHtS/IINQ2j8nygHomvpFAJsRj7/mvKIEHrEnMn+5b7lkU3QQStdhv/wRz8yRm/dQ+xm6TPwWB
XXUpRb56kPMr+CZc8CALhsUohkA6FKRGepIdyaL+jAY9H7WQlf1NaKqwKaObwKA5E4CMof+sNxgW
tEvUa7FWx3GdUOTJ4pnV+bc11P/ra2yedvq2veIoccbJWrXCXAF0ltsuXd8nIA5idpSHfxwpqk4Z
RQUfcuUn8pK7ME7sC3NIZ/bEzUE3qz93WE6l6qPMeV2zLPjlpKoA+mla8PcTxkuk1fIS2k0E7NoT
2bEW5sJa+33NJhNWb0BZRY4oNRs76r7yW/Mf1nkqZzeHwHgInwMm22WuMi+CbXCtO7zcWy9V5qLw
qaDmFpDOj6iH2tWF23tIQ19amdF6qQfZh+MrFpGQ+z9vqYCgDKINNQ9yLD3KQ50YRWzvZmjdJbC9
Sj2x1ica17Cri89Gi3XeL6pV1VwycOgEDdTFvhe6EOb759S1WKUorxw2eGSkiyUWWrysuSnJvcEP
34sop0m+wdGc8Xf0YO6bKTs/dayxPyzSXgf6hf8tOueSrCSecBk6t/vT5mzculr1aPwDrYePBPOn
IczPp6K2c6bBHPgI+5052FLGSj5Nh5JzbPfIMGh3CBvi5kk0Y0+YSTOBQ/elytUMAwORsBlQWmsX
8I75hMJl7g+ZCizXXuEjyw7lJ5FNHzl/jaXF5HkEH/7rPVRdFA3/kpIgyMOdD8QAlWWokKltyHAC
LSTLWW/Y5cjNi6mJMPZNXkFfLw+BIa4eHH/fYEoQjAKzXgyG0QjmHdnQc584NMGu6HR0LUgcf8P8
e08D1Cru1qeY3dRaFmMUHt7WUTDA2ArYCOGI76QxZO4xKoqoQuqhTR2j1RyMMVrCHbhuOsCkb4Mu
+vAs8Lvd/9+37WzukTtAHJHJdwBNgvcl0dZxJiKW5sx/RXYnZoQ0HRibl/WAVwr71GtdHviv8DZL
HFH7OvAs9fkyadyeisLtbQShBbf69sq4PUs/EQ2S4PITrLlZRfpi/0rWYNWD/oUfABQzBTogv/uu
FlOx43UcSHACUtbIYooaMe3chA2x+6ZxcsllLVqh0q7FG7F1jnXvEE2yp/IoxnqySRl9Ue3cf7S+
i9oe8raZ3+vUTpFpJ+NlvvV1u3uN5QWLCp0bbw3yGHzbTHcR3yYMGJ28rMDGuIhLkBfbJ+SUyzF0
S+h3tQaUHiaP85So7U2+KAFKKRXn3q078w3a6KNPvSWxy2X/qJSdAUbsgmmRUjNrz5/auwXROMvJ
aeGiutihrrbaD8hZSvyJKZAmtbRZAXr0K60I4a/0Bf2eWlf81eQd1o5D7CYBNG1gA1+5kRu1lG21
olk3BM2daKwW3b5WCugfJhoyuEwOxkhjA7R8RlK6r9bJfzYCmlrNdev6H98C+0ae4gTTskxt+SPr
xnr3KMhvP4XW1y4W6w3QnDhA/p3in/HDrdciRvwy55kaaNwd4eKLQzAC0TQwBKFPhtzZMbk2dE7c
oPhcbojzwDH6RIaeVIggGo8F5RZIYjaZ9N5fFyRR2JoCSpi/H9xSQbJiynsE/EZK/S5mAyhzBgjH
uGbw88gp0AluZaeN3q9ouJDe8o2+l6yPa9UwILGY+NNtZy3dWujnMdtJ814TmpN2KOFQ122u/nN+
ZKKSN+oo/o6wHVmHuPk2ZeZpVbBsSvJDLk0IPi+2Gji2z5tepvntm9O81xqoLbKG6PSE9YlU10+p
QDFIFEI531gxkgDfRNhiscFmOh7k2/xEeYsSAiYAA72qy0Tnl9U+58t2/suUARPXFqsa6+d5lCck
ltj9Aios084lhvt3bIUip133mU8N+DkEFQ3naAaAC8AdCg+R9YwI2TpFfF9r/Zjy5AYAAivvMg8g
9Tu+izTuoL/7pEgXcg0qmp1sqMxMAnN6PN7ETrAW+3WmSjjDC1aeNW6+FKlLLAH5Vf47x81+jqiB
0nMCbDDBzfoU/9hCK3NhmhmXG9mQl/Mj9rOaI2FlUVQqpyaIPmYmt+YfZ+pA7Lz5WAMXCj8HScF0
u8F//5pfhFSVhDLbNJL0xanKYMovVuQ8gPm0wx0ROcabfIxYSEnihqu2u2uRA7PTQHODxz38Dt42
BnZ9+l78+6jug+Th3GmHeIm7qstqbgoLzoIAsV6hmYQSdY0vGEfLtqjU442Pok5X87ZPttZ//Uqo
mEpwybF5LXMhl/Y+L5Sm2CTeX36iAlh/qEROVQKqgt8wRhcij92WOKHkdClCXhx++RrPU1s68vmm
dk2tKRxa8k6XOwWC+Yi3TtyyiLPWIOVsU2N/Fr8SnfbHChicr6xcLJF95IMfsNNUNZ9ArxEsyWTh
D3CEC5TS4ZBn4RBGsOHGVDad/BRY3d5oL1+Rj649JmGQFai7smraNxGLsrHd5Grv1EXMMASynk5Q
cRhmpdxwbZY8FulHkCQc7anU2sOh0VGBJsOFewtpjRyepjU6m7kR+tLStg6gQt1G7cMAXZlDgDya
es1fdph2mOxMKVIVFLLPHBkw2MQR/4fEMpAC0irA1yTxCZiOr1rHCBOpKp+83BA5MaWK4w8C3aLA
o1SkZHpH4beahhwSofYUO4x3jz0Yw7FSZy2wgtQ2nzx9jWazhIuzZmavBe5SYkyrroNFScvSTsXq
5KY9ppu62sdgGN8QMR+ee2noi31RY85PYJJfGtZ/5qPTRwZXQdE8z/QUIXB14y/iakCXDiBGj+mp
w9M47EnP8RIVHTMlFcLuZpVd8pLhQR7+h+3YLuaq3mNolVETTp5YlEDj8Z0y6BcE/Ai580h6mePe
omG6HvdFyIpbsdJYQjieLgCZuhI15vXa0ff6k10HDB923y669RSOPICqFaRAyor4S5uKyWNIdNpW
d/MQavhvMZrRfEkR9Gn7LGkkPSDoHPvpsBOI7giK6C5dxR7s89rpvuSMrwIo1vpc1uILcb+h6sL8
0eqBnbZgQXy9/I55GFqzdFe+nr8lW1OwYIANj6m0E0/WPLurRa/2+JwE6y3tEMmcWNG+k4lnp0Q8
khqnnEUloDvW4f3ok4vHwPFCvnr2wHJG01pNhWoTNVgO5flQAOL/lvWC5MjTuySn/8A7T+da/IjG
6GYOizCmS3msnskSp3z4HcoocXUSziTiWHiV/O3KbUxwCdCqhwskBUl1jPzunz93V8ndZnUOL0KA
SIraV6icd4eyfZsnxauTq+wkrMjBOE67hFqWQ1+d9ZlsPRVM4zwNTOy4zhA9zSVCfsAHrOLEitzn
1gM3hCmo6x3A/rmRls4TordVQl8i8o8oy7hwY/7may9UsWuDinyARSmSW+GQlG513AnXwahXurhw
IoJX2NSj5hP2DUa2E8v5fjWjwuuWZYF6ou7Y3DEhngOy2H8QVhZ60PLHXEwKMN3vTeXvApvhx8Z1
ohf4zZonA/DccD8QAipo3s1MXP8T7TBvKDSpBggPnGc9u4ZJQewc41+By3HbpRrMu7Z0s/sqf8IT
xyO8wNbnzywx8hrXRrqLrq6v86MT3/4UDvJwzfEc/OlpPSpzHRTuW4Y/6Gd3JnohxrTqaDyr+8Gm
30BEXS3idZmgqWJQpJXMiQXHH7Iv505ObcBawOE6Ut8wO6v/jiSqYZftRzn7zzhuTQex4QT9lBB+
4Tj03ntz2fl05Q+feNGAKyIG3WZmWIqeHN3f2eNmOWP/ijuvQSx1R83Q1JSHwHTKSv2DUhH6bYlI
fnE8KpUrJVk6v+93qqIYeUQVTPj9x6PmEY/yp8TJtl/z1fmqtO2G1IBFKKpYKfdEDP5qqX948YDT
c8UL0HxJHD8r439boobrNvnbQS5s/iN9E9zpsYCMZCNdTOYlplEUsuxkDtChtlF37wkwkmupq3Wd
85c/8RZkIhvIzZtz7jY9xAQXdYaz1tdCk1VTpLRUlfH2QWJT7NFFk37NL9diIJXPVodZH41UBFsz
2dqhpEWTUN1BQsEC+IMnFgjLeSkHYy6M1ToInVqmT0+IclzyyD+VEVrmW81LZmOyu9WknXMCTO/b
WlNHIzQs1c45uch2ggmXCM5brhGqcXn/fMtI9aAxuLG84ESfKoXPdozOPun4/izYAPxxahOiOjVF
rDVNGwnI/3/ukLxcZUZE6PEBzcsJblxcOrqKx8DDR/dvp5fzHI/adNYnDJkHCNzXHVoqaTQNGYNv
K/WXHLQym6KhW27rSsQMFK6/N3zCaTOtgAtEBg7uRVFVDpriW84xpyVbFe1VcdAE+taj2Cvk0pgb
6xcBDz7+bXftBYJEXyVwu8cEHSb9Zmdm481XcirmcoaRgcMe1YQHG2q1gievyhqlTWckINagtLsk
8IRD1ovuraYSVQ4s5rIMGkjvSVM4K4ZCyaKbLbXq/bK6kfO7JCQ9WK39Nn5wpJoePiL6V43iEGBC
Wli/9eWT/6IRp8uf4sxooeQJWAPlqm3gTaddQ7YW1BuCabtZCFKuksRYJWh15DqgTBIphXYHZcZL
cus39boy3R3dnLlp51bpaX9RcXFDhLBM7nwD1XQ/0MXDorPFCR0q2h7KYQD4xoYFkbEQk3TMNfAA
dTxnrABwzk119sXcKEFNCyVUpIjBOyllTe87XSdtC12M8obAzlcuVGpaOQ8kdgYW5nZ9PzysNhme
+Hqp2u/7ZKy6XQ/0rC8q1Fm8ofC/x3MKcgm5mvPMyfTgiw3cqMTN8421TaSXpu8Vu3PjFbPyj+kn
dmoD164azXi/dUwUfSyMirxnT6FH8vNlOGNtp8SnJ0TLlBXPL+0ydV0ieNGBTIcjr26ix/npeITU
AP1yleLybe7wL+txd89JWPe7vav/oFSpeU1CLvCN4vPrhITuXPQzrDtK0ullLuqDPho3QuFKlQzI
IVSOJZDltecGI4c7S6IudpQmGJLhz2GjKhx/e1NKEwMuvivm8Zja4kkeePYznJX2C1oe6byaHzvz
YB7M2SwYdhdA7IRFbNlszXtqAs2YQJGFWUqdSoO0/JchD/BkOK5gFuGcBAztF+Q40kmPv8mgFIR5
QdqVXKGXZGe5SEfl7Z6LHSvEIdKm7/GhGQrU34/vZIpilcIlB8Gd+QNbIWObNjC6AIC5PPb5cych
zwmHp1GGP2J8FMsNyOIAht2m8gDbUDIqmHqgo5/ENUg4NC08HGAmdLr/WwecNL88CS9bwdx2jY70
tt0WScGh+mXaSHylBjWvoB5yV5Pfkv6EnjFZmdq37ZCwc2wGNar4fK75OnGWPW9kCrCffFSadDXO
T2H4BcevPE7NghXLIk/l8NX7sVWMRHBp+k5INCFDqg4j6sVKBhJygbHwdF/v9bAaRPRn7qmoAo2+
Q/WD7tqIHQORNbmVduSVSNgKc7HRcRdArvNt96AuwBcdhgbm5HlURg/Oe/uBm4kWvLJrGfmS/QfX
XFqoZ8Nj3J3F0L4PCuMx2/cJJDmZC/ccTzALhJ4bFzNEHlOiqQuv2LkcJ+TeL4PVpJ8QUFqq2nrk
ZZj6Hy4oueMomXJ4+7xsNx/YHMI8gl1QXF72hmfJnUzOXr7Fb6QRkVvRv3D9f/JNSitqB/G/bhON
ypYL5mST9htOhNOsa1vUlz3hYilMqYzX8wO+Gn99VWooikfVYoR1ibJVtkIIodZgoUq+utXQD7Za
iiRcRmhKMHeANvMuJtybrfM4ePRXkkJsikmvxVV9TeXJCS779gQkWKWJAxLVq9v6/X3GR6sjQOTP
hmDRx+MVaX+p3W35livSsLVZ54o0yZIDWQch4XOCDnjXpz9RYj2e+Tjkuz0+IIeo5E8Ez798h4W+
xD/6LtHXr0K1zyvkF+kOu90nvNFOfFXTsnROGw4nmCaZaFY+8YhZwMcLS4FNKEyV8t4Eu3r8Kvl7
tbqDKTFu8w+gNgx/fGznkdpQbnqMEwPdyoVHx90STugbRDerQjeJu2ouYxBcnoGy29hukHX/xyBN
jQpsE3wp3HJwNckSQ0y5E1GJ8c9YoLFEBdUzkHXBxJzAjyHM++WoxXQd3nOb498fpX9ovHQnPvmF
dB76PvCGOYw4u8/5viG13AVn7hrN0r0p2EPme9nYYAZztBky+hpzI9LxraQI5eG4cIFhGZSGpWQs
t3i5deXTmndRLB9/3o5JhojUIdWCRsOvUmnWZeETskwaBrC3BTRYnwT13qsGLYSFJHKoAaubPYQU
1P6MMPC3XuO4A+l2QRQcvH/V2/qoDWSz3YhYVxJVsLd6JIrmWaj0f/TVE8TMZNv7kCCSv1WWleqF
n3SJbpLaGR1Z6qzI4DN2jT26MFNHBhS75pkvsqzvdWozb183xCnzOY1EBiu6dipw4wAca/D9Zgi2
yAA5FTMyReAK4XL+UQcpdfQlZPwQzg6jOO3JcZSZwbtpgytIniARPi0hqAY8ABspwWBlb8VZURXT
j1oY+SjEwHTphcTU3Upxj2voFNfoO9+8kOlS/d7Kqyms2UTtdtuvrgDxYtERFFfthV3J+6AM8FZ4
zM5SR7GR53Y6m7suzSnJh87CdhpfVqCrhprPrzjWZ4GdxeCsfAOKmIvKgdTEsEtqv9DMqkYJArWj
rTpBZUnJT0cePloM1gYBDG7VPO/bgl51DAflChaJzOYZ5/uwLurIgwaQ9z510blzfOIAnDeFyWBs
sC7LiagI3LbL0Cxwl3mBFfnKLL/9NNmixqtDSAFhMfptj2gIlnioCSzTIDshnujiGwdc/S8Z9jY2
4pSIXm+qGR12+8sKa37FQavWaStUqYfm8hrt3BfUN98nsM77z+J6CpxkVdYppiG4fsReY8n34gGj
L6AOM0ZcvPX0TfOiReaJAiojA5zsqtn1mMQseQp7i3V1MAG65VeCldQpLuhxY0vCW1b2XfGvnJ0t
g8N8J56qiGG3ts5UAqge4Drb+odXamXpxzeGMb5oUZKPtZih+Lpq6JNcq8vNrkb1BepoJYoIJBap
xAWswERa0z7zIhIvpi/7qMR//wINy4CoGQer7ddQGiT9T7pWwdXlF1E+clRZ1qrYAi3jVpqYa36C
nRVdFHqMOgjPxOjbKutZlODBM4ZWiVcm3MsBse4MrxhCOjqq6JSiM+WiDx22LiX6Dkg3uDacx92S
Yj4R3VLcOQ4FprCdTrirH2bWRrU3aFsMGb7cUQ0PA1RwIRUSNyU/fXY4IRtitSh/nuugWh2eUan3
0z8cfkYgXqDSqDlhVTOzr3IRXt5DDu+xXOPQQjHcYtrl2p4QmAARkG92ykNy6BvEU+ORQ/1gt+24
fOPqCMGHSQOVj880MZ4uG2O8+gyhvtdkM3wjty8/8oxCQBtkyQdH1vh+Dbg6CICAJXj5t3rz4/n1
oD9d8cPTEXSDlxNAL8+FGa6x7H+aViIcA2nxeR7NqCNDGYV57oyDtdA8VkIWBmGw3g50m+3/vWLl
7ldIm0XCJTrUD13BXIx/Q5QZZ/7bQ8WXnlLqvqsokde4uR4NM5IEaH9QfCo1wjtG11bPlc0HJHAF
DpHqxcilRlnMcEt14YPuGEiz8Ar1sIDxcZJMevd2h1wEkCkzccIr+uQ1OzclJysZnKAcGDozh04D
Q6jG5mwqpaPXMOVYwH8mlKGdhPls4eMvflElc2Qf9D5o7aGhd/+DzPPDL9PlyWjL6Qs65NUnuY+f
3ATPi/mt72qQB+LeqAQbpwAjgFXpGEWnoHi7xO/KBLUz6C1UD2sVJXEPEoFofMa2dKDlqWeIuwpd
+ZlDkzHGfH4eCfKjyP78IZOdodeJx29f9J46Op4uSy+aAhz4VvkAgR7A7FWY59o90cM21OdTSWh/
UBHkCDhX7jPH1IEAnD4/pt3HTH96SqIF+rFd9VmSMq0JIhm1Ajw5AVGQJFx42YfdntcqnxG2sjl6
RbzAZ6Cypi9/5HsVvmDIUXSKHWJAWOJ01GVD1rPdup6ib9+xBo6khWBSGCxJaqkLPL3nvEHQDpVp
tk5ZM/RQW0LgFamXoZea5FDblrynf72CmdaAF6Df3b18PdEVLywAH2n3kRkk8vpMRIMPMl235pV6
jaUG1uljnSQTEJWBGP7yMOhP+Y48SN92NM+t603gKgBImDEoM0iD98XHViB/74GyLnC+9RO2QL6y
DkHd+UOGqHZgnIhq1kjzXe+RC3dd59GbZ569PdqTj+uXmWkaF3L+zDQkWEBhE3xlPOfTwwM7h7Xj
yvRBDC3gAIKPs15/7JHxkiHQv+MeoViLAY6pw1XJwnxpQgU0r1n8sUYJkHDFldlPEKxl1hcT8nUV
RKbAM2bwthF9sjjYN3g6Eh+QLsibGU4yj/q00MN4LNN9c3HbKNTQLjD1lw1zC8RAnWEGgrpw33Kz
fnSw2xjIuV0s9JcG9jKzh33yDOHarbBvQcftgFqTAb+1Ys7Zs81SrI+YKQKBobUhj0UEH9PepmtB
9n3AVxGTZsQ2ukr64ZxrqoFB329zkV/2zZy4v4baF8E4K1Yhnm37s2yQLVgRx6Nn/g9t7V/RVHGg
jsjXnlxT60iWMHonCnjvxMSbmmLGV5QJ9xW+YzVyEIfLgULMEzIkjkGpqxJbJCQue03u8Dsobqum
vk6gyjf6EHuW2yZrbwcZdDRYcoASE9qW+Y1k/pKErpopVOcfyAmq7S2da/7wyYDoi9OXVhPVEQLO
5dvHO6sVp/Lh4EZaudvGi+0/HrjWCFOWTVioDUbV6upZzru9fUVvamlIERfOm0xVPwJ6TL1Z//hp
K9i4Yd+/hrmIkZgCMM2ppWarM3sgSYlQhWvoPib0UA4pJGBOaVPUhph5kXdU4wGYPS53B/a09tqC
reEzQHXTCi4YO6Lj4IqdA/qFZjCIjAXdmRBaruXqFDyCQX4EjB7SGFopovGBPYp0cP+/1CvxCbLH
VstEQ/AH7sU491Tjz8dmH4VCVyP8dPR/L0wJI0/13oXdZGAtYzOjAslLy9+mqDpH8aYtqo89CZCE
I01B3ywtiPo+4kQvOivnlP6OcJOrNe8vJM1kog1AZmXmJFKdY6UnJbnhhwM5zUStN4T+e19lQAvJ
a/E0zCe0zCGSKHNm6uT9h2XDgnvqQdUaWOOKyiA1oTBAaZsSRt4clSaGzwFWQUXJwcDPVvfSLTHN
oxBwJ+cGicUM0rnxJKuNt+kUSCgRgLsQ6RA09vBVV7/mjJ4ID9XNW+5AFys3OXgvnuaPxoN4P1bB
tU+G98KzYkjkNRpviwsZSSsJ3dLcs0uVyGYR4e+5g/Bw09R02W0yOY1pnz4iFPMJkv0e0RJCnbNq
uY+7H2n/Ep8wVW5FnxufU7GKD0LvtHp68zpUIeGXAiIk8n/gGRFGKQ+tC2CZ/zm6eeIwQjuihB+I
7P8SOeQKw9y50YJedxSfoxAgQ8fY6axxfQrF4esFZiD8zQUVd2bM/+Nj1IKrlgNuX8mCJ6nrSvbX
zi8t9oQk0LA+A1k8/9xS6+ZDwdNkXZIHfmDecnpHVM6axGzNOvIQpsiQ88J8m91ZpyYjl+tVUfcy
z28o13gkQnrn+4TjXPekrZeximnLhT4gmxgD0kDYLV+2wWy/lLHz4yfHMoHgNmnxKfogCtKQdIz8
lX0aWYTO/r2m7sgtfCEfpAOwyMiawqVSoJd0lEZTOZwznxjMQ24vwxxO3383dL3YDRa8+kzaIuDs
zIT4b9fM0ZdKCVVs/5XWeczKKkSRWkmAin2dElXy0KNIPHr+Xd1uvOQx7R/e38dDwHsLkk6rCQ9K
6BsfOykXgnEIpenlTaGYHwZucksvwgpqAhyQvPgUT/Y0+dWuhLhS/Oz6/QdC+gphIoNa0HYVB5PY
Cy9O/g1M75o/7msJ0JrNWIOSo5CEk1s3p1ZH8TuPsQQWqBUz7VLJvgIxKblQUwiy7TvN3TNxFh+0
e33S/04tMzcpBMS4Dh018I+PBbAPrrAVq7DK8wgBP5maNAqy+xV12qi/eGQXjvPDuP0PEisOtmH8
42hYMD09GDjLhSKwk+Abl3Kgk+3FmTsb3JgF5cdZNH3Y/uisarISYlu8AvDNLhMDLFrmzbY3QlLS
yQgJdAjhXZ01+C7GKxq6yS0A0Uzyk9CeBYZ2qE9lAkrAYj8s5ID4Z07LwbKlIoXUM8gVISwDlmlm
W99DtA/V5nbOY9kuH23Pq4ovcv+b9Qnt+loJskIxLNJO8cUDQ1SVEVMLVb/PYLX/EOEVW74DO3oy
coqr985zAZlN4ymT9j7/AbOZlGDlaxlCMjho6enefDexf9I0wTRglzKST8M/GmcyQGfCZ5mM90RE
oYIS+xI3Fe3KD6mom+v23CfenWVhMcHW1HXUCQZqwTi9XAqPmskpMExnYXUWpWwjH50pPutn6Fpe
DQWfYLNGJz+MwRo5FtDcJFrIOzosCVBpPlpu8m6grIIYODE4SxF2uiP6leWyTyfnY8hIU6QsRyvN
oFmANX59ylZXywJaDMvKkOzCMIFi2yUz9IXcfTSAvZ/H2Iku/8g/bHsNo88PDPLBe7yKpvwuJVIi
B2t5ouYCOiCV8lfpjU98EQwzG+6bhZVu3mu6jfE9czk7qvPvcAAQZajr7QAe7QMQkxy03bwMX+z9
FIwwgolMhj3j+61UstIK0BUPduWyc8MRCN/2gKVn5jsjP4TDGaDGDv+zjd2Gw6LazAextneuBHwx
PBWL7ekBhxlhFDuFf4lvhbebnuj9fI7+3cYCeq6QGaaTsVx2pIIT+Y4R48Sg5UfZn5ce6AG5K3Xz
EeCzHXijdmnbzY7JbTOziIV42aPZd+MwNK3OX9lCCjFAdyblfmjTS3Szm5uhybOdgNwTgLubryqW
FfTZfMxZD6oN0Ufuul8ygKWzh0zCfXPqInsx/8GyvZ3yb77e6N+UmcvuexCH99EZnrEa8CmccOWy
kA0Otd8DXz7ZLEnWBUFW2Q/RNYVO9CpEUorXKIvrsfFoYiwNZV4chAXLY8R0MeUsxdph2jEEIsKG
72tCMMK3dDhGDwReC9SbakYY9QNHMseRUUXYacKpNMPCNyTFeOGKcGxrsedERKr1vi2iyxNsidsk
/en70+lXgh0AUA/857pkE7Rydl8QSyACzlt2GhswIcdHMi3IzjwGsOz2iT3skFZ4CdExpgeEudhm
ShMqEUYQUoA+ZOWq4w0FCbn3h6odpeC7Ejhoh580jGwZzaotiF3kP3NbXMLF7U0dDpxSfOPtjnT4
3OnjEF/lyEpJPycvK9arbQMuBGwk3MU3kPppVOc3WxGlTk7FIvmD3RLSnpIMxIe2f9roC8u9zae7
/zK3WbjxwdG7pI38rDmWjS9A1HwlcaXTOgn6asa9yHSzxGmJiX2b4jNI+N9PwqB/nbIWq9SI91kL
HVMtS/En4LK2GwGQOLLrNpOVeKMhUcz/tkQMP9gqirF7RZJURxSRpCYD6fCwrXdV622rWhMU+D4F
DxkE1EI1FwtYqsTpGWZNB2aBBXZ/80zXsC8w53myxbyFlAsUh3chc04fNG988+2tRyiaEmmrqQ0X
fUoGolbP2K11+ChoxDim8d2NPGDI5yCMU3YNW8xoEM2i8jWUAf9jtBSpIQvq4/1nsBC0YcY7leeS
m3wTrkiyVFjttz+cyF4zIRhxLXYWaagfqXfypWQYBso8FIinhje50a9zSI6VVipZ3O447P/92cK4
pUS4eA6jpjNF+hsjuLIyFCAKBz/N4XO7mzmofcgvRPjb7StZ9hqxZ8FKduZ0Qu+1Gxu8GSXOYwb5
6SFk4qnGY9nopIeWfvPFl3i1N0EEz0Li0Rv760PkmQq1FeO/Subl7l8nm6EN+QB885Sc2I826xFG
3SSz0RgQe7KrYtBSPu6bRsGhjlVAIeW/RH4aq+2ZnyVcLMDvOaJk3KpEmLrk4yd8BpnValxiJBKW
RU6MKHIsTvn6+pkAyqAYtjKGwr4YJin7te4QZmJce/ctm2nU1S9vy2uYQ//ZksJCL92Lh32l6w8L
RPd4LvRpp4Bru0ieiy1vhJqhsjbDSKmIBkWL9tUTvCKsLo62F3VZhhhxVi8/LihLsoebCQUyeNCw
jQLpqdwCspTJKsLpAEvZ0RdF90L6iUYVpDeUD2aK2qjO0SHJzSonh6kKSlUmRHNulDQdS7K7Ae3E
6dD1WASfyLyroDEFAOiR1Xs8UezYwsLI3ykWsHJ9LhOZN6TmaTLvatmqLPJhVq+kXXXegPJoI+zj
fQctgnmclQK6f2il1fqpTfIGVc0leHaIoeNHotJeV1LZFPO8SSDcsYErO5Echm5kqbyuceCjJFac
ALT4NOJIgHWerjnRsfhdtmSAwcq7Jat7oep4BsaTThOuEKAV+fYLmHDoHWfK5vEj417ZRwYoL352
U9v5yuU55EXbG3cwKJhN24uLqszAxmJZT3UNUQadbHtPJohuiHenkvw7AYHc9FFKLIqJQPUtotBP
crW9gODDg+PrBBEo62eJBw/fHQHTHFisgYf56nPqCFHvnLumhVCwRTht4bl0MI/c8wLqwwzFem0o
ln7+c6b/FCrjrJb8lID59ZrkAd+0UHC0gzxVY/pQ6Xcw85caMpO5+8MFneehkGNUtfJWIJU30tUk
MIxBm3Wgxj3evDh+84CEDIE1YQTlxwNFDSGa+tpwRdbZ7u93vZgpYCIB3QqXpdwSbizYgo3CcWXZ
I/lozkLH1WB4Vj+IEEvShrYNIjCTEAQnAd+QC7LPFhbD6A4PinIviqpdoLe/9VKGwI53dapoejVr
amDuoEszEL0/M/Na2pmGo9EfEs8NMxIWDOIoUmZusWEWg/KPVGwysiqe0sYjEzzSy3HugiZugG9X
BzlcBhtIsdjnfOnkqKm5EKWJyFB6pphtmhH1gYuo5yoDPHM/KoH5wYBBXxBNXJzzE1RtJ93qVcEy
nd2D1vrJX+0YvwR/eKtRrVOwryPv28+UZ6qcEznsUX6dnGWtQ0wbDskOoMoCk0dIc3t4R1LzMsp7
2YOdXpbNeS+wEesRpn2XLqogfqw+VWpHa8MDeccltGtqftXb6cE3mj/+43ERXdfTndaQGZGCapWw
1862uTXTto+/HUrXqdVZdPqINpoVxHS6VZGh+5w+vplNOodKsJIk5ETuiI6iy57iU1RzSewjEHYJ
1WXDnQXGxwlIqcB6hrDLAtuJPtYaD9Ng2gcHOT3NfMXHfPEIF4k8BPzxB1MpdntDMUCZaXop6lVh
0EMJomDphrtVhk5vcrzjPiYqkpOGv9mL/mfCAipLgZgvZPI6i4eUtm/kogmzGmvE9b15LxlOmuHZ
xyRFujW6ZaOLTHwYIb+JdS/7hdZJskFwQXSmpjeXiyeTHElz4OPlak4REbLBMKR8LAeZOHD8/Pzb
/HwIOk41xz7mVpAplhhic/dYpOV5ie+9COJt84kOGjW7IL9iazh4KdEaPB6AAO32h0DI03th4kZ6
urL6inAAKyBmhL1iX3Kw/Er0QltYYrAT0IfDxcyfBAMnakEuEEbcxDs24UP2Bo9akQHWJ56nMMl7
KCGgpUAhEtXUhIz9yiR/XZiKMnsvxxeQdJGxIPFObOYAhimFvVI53lh7Wc+2RbPli3DbvTtZvJGF
IiGpeoySu/IR+3lxXZS3KLfNdtZdfolOazRc4rX5GcGoLw3aWCDPCGTZMIS4/x4MQj+OyRE/fTEx
W2qVN7fGb0E4r/BjtVRPKR2niFZ263GSID2dW8e76YdsZhCJ1n7JLDngIYN/qhMx2/NA+V1U5JTL
fR65gfGpToM9tuyJ2UCXn22+9wufufUPDGs6JznBugLNMmJqVTacCheEFScyB/rwxtGulA25g3VG
QUgnhuXL7PKF2bf9RLYYC48oZtzdSqnslANF7TT5utzdeUttqtp2c6dGxHikKUUWhJWZSGiLN5HI
WreO9jCJZABt4GPHoriPsVbx0dfSktMXkQKZQCEfPJy9uLvBBJCR0RxS91osNBfTg6JljEyQSJC0
4g5R13LMz8J6iyCjj+zsFk+Kgad0TY55XD7cr54GrfJGMgpK9qZKQqRYFDg8dXnpwSM7QPQHl/pr
4smy/srGYXhXTQvjrNOeJq1yTQ1sO9XtPl6Dbpub3CmJ0VZHunY922jog2Z3SIvNmCEAmVp9dHNH
Y/L+4xIpyM0TFfD6MQgNjr0pf/bckqXzz4iCGCv/GdSQ5Ipixoz+V0kd+K/uehzwjsC7j0a30Iou
S5vt83QEwdejvlWkpCDltguXdxgOs5TlFEAc5ihLZmmoA3oHxLWxh2ET+OEUywsMFOcfpKokUKpZ
c2S2Q/ZjgstB6f7uTOscI5pAq7GopvVc8gNOCWiBDtgO1Z8mZ49J/fYscxM30bR8dElKmYRXtJ0T
gl1SJ2IgW9+ES1WTqz0mg4bc/RT7K2fiElzN+eTr2Qe9uwO2gbAm+9gMzP33dxkP19hj/1uLRHsQ
9lie9L2T7Cn0E0AkmNXai/i10NMSQrfDH7AR7qplbm7JyQD8L0j+hOqaFmT5EB/I4ieB5vTYC7ja
qEirc+7+/E8YsQZB/HaHrFK6w3EEaw7RJS56vW/6y5uWHU4WGUCjbCdCXcuFK611TOs0yORFDXLe
cdiAaJhiAOXzQqBo3yVKjxVhDQ9FwtnGVORODsIfwBsFBr8GJA7c6Wo/aT7+9Pb9hLUxkYAHBAwO
L6KAgcMUaHUBec2swgz2qmp+pAj05TVUonKBntkKdi+vbHBQ9pmZeNLaQYz/ISWRXVAMmy5kjF0Y
znF0jdTVln94EWT9Bzs0U8rgSp4xGVKJGfpNzZm3CyBIznXVMaf4ybJch45ZLD2Ut4QPNA+KIH3o
vv3EW00314SnmBlDJVlP4a/VXBz/ViZHcpWDF9gBCpRiGjP6qE0Jtcj86TPkl45BctOWIVsKzbwc
Uy6xVCNAI8FmZHCongO7sNBPF9MWDc/ujgtvKoqt0ecxctaiMDcyZ7NbHalK9HqxY0uvOO5RWbad
nTPgqZ/eEWkx7HuRlXxFULl3M5bUQz7UiOuSbGdx7IfdM6r51QPbiBQtOn/Ndvw7NB/SPlWeVtKe
vwSgapGwRmfCbgytckfiTNoClXe4EFryjFX2I+fBC6+/M06whqBzjQuotUvZnQIcB9PA6onXgHfp
KKE83D/yoqkK0NKNOU7l8CO+5zfFStpKfSKzQQPavtH79fmIt/CXeDwoYQA8Ws8yVog+aa6JdGZ6
CTy1NZY7jqa9gXE4g8CyJ6ByDJFRbun2ejUiyfRef0GQm3DuKk3HtycfAyOi7OnS0SEDBxM/U+Ue
N6JU0vimjgaQ60CuVnMNaGYRnBcu8omugvcVA+bCxVH+WJfUCjA7vWBGqVLNLk/1wQQyuEaud+Bq
RVoz62EuWNCj2zzBSrJSvAb7o2rieE/RFfWlqN22OMpl5UPlYe3qR4mkhnrEPkhFxc39zYB4P3Qk
GDy9WxXFc8tRDUvI2JwEO4US23uaBpYCW5CU7BTr3icDr1yRcnAucduFOpUkKR4q5Zg9rQK8femH
oOWSBI6pmKYbDsPiaVpnZOOGLEqEWbjvOOBnUbJlfwel1cLtLfWcgFPbmlrV/LIZ154miaqGj2/f
19uBr0PeWg4Gw77O50Pv5teN4UYIurom8gcnjWE/SbEFAsXiJcdkXirK+M2u4HCoBnGBT014GKYy
F+a1YuC/jXXAQv9EbL5HMatVIz2YOnKgJtLXt0zzFaOc8xi0S5VDpVIO246aXAv+ApM0KbsbluTm
XWpDtDUcxaxrqtu9pYf42kJ/QhE+0wGKQ9nT7QeedE923ppGY2rNiamG25VJWT/R1+HgTuzJJTpx
XB7AJlkWpPJCyEaiDnu3eCPBNfNxNa+TDj7TlHzGRiDepb36j6mD9Hx8UYGtWALlhUxGVzZ7PXew
pbDHqCk23tjrnKEbxeDx7ts/NRmMcPTUCHzSU6TP/rlTiFYlepLsJtXfCSfHg3dvUvPb45GFY8B0
QXa4DBwyY1NUAdoGNfkbDMcIkJ0OfCCe1wllNocDN9OlB/aEX8ptSWdG6HVfWavJ2sBZmdealsUe
Bv6vMpAOW0SPrw6pJ2O/JW9Tma5wzXf65XsP5e5dErO/KAa0K+ZdIHA2EaLc/6aAi+WAOxp/C6Gx
fRoUtmJ01Y6yDqTZbcfhucKdhLjaMtVdrUWHYPmV/45fQfqIICuUQYgj2/92f5j0g8Xnc6OomQVT
JPEIZWNcTuuuizn3z4/hOhGMlDACJdgypTXhnzYMCy+FiBd2tPwwKQTdxp0Su8s7OWRZj2lqFeUe
5YcgJGAz5CcOagyRZCpOwjajVo4T0gravkv2AwomOFIyQu/WiL785hY+Xoc1hOHE91hP3OMYPscj
mO0qliz9ZtQ+QFC9mx4y9tzFIPjpmqOo0ICzTdA5LaafqfrfgixZBkbvFcKbgp1pk+Mf6T9wibPJ
BK4O3+u+22i35AXeohmk8C9Oum96bPtHfubEGLUTYFsRBw8scELT3YRmUyTlu3ISrp5B92h+OKxl
ICmhRKPpTaWbauaKUpox4l0sIEwP10qjT88YpUiGNiF5g8gLop0ONp19pdJN47pDkjUPrT2E41uj
VQdZ9EWbspUAANemTX+pSdxLmxfSKIvWkI8APAeQapc0zAng0ZTb1nKqeUVawtHfGyK5RHeIsqrF
1p22BgvMugK+NaXMGEMYmZ/JsyYIWfXX5zW4VURurvBJKDVzBuqvYep+rtMtdnQKWC58ka8kkgwS
bcVmWlWN8jNCscA8y8a+lfniwvYQkgfpXIwW2Y7mMvwEVHlIhZ2+YfFTtt+3SkTkmgPzUeMNZET9
qeL8vNcEqKSpM3DKUsjCOQBo6uOkLdoXOKHMpeUB2H88EsIGKHPGam7Wn8Ck6Clf5WA2fuZp4768
r0LSiS0+0ADoYmrXycz5SzPO57xoMJR19dSPUVDR8hnlfCxP1R7G5m0sGfBVrKMLGoJ8TtY6o0on
I0mVUbP9mMpmks9Snq+dvkTyP1Qm5duWrG3hO2nWGChOYHSFM1T1zEHv5JdcAwjYCJMsdeTpM+or
zU/Q8OKQhoqOOa0/ifJo/ziqvXLSFnHa0zTvONrloEaPGoH6w0DeUwdJV//U7nui25yFkoSJsm0T
isWy4qgTCsIfWzOTjg4tcvbs/k9XiIYzopBsuLO6GHNT5jxXE3vpIuUrlG4vGJ+XWcBE5WfUSBEi
Y79/EoPA5Pzxmh/BvTkhMubUWmcgC9zjLU9nqqbZGkKah2qZ6obzV6YIkU0T4WtPtZNMee8KDTLa
5GskDJf3hxtpceb8g5/IgUicsfiYNI9AscGA70fU3tf3OPGq4+77Q90FHgWfvxQHGKqQG5af/P0s
CaJdyfpm24gLT50XD0xAJmwmjVExkT8Hp94RXVPJTy4bF+HAtIINqdxX7QMRK7RAh9JMZmPeSrzb
3+Wh6lWVQgPXpIc45roXRXk+8jCLnmZG8KXbBRiBJ6QF4ai49VvEJ9qka3FHNtUpeYr6GDd6cbCt
TUwRo99uvU6fH7RTp3CC0hT/6lVTdX8Fb3E7CHg21w5zCa2USeMlYK8URWoI8Ht7uASNWeqTSwii
wOcKUXxsoxhTTbjjcwWcixbTdXuzF3Ho6fWzUaC0Ag1Dm29QZnD5v8WYXIQc6TQLbe/iEH5oCuSv
jd1FesCz8EMKDFYM9j+ZtW6QChewNHPrPTeWyaqQvyQloCm0NaiD3eA6lcK0L1fCjH/vfCGDe46u
B48H9Cx5a/rqc1YL9fcAcpoP5fhkKTZEkMe9Ak3V1Yh0gpXY9fSQYqjsDRwOhl7LDom34L4/VGzR
DLzrel8SzRk33K1JVXFHWh1IWEp1oLQoBdtF4VI34kNIYm7uvIlKOr2yzZ8clEyB6jQA++h/HZPt
ZE1r6jl4CaGrQy2OLqsOyHbSO3jXrPeBXWVg45A22HVmX/Kv5rXV9ViyfHX8ML1WuX2SkOi0Hxnn
Pgiv6SOFNwy7ypwcq7mPLQN6Zjp9mNKruU0EM9NhI880DnH735TbqjNFl1Y0HkBw1blJjD7SKmzN
T80ugXs5Ocj1NP1ylTNDQkm67Nw+xQ3SmvjgiVOE1g6pSHmKLZykheTos3kNzw7lk6ie6v56963+
g5HKTuJAEbU4+ExL9nIIsRlKJXH3ZkJhpBJmB8+NEXKPG8S8y2IEH8SyTSuZjfks26+XzTao0oIe
daYxFFNOx/2i4Tq1CBG3fYWAa55/0GkvcHPcg+cJrFLD3Z91pVZKX57Pd3a+c8FHZgNvYUncY9Og
4QWrqLqrbgfY0VyS2GD7e0SDCKATI2Jq7hINEirllguQ4Gaz48BZjHk4EU40l3bwixkjuYXhCaZc
42r9/+rFIGqdbjwyuV1HfYpZAkS9Aj7ps3jZ4fi1bSVZNTiWyhBu0WgqDbL1saIcy28WBEt8gpm5
iHmhyhoQzL17cMRTwSIWZqSrlVEpbn/uKT1CSVTiAxJ/3ARJ/RUXigOrtNzdWSJ937H1OAM29kho
w3OnN/lWZHolACOg2v5n0LfHHN3mJ9zWxEe7CIAYT82nyFnpN0JjCnhkszPC2lAesw8DABdu+l9l
EZ/y/IbIk7VJDq6jiV0V3JHI5+7IvGQhqnGj5QY4haybuXL4wWFwWBgDDyU75pFnAULivgTJZoaU
yqJUGRtbkULKCyAB/x/8/8i10HMdbnnjiY/8TOV/9ZMbTzdpgfY7nUX2BwxnokMJULOHcd5Xo6yR
MXe99uMcU64NGZ3xvUr7rLIprSvp5AgFBl0x7BFduBeGugILdCwca2x6yh6Y+IIzmC2IJ1QSckqq
8V04A7EbNeJsJfjHQHbB17dNPTL+ChHOv/PoZLFxh/fqOnxlJocV0N/+qkcpYmhZ0DEz3P8GsLxP
mAZiu2SyYQs4sRrM28PNFvCD084vTlOKlaiS3Sr1ZDZFhYOGamkiieA3geXE4LB9kkHO8n0qjTjk
uXrWOSCw8U4/0lLZu3ALSND4OT8qLklR4F5pdkNIKSQIdPZPJqDQHrAusgATU1O7U7QaKpe1QD9h
sPFONhKHHIw9Bt4nQNFtPg8PzX1sXrkXWHa1vht30J5YoqwAjfOnVL46Evtuzb4qkBYAHWATmhRP
dmr5IZIh+0TknN9aUPCGVkq+qPtsY1wlgvEdiVYGHwvV0HxJyHwjgOqRbR3zphW1o9UFRWPZ7Mwt
JkoBuysYbBLzOmxlK0UD0UPbO8FyzTEmDGSh87C4EXQeaBBDfTLLWZTxamZhr8hkD92P7isnAPnQ
KsbPZ/3Oo4dE3qtmYJpFDkAKgQF6dIuokrSJLUmCQEpQ0lDLtKP107xjA4daNhwwvABMBXbsD5wo
/UizjW5hUNigDMsn6t3DTSlSj07SME6cQbuZzdbiNN4FcPBLizqBKV2wS2+uFPqjFLXFwU8i+1G+
LnrIDs4xs5zHZhqkdpt8wIs62uHX9yJ4dX+1hI1QpVcsjZ2begxhgHfRu++Un1ohsiOKXoXtt3Vi
5UtUegsyBTnMhcwSgr+/+SF9b5mvE3caft6BIR58+bIxKsuZsH/4IWSo4xikynhqRfbtqrplfCLV
6HsFAYYhFVc7wJOwfGMDnIWZ9q9LPse0C0FY8aYUAM7s/vJhsyz5Ez+ji6z/1pizOV6h+PS/m74G
ZV7rE8svz3DZYR4rVy1s8E0ZistJSI+a4Lm//mW/H3BsI1VDffZWH4KQ+BnwwMQQHVjIdwSVrf4F
/NYY1ZqP7XMj7SUbZzdV6BpMjRSBvSZA8I/g8yXuVQncUxa8SlIFgyo0SHZnMEK8jHxFgQnrHy1J
YldqkNBQoIGuJYqTMa4Q1mBXTP72SJFjftEiUgEd/GM4psKTa74bB4fMbEwMrfbgLDfFrLxT4vom
xGwT9qWWr92MQ/AxCYVgFsXmH2zRWbUsqlKOJd8bHe+IYvxB2TMVKOcGz35zIrJeKighdYIcEbzk
fCFf5jesk4yRoagOkXsQGQbkbVQUVSd1MGXpGHuR2nCJitF8/Ubq4a2Tqo6xZW6adpl1rmdJJFOl
SatH+DRrvQwIaBJ2YUSL8+T7hGWwueEdwH5S7R3Y9Qlnjf/QgeBYX79tOEVx+W3Y3yOR9slskGjt
d80jtVAbT5pKknfnj+/9VwxnyhUu0yiF48Ghm7AcxnKYFhU2cNx71VdaW5CjbHsC2KFBqD+/zXNI
Q2cX+s882BueVoiZh4NRmd+IURf6ju9G41Cem2yE/eV28aI5idsfU+EEClCEZUYoh765c3iMvmN9
gJmg1elcxHCDfhZbE7zztUlh9a8aQW7PkQ8bsVGh6Y+MoeGtW5ua4V/grJ/rrJJy3r5l6KEKU1Rq
qMlfnbqoOt/+f1K3Rf0fp4AE2Q9/Zhja4q9kaWxkWES+wgqK2gJibMufmTUovIBHB2xOr7bBXcg2
dCSHwJGCoH4iEY0CROh0dl8fMQoocs5FCwQAltEUboFpCHHELhNrvL37uT+lWQjYAZ+DpVjsmQ2T
engVkbiZk+xVGTMGhvH10jqOkdpoixumIrDinjbEoQ+zQD28V4ZDHbYfp/4rO/0tEtg6PsPCdgws
xCKtl9JWvLaEUWfqHq7oghncwAHHHUXumYIHLCJIsc96cvXfyMyr94CZkjiG3Ma3m49MZcgYgz2R
+HUkdntVT4eBqgcw1r1DtsY/7TNK70j8ZZYmcXf4PyxJAGcqB/oQ40yyynmVrTo3HrQqVzgskPQo
IvGq7moPigtdxl+7xG1SspnVH7Y9zBPd4OZUUFF3t3/vwfj1k5LJovwkLOVhewtJ4vAE0RncTLEU
JtLCcif9971uRaETR/UFfcP2gjFjXbAYp1o4JwlUgSZmd4TNodAonTEKVcDIs5wLQxg8kVZdQlvr
o+SMFiuhMNug1eGiNC+XFK+1AIxZGIRuW9Gw1KJCcUPTcCEnJss7Yu++1xMMCO1/9g6WdjZoiAKr
koGWmxGeMuAiZZJi5X2sSUeSm3UBzyHAowAkk+3T72hj8/cYMutoG5VCsDM6HPAFbB+RaZY6V8N+
jthkOC/DCw2VSWrvD0DL1TT69NGLjGRjYWFzqPYEEUcKy98KTtWqJmJLjSN/xgFKTT3hk/ULdH8y
Zvbs7FOtrQVW7E/4/+JTcuDuGKDxcrFdSEILRV4jIUTfEua4U8/V7jzLeb6s0Kt/AqOcN2DdUeHs
WObiOErT8kuykaT1TA0YMJ7NUptInTd98+U+Q3BK0+gLpgvQ83TnQZucrAO6OjMPg5z1X3SNWhXt
QSKUIutPea7WhfmD8ShWFBcXBeOViSljtAEsc4BLyJDPJ+lsb/o7Lp7lNoC0UzwTQseyRQaG1tMV
eHazGG2aGe3bMmF0DYXY79nD4RBMxqTg6LzBqHGPjivuhZsK4dPPtAqHl+Kuw/dsrvamfF5lu0M7
hppKkvQROig/a0/1EHTD820R5YgRdjBTPcNyj4u/7+/9f94yJEghWzQKZ57ktwSHwpQVVJU+6LQv
//Qn9Widkjk1FlgOu1nF05XEARCDk7WhZbnqr9K51a3mJLNqYyjWz7gzSEMDij9q+w6RzoogBTFf
9uiA01dqC8iQT5uVPXDAAKwr8TAubSDI9WemLgAY6PqtE48TjMIY3QSvQLMDZDc2H0cV0lalS/xd
W6FO72AfrQpBfO+uaFBX4yoah8yN3yEjR1gls8ejsgFh94YK0bGDwIJK7f9dCUyDuQrJg7TosmpZ
FPvuZarltWINRgqyVuRWnLzKeAQG3W1eFIaE1ih6SA4Im84l4FB6lr2Wrh8yq4AxbomkBhsbmElv
yhAvjaKJ3AKaWyeZ3A+x67QJ4OKrLg6pMLQ98/fPUvGDVvu9q/d0dHdmL/PgtZTHkRiR3tMshoDc
8OU1mifw1jBwTgVVfbT3b+oRcjv8E1Ba3g/bPwJp5pmF6leEFQNu97IDdTaPH3/dREfhOCLyjS30
NtAmQJFMPjve4IZgMS+WgVUot22nDpKr0S/7be209cEIYg2cFiGDma3QUIgOUxd3DBVafX1dc56S
Y41KuNO4R3MlgJA5jslb2qFKflDUc7Agu2XtRKQoTvrh2nofYo5EB24y2bkQ4hq6VhD/w+Ry6c6E
VY0gclNwQDGum1vuRwCv7qvFpkgL2kvQrvI507f5yw/va7W3HiN6XPPacKw8+pvCu5M5MSMlBKXH
I/BCJfdkVZLhUXmAE9nzKxM8Hmpb+UwtmdAITIM2+xsMS40KIjsvoZcT1BLVBhWWMVTKzo5eaLt6
sck+/mQNvlS3V4FTOSR8IxmwXKDJ+s3KdwlZIvVYOSfDj7DibdNFwuV2NaAamO1wf6PZF1gOFMUr
gy5gMipszNUfpCwEinztOkJBZvYfrN7f7ZDl8NFihs5Vb+vLqngjw5hhHvEVI2gnGzQMx8JE8xtS
/1WwP3mEUwsz0ikYQKss5UuVB728xB3UuILCiZnNdC6LE37Xa3vBKrxHpYjaja2oVdTcKW2FhJVI
zZE9cIMJKXprQ8j5jF5fsaOnA2js5vWvyOgkHto622dbdlYQnpcS3zzBk/53/FV5XsLMrftFK15n
XYY24chcS9ppWeboQ4lnxpIkluRbIEYxdYFc7lay4gwVeoIAER4TnEdQXKHP/9iObtt5fJA4ky0B
Tb0/NOFXDpxX1ecqfqucVw+bxNihBx4SvEpqaCp/lvi/s9rbDM/XZeFbrVoru0sx4dAZe4YUbEnC
2RJL/6fxivHvtPDDpaYvEL3X8TYT3DMckUZmgJnPNcEJzX47JnHNvu0TM2CEc4GZyBvvy5xal0/O
I67Bc3J5gvShINmRnefSw/blfEFmgBVmqPmOhBS+8nQS/Sp1UZ4pW+cbyVEzBWEWUY1rA0LwtuhR
44E2zMjXVF6qLCFazqNRJcNV1wSrOUSyXiq1iASN/JbPLAzfd75kXSsEJwJU2KS0ZICNWRtep9yD
WauQXfKEjDxtM8xIh0KzcR3zLrLiEIVP0DojY3f+rQvOGmD1JpAp0JNt6X/rdKbBBL6/3ewW6geB
SnwG9ZU0zBMbQM9nMj8+sEg3pvRO2s/aujh0BX8emRwEcw0HK+bCQv/OXwnsGaURzW6FvjR6kc2a
J1t5hXvFM6kuS+wIfg8rCd3DC7ow4KT3zjhQN6urY/D+6wwDqGE4aiJJjtOeElglOY6MHgmwTcYj
YYbL+k8uHBfR0jACnH21ScvTUsnAtR1RbgI9g0xXKDnznr2pCwYprIqul0tvmk8gjy3tpFDjlgR9
QNd94YModDiYy4yqIQeSqnz/VHUE4LncEHSRzT6A3j/W05AsV6hAtNm7RPHLW9Fa/PEnj8g9epJd
jIEiJoYLVeIFSLNRNbVuoXQgMczgsUzUukCopljv0avkXkToX3HeaYhmyFariaTsWDNU4FYZZr2h
T59WVN0FcNXve7M6zOvqVVeeabBg9i2haIAGN6aClAtdG46KjYzrGIP65KT8Zw985IkClPLyj9Ps
Cb9T+P/8zd/ivAdnduX36C5imtlM+gn5Q9J7a09FcXqMCfGknmtf2jeOZxfoWJPLLHRsk4Mcq9T7
bP9HDnw32PHBFkW7FirdAFPLTZCFV3UMpA1QiPryP0+DK5gvxEpIzRhZ/V8aEqzvwXdv2TZX0KIl
BWc4sNPO5aWnlshGXnMBtdYbptD711IoCh4Wb+/6BVBqOmnE+J8NmV8hCHFdcRjtZboOI0rod9zG
6IAz3h+A7hbmUl8XzfZFYyB15f27E48hu/AUn5rT0EV0vXQ47pTHDVqLsSUVpy2lCTOpBqAQFvFB
BJ6FIXiL5OihiNNhWXpdF2eUIpw9/N+1q3fcFO6Fmyk8hF/oea1N3yOo5L3Va7ll8yPTcoFAyn6Q
ULvcjsAi8XRyREwcGg9FgCl48BGgCztVe1usvYy6anVZTtLNbux/UAi5hAULYHTn0FADfK5CtQH4
QCDhPgJAwZ7czk5anR5rpFIPOOYccXlmOfBuTf4wP8JkSOHKc7fwhz12uqnb7F4/IYYZ65rQ7KJ7
ZxH33TFc0tQet6gl2yKQ5zx0qLw9bzOD+hClXCIUCXAS1ljzf5GWNV1BgRMEwSE+p6GFzS/pkRuq
kGIQMjyz4T8ZNinjEi2AlmzRLdkUSZI7AqBkhiZfEiLrpsgq8G0+WOaSOMgPYE5ojAnbc8mi1aSG
S32Gjguh+EK6OAhbxgw/AJQlKKX1p3gEWA4+oPIWBvJzt2At2jgaIGABuzru4c34xA5m42iGcrMh
wolmLFlx2zzvK8fFiOt7zDdzPou32nSUjCi+801eBk0WSOLevffeLwp+7xbV2hqRzo+hkZ7hGO8f
3f+1h9loMsuRezPPG3OzCH4E+xeb4FQFdQvFBYJWNMc5EC5bsUZvHv/xxaKnODSUi9hV8bEvjlaD
wHbZD4/XtFB3ctnEaoNGw3llV0qz6FhNyjSZWn1Z5PCEIc8EyO7DRjc435BtuhueuSLKszYeLvbR
zAHk0PCYCJtjZE1cQthVuNaTjkxZtEz/+94gGtUfY8cNb7zMrGpVqaqiaU/i4x77pFg6Whf0X3GP
aFazXl6o9MdqqZfiAri4js2Ap+rmghc1TgWQtPmDNq1ZZnJsXuRnhfFe/03e8P88wKY6QmbkdMIT
XmPcH7lZTmi6R66AGDbEokxPyNo3dFJ93vkPFaatLazUw7exM1Qs/RZJvgXhat9foW+uObKmTtpm
imQk/1cAaV4W3ccMdPHrMdX74o/IBRmrJl1n/gSz3VKSU2QqyYpVgDCvpJfMp22ddXX3B2NoJGFe
1Zpg/Gz0gElUiLFfcIkL4NUnxlzF5uG4HKrOxSyW7GFp8LnhTIalKyOd2pOFromUZAIYEKLMr7qr
PAQM1yTX8Ly3aIiKBAmAdVKdl4V8Ivka+L9sG2wCmDum7uuaDZal47rhWIgE3wc5/H68JWeGLZ6i
rhGYbIs4UQ95TlVNcUxHksbsnlUOJ7ZNhjF1RZ1t0QQ2nxnJkK5i84ixWHA+pA4Evosx/bcw21DO
OkbJpmGv3Cr4gSIJdlGnisB6/aWrjo9IuOzRk9zDN20wIEAg+1/GSn/TY4WLI9U5FSfsJAcNbnEy
/5jai7bGBotgQMxS4wLDQh+C9yFlme7lKwZuFzt1rIUHBk/emXQo1PgZZVKzMzXW221W3g6AtxKD
fGAd8Ln4ZeAiERyn+cqOL/MsosrVHm3LipPoT8U5TihXkT6ZG3y0ZP8jKVQGInbOtd2PY6FLRw5Y
0U1ni0t4FOWXGKhAvMMYYOaE60J3LVNZUPSA8jcf5xAZFroGVVc9wq9bu6lfPolWN7afZg1jzEo7
U2YMKIFpOaiSNnAFiTkr24fuHMXKFrmhtwZCMA0H1xB7Y+7JpYXb2toWNZ2WJnq4D/30sCovDISo
aB2mPe6Zu8SK7DFvAjgng+zDmdl58DoeZzSOE3Atw4RWvgEbfC5MkelGmOHzktv/ar3RLqw4EvNs
xCWf1xqYJLs+MGG3QFKt3mAkiywH3DRZetZR+xrcmybeq5uWI7QvNVgdJrBui4VMVFuwZsvigl0U
bwYWNN50Jw52T/usgXz0ygZKSbyhDSrdnOFG40LJ6X6+Ktb+Zh9aHAIO+rdkjaPslGic/RNuTww1
mDTDWXFxT4vDdqLmni7CpEyHTV5iGwOqM7YnLb5Gk/+OWjU14Cn2wGR3+BPrL5F25oAr90g/QYEG
IEJxDwPiqVE9xs2IS/UaFDb9aGW86kYxCBa2LPgSySUdi4PyX9tcfNjgR6ye+7EBjtjStJ9FNU8Z
InRlP6hCo6fVG/OaPFCR1inXFu2csA9ex41iHPVEZThdOQB4oHapApRkaziXypPnN/V7gKsRLfYJ
3U+rlZHXYuvVxDdCIhf2YtAOosmQLfP1tcJnZ1+7LgIQKjEDKcFH5BHSv0sVaU1VI1t4tsStHDw7
iOMphmrc/8y9TEHKnSvZJWmGrm8gJSazMLVTkasE1YSIxGKS7vRq5CZJUe3/UAh+owJyXEuCpJQt
jUt0ha/sihfrNBaDUNnh8T0OoLfGNU7sJeV9iwcKT/FSIReHoeqJk/CM0BSt6PVKfa8sfFm51mVz
1XPved7UEkrDSrmfLUP/LppnaR4E/UzrC9bK4YxjRqNZrB1AtEwpGpi51w/eJ8iuObunnLz8vP8l
J6a+zfLyV3b8ge4TU1FDdEd7ZOYdG17zrXk7rP+XKsu8hgnDIFge2qP3za4jMg8Dqi/ZlC/CE13A
RIAZFuyBpW87xsQGr49NEIdR2bmqRFhfTDuIqNjCENKgz5DH1wEIc30787FVj3pGmSxiDjYxkAVK
QvkL7WVYtmX0ucw/kr98ITHxdP5C4V1liDaXbGIki/8ulC1/twgOIk8vetFr1TzIe5faY0x1UyuN
Y0SHCE9SEpzlZvMUlsM+Pw1z3OWvVWpra2a4r1WikLR3JVyI/hkSw2xo2dNurzT3SL1iT0SZAvqJ
8A3/QT0fqL6NfywdK2ULGw/uZ3o/ljS4O0INCrOJXU/X+ZAC7n5NoB8ysqO7AM5WsSCi5K+oMVnk
tFyVhZDp+mUoNmDoLvQOSQ0/QDduBRU9f02Cr2RCY+AizSK1B1HJ/V5p7TEWst3wNjJbmybD9t7Q
BkgTfrmR2UunDA65ZkmBS+Ie+8UMUdXKX2G3Uqe0aazneEaJ46OGG7HDw3ij5iQBfJHv/5AGaMXk
vOw/2bGFXDvPog4CJVAHFrri/EMYJvzXnrfJ01gr9o8TlGGPSN/SXIxwtnWcudlxzpBWcsa2wCN7
aGlCwh3bqHy0nn7N4ih/KqiWPAWKnbsGqrsgtvx8+IoK4x4v+lgx0Doon7Uk4T3nGT/VyAGplx2J
KLR6PYnpWBxRZdB9expYS4XsfF1oucAHLH/5Aka1dwswN5rnf1XR1qzKPYF+Sspj7ud0hyWoxc12
JDYyQxyN4jh2Xj7nqtj0vohK164mtMlMzDXjbRqpHakgI2dBI64AyDqZUEqMFQXlBCdFOxPqT2lR
dFM28lgkLLLSqwv/E6U6BJ8Xm4vSXjOO+qK0794gh3Dh/nvSh3mHdUkM++X5LOvPuIzbg0kZNwfN
XstlqBmV312qsZ1Px1b5cWqxs04XV2p9u2XDoFId/QSDAobXP7vC74vrZ6E1TIseuOCzKk90WK0y
p3o1KVuRppN3hKX/IlXtIUJDQYW6R5u04uCEqY+s0vN6FL0bUn6U0G0V320+28VRx531hajw3EcY
vfn5ZGoqceyFhgv62V5ssuR/Pa9PDevwOAyiw+iv//IkmShILNNktcnqvnhrhMOJpaMCMzP1USIh
T1rk/OJ2h9K4H1y3ceVWKHgOIx9jTA1pAhr3C3rnoWFezEDZD2GUsY4xPWlDqWTrX3Nk6bjRPDPf
11S0AdgimB1gwCfyJ4a10tOlWh3ZTMjw60P91aDs6ic/rGpQKBRw5m5xe1lVI30sI5Uv0Z2UnjHq
Bv1gr2C/gazm/9W3mvlz3uqga/snXXh1oANy9xWv7jQheYxrFP0yHKkbZvlulXSfY6U9Ksvw8JHY
BNe5DXdPqPTgKXb7X/rGejq5Z9mMtASYmqKE35iA/W5iTp5KCbHAcfv2+BXK26hE0FICks7+1yZT
vA5OWZFB42e1wnUexjocyZjEPP3STWOA7ktJlherQ5l3Se5/TU96o41h5hRDwsQxjkFJSf9f1sVh
Vlne3clatnrVh2VXIBwhyEnbKxuXSA85tDeiM8l4PYOVVy2ZhzRv/I88dj4YJ9RLJ2jJs9eSF+XQ
yBUAsay4ZVsgKTkV1bzaWRsvA9dq0BPZyDtUcC1GJ2Cn1Ld9xc9I2mcSJF4awUJAnB8FhbIvOlDj
1T3vM0XzPEj+68691uygaVkRAbf35CNhP4OzL8m4MF6qW3IP7jzKE545yJekmdroIi9nSgkAQ6e6
AtZsox3l902WxOO5/dYKYHY7pXX7SSsVz2WzB3zfkZy4qmeZyiyzOG/mQmsj/0pmlKQwyCw6BjAz
EKfbVMY48SoC2FXTDMp3opNCRfdxdgqcGW4XpIshgQZ7XGJBnmI0RwBLlYFb1/eySAtalR3PJimS
gq+9LiTPTM+gQA+dB6S55Mfw48jBBIHFJ9/DB2alMtKgNAJev2/H8mo+E0c1zwJFyyEZt7b2ZF8y
bbWiLF9wJd/0Vb6n+ua/QY46vxAX5tRjLaU06Edg4YYyd1wOrL08Y3ihDEfsA1E/SUI9DWaweJ33
YusoAns3fy3xha2moBewtoL6fCL+xEtkq7yENtmBsSYx3MRkzjnEmThlhf34+0jTqtl8gWeyJaK4
SqREYYeTQ5IoansQpZXWekRKzOC345GZt9/JqodWHgHOc9Mpm6MKgMlLncQsSpCQ6LvtR+gJKuCw
6K/KsPy3IpoOiegAYUS/uqxJND+fDwP4A+q0k6HffYUlrgLmEwtsd+OjFuoCJRPXwuRYTYt8/67E
pfRtF+tGvFRWuOIkY5AC2F4VBKOxy4wL2R9f6P5EYyUbFCn9grxzC7r6k5e2dY2REQ/7yvn/DCqT
JRQeAdosigzETbT1FaAp3ikYLAcN66trgWHRllkLBDxZ3cAXwQPveh3v3WDme8sJHQFyIxtPzIRi
EvSw5uszFhozfnVizGb9VkLipcnft01zctmAiCkp3DWtrPE0iXwt/mUAOgO6fQyTd3ps6x8K3A7O
RLMj40k8ayIAq9x13+WVxu/zHGK+zBnDQpTn+0FFzDeAGQS87kk2p6GUvT+06KdYW/Ie4plnHcoJ
m3FOOIdNPlhnX2RJKbwA/jrfJxF7Mjr+/HOPH53L7MiXt/HrNXpKqR/by1KRsB5HnoUdZkFccR5V
pIBVNJ1Zi8Hec4TcxwoyWrT3hJRk5GBinAHkBsbBz7lXqbgbVmaFbaismzLuZEwwJQcqc3hkOTwo
X4RM1QCY64tDJjWZEgBx3+AWAolL6Ac/RQu/5yiuC/DbdNMc+Lc6hD84VsRADFQbTUO7/TScEl0m
Aih1v2MTIxrhIrBjKDGtGkFLtuOfyiDfnWplpv+oVLTefji0mMIv4BjErssY40dO+0Jva7bk0HCE
SqYKRW0yvtUKz4ZTg4xmD1fxNmJ+2wRBivIY0rn0WEgIGkkfn56C5elLo5hTDZPRa4gSy6OdE8Vr
LCeLMvE12eKGobs1CZPZxYf9e3FqBN6ecCiFX6hZYI1we7beZ18aW5Q6j2cFg5e7pJkxEa2Q72nF
BZU/aHL2GkXD/oRChdma28NzGdIXTC/L/C9KnEF3SibJc+7BDM7qadoytfkkKPasJnwJNRz4ZpUS
O++SR6JoQZTPp3rP5VNgSsTU/KdEF3MyVLe9M5lRROjPBWQdbYmcWVgrqp/Qxo+jC/q6qcDLSVRt
2K1UzmBlPJVIy7C3CQIeVgJYpmepxsnDR0TmFefqMHj9JWi1J4l6t9tnLkk3UeeXgbfNpbyyIOv0
KKCIJuXoad4ix4ciks+DuhMh3SuQUhcpwAdKACV/PpwzlfYC4esBTDW6LSMlGMTfGKDyXjpnZH9w
ssy/qK2ltmAAQz7dWpwfhaY535Ek3o0ZQ5vx9+RvBPdO07i+slanbi0LJKXSEWAzUalKYh542X0W
3EjiOAP1PMCMI4mrdWecVOIXs+gza2P8ZF2WST83aK2U7owObF+C80KBT3KAIztGhHH+8cye6mfW
xfZprbfuZOxLd9x9/KLFsKUOLbuk7mPP2cbtZzugNE8rD7BmTIYyym/AKg5jstQHTRHzIZeMpW8C
jStpTbQ6JKTrryqkCDuYuNsB8wYamLdZ7pkRkInmR5r9p89O9IRlOe7lqWFA5+Zwpix4dYtLJO1T
eV+yXhP/4d+4dg5cXJOs4UFuyxT5+GukFoiJ0ce0W1+qCtqVuhCvpkq8QV42wEI0AbNxGSb/rx6D
zm2Qt1phnKrAZS5S+Dgmu/b/wB5j0q3a3P+FfL9rinrvXlZuwEt9uvHLl2TG8w2Dr/T97Mb8CWPr
/l0iVdPInIKgG3DXD8S8B74FRy9POw7gVv2gEME+EQ0B25hPz/w47Uzb1C6U5okR5ut+r+iVTkFa
UVaTAlMvDTTTSJipl8upFLHFobVceoSlZOldEORflFOTQ9IN/t2g0sVxMyWqSDUChuIGgYXjYprz
hx4QTu4Bcs7NwNe0kLLY7kBM1YQHO6WndsbikX1NiKxA8VtpOGkmafTbvaDfFMiCkGEntNR+LsZU
0aa5toJTvE7DCfWmDlqk7jNwhf+XXPoXntSCYbfPu022978/sy2Jdmbh9dSZvcroL7tMyqfNOnfg
CcJzH8WXP15Ze7EtzCv81KxKqxLTqwoTZecRb6LP2CrAwiX4S1q12O+UUYsfL+2/hkK0mwEsWadc
x7InxQnNsvnV+3aj3+84hblsgW4DUKyf32qwIVVRP8j0KvjqiePPBjlbCTYPDBNabdXAgRd7XpbP
298RnkQF/wyJ/oxnf+BHbENv6WRrcEFwGbak2iAVkyqTkIWK91OgncxO+2tRA6RzKWhON5xGSzyu
InX9fdqcsi1tZ1TsiwW5nKJvuYOHRezf4td7cBf13C3lZWhiFf024HFygF9vDmNVYhSjBfb4+dLI
hii3nofq0YpcaFa0iCKBrFTV5VYo6qOX6wnNUDD+2+liAUJ46e01LNIG9hLVuVLwF2JFf/t8IZW2
pNL2oGClve0NRCX84q4dYhKXG02XxbigKQsHyXLMYmduWczBB1VuFdp/qEsugK5/AziXWAUVTgD7
OJNySU0H/DYUo1FjKuhInAIGuZKXJ4M9SSjdLHwk/GfqQN7Cy76ca+Wxd/LrIg7XwRdQN0ieeqT5
3vhNt+dNpc00hfWksN03AhZVfi4CRNalqrU5QDAVO//AN81lIQ++nXRZrE1ILiJVsP7jx5LYMJeR
hqxXTYRkCPzmB/J+j2xrLYkrxBCxell9K6CGR++0bOXNPvP70DoBADXh84zllmGrmGI/osFD2UlF
5VdvsRwbsRSoV+QZj9rj/GbrZ5HgAXprjXMUpA+qJaYx0M+q7oPNcqz7A5dXlVNd8UREkOW8nFk5
nMKVjC3M2EW/8TH74obNO5Lc9IKJwMqnIBCKhoLn5GSC4QvG2F36coTgxAGZccwX4dWyBlVN2VdP
2M6Tblo7tAhkHz9NDiuTji65DpXnMt9jzOiN4iK0UT5/Stb6coG8zvGJOfLDPovdSSwo3eT0iHqH
ikTllFgoTsXoNDVguRf1iKSmldYpBRXqZ4tFnPVHimfoYn14I5pMR53hzFV7gyQmdVy1z/07z0V9
VxhMFnumE5sPhp66XTm3x2LAeXlp2qt4aLAy6fYyTsJIUQrCVBvGNBO3CRWNE8UXGsLtYP9oasTk
VFaE4vX8HW9UiCn9sM7DvyDfrLw7wjtqToFsoWsmdk44M1gpsXV+XLp/CxliAJQ03S7790rcpaP7
ME9u6EHRfqGXGSvId5Q09+TXe74fPJDRxkbKJLvlnKS+UmxHg1EBG0U2Zjsfeqbm7qtLT4FwF58g
BBO+PIFZnQSsodbZgvq2vNMpG5TBC2O+vTlCwdzPBCcPSXcCANQAsijErxrdgoy+vKkA5UKyURDw
6E1Sa4T7xpqvg8BDDxThyVfkwheqk7bu6i3UxwXbA4Q22XEPR/RMZo3oil+81gHG0vVTT4Z0lmCZ
oD4ITcjNN2Gpe6fjmUmFcG85zEpN8VRIbFSsjqmwL375TrJAbxYeSiotrrVL53u+vCGNmpLNxX0R
pFSUVzsIbKSDdTHVY/deSWyrgoWSEKDjpTPh3sLUwk05BVAeaYKZikTzFhJYDXZH+DVRpdlSCVak
H9wbWtpzMML2YTMsXQWmKOZKduj3mUVm6YzoeQmCJHHxWB55Sx5yAuRJIka6X9HVAWaN/J01C8Qp
UzMtwr4dnZfVJuWDOW23SutVhGgAV/w5x0DLlGYzs87mM9HuM3Xfd0W+o3xHHvwbhMpHZPBFw1CR
zzPUHLzYsSPB7fvA92t+1U6Cn8BHVSVQTVSYDjjcSLz/9KEt0s34oB1/UF95DumKtFzDzQc7m1ya
r4dbOMX2hAl708cUiSJpGZrf2xbVCkHWnZE1slFKdh6/DKL+79qEERCUF09FSVhOo1Pltm11/5fK
IJZVEo46svaV2u2EAfH71as1Y0zGAuhYzhd7xJevQ2pYJyN8LnAaHIsNXG8VWIgKT1JK9RArIPCj
+xI5EYxtBicovjNM4ryhzHn8Hy1zUPK/8mLVYFV1iHt8f4/XQKZLHiOzpCOj/igeZa2cj5fOwUA+
9QeT9JlDqN/kOTVI3eQFUiwkvRki0J9io40AuRkxw4xTc6RVpX53YducpmmAunEsBVryaLqiJe00
SG3D2tCUVvLdnMG8tFMMML7q1iLIf7V69AQADZBENwuEi59fbUEh574dXA4bk1I3vEEe1OndwEiY
/wDPFHrOxIpvmeFBVHvKoThPI9JPJOuFBUiTsfW/uSYUfGBdeuVAs+hKMFb9A4+EzyCsKbtF4d22
djLktaFGxsM6BsOu1tPXCKe9KfLi0iLddWAfvyiPIgREIjadvsLkOZOxsnuRaPsUvaXIb8EJX+RU
4zT2oksiDk/tXGUqAxmZ8trdgLjcCKLOgMbdhc7gdSkGW6BirSSMG/rIXNQmKT8Yut28Rm/fqUeM
yyQi01sekURF4k5JZ9mjyEWCFMq4JG6E4dfsbnKMGwteroTMLZJagEDEyWwqTWv53vlyiYzeDnt+
7V8cuSz28ivnuT1EUNoV+08WFyLF79TosW7J2q1Rm+T4NcWx5sDd6UXIGuW8ylsvpXBCoYEI/Gvx
g7YUGQg2kF/Rw/z1tNZFsqlIZQXiGtf55LeEQyHMAQ7QLCvvtj05WQR0GASOZQk9nHNbP/64A6d7
08G1UHePazGzRw5HRmW8goZCMUE/xbKNr7U0Uug5yX15L1gIHDke16b32yEaYAJqvn47dKadveab
aG/x3Uf/50VIwndr3VfAQUWjlaqZdTPTw+pBOBH5Hm0aKHp2O6RBYn884FxHwzdYtcnnr+9EBDUz
yvbNjledTprgsUT68s3JRhMZjZldgbTIpIXSbXzp8Aaqlv6KAE/xx8xKXPeC1TxbrPG5Uihez74z
N7eXnlJGBzzxMrdbYRQu0a0woGxAs6wRNouEGu0xFGgGrVmcnDF9jDyu/3JV2ClMk+0HEfiwyS9e
O2ZTmLLn5GYbX1ZLcAnqR2rozhrwN4kpEEHn9ZgXcoIr78k18TwZ/yqTyaPyBbi+dy/0Wv+oerc5
ZOjWDnP6fKJrgFFGL6T5JjrlIcqjbzPnGG8QrooFUwTikvucSrU0ejau3OtlM9g/HQA28HE9nceM
L7YJEbt2KCmiFbPJndYD2MDvTd9/7dZ6Twoq8h/7EeIxlkzelZwlGQRXu/lPJHHA/A/k+GiTgAMQ
0CCA19qe3ZrLv8afvF6CkfLi8SSJBVs9ysYPxPe6LD21rUo1HvfFj0ZPdui5ivq0ul/yLkTi/PCp
kCeSY0OJ/rQceNfNa/GevvuM8lIWcm4MRUyXtUQxXzcEvGLbjp5NcBur9lY4PDOMRy8dAkueknxt
2RdjyRwRYx5zmBgYUU3aCavEiTnqSNrLaqTSEY0ds1LtWhqof7TzG0ozlaa16e9+3UeBGCWwyB6p
MbU4E4/7xtUaH00S13W6Hk9U48/XzD73Ip941hClfOU/XslIPKG0Tg3Zm7DpbMiR5IUPgdOG7Pj6
Au55mtkkgxv6QiJOwI3DrQzQp1VJmnRpdUIspmUS9ZZowdkKsmMG6vUxv166+QJodqp5YsNGI9bK
MnN84UFTM1dsGsZW16zLn9biJ4aQYRw8cy6OaFnPFJYlxJ84/ldnm9Gd3c1kjVGF3gjXzMCkxw36
INSUCOsNXab884Wfh/Tq/Gr9zXiOOL7asbscm2r0r3zOHezlcl9cvXUgKJcASmFvsMRwIcDgw6Wi
yKa5oMI6dHS7HMghPeTMWVkG6i/U0CU6OuxNvl8m0+nlE8TmTv6dN0P4WhqQuRQXJbaWWRf/00EW
Bapds1O/60pwdJkVzMFMcmJDdXjZ49OiLM0e9jOBzKqlaxjyxt9E8n5BmFJvGuBGZVy9AYC2/T6j
1V6AE2guz+gs4sfJjzg/AmxALV+YfpE3ijJqhnO59pEFYF6tyjY3UJkyMWx+mqaetPOVxUFfXyMb
xfGUuxLb1sBFNXw3fmDUDgNk2wgv3Bujy/GvakGH8wVcFOYIx7W9yPy7FVRQr4OvHP+Snz//ciU2
ixRvBR+CtZlu17ZSnYgVxGEcxaj5L7qsUPFWOX8mJPmVKLDxwvwXAdWPwWklsXP9AmBQjmvdof6g
YeEU8kh0kP153j5gv1OclAOxhu/wx+3UDNdeaRCJogFEGZaVDfwEupXblZNJ1cBdq55iJrY1W7xt
i2wvAfz2+/LSKRw84Ndbt1w2WYOC0NUiW7HMXRU2XQRxcj081S+EIJ2hdwgxK1UDviQ9wSrpwl7l
qZK4GMxHnjWg3ANBIbNChUYgDS97FSanPhErq+14OMsfd/tM+PvOLaeLLTpXkWKhkoZJ2ezOq6/V
3LJnzBq+c54bCUSFrACqCDb18JrxAwHeCAtpfNd3oFGhdK4gUci+1JAG4aV01N4ZMURn7QD7Gcu9
MDEQJfJYAbQDeWIZ/zmBzifClRKSoGc1ystyzzE0dZ0WiUOEkYi9RSEb1f8v0sX0TywlzJGZjQQu
x+GVaKZHAs6iLChfqVg32r3msTqbwFwm1eHwnpMyWpurAD3+TeR+QzE1gz+qNfXtNvFHtdkfcsEl
sXdewEcPRFLKWdDlav9HxPM5uEdur/6avycUu9LpNmqD6/0H6mAzJpLCPc1tEgxBq0pSQRWBOWK8
6vZbFFcrwr8aKCx6JbQi7Ud/IfQzdyDO7Ox1Bc+9mNKpN4CQXDPHm1AG+4pzGFkYRRYjTvCOAik3
LGbT2qqdz6OLzrOktjW9W+l+qmmoJkes/WsfecnvrEZe82rNt0Rhyp5b7j5o6s811OOoN9PUlpgA
IkCHsMXZGYQcA/eGmL1nUBm+OnckGrZz1nYmZouaxLBRE9SfkwSZorlIx99py/XNyac+V2KUt6/1
FEKS3ma305RUv0dc1qxLmzN6O9Qgoem9SqSD0GnFJdZcBeHx8CKFjjILPuCoV6djubA7aqTWIyZh
Jm7XND+dV7a5XFQK/Z/oiTbA9OGKhjbifQSNkW8U9pDrw1ELskOD71bxjyb6q5XHbyvSfO1mSe5a
HE0gwTz5zAc0bTAfX6uRXrMxbZWPh28yI5CcZoX5V+e9kfna/JUelfDTEQ6nM6O7cNeMbERmNpGy
h675xmpYUB2qONbRB/GJ5g2qF2ppgnnAC7Fa/AY8O2cdtoOc7DbCSqM04H1aUhtcsyf0/20zmNJZ
2OSuYYCq//ur6KGrEOjDllh+sBvhfieU90GgqdOzSZy9ThTjUFIhEyR2ln8tHaa4WxeBrouhLaL/
2wDYUfcOVdU9hZWD+qHX2awUqkCF/rnd7b7xLYyem/lbW2YthamIquL9r4EeB5jsQb/Bs38DKcla
hv8RuX+RBrkp06EVfCeqbKLg2mGSNTZR1NZNkTlZQqdqIgSBVl77A3P4giZn0yyU3a7YcgTjziAs
o5B1JAAPFqDAZ6pl+g/G1M8pHDGaMp6/OIFXGN9VNgLlLVUfdlSOmYMh0yylaFJ0wsx9bz7/NKS1
SFFLDnBv1xrNLt6n32F1OROWDX2q8VnEiY4PIPFQM9h4eAGl4NFRCp5t2pp/m+foT9fIEco7R/fY
6+M7R2zcAfyGVh39OQGco2k8325hOouJ/73n4uQkm0rB9DO8Bf8iPTripR/VyOAapZ0wNZiGkJES
cR93EX9Q/LLuQ/qaDPo79SuF+dzmKaDSLzSxsjC24Xz/+WcbkhuqLqa3haObu5bYpqrfCDB9+X+U
bP3huEOoLykp9pX99Id6GNaoSMLTW+vqkEaSGi1/CCUm4IUD9UG1vDohFgdPc4qlXszb9utL3vi0
WikfAh87aEzYQGYWoVXFwA6J5HGXfymOACSG6LpJx0O28hYvtHDdamrs043dN8UwmTQVZ+KSYprl
AglCuc4FtkJYiRFk2qwZZg5LWlPvv4Si2zA20u+1UhD2h6bCaC4H93fhjrKPKltm6Zm0k5MVTGv7
0SCSYYerySFB5CZB8UZWsljUk+57c7xqVgHXwF90LfFI1PD9AYa0CZUl473F2GBnlDw7QQpwGWEJ
qZ8eAWJq4qAqNtXOF+XXowGZc5vbf4VEh0XHJ0aveG1MWYYsLuopoUOS+Zutf+tQeUl8CiHFMlFu
DAhfJUzXp45i98/09V3YEcF+RHp1BbzBZZKBWx06k/T2fCWWnHIV2Pl5IAHHNsWoUDHmg+rRgelE
VAeoJqwuhzV9fwNIqW/NtLY5nDJ2fsTiOXtFFmjBkwrcG6wPc9PcpCafJpy2P+IIOtyqLrZOojF/
YCdiQ7I8hpZpQjdx0Q4IlkaFp42HldbCGNLUZj9d5BZFCzseJ+dfCib4M7BVEZV/96f/egelQRXJ
tKlJI4FpZPv/ND5sorOLj0vnDmTCDCOnVcm9nXRiXe7mxINjJ2RJ14Sgq09ldsdkYJg+OdQaN1E3
vQIDO4i2OpMbxGHPU4rAm0sG17F6ga5j/m01j5motpK9rNMIa/VVCOdniPmlumYsXFLTap8KwTU3
Mot0DqQXV7zQrMQ9WHkxYFPdhZIGk4eIfTd16srzpKOeyqYAXImHgl19pQzXfHBb7kBlOS8BcyH+
Fa2ZHpNXUjIKqiVxyirg7feMMu8P4gsTCtzBIHHFvUiV5PzVDX6rEno1n3C9lBHLNG0LRreTClVK
SO7MyenShADyid1rvED4NMR2X2FQ98wE0bl7WEzWmV2TPYBt348mcHKyc7s3l3DMFGDK/F7/i7js
Rykh/Umo4DwgBct7186DDIJfz7tAgl2tOIPjnovwWDsSdmEJxgX3yGx51pgDnDkMbDv47HH6Hi4v
AjJjJFNy6pORZyg3VbXkV1L32/QyzdDJQ7ZbJI1TUEJ8Oi9Uk3udanYbsTOxf3EkSfYX/S84fHVn
zXja9h4d3MkIs7Xv39IAUMoX/RrTH34IRsknx4joLBADrstP4LKbhnudUrTUEUZF7CKZ6S6v8vZZ
9YG5yDMVZwS/Uc3mQXrji7MbnxW17SBmeQT/aj9C4P50QSGnNv61IuzOXIsshnZMbX1I89MrixWy
RVQUqVxvnt/+I55din/9cYI1vRDSI9NuMzOwtdoZyeNGqRwS3PPD1NnGONqUMi2kvU/2PEcUMn/q
ZwiTHxpW1ZMaLj6NLjeTGQCIpWuxJVmKut/jjU0eUWAxdtTv9uK8s8YiJrSfQikw9FpPHBw1h1vt
yR6EAOlhPHvw8BRwVEODNntiEd38CIXZnRC7AwV8tSqzADX2tSkrnMpbl/tUeaD1fYKSa70DFW4D
RQnUnzZyr2OlBTUCizIFFAHHdInoporaRUxklBUyeGAzTT4txhdqyQINVo/Klz5P67y8SE+2y8XH
kSfSOBgf0C5DbdyCmW+jJegSmZuBaH516EaG/K1aEyQCzE2cKXCyV/h7hafwUW7geZPkR7resygt
H35pcil+QyhNDdahBL4ri9VGdEZNpcj7hD+qJ3e7Bd5zqBXbLeVTZkXFVUd7rqbM5HWMpVmAHXW6
n0E9OOItqAG433mJ/yOTPyH4WVJz38QiEDHggpTgMGs/YQVzV/m4/K43l/fBkvUkcOqJ4z7s03SY
U8R8DOLFMj81lHHEAIZkoIxjHLG+Hj+ImdKumBsp2AFRPPc2BAm+nIEwMgjFahz7ww7INcMse0Rk
I2vErdgC4MY9+G4vmQNlV37LLF8CUkdqsu6KDyk6jng7rxzOcqC3RfwNyWHQHZODAh5tTco8YaNx
E3oaj+B+Ycdm4cos35qePcyOW0T174i5/VBT2VfgdFQHUKIK0jyDJqA1Z7bzi6p6ZknwwgAAx8W/
FNjBZaXvkjd3AFG7if7diJa0IIlzrdbURq2o/cLxNDLF+6WIclYv8W2OyhcIuO9kLDjTj84Vfuv6
z/Q/BZ6p4y16XZRDtQZV2mjF+J0DSvLxfoDau2o8ZfnNL4dbJe6pZLl3D4ddi/u76rsjsvEQAUbM
aQlrChcEuSKKNSCrRpBwYIFfzna21sgkwiSw+C0FwGRihHZM6zpLLJougBFrvVm9D721cN355UzD
L4Bs6ffMYJLUwm0h2M/F1yVO8gJWG4JzNUFvv5ePTo0FeF2Rkx+6fktSDply39ZmwnsI/sgHvSd7
EqqMZL0RJXLjkmrp+zdVMXaX5QDZ5yq0Yd0xclrGz4kEfNLo6Dg/bgPto6xkECSeiyW4bh1tUmbY
yQW+KvC2BHa4CBB+MkPvqtP+x9aVbXJH3O34S/hxGARensf9i0EOlGT+99Zfx2WRF9shlK3LyxlI
6QHLjcicpxJ/QHCAc2HWZtmjsPmajDA3RgjZZz8nuDLq2gxeYjbrIZegf0odDAIeZEvWMFygvMTX
W1AwV3JgOMtV6oNzLKbaOu3fCc3mwwekM7Ly8T/L1ZWNm4hlmA8Dv7kAsD4e/SK2HSl2FUobrGcw
qMlSuUrbyrPouphc+N9kt6tPrDUkI9feHRNcP8TvgtMTVNVdmQ0NEXOk6/gkRSeETce0D1BIFrh4
ZT+R+PMEuySxeKtqmmwyCK6ebgshaNbvvhhfL+krwEP1EhpWhAG8OHlC2bAz24xe4lMCkYuXo2iU
4pocfNCDe7icNI1VIqsTQsvJh2pnBLQWICTtBnqaKoYcGoWsC/18feSdp9xFBi7qgkFK6muFpKq4
DmUY7pKkpt2rgZEkX3f9bjNNHc7686yXYiZCwc0fGUjGC+SBqkbiX7CuNT3xOFhKtxvGgftQla+H
9141+opsgCEh/R1l584O0BGqmq0cVHsPGfVGY3pXht1WlRP/Vbcna1boqCGpEHiMhesC3lAsdfZh
rGoMbUL5nnmy+ofKCBr3B+qwzilXnVR8zifERQTPgzjpQFhNu+yzuHy0UpxSf3iytmHvCZbRGew3
khp7e8pHR7nUJWeak5Ek2cL0ydTKSb92Mz3KzIGQTgmkJYQvuKSI8NAV+bmewkFSGIchZn6Go0dm
fKrbaYZPhELY1leL2mkA9x6Zw07pFUGrRgkNNMrEsrTFteylRxmLr81lUjqCyZmF5gRF6OTLiO1P
E5C+O+hXohoE+cpi244Rp3p4baoi92nXFU7tF6SGupPCJkpB5SW/kJ7W3fN4P9k2PNfrniBaXc/U
Aa1z/WHZgGS6csnbp0lMrYVwpS+zKpG84U2TtnGwgUNAMAEQK9aMnFXIw1BKM2read5OKkcoZG6r
vR8tRhq/lAZkL9STx5u+QugIH20/gaguEBknuvXRGmO3ieu9Fq+fJTqw1fy01d5Sx/BPB0AjXG7m
cMnf2hS/j7Td4td0Se1qCY46ISE7Sr1pbZzp8xDY32elptLO1w5Nwk+uX1H3C2CDKtEUVG0qle9i
BVl7O32NCNB4MWd7I1DnEMdynuD+D1vaDtaI6qemIblS+NawXlgxiu3c20Hk66wnXjGfiAdRlD6T
wDbTT1s7hXCoNYC6m0ZSovbsdqSnU+uCPSnEM1M6zIYd5RnDpIbsYBC8wMIu6pknxxOhlBTV4Y9j
0wameVdcKJdTCK0V0lx0cWovte5ZHK+vvHZplHpOnv9mrDdWNsBcyJW7PofSJfEkTiW3nfHhnUr3
S7lfE26dCfj1VRUpdq5F1NIZgDT1dZHlrM9QYbMrJGVPNw3uQ7wWyYU84ExzGPlc8Qv3jjhI7Z9o
6y9+3iPKqyNxlCQsCtrhhzGIjjgWo3i9cBIlGSqsfjYw4cGuWJz113s53IuQC7Zaa+ZtJytou0If
Y62pbXXJDjgWv0krD9PImtlJrIayJ4XWkONRnJ8fHBBLqLCqqdTFJ1mzJ5xOw43VLnamzhfpEBMI
sqO1mYFBFzQDii5qgO/iszS+scdLolV7XEY3FjVKJW/e1q0j1HHn1KOjXHvEXckANVNkTuGX9TwB
+Tk0sZL9OXnYcAW2QKOH2xkLEDCVpx9ywohlO1ctunMS1aNtQj/LPYBiX85ibWUopjkNdu5cBeJ0
n8pZ5sx3QW9oO3I6LhY4gGXmudQYKx2yBHnsehyFiLHHmQ2d1iObp80cmrLA1nkgGOn/rjqEEg+0
3dHd+0qN36MG/Ilyx+79KKUBTsns0AVH2aQvznAwetoLf5EhYAg/au2Z+fS/pJmbwSKUmm4gRAWA
5c3qkpQJFUm4rbmU71gZaLejQLJpEh5cTb7iPvJoxWRPStRgG8hW1hySylxoCTOAeavwLoKipD0d
7Kvz1P6UfYvAySesWU0Sv7mB8wWoBWssAs5niBZIhNSkx1J58hEk+2RQWrRE/WqZdcnJzdQ75G0r
olOtY7RhuDKcySE1+ONrI2AXIIJlN1NZTfzwL7kjh/rx5U/50Npi92RTRKpzufI8jPtJuF3wmlUJ
TToT2bzhCMjyzU30R+id/dBgLpbIchPhRmOOqrci8hsl+g4ETI6yvDxYr/iGzeEa5mP/sffM42n2
xNWEdNci0T70R0o8SsetGzXEfIKeLwYkC3O9ngXOJzgg76t+r5qNXFyOc3pAJEAK3srIyeHNthdo
T4V1/Yq8mrxecq9ewGdFyXgncoq9xRLdfLY0PanWWr2/p264Gjj+qV8G6zK1OO2gfqkgJ2XuOTw3
r5W+6M9+bOoj4emxOTt4XMsm7sRYlspcNC9+Nq8+xeCCNjD4iO3UmMkNz6obQp6OKVKZA3WW2BTx
IRuoqERUqnNdrfhGALUa9e+06rP4gUYzfypFfD6jgLj5hzyeEEpk0o4WFizSIiEjKVSm8g8x0jDv
rxhDOz6mX7yNRX589PA8/SQolIpmubB/6yrhCuyPEFWI3iBgso6nCrS2UYFx9ZACTBhTug+hG2TD
w/WY7XVBwuheZzIZA2eCnD2PXe4LtZwKjeM9MZfFepCI7PoqQJBAiq6bRNyAivi3BNqMLS5hyxO9
ODdNGEDr+63HIxuz4fKUBgWjoDhfoQo9Py/6F7BaIbsdpm46FX5Di9DRyKhXkcfbnse6Cto10tmo
wbJr5JLRGZ6ScVj+WkaKlqhJewzpM9OermmABRtRMd/S3BD2HPMOG2XZOuTV6/brULgHhAPsBmMK
o2ngV2kc2fHWXbx72QrAtsf5UmVCE+LnLnuiviFqNMiyh/+rqzUqPLeEglsudIl1k1NajwzwVAwo
WUTa15lc6YkjMqNo34BDr9DApzWfxz/QddfyF2JwAQRGk7TdsUN4wNrV98qSb/W+Wfh8w4C7uyFe
VNe50GP/LS7xK6HbW4awxnjoec3OCebEqcAGP6TTEAiISzh7m6kMrWDT7qkjAUnibwfRUgn6tDiO
ICaCUoj4D9+TXm8k9qF17iBTFLQcdzEkeoy/6uRL9pirgOr7LAlRp+fiDdsLi6brV/bx7/k6FEmK
NUuFFI3k92jsuoRCQkHjpSvIjm3TVNBTAymOCqginDRw/H4o8tO/fNhjvNxblkExDvWl+0khhiDI
b4xpabEEwvDEFt/bbNr5Jod4IzMD7dzjYxiVuJDqGsibsrEyv/KtkKeFdmuky5xcWQP3J0DU3T2i
O+sFo7tK13sSn00Wi5vYyPktIeRJwIdQCUdKWB5js+EUe5X7fhBaStADckDJoz0MEromGGBlovlL
vL5vcaOrvq2SmMkLsq9SjXiXt1CvhYGi8HYSC+KX/mOjk96fkbReS60JPdD9PaHfrpqFuc2Vswws
1P+9RNrd+iNCawSNktVZSrTXpa6aTW0E5DqhfHpO1IPxLoSwiltrgYvdOdYYD8rXDCqXBbFiOtl0
F3RJSj0III4wC5kG0RjYNsRfuAY0bKY5sdooSHWrPfHcRDrAw1OvtgcCFHkSSEUR+9dEry8ktBj7
QzCa3knxGdyp7lmoh4Upvgv3P7HrCfAQ/m2UHUS4ZjmfNPCSJweWZfjw3n9SErdgi7jjhyqIjeT2
UwwJNFbOduAyl3FFyvQS5IUq3bnzpurCBvxJ4+QYyUZOPWMPmeNotrCg59p40+nUH4yAmbi1IddN
OWzeESNh4ZllnhF6E360eME3mUShXcBvNZ2rzNdnk68FghWJdOO/bk4+BCcdNZipleJESSShEgqi
jnRcq5JB7BCFfwI03+aWU7KwqGynuOuece6qWbddMRgTlfUdlwL8pvxgJ+eMhWE7YlGdrRgY6bXP
DQCAL5v6UktRnZscWvhgHcv+My6iEO5V9ZUqOb1J1FHp/7a1SIGd4v7qjcIB4hTST3Ip6/JlEmj9
ibzuIGBZNXI7x2+lg1psceXlMdE0/MeRWAZKh4joUX8mg6NuWWc6/feX3bfHk69kgsJU9d1Zpj0h
9cULWNV7Dpc69WK6ujsVZlu7k7WOW6YxdzMLIC4ZkScn/NofPnz4SQRflDda/xBVLtm7PoNUrVzG
n9QR/GZhy5oCcQd1tQgwYTXwv3SQIw65CShwR7VLoRlaOTXnCaPZ2XHDbRHI0HEXyMPFo9vzipV2
difADldkXq1XnxUTopYSHr57o/3RfcM9dcgTBwUvfhVCOEb+MzqnGevYaTXdlJY0ijVax4ExS2Ay
KvR3uJN+9VZWkGkuHkodp8H0DK0fJSHp4HkJBogeSuC5Ed0I33DIQi/zPApRvaT/r0sgt9TjuSTP
1+OuQLSzZqpemjvm5zWRtibXtFyhAjW66mPZE7KNNA9avKbVZNX10WE4BwP4CGINUqUMenkMuMvi
HdZQNd2Tj1Asa6phF0917wjB7r6vXi0BRsUoPWH2M5sw0SSp/3WwxIbtvSlRNQorV3OWr0QiN1v+
BVrTtauAAlOoECvQ/qoD9Q7U6IW2inQ7eMvjyKvwK4w5QMsknExW3hxupaTdCQVPC5xyW528kQHx
5f8bEnlnNNGTeHmUMQvGDNA8m3YouV2jGXqP+kKSBPK7BMAvlsKUxSysCO3+xvw+WP3mIoa2Q2Ib
CWS1/fttNnemwcQlBQpdbpH/hgQ4ATvvU4lQKsqH2+fnpJYPZMAjV3/sPmNZKTaPbnMywqvr1Q0l
pyo+4Qd6Duy00ELYybzK243vpdbMB8ITEDbWc2hxGnyV6lP6n0/ioT4fWSsFGxgm9n9uF2AbF9lw
MNKX7ha2MNj5AfzGnnrcJSDyVwTP6XmF+hci0RrdnHXPLeP5BtKnPOw2IrJuut2CUj0HmgXRaDwx
ftWrYOYBCV8GLoZT/CHbTARKNzhvB478igbynoKwX9c5VSyHag06VdJh1kwQs5vVOxdzkvvzHnhd
gBJUSGBhpxaC/OiUVX9BhWVnEXfBwOFG0vuM1N3Gof5XQii5ysFFoQE0NtRM/6vPUy+JxtyjJTgm
J1IYDHkNyrDVcngrJUc5nDCMk/a28919AjFUKyKrmQ+9JPpq4n/0XHrw6QUl9xqD72Nhn/nEATX/
pVHyoljK15+CpfoiKqEgVSy1TtqlP8HzMpaEokhCNke2L0rDMNnlrgTYPNMOzl/rAH8azHD6g+Qc
PLvAPaj2nCS/uNmNd9MV3+JkIWN2gS0ff2SRwDt4KMQFxcOifJSC5pwy4IttdpfWm8yNivK81zQe
cP23VjkX59PU4uqSJ0MFSVGrgQBoEljNNoP+1omNQNaLcBt8mcn728jhhG9klWmENmBHy5OrZ3ex
NII3HWmYQRHRJxBX/xAUK5Wd70JcASDejIG3E04AkdlKIVvI+4AIlvCsYjzUjthpNdO2qnPJHp8L
TgH+b6qGTCXI3hzfXb176zgoG2XTmu2sQfzrLovokClQQ1vd+/zwSHfo+KVOh4Pm5D+PvHkHlegb
jnrc7O8RheHx7PmgsU8pxYHJQliQpO9gZ8h01ln7XVgjD8SxpdeIBqrIWcbxPkdea4nkb04VklgF
x86M+4xkrMnBivepPJnuhxaawykNT7NGV4/GFIh2c+WzhZMqQGlgPkg/RgfqgO0CsD7kwFbgxbhO
tH/g58RbCGKRYk6oclp9OYpys5YubGiZE8KwBV0oxkZHeFzHhFgq0ewkQWgnAEobnX0ZA5nRpQ/g
kzvBrw0QZxPLUePmuhkapaWCn37NR8tXZo7xIIWQxk8TKBdk/D32XD1/ifupiCEVC4Wo7r0HzvVo
dDTTQoVgQT7kXt3jB4YJjWES9nF6UmBHsuZhBqLh/d6RHWJwmQusaOxdnDAU9yctKRFtWTCG0uWS
MCEvvD4dplyNYGmAWm9N3iVBA8Y5zs5BpCWDHX6Dxpkv7yX3qSUb+W/6dWRyMASf0BS5K93YTsP7
NOHGnwUlTIzJWEihhMFgw/jbPO4TTDYyNWac2imMZRi51v7Y3J7uEEKahEklmXUJl2pytFDkSw0y
TT3tvOpMvnkuuBrs6qwgu6iqHVUA8GB+5N13qBCAWM9KkwH0IBWFQEXNrn5NNLngzSAyHZ0VWAgF
39fa5mNWoP7DaMeG5GUzRlUwpVxEMshXCe2PCFhzvj6dkY81R2SX2FvTpgkQ2nfg05/Yq89Qlgz1
ocJ3KfqGx0Id3tEeDLH3NVFLZL2ZX6f4/OrHN2dRIWthb1dcSeZMXYpJsaTjjBTNI653JAZT+BrI
vv/A/aXsN+kSMtP+t3JrLo90fN1jesXSm8c8L7vNG4ZYl+VfyIcbjYz9SiOOH9Rx+/OFqYaJ2iVM
ZLpu2SHzMJPMYOgWg/ZgEhqAoZcxlFmSeQZz2PxIuoLf7RJPrG4g2O87+GNfx6+5TKf32iVFp/Tb
Uh1aBBXHtQ82XkPeSZaLTJbP2cuLmv8kUNj2ia8aoMryRuxCeYGMBSMVwXPgw6W1Qsr8/cAujUVy
WbrmVNQxKLqMRgO7vo9ZM84LGfsy5KGQ5QrKzvY2gzSFkDBTvrms0dkotfvTlFbvC4G401oghFGX
YZNPKNBx3Q0sW7D7e0BaSX++uO2MWTgyF+zcVazeBbjih6PiKdMHCl+rfab5Qi7lAyBZnA5qZuaT
BHyO4jFAioUEkqIZfnl1j+kpS22J6rSmDVW0xFRXH1GZJ09uh/2RNcMrIHvt7ro53ge+Enx0rYmh
GMrP7gopMTyYfHjPz/o2eizgkB0Qzg6omNKOQIgy4Ul76bWn9MtZOtwSyvqVI1NeUDyRDgRA9uOJ
CzRy2zQI4/5UjD4EhFeUvsYNo/PQnJcc2W83RKYWh7gTReMZjQBBiBEWOzJqbOsVyWHuziZyvuD/
D16I+S5g5sUT9g0cnyOobo6bkIeLangOlWkmRNvngEvvj7wgr7llmPjhp/Cu0zhIle4Lvs4VLwkF
cbOhHmIuY79sLboApVYnijy5yu+C7sECnbDGe0IYHwWXb/qfbPymLA/ImU26asD8kEUA7bVjPG+S
Lqll1TdTt/lUftdPIVYmCeWS6/DWi/F6YHAGI7eIfSsy+3FsdjgopK574NZb8G6sEStwg3MRq91L
lHKIN3xV71T649rEROouuVcm73meij4c0w3FkLph9EZuDv3nEqK9Iev7eTy2YNgAxLO0TtFMnPcB
LtH7sfGXCBuoezJhNhRMqbZVcq4q/FdzBK3hXNBWQ1TRyxzI3qGpSMB+myEx6eEhWEZ9Hm6DT8JK
NQ+ps5Jo5V1OVGG4vbLU7F/bvmrFbJMBWWjrfDEJpM89prSmGvrwN/3Omb5MQxQNt9k9ird6BzCM
qGhQwpgq66pVPutKdVdymMeazXmQ5obUaJeHFrxjKSLa+OrB967vRpSg42IMIZDDvEYayR/nbu9w
UyqY40dpK0r1bJF8CDUH7ZONosgrpJ+GBwyaLW4p1Ttl6SfcBtzxKtxMpks/OiAXo/k7dQEUpkQH
hac9y99XmZo30+cbuIJn7nZcKiH9IroJwZe5MaOHbwhcA2tgJCCpRP69uNSsR4lBVUxL0L79t0AD
TQa3xBXAwQfZVgmkdS+82jnKYdMk/1II9Hcyz6njNZHbCSdwHKawB+NykOtbnub/bmFMwiO73msY
CF641oy7SMMXi7omDJ6mpbbL9pok+I3XCMWsQfJmy9E8IPE+0D9+oY2rfsVUCQBRVWlJHmFAJLLQ
d9xLx+zEVzj28Pofriip9lQsw5+don2vJJ/rJbbL1Bo3fLJN+3toJo9/Yd60RrOFkXkDA1CUERNU
xe+lCLrczj4tJuAN39vN2J44O13ppOzWIyxSmpPx5qX1G79QLan+MryD1OqoYdfUrs1a5Zc8zg1K
QaDrH/nsnUtOKaM4ZdvZu8GCzfzJiY54GuOXmubFRPc69dE8ZUBAvvnje5vq8JapBoj7tIKPSOVf
h+MbxkmJl5ahNdKCFGqnTSIId+vKiaKfqi0XnYf7RmKchqFMRGVpB6xQVJKXJap+WnRG1OQnfZPZ
YpDYNRJNYUCVUm42uMoqQi/a8n0d5pAlEZY1qG248opnja5r1nDeCbuZaK610oKrQ0DZ1JrCJwl3
Df+Z5aqlxe6KDakQFCHNZQEUBJB9CEXULjvwDHmbo9cTHT/N5Z4LnCQrxzMTRWQ3Vhc/7H3xLBed
C+db7sirXEl7RIF/kXeM+G6flFv6/6kxa7IGD2aQpZPTkOt39nbNO9wxUECtnJhVqLTo0LnZKmqp
qioN3pX35APqRbYnEJWAqKti1NzX33sjzfcR057DuOtjmGdoiDML+h22OSrsgGk1xApslOlY4K8a
OggHbL+MpAr7RGrY845n1dQw7CqM0AqYF5XkJxuj28n88f9UN8TuT0hcNsmyi0/YoYA8cMvvLFmD
u8AhFawy4pxqGUev4YNySRdln7Bns5DQrx3XgJVB16ZbdiO3BSQdIF/oQY/wRWl+Jpg6AG91/Jy4
e67mLAmpqHCczzporVhNOtxqDscmKWOJJMdfC5FQV5f5wHibmoFidz7B/z0bdDloQgDOELzUnHeW
7Eiy5UgDGvhCsoJvm62tdhfJdTdQxhTZZBB+RAN45uQOmlZKKXeNA5P0ixagRCc517VJLabEimqy
Gvr/GxQ/+WVQg40Y5XlUdzgpB2UNpaiZRAUyMs1HDezsATSj6vlFhHxcECc97lbMWXKeKf0dt38h
bqSZRlrHhBfTRQaB22gfME0E3QhtreCVuq0H/yQWZY94FEF1NpHpayoDR+eFnQZhUzdERhqlCgGU
MqOUZ9TgiBjf/vOxSk4I3sAWkIKtI7tZnl6oAdpVjGgD94Di5Bksmi43gUGcpaKMGFGQBVpqk/Jq
J66YAKRWS99zDzloM4b4u1veJ2IUycPhAHnfFaMj8xkxNCrSxNJDCGcdgGzFBHWEqMuPrP2lW5FN
ZVQ6cQd/G/5ml7yS0rruESMzFFjmIN4KwA9Zx1+Iw+HpE+d5O1pO0avMCny9Y+3X+gtn2DNv0xQs
UXoc8kP185oUT2pYQHQoiGfnyTlYeJ+x9k3YxXQX6hxoUb7UEqp7DOeXQEhLNFHG/R5pvzSngB38
indrAuIw+9hgVy8ucHKwWilUG7fDwKT5gbmVIoIIqJyNzBfdHknzCAFYZSTA6MpIM3yCgGw7WHsv
jRULcOyFqWiOqjrk7pvFYyxPfFmcW7Eo1HWmmWTPQqYqVOKf9HB87HuCaD1f/nVKTvGb5uTQdWod
+LwVoXF5Omao+yfp/nSHlozaOZy3b9OiasjCkaa3gnX0wpNoVEQBPQCjcVEC+LTIks33xzexrqCa
/uS8+gzMSg/QYDwptIOGbHQdeZNaGTzCiuk1YkmBoLDq1qXOYBjMftvAA4jbo8c628n45tufINt+
TuT9BC6fIAYyxjUqs1pNDKBYfBWUCMPHiqreWjZa0zUFDAG/lvrvzo0+zVI8nkLZGzCWxhDDuuwI
KWJGKExj+u2JISKZWMROwGNMr30o0WTf6UKQyOMKpS3v320YrRRtGFAwsPuq0jGA2BEEmMvyL2eE
4fE4zPQ7rFhVCL6qviDj8M5Drp1Xicq8ZZ++eOIbvjgue0eksPTKaJHawVtzLKlsNQPLKUivSP2S
CnPx054zR1GrIvTdbRV3/eqLqO2U5yUBsdWAB8kOL+nLTe9406sruWBVz56qfCBdHBT71OsUYr+6
UJ/AL7tr6K2KTAn0d5aFRjGoriYUeBRDxMiTG16FQ2BVNvys8cNj8ayoNLanuYChgfZtaTX5QkSW
0a3Am+H3BpbKMFpZdDa7esHwr06QpQIfOIeE9thLYRBYAb2qn9BCG0wFg6voM7N8IH8DOfBdpsNr
070gE3Y1d++1WdShooLiREeefSrmpP5L0t19Qhb5Gji6OnrjcobL7AXUobx0bNRFrRiZ29Ajg+ps
LC7nPLxMH1sCFSvejjnvGBDKINFpUMhhvUkintGdJWtseNyqxjDOIAg0j+LUFRZfTOgHFhgyuHVc
UgB0lorWa0L79YNJx0utXGxJV9a4HrVikaCVYxY0v6YhTej5qqkcH4dDJzFs7V6TKUvdv+xv2gXR
n3nvbI5wQ/Gl/K4XTgumX7GeH5tzrTC5m2aP3AGia7WDp/hCWJ1DW2/Crcbdb0fbUcgFBWdKonBK
lqiDOOJIlML/AboRbyfMCIWbKjdAAzKoxWDfKF8LKsXYRG/DvpplZOcPNxZQ3fK2YRmzlguxWmBY
NZKohz+duZSLed59hlw3yDZO/3cIqsTbo3SidDbUjvSynwr5uTSbhMx+LGEl17FBWwWjcwKmNo57
72kzv5twYI0Y32hoLyIkrgNHGPlWoNKky1y/xTOxSjKZ5GOO1XwUMJQIWSJKuXiIK3UsXpsNbOdr
MGxXTEcRBfwwGhrtMfUbdJ0O22F6uU+FuzZorrfDPtprvYQREz0WmLJSdMVrMMVS/Jo4JKLkcqIJ
TwZvkZ9NWVpiX0i+1LA+lqao9qx/f1e0j8F3i5bHQWaelgFy2BHQkbcfSpL1SolPz6N6ILkjMlb1
87jfy/EKvhghSTjOzimniZODK9BL3ZBmkoGVR/yXLKX2x1+JCrrJ3uiUOtWoMLbi7wD2skv+VUTG
xYngGeJjInDBgwrFKcsxsihxxMI5OeSCkmCMfpPJ05i8LdxwGlGHtagjZJ8iwsUyXVvPH+QBC/8C
76bbFdq/e9+eKZYXE1BKAt7gO1BigqVioNY+sRzVVS9MX/5ke4x6AMfeGUmNWisxfCsPbKRGP/K9
QsSH6CEvV2G0+qlYYMZUJxke/Ci9TQDXEOJtFB40l2EcsSYKbUY106Uik67eQhYJzpwezaMcTQFD
3w8rfkL5Pm2iE6Rm6XV0jOdO//ckpHcm+YfDlj2nLQ8a044rb4qAKbNyZJ6aogd5+uVNjxU1vBcE
FvxLFq4EIwxrNj9DJUWQnBrsUZ6TDF8+QpjWegKUot5DhxpkkDao2eL0BXmRJhCR9XJHO9Dwr5ZH
AiU2+xCPj7JGeMAl6h8ltkDJZ9qm0oUJMlfJhwC491mlKAPPvbEr6y/DoXemBSqLmD2D8jPeIYEn
9oof/q+Aawg8+Ac4L+NQpNczqY50EWSJmHP1WsnE3VmBosHYx66YLoVN71MvekO4hypiw2SBWyMN
OLjKE3npYM6RdTZxhXF3yw6ioCKM63prsAz/Fr1LOw1pjq/toNldxWXDYAsx8meZ47Ygo9/u6ivW
uyD1ZWWNCS56ny850BSOII7gBEqVacHB7+fVew6ijb4W4eKyByG+fEJlY+aOTVx0v7CRM3cKf4IN
zz5ASeiXrDJCuKM77bUgy2D1kO+9sQcpBfjEGafZdjlmMZyXlyEInl8r9idO50wrOHca333HbjJ5
HTPfrV37hTapjNkuycWBjA2e91A/Yb0Bz6QZIy+5ulCXyPM1KVaWNJvvPxphB2jhFSbz1UFzuVTf
U32H8DM8F+a5hiExWHytZq7On1dP+jYQ0LHiwNTlS82w/20xhuw+f85TKCDxxYP2DGFSjTRCEVwZ
f7IMVhNI9yHwgUOnX1X/L29ZLw4CuPmTWVRR93wUc8mtuTTaDBGx4wVeTgAemuvaCaTbJKTxhH/X
CtKZmvcob+GfRQWNURwFU57hd4lT1uehNLlIAQ1tekaVWC0q82HazSUvrx1NzZ87wwE+eg8IwT1b
6xzq/CIs9mjBJZLPu4DdmUgpDb2kVrdtG7ibsddOp6JGp5Oh0fzP+9+wcHqszeEqubLwptk1hiAf
iEoznb1W1EzwDqTbFViWtQhw1CvzuAXavWKBpJE0cPRW2+RJp3fi4+2B6tyjW8nnNdBax0TIlkeJ
1+NuBDhHw3VNzrZdGQIeOlarrOw+QLY0X2/lZtFs7E8bP933DoJ/t8m0pAheHeZLFU2sMtUadOfy
WLSEtsG7FO3+v0eisDSMZNCZB1JseyEmpP3GdUSqjOsrMPNqW8D8QdxlmQm7lo3T/s6r9U8hPFkf
J6mmAQRYXTl6hQV9hflSPxzpEfqDM/NCY5i6Ut6+UmpTEbQSptZoIUtzj3cF+jnlSpz4JxNMtW9V
T/BeoRS4dGge25jaq5FdUbrv+MEvVGpFoVmWtgLNEWDLnFoKHZWWEyD3QW2GOlsKVScp/dATe4+Z
q29or6+u6uvj9KwSUkMhlBFkiH8CkNvTM/hOG5tHdn1YIveojVlgl64eX+1FDfFSB/bh5w8DzFcx
1z/x9vFwqMcZo99mCXFhUGJ5Iu4mG7utvpmJkAIPbLuoCr40N7HGiVpJ/eKICW4Vj9RKmEv8w/9J
hJ6lEUnVFfByeLmHbh92I6w8YYYYOSUlfH6Hv+THDMkYzBeYjxxNmIj4AIwCO7dUmXzIDa9U+Ykq
FM0ne80pSqEYuNO1IN2T/bwldD0S4sRrk5tj+kEi/4KQ7PPm45utRibjIM3DkL4Fw2CQcUgtTCyn
R2dh3K0z1f8fl/cM34t5Rg+hcPTxJR/S6PYTc491yDuyf1QXV5+FXz77qJ0j4BKL5N9LpO/4V03Q
Ryzazm2vyDQCsQTCyHnhddwhvYOt/qj4wo7Ydi+oum6sjmBv12HD/5vEDWzHtSu0Ax6hJ55EOhTJ
6iZuMmDiv9EoqgIhSp9o3lRCSzSvtY3OzWpIu2kx4GSnDOqxeCTAanQKZMrjUip4VvW/SIlkt+vB
ZQ6jUa7mtwzjyU7gGFAKLulTVhobUExmrw8tdIG9TYUQZlpkKiuIb9sZZu4P/vESi6xaqHtT2n+W
iNSeGzOR0NDO6t9lUTv3F2jJJlOgwPgDzRq3ZSidEqxvpPnLJZdJ6cSg1/uk33lsSJWiVe5PKLzQ
fsINonB/uTZloPbFzU92EU4Ywt5UOWe+/3HNKqFJIdixZRIGZDTDUlGJyY3dY9WsjvquJ8/ZiUZ2
09JaA7FGeafG+212AhX0OnpFXZ+LaXTmOF56uOcqSkH5K/EQqP08yKrwuL6eSFdFEWykQx4ucPVu
ZJORlAqBT1D1go+xCo8kiTbwA6JhtC2HS3+y/qEs5WcrevzLB5R5mntw/IhHl0eCNUbyYqCnbpN/
s1dPkYM/pXyLFJx3yCr7ahb0mzRfSJ0OsnNOjuTQPnW5HiCj5M07qdJrnGMaFgPzE1Mp0U/pziMw
hmbQ9MmAC8IJAaggZ8PrfyiAvSbqR46r/PjQ7MKtor4j1BLFWtBEJ5dA2DLyWDsn0sW3Oo3JXF/3
cwGzn5DdPWr3HkZqgeM4sUA8crP90hqG4dJ3LMeYusqpUQKp8k47oPqRBZUWLfTs1zPgjgJusDSv
UavXhrozI4zfNY8NJ0fFhY/x8kusFPREjI80Ui+10P6mT3KCzwlO9ZQgaobf54BPg/d/jD9hdwn0
sRdnNCrRLiI3kwGctqvSTf5uxGNdQ+JxvMHcjWQHCZe+hytzTfl15IJt53iO/v8iShS4SW3Q9umr
xe/koUmBbI7h+cMgPMU0NvmBfXjgTrGCCvXlA6F3BcwwL6u0AMgV2TNt0mn5f06IyDNWyEkdwR+o
4Edi7hVDRGTDYpoNlP4B9uftHoy7RvTZgHmMjoYeI259ndXiuDCLUXdQ3oHFWNL3U0Pn6J7DZzNW
KZrEhDTK0xCYlg33sljqawSg2KXGI441M90NT9ofNOoHiEkQPJiqgp1msWvyTNPnM0t4Ik/aLNUQ
YWqK8PzaqCWTBKRd/2LRCHBVIR8DbkJLagWuOpIncG2fXaH/pKEZTgEpUX9KbpybnLFo9B9SOYqN
TQ/+9z0MoApqV0Nm/nsMC84UDZDATnAcJtppwJquRsoar8JqVh37RAnQuwvJNq0JwkvPYbUvmv0K
KQL45HZMlN3Sr2/MdwJftMLodq6PKDQCPbbIbunoq4KkuZgYw/giOehcDkoCtr6RFelT+LUfQb4J
2FfHCwa/Hgo10qYa/07uxkMO9gw+BZXUOtLNHIStCl+KhPm7ofv9T9VcmRtSXNPVqIPFkSdKxgtS
UD8jT/7gGRNQa1ar+rdvEUD4LaOuEa+1sdUtZHq/ipux4PC3jXYvXQ+CJgvVcB3RBC3av00/TK8l
NZ/pzWnpyzJYs/MiVHK5KYEC1yM3zauXramJM79dm4meeFAJ62Dg14QxnAYNM4KsQI3wMwwSm9+v
vqjyEhmlfq8ll+jC3LUpk2FLkODZbDTms1P5nDlyF4JGKVlD94l89tVHXtjhQ+w/O7gjEx87RkPi
Qsulm52QT5dLTQm/XEqGEXIUauk059nT2hUkImcVoEadN4hr8AA8eY8K4FuFoS3UE1sCgrASXEpX
mp/oxx5WcelASCCGi6CZPIQ9Xsa4cFNmSI11EJ4Rcl3i032pfaA9DJoc6pSaDHu1Hxg9vWTqiGHd
X1oGYHnpQjpqDDNfzh6JWCOE6mHEWi99u0Si5uhPx89yYhS4POUDQiNQ7gIO2mw1yMnOAHiDi88r
3HROgyyb3CpIbh6bVa/eOyVoRy7yrf9pm7UlVeVpUYrXBEZpyFPb4ONbr9M2d92GbAF0pgvisp1h
U/IZ27j8xPv887Z0KQjIZqOJXBbjLTHzy0VM1wMYsTMSGT+fSjG6cvPiHzQItW2Zrtxj5mMzdmI2
MqkH4/LH20yYI7rcjYp/1MXnqW4/8HJgFVcIDRyvUVHZj8Yw2fgX2a3u08o08La3a6J7syYN9nH1
KKDW+o68Eg4vH7nnf/8n662lEkwBOSIhy8F9mM21OOejq2uC9wd/g+dKpRKA3kPo9G9QW1JfE2LT
F4dKjb+lxwHvTy4NT6sRcjiQI6yj5/XlCboWbv20GBrc9XARfVt7AHJr3iQZvEse7SXztfft05cF
kgG3QClCNzFeqTdTRaGCsqZ6YJSNCcTeLFuzVSRxCnCteRUbbjpSapRL8Ll9Z3wBottQ+HtI8a7I
C2Vn7IHpCT4Q7IsZT/Gf/AMIL3BL154VBQ65sCNF13v7uhkNasp0CeWOa4c7FL6Zb8ZkohAVvjzI
2bpYaGkihecRN1vK0w7ZLmgt2dduoWFoEw7TnRcvbNQqjpGNEDWbci9LvQTZlAwdAg6FjwPh1NqA
PrIitwdNWRfNs+INTgJ3b1Ta+rtusZazwmi2Lq1lzhzsDXPibMnyXWIpkluqWg++yCaWFps7yYyC
MOfu8wxjWgNiH5OkRhSLEfeReL5nTR/d85NRFL0JL119sr5b+J84DFdT6L7RTWVZ50dLBhaphV/E
tmAzNi0+KSi+/5YAMd1I28jSB4g2kM6IUPetTwx4NvdmNid+30m1IvU788DNhNzZYcq1t4r831H8
ue+hJlMHscT3o2NbX5bvzib8yvM+fMasLxnPJJgYJNskusoc/hJ687MaZdAh+SmJ/JceDk6hkfQ/
N7eLMLtnqqo+jnm7ZmXwwU5m2mWD49uCwWYuE6YVz6xIhtbVhAKhmt/LEiFJR1MzsHb0OWVwYGFB
JGC0Z0E8YoBJox/A7nTIulrm8ZXhCFv0LxQXpaBA6r+aioNQAVqswf8MFNewV/htHsRijT0syMll
QH+pDS5PLdJqsir4J6vZeXHZjZ2cPxgUXe/oOzs2mu+Vg4rZQGV5vkRKut/b9kQLcRTjDVMCBAX4
GjtBfguCdxP2msYpdM+FAxUlBa70PeL2/zyQOUPfhkOL+G/qPFEQvbTvfs8gjJIjdaaPUfojq65H
y/Tskh2xO2a1ByhjW0s0ry7d8Fopt2ub+GKoj1K2Bq4d4KwTYgti2Y9XGA5n/Cy6pxeFp8pe3htq
rPhWEzBy50QaUnYKTDJAsZW7RG/zCkNog1SHlO6iiVSyo98GuwF1DrAt9KFYx2a2gshaYuq5i4GK
Kroh9JyIw9AzLngEEu01VyU7XE72XYSP45ZCPDvYN1ZBT/LDY0kTkfxOC4bUy3+ZtHxJGPKJ9C3N
Kmwx5/ZgRwVyliZlrvDa0gJrmwzEYOPq3UevBKx3DGH+ThQTeULU9zS3LYWyHJX4dAKdUFnu3Wrm
5Ex7kT4Q2BkAt0ae1Z9MHptzpN0ICiLhZ4Ab++51oPuW1cTB7/CXmwer+V5U4kcTj0EQ3tu2YcWO
HsY0Q7R2BT0hB3V8FxbwYN2J3FQoJI/g+7oNTWbD4vEd/TzRoKHgjcEeZN1T88dJAEkvgtM+VctK
HcYlRGxlF5Ua6ZOw93bdds71v9vkYgzAJIJKg+9dYQz6I2iD2WR9KNWoowtFbDolJO8bw8V9Nthl
lbzdUi2DqYQhPLSMKMsFS6zHGluETf3NVnigSyM1mAw0AYhyE9Lx4QEaOuGvBdjFrbxtRdlEoyqO
y7uZQ1SHrhlHV9aD5PHqAmxm9JK5fjxXzPO2ngf1H5zxeNzppXfFNYBtbjYD3KGbdo0YL63TKgQz
UM805/8+fynuj0FQ6jK3CoRWH8cyUgm4qNFF389Sk/9TJM3KGHdl38pMjUQJJps9bRL6RbIRcK/z
/9ei0+FFvyyUI6QuFN1Y7QgatxfZbc//LHtuFc04J2K1s4A38XC350bE/ucCWvUfJBcJWIskp1K5
ni+dIzcf7wWZCEZiBiLnDPeoYxamAnCEaVUN8RHVgCyDN0l8SDGyqxySlqNSrDQdLFp0lMKjVoRy
mIztDkSXLgT7Zt11JOjrKIc5FobUMlGJWdvO6132aUnH2Zfas2EgWWh+Puv08l++pKSI/Zhe5JP2
RIR7k7RBCySnfWHM+tU9kIPssD2vSzjLdlcNgQVVxXtvDDLqm4+JDDiB0Xe7qKGhDhirhb0JNCCO
3Ggk5SkywED5fS1A7+f4INj95NdvttyLuDizFU9vou4i0d+2pYIKAVkcGXmG36NCK+ZzvP1AgzV5
qpMU1Kn8qecg0xzpCMUtYbvOk9qQsvmJ5W89wg78RAY02CWycGjrJMHLQfcFt9j+m0mbMOtSbLGX
uJHawcyD9tyzOMJB0spzhCYqZHadnldbzuYFwdaz9Nb5qCzA/nxPI8pv8IKYUzTw34sdHdFjBt2v
hJTwKLOEYBZptnETX4NZmxCwKhOBzWb5CfsKQ4gMfBq8P217ovErZBarI+0bC3nuBFOC+jXiGVnj
Wbbm7aWwkJf43MjB8cy8gKb/m7Zr7UxXjI1LmigNr42TvxF2V8LKZOdPK8gMqXr6pNMieWBwpWMm
YGtqcu+fNP5bym5ueIIMPis3bTx6nFo1Kcv/nINBsQhqNkCapXRo7f0o5jUVakgpM2zHn2dcCvMl
pD/RCPbbueSLkqluO5nnqiY1XsL9b5wT/2Q7AthbullTbkGlfa9IaI78jlHvsoeFX5nquFAdrOrb
sJzNAjq28DPrry+7EzEmBkWDFbGU1rssOgFXSpBxb1ZeRmEjTV/6ZQ2/ceEckBAtjwwk3ktcLu1c
WXwaMMLxAv1YkmpjUeVuixEarMrOsmeY5W1hOuK7xZl57/dcfY5UD14nrBEOkrvoT6qbY3P3wibC
RVJLQF4zx68CRNvha5b/FRFeLRHmrB8xqchBtrYA7OawiaLyaiylBCsEJ5/qOVRg8Oj5T3OuZs0z
aIS5/zbeFc2qy1btzenrRNRRruxqK0hQybdYM07gmbf4dZUfhgN+RZzAArVHnHnr1xR0yLCZmGJu
al9e9SS8qAtksaF9dzLyah0uaAFqu7YDX7b+or8wpDvSDarM/nDtKigZwJs7RvB0VQcel+DxGMxG
V3VdfPUoHor6uT/OjZ22gt+plu6Uel41lN41EK+99YKRrrqdVQ2MPpxlOKkdHuqdPuMm3/99kKQy
fmgS60syOvgoCg8YmJgLJTexiPVLDIlA1GLA8/j7wUgdC1qXYPU/lEEfeiAI9kKRCDHD+2+73jsG
7SmGs3hXuJLhVAyLRno1OvjEyi707tE6NIKMcSWua96au+ZyTkiFxMKUyBeKK+dDrc+5bSKboz2N
eJF9wLjFO/luSwDSBRleRvkIHIyFp8exa6jIueX4tzEdCCXiGcLrQ8D1CQkkzMpmLrjiRk0i2grc
WxCVOrSzVAWic80hWgFz1SV4IIWPivkIfw7vNe1nQd1W83UJr/mD6j8cD/e9Js9lHAl8Lnv5LOYJ
AdxOIgsGb4AdqIWtofVnUI5ZZ+7ygFnjQ8dtHFcP3blUypnBefql1896xjjnqEiPPHAt41VL/FX8
VnBB9Y0ZFVeUFS5iubjb0j2Dc0+rp88WCCQbYSMNaXgT4KV1QatP39jc8XT+yyD2NgxYzx0r4kIR
CohZObxg16b4d/rkAqyMRCjYic3m37w2nVZJVfr4tAaJ30G4cg6Wp72rUHikKQLeoVtYu80Lfv9A
CdJyxJufHsrMsRVY3wuNtWm0q9cOKsnWQAEJ5XsZR8934h/QNOXEHFbFMXC/luNt6wwWqeoRhsa4
HdI8Ui45ClEsbZ+BnbkGLy0PRpdOG5OzteK2Y7Ml56WX68AYtb/PvokH4K1N57O1jRFG2TzzBtjk
TCdzRGhVTY9zQ+3fxk+XzumidEWJkRtz5w4JU0HhswK2vuxGUCjM9l71iu7kJkVBB7EImdebbjBb
HMEmNjTci/I/cUOFE25jycbmtI9/SHNlOmzZtDCyEEtxizoTIzngsEZEs6Cm2FPYQQ4H81DZPbkK
TbvG3qWteBV71g+txuJT+retLOBsDLBdyiVxCPMJW6lNiZZlyjfTPGr6frX7QvCzTMSX8nvlp4Vv
dj37cj1bx9I2Q7syu54KJS05hjIHP5fb7Oav4SfAPQXgU221SscqAEvxbaTfeySPhnM+IGZDboZy
vCEKMVNsM3GR82Eikx2F6nToNwI5mYrjl5H3LG/II5JHAGoMye1xCoKJtSTnqePcbMZ2GM0tbbnr
dKMG5hDDxOgO0V5pY1KGFWvZYI6we/XcSw3i3bBFX4gX21mpdcox12ejYmWhapzpe0L92Ebg/7Es
BbIz3ZZHuaYoR7BY+KzraAbDksHfQaz/rZGCxU85ela/FbKRFL+Rs/mLg2oX9hsHkCR9WjyXwpzS
my5Cn7pDbRjpUKY2q+CghoHumHG+pHusI+kR8qCchranYGN3QB+hn42ZKAsCHEr2njRXt6LfXIWq
C1qDzy1wJeJ1m2UkRvJeUTqus01l1p4wtnZlt9tOCopWKYucYNg7RS1iZprre69cYTW1eKVGIayf
jWaydYlEVOlyLcCJp9+Et+NK84VOmJ+EmWElmrbO/DWOS/nli0kkVXl/uc6fv+0HSWpuvFvaqDuj
PrmBFzcupaF1VR9418NlAAlcM6aQG/F/z+rsO+u+NT177XOyQWGZCATMnf3hO8qoDymrbAgBwAFA
ZayjmdCtQnmKUOuDqiEC/WHX77RYfB8S1bGC25FBfY6cdc15Y+4nNFiOSx3twjTLwim2B9a2tu4W
SLuaUdm6HPcUIg8vYBEoxMarDCPekLGkCw/8gmvWIcngRH/TiubD259veLIVRbRkadbKGHvgrqT9
vHI0L9nIwBaQqrrmFe76qxZEIYzMjbZ2AF7yQrcDy64yZkOTzzPEYJw5lwnPnMaC9RqEXXewy/lH
HIX1ol1qvVySRhzdZNGPn7BCr76MrxMLmbwrg0YxVF1uRhYpeURDssxeOSMAoPz9qy9zadhU2Stw
yA383jfrCkWJnJwo5EgxynYl1CxxAaKNGqUIXvNMidg88O1FGyiyK0v+m+kinjLaejaFMN/mltAi
avvNO3BDRVFYlEpb2QdSLPveXOUqVB4ZVPxfnY48F78PmS8HxrmeNQmvB5PNyD7jDIM54DQLiS09
SfuwsY4iTLd1Ns9tMzlRmb6ti7bvuMpHnBiuIuAxtQGEjpQHdFQQZGJsyvVkgRW8CoaL6kCQ8JNf
zK5EAed+LM2Ps25bHxvLnIAWBMPMH9j1GKE4NSA1bzSkJU8WLUcpZqfKEvLxRt2ycUuywURYGKUF
LivuNUV1ipuCkQBp+uJiilQkfzPkgU7RVmqxBHcDYqrDJshm6HKekPPArTuNcsWaQyMPYSWjXeM0
XHktEFbEKgqJsOrF2ax4ISOF+ffHSpwsKztZXuU8DrSxwVT2G9KZO95j3tfessfioClodkmbYbSz
wZNUt3dmuRaGKNfKaNXTISxZX20R9BKqsidtodvwf2a5MVkzp/aQg7pnWDZMt5++swJctpIVzDe+
Szar5hXdj6ZLrBiG/Mb3cyW5V/irW2C2AQWdAz5HlAN4i6gdYxVp7W+mKZeKJR3xjSSPUdooxbzE
q0LMGWLcEHwHQvLBSqh0vUTpJKso73SNmh2iUd8zrQuLsBlfWn8hssaRA5AYfQS8fOOOT7+tgHYZ
v4R1Sxv35z6YptWk75TPzF6MY43NM5u0G5s6/7Wyq6s9byP5e/JONReNBmpTkN2apQWQnMNeU1lw
K18PMFpiugFExEmpD0/SXnmsfVQ/YTCfJ/7ry4F4mtwYa2xaKzyMqN+OasU59G2zABhojx5Y5V8s
OJDhXBLb4+fJvbWmto0N2j/ccYJZ5v29dNXAfCN1Rrf3VXnRc9Q+SMGBTWQMO/jlKwcrN7+xMdFk
IXZIOVMfqmabIHgOXfzbOjYfzu+nVxW9gLU2RWTnM/pyqx2IWHBrCFTiz/U4Tc2tlOg+G35mJnoj
QohoT4ym8KxUd/OjuxDBQ9dlqgjdkmoalkO1ifcpXn9ULg9JA9IFQ86lv84MHdq8qxSM5viFd9ZO
IuvWxUMeKDbbOytagrNDBKkP95zn3BNDjIRAiihLUlqRUEigtOHo115nGOSSgVDljEMAPtyV3Mng
ALBSCgkqlF/UtMQ90+JsL9r2jNd6p0WQjjZeX4uQe8sTp1MoKrvORGMoXFWergQ2KHnqEPGpAk6+
C2+scSVdRrkxBpcg0025XTzc00za3JqWKaz6c7K/3Eodrm1UfC3+R8HOV1iNTRsYaZzey6o3g3P3
g7iqit79pHDyTc055zQUQsvKSah1Q3j9OVcd2HXQJU/upurTKABRm3rZP8kl8gmCddiyekNi1gum
H+tUG9G8ToZ9dAFGbnhOl6C1jaHE8dwpntcD8mn9gMB+UH0KicxMLMweVQPnt0dv0E+QnEEMQjFh
axBl4gZPXkPNUEuQc8aOmumZ6A8JoKRh7UMpnFL2aNqoQnwyuPxp+F6+qeWiNrCWvlVZ9bMQY1wO
MGA/lGA7hXVVXJKzxBOoAofoSaTh8PXr/4grvNbt7Ah1L4ER/Qa6a7XuztBcDjk2UlUhsP1cYV6N
H5oGdktIl0XYR9hMWbDGyX/kd7hELZPK3bxwtO/wesZ5AmZRnrtl9RMN7ea6EgvNFcqk7nn14dtk
Pr1YhYJiSp5bMWtTbuJtVSIAfBa8hJVgdA9UTMERll3xqddD4gL/bKq3xnEERqCcB83TxOfR8Xbd
64TtDqcAQe3+sfoMs1Hktr3X46lvKj6TA75jvfBey/tG8fN7yws8iUDC/lnGTnt0u6W92W8l7iKJ
deudxZwvuyi2VF/VuMSoum97Hj2ZOzksNLMDvcgDNZpDq9jbU8ScocVn+Nch1tUhipQ/KBMpJT8O
9mElMnpIfRpqPDJPeQuBxXi0Ooc/UJnjNjNFtHraDrVZ20mtfEUKVn943RlNo6s6j3MjLbGpyvZP
NKFDgE6wP1U02dhoNsmPt9O03wfGG6kJRIJT0dF1dTKOSc+VCR/RX1HACvhxss5rUbK4voFR3m3p
oYW/oCFnLE5PtuBGas30RP8Var1uHLIFdIEgoEfRjTY6PNG4yRmJ/qFFNKMvpfkAkvwMTLxg+q1l
QosoKGcjg57pEmfvczyVp2wr5bd/wAtWwEeGD2LkcWb7wFyMZfoPIoZ5jNY2DJt3DrPbk0FpyP0S
82u01NGGoM2GZPD0S9bE3CpzRhLWpK94YCrcz0jATHyncKjCZGxdhwpuIbK3kHyY8g5Mug0s7+bA
YiMRB5Jx0eY2C5y3VW6lu5TgYCHhS5V6YTPUXj2VVSQ8WrKW9mYZN/EmY2yWZ8aoOpRxen7znniG
3OhBbXeye5hDJdwgtKTIjci6widE05UAmZgCjxMaZPpLDSXVnwbpueFUm7HNDlS1DskhynL2Z0An
d/FjCaXDKhMmQ/Y6/Z01MXdBzgp61+dmeDX4gxqgZuKrjttWSOMQ4vVkluiNFyqWLhtZ9TVzAiLw
OX21bFiJqo+qAHx3EnuOFnK3irQicUsGwx9FDcNMoJcL251aqIZ+RPgONY38WaeiEKFvjuu21jIr
Qg3tjyDxi8B/uDGnqKMwCrciqYbGPsCL5FB4eDWzO1qtuC3jHneEhX8AKmZSdDUaiiFmHhHqT9j8
OpLYjnSeKjUgNNdiIhmB9lUrfn7JL/g8I8uxgaiOwlLFck7wt8rVeM81CtxDL7D0qqWaENM/a27G
ABdGvKtS66Hw2c8GzQHZGkMU59rJg7mB2mT1JvICOZOvh12egsp1ycUxJ7WBCGz0Z4UjnVhkX+vu
8K4ir4HbrwK9KLp0O4cVBQah8W2tMagQfj/dXZG/PCCe3NlN/k3dOcDpeo5IhYdHnWcWhOiJKaLM
adxCqeB1t1F5tpdhzrmvehvzf76SFgKivjQ58WSDTJPGm2rY6zmk7bm1gpHbCPkBWFoaHbPxBEt9
NRmgYXKpLGXdorAl12EkuAILaVktQI5QGk0aUMEpudHh4qK0aLxxbXMRMvJuDFdZQh1HkizP/mgx
mMdcgm8/HSVKlATftlNtiu/f7RS8/VM8Y7Y3QcaeWBrNM0Qd1G58QLxSCqPoql+mJ7SVdsXAcPPI
qrm06HA+ExCYTD7upO/NRxSTMLMcKd8oNnze6N5RNB16UknciqHr+0qz7dEwOZYR6PujUSYemfuf
cDZFGD9TVLZb5JHktoY1kY//U7rSOSzuLwj5K5Vwi5nItBMl5XKvr80+G4VtsPGlvsL9wBs3G+hj
NQKi0o5opRudavgQDqwhx/5BygXqYKDLjgcNg1TvCv5LyS6QcnHR+Ycfp7gbl3tgjHgi1g2jPqoC
5LFLHl0XmDXcor7fX0SPYs+CkVFqLEHBOMnOBieJMhNMze7f3saOXMwATrU0FYd+UvY1sCSCxNnZ
xbvKHnUof/uwbu+BH5Cr4xy9ON2LUfQqfd4k0pHPJuEYVOyBDmgb2/TKa45s0oeEAaZb8fWSQwLz
+4PlKG0fs2u2MAm2qQ2jZGEEdKDMJrj4qHXxomv/NeUSZP9ktt/pAZIUEKfZ5f7xzq1LbhB0PN7j
l/rSQ4pYgMMW4rs6JKxWkDDuVNvrnW5W3lKdwV40Bsgid8S0dkIUl5meo4FaRr1ZEqR1vFIViNYs
3H5f7QPOzPigHVuJjdQQUSd/E/5DjLvLRK5AtKCal2g5GzlSVPiKxVZm5D6rg9Ew5PHue7kd5Rs3
uRvSdQiak2tIpGhGhqf4MUGoSJ4+maQAjuITaX4fB9tm4ofMaFFWbBIkwqgN7povGVxLnmRBQn2m
ttkQIXmI6T2dwdDabai/xG3XrYBvYHdZZDr4PRpJhqed/gztYTr41aNF47249SjnwBPQo3TdvMeT
IitJiq+Y91x2kmyVJdCjKJgR4ICgQFwJVI+RB0vF+AH8wIIeXawMGKWH2ht9NyBTR6OzEREJvH2p
jxX+OxSAS2/U0wpoWj/NtVLTa/YBLXJLyyqsfImWgDclu7L9E3ngMTkYUQxumdZ6nGmM/Kn2wt1q
l0TUc9U8ZAamL+9M2qcBAV80ZaC81F+MvKt3zXNWtOzgNt6jsAU2QFccvIztewNAp0nn4rp/s+AK
F4PGKDm+qaFJKcRtS0O2y30fdh9U0d4Qaaz3pfvIeHWhfAzJOAenuaOTdYsM5u+HrOfRx9SJSpWH
GFzYEFxBHb+bAXM01xHBshGCYdwddCVi7X6yei9R5xCsYvN+kVKo18j69L1J3SQSAIUiC158Wnj2
Pez26yKBc+3dP/e9h3sFh7xSxXvD6rEqeTrdTOS/jKNXdpN9hekmK4QOtZrJcIWTtNjF6rFFnS0Y
s8/5MS16irY3wQ+4Ug6Zc+Hv7OhXPJ2pxoFdmT4PVnanqN7icu9blliHoJUtR8xkw74P3C4HLrZ2
bTxPXhScdXYS5t/OF6e7BFGu7vaShULt4VSQtETi26JaBYtv7kqLMBgHJqlixWqh5kVwi1obXVwn
PvrODcbl9DA+gH6Hc1QuF92e+Nt3cyrzi/g4apbZUmXAca4IYkaQtjyNETjUTEi1wcEDFwlChZdX
ih+AET3o3Q8hko4R61fBj3IIrxEbmO9xb04Wx9Zco4Rymlv9qk7Q7MwR5s7fJf3hbWIOLLmEFG3b
82alNchdVeHRGDOgNo/kNPc7xVzFPIs72bEXc3zqKT4oybuFd4WeiFDNY0lbBFif/pX04eODEt70
S/GAcnwL2+nuqtI/zsLVSz2cWJLap7GioQJXsbGnB85HMQNaZaAohKVdz6eRl1RbCdWZO3IzJWx1
rE3pBseioJ+o6B+QCrbwaEnEBlvoLWgRJA5AbjPIBrJaUC9UPgKkevz8/3qUhE3LSzC6mmfdRiNq
ygNxFebAvxEGM2vhS+bZCQLxqlKfk7fqAmLEf0B5YfhdYsMTMPzyERoOtFXkEZ+koIqVfunzOafd
wkf0k4V3IAQtT0ITEKO/L1YWYCesf3eWDGJ/7pFzA2mMCKmUdJTyYba+luiJkmG1Z3q5XmtaMVWo
GgfrSBuCe/2OpGCRG+fRL4LsA4zBIOjolzc1zMGLbBFe7bfaLRc+U7WOwFByTkhg8CmOGwhR8/ex
D6YW6rg4Cfv99hUyZXRY54t+1Zr6KSUW2iqqyLprPaPx+Jys3IIfyP9RkxEdBc7eIi2DBpAfJRNL
TyfYWe8zkacSIhFP3X5ZTVGLuPMgbtrMCd8F6uqtY02ETPGpHIpIpDMBt2brYVRo+qS26y9NRIn9
mmIlEsZo6BEmL8tc1NZ6XXnaZSQip4WjL6I7dSz7d3QNc2ZnQrlnkxzcOmL+4WGtp1/PVVCF2Og/
dQUCTpv3OMRTDbVAPp0yoRHksnIJLyoWpuCV5zYc+UKCXjvnRxnrzD/chzXIR3GiKtF2Q1KdH4l8
/FvXfoP4cWwStZaU2hqBAFOmwKhJK9V5ySiIDxSijScF1UjQ2rWYqfkk2y32hJvvaXJBU6tgaBAM
S9UG2CR7TZYMHlivgJSasuI1mQ/EvhihiJPHwYTDDWq2oxxPoGV0dDwBINuyyf4G34OiAv7p0zHF
l5EosC33sCCgM59y6gzkTd3xpPy+tlgnH2i8zbIUsgRASkk/CRqJsw7AE2zQ+jYCqK8flg99kqaX
zzEbID0bVtdyP9zjRpl+pikBLodlAttwzNFssJjVfnRgB3D1oXV2txb3EFHHoO/IcsWCcIuWzSVF
BqPHrVWTRJfjJawiZZszGiGRKdg84i7Bvglcb4qZhiAU74VRF041ItsqSxxmB050bn0ZYHgFwbYG
3i1l0A1/GDOUGROEbGOEuNT5vLzU32s7Ppo7VqPxLYeAh7wwkfx2otT8YjwRWynkYZHXmrmTa1EY
cb+urypj7b9rCeXtUGmEZtBzypzqK6WspyrLlQy/hmh25oCeBl+Q6lo0FJbOmp3l/6EOr/v3u6nJ
26bySsHZRCK7U+ubtZ+lLsaLhsse0PQLJ4eDwFhaFMA7BBpDj4IdvR0hOIEoQlzbzJOSTJb+OLhn
7jByG8CzFJI9/K4VI729OP+4T7Ro/ypQ7xYBACA2JnNhHnD+aUbBdKVUy36Tl4MVbG5scl27gWMV
f/JTLrxl6TVRcalx4OtA3VnMv+0dm3asnnBbZBcveAlwy9Oa7YRefYGt2WaUl2WqNox7zDY/4UMU
klJO4iDacKol3spPANh0PC7J3LJnBnZUhi8ZjTsRGA29SYKB6SyHNhCWfWGVsV2kS62lNDd50mfN
xiyHJMPMZbsUAF0KKVBrRhRWPRx89TSdn1cEv/Cud6FI5CnSKj96kbyCuyoHLkEdQDrsLgwp84FO
446f7OjkCyaIJJ1bpbqzOodnABkLUD4fVLnngkTtE5z59wPyPBIxVp9FPa/XY5ThYviNS/y9EDWb
GH15U/Avc6+C213CTqv6QiSC0t+UY8RynB+iIrmgPtxnbYlYuebW7pnsuxJm/KFbAagCEi9sj2ji
DzB16GPMRU/YusVvl2KnISIYv18ujHy03/w0wpPragtjtUfN4pOhTWyCUlMOHt0/bvetl62wPkOD
jtSFqBnU4KzQJVawz7JxU+4eN1Xq/ju8R3uBsBpCW32vXU+SQ2olNrh/BNW6tal23FPVtYTKwUc7
430Vp+htnlrDA/qrVFPkdvjitD8WcaubrS/r/Z1yr6FheYseUX8Q3H/W6bIE474gV94tISDzo2xu
C6km7VZuWWnHClUGtJnTgluIVEb8mxvg7jPOLOtSMZ25OJLETaQWwUlqFl8Ly8OjpGZxVVnj9hxF
SNeIcuvlxIPd3Xu3Gg6pV+37qZZEJAeouoM4VUoMSdQSy9+zAHu1l6E6ye2rEWXAC++m3bCvuPBx
U4MZcGhSo5KTdk1FcmUm/oXjXf5i+T/O6YWV+sgDItqfyujyOCFSDUnk8nnX15E2Kuaki2mBz39v
KxYiGsjGz09Hq2rZRRBMSLqKy+WDrIoWRM0f04Bd5r/XLo3KviodtbE3bJFbAC2/J02RYhHThScb
r/V/kE1PnQxfE6KY8ZyjuRWShuznW4rJVVqZ0D2AzqWTan2pc78wSEbebtT1Djhnb6TKvTMhMVst
tNohqhyuGGCAeBV9xOTE9p74ap0v7dUD7A4wIS6a+sfcj0ajVW0xIGCAtc9ROeVAFIhRSCC9CX9f
2XSuW+29wT1YsoWFQAmaeFt6dH7Cj0nWC53FklgHpuTg3DwE9oc4fQqiVGGuWILPDWO26H4KF/z6
+tSTTST/bulSsgDVXvZ5z/UdLAk+yVWMUrW27jj1Lj3cKvtjdZio1untCqNIY+gPl1EgD1eq49Mb
aqWoozi+4AoHE9SiTFsA7R5fjDGrChj9BIjn0G9oo+PIo9Kkve1bgRqynivP8D4R1mWYdQZuMHS6
iCaqyEgCGqr0muHfzxnZEFjEbwgsuPg2mq9CJNyZvauTjx+RGclOU8saPgFvMeIs2aMuNeE6Yj2W
RKyihTqc8JTo3P4qqNrh4LycqP1HTOFvyuZZ7gBcdoisBqTdWtYzC6B7oDn2T7f1rjSoHP8LlC2D
QScKPPdcBhxG3cqA10+cxPJbqnKWQEuzPQU/Z0MQkLn5O0zSl7smNn2/XNb1YqJoLrc2w+9SudYP
zcaXhSUPMriaZD1vDJPE/ehhoAo4pxoFsfJaBE24Lh5fyFjv7ieFpKjKz8ojHISTdUEBhlCmO9Rd
kiGBDrlAMgjw56fqyqDQ4zKwQGC/qw3+PtnVbaHPXgS5bNZIjZtfBwCx3IyB/s20nZb61ilpsI1v
JcBqqeQB5SOw05K0IJjkuQM8IfO6TQIE8wdfLdA3FVf/y8VgNJ+DKA2Vn9vlqKFSv4gGZ0JcM45V
USQS12xHbJl2NXisohSnP6dQJ3KZIRvHIt9CKoiM3jqaDA9dGbi8MXrVkUzpSlkO431K3Co/p6g8
jpf8WHPGI2n2BDytrbRRKTFjcGZ8Vvbm5uIByQohu2D902+6xRJoi2njvQE0xY9q6ZsvfF1a3Bf5
G1ZQ91ZOCXUUGkll/HMF9RmmjWdR0ebNNMxeZbopb3haLDxWgSClVvp0189yn3Tt5QSH14jGIDEH
po5q2iC03ewjDWf8bw2qPwdE7G1+zblOVilAHkS3ElJdCxtyigq5mzj3SfsPG9UfOCb97egJFvfq
YftcYsJqL8WINMt3DpyMcqgeKTRXG2SSIFQe0yHvQ54csue6Ox3+YUZJ1ox94djIapvAQ8hReo/9
+Q7oM8JmueaNmi4Ak3Tp3yod9F2aorVFa6H0coiP/PLSHZBAhX5dT7Ii1qzZpXsHB0tJ02rRBylB
Wx9Dw3Prar5yINYzjDKL7eu8MN62QsWmh6l8QG1yEz5VuLezBKfYvNi6oXj07al2Ikb6egSNLnpB
hvs5lI+ybQbbO6P5f2A2BpN1Qbt59WP3ha+VqNxaLJXpLNRCtDt9jvc6Qa+gPjIChnJ2vIFR0IeC
v33o1t7HjX0pGz28hE/aUD4tu4zEu95oJRmuvewZWiXIUsyLSnvRjvhjMdebK6PvxjwtNHCsKRz9
GRAkxsmbBHuQUr0M0Z2WJcPxnm4yEnaO5yYby5oEFVmhu6r68tDJwwJ2OhOAYW6puRN3nhI0U4+i
c0kQMAyieaT2lGTvqo3jTOo42LdrdeCgjqPjS+GUTEh0Kiu0WNt0yJIqlVR7FFF/jIvGKe4NyoqE
/1EdUaSkV5BTlFVO4HeuAQmrUBHhvKNI3IxzuJDcGDCkwRC/jA929OYaJlXWnIelJ8QhKjIRtahV
uZeew8A8tewP+BObQYoRFijmV2CPZdc5zWuGQ0YBJnIN95DqDFGTVt3n/7AN8qwSuGvC/HOnZv4l
Asm9aMM7RtIo5XDYBatx2Ib3R8FasirluEOu89fYzHlxls/K9EAPYLpQghbDJdgtK/YHqJumJShL
JXlqggSqvw9iwVO75A3f32Fsf3fc6jmHYXJNhyVF/H3Z9WKDjgm0KhkYwv9d+Utbq2c01EBjH7Dq
SanWhqPhr9Rt6cAibhXT/ETScDvxzKAnFtOIIbnn8tlL28PWjvCCEyNDzjegEUYCmmYEt/zHMMBi
y3e7CTixh9hmPPIDKWCWTGTJNi9LRIN7iVsjBTDXGlpmWx4wRO/NW1QDiduJO+wOUojEeDPnP4GF
+Nc9bcs9/xvjyAwB0iP56e0r9JHwjThZroOuq5y2eEedntQ+nJKrOGrbIvs1VA1SEfo99E1UzMpO
4GceXIDF0RkNqLEWg/wqt69PGgQ6lZugGIobJ0asQ2r1RIC/Dx/bgRIOZDCG6a61oXUO5Y+BnT3Q
AM43sDAvCCUP7JPPRbsBCmSyjaMtS3+ZiUDuwHyLu7BWaBhj7FRruh456sSdalkbM3sbgj/7LsgC
HV4TcxNkRXjgK30LZ9VomLtLnSgWL/oPV0LhMqTbS7v2ELXEThjb7PjMGZb2jew41201xJEuguUH
NMeSBlQuLTrc2jVkXODzX2pnFj+F2OpRUYXe1KT0lDEFby0rofwVy5dlivoLBG6ycZJhOFLWddl7
SLZ8EauhtzBX9Sj3gnjdH9FTTESx3TwxCKociJm+2j615IVkiMINb1iKU/lMcnWmQff07rAUGIuR
VmA+sdk4FfsiIPXtOGkG9SyT21oVY5FR+zskylZd7Qlcus3a+vAcZAPlYUlPdYyEQEvdggfTMKoE
a3DxSW03L7efIxbEpi3ZY9D18NsQ4aVYUU1+EulYGwrUT/8F2UO3bnFcB+UU8nETPjnWfMLkOGbL
fH3JxJiWfK1UnQwHRZQLCu4oxUcuQUXMeSsCMT3eIDOu5lFWbjlgZPAMefuI5fs8ow2DIWLCf/GY
clDOfsYml/v8f0aw7G17TZfnfBwLjNZC6GM1YZqqGaOKoRmtRnSmjw00LmK0iXJUyqs1QMcBZQY3
MDxfcEWGB0qgg8O5iUdDC8BuQ2JBGFD/RiOWzyxzAsakjIvu9PXXQVwXI2RoNmpYYP4dRL1OyI9/
b6GiIwURPVGRPIoSX3tevX4Gxq7RXJDVeE0+qXB2Crx0GEvbdAn/7QmWzF5yrefPuJx1+f9TUId2
1elfcFmlwgSNcpUATLgvJSLwwjNnZUkdRJ0+aKAFZfN9hLL44TEkegM3rwuguSJpLVtza6Wd86sU
u86cxnN2fS3hmn8MkvsTK1zkGntMUB4ItFdK07KzxaR4JFreiqJcLgVRLbNe6PQO+L/inasEzrRJ
SuyPY0NHPUSlGdSrg1JbqyFMrqeJRx2mmsN9X9PeLRn59sVXdfgdVMvFTj3hUPhzJTX9y1zqaIL2
PyYaxSwZEVJ6iwxujR6maWWG2UGMz9hs9hGng/5/Y1MYOC+FpkojspYS+Nzz2uVFdaEf/cL91tE6
y10x+ca2x9kTbMOSS8SZH8jCx6lbTb9ANXfCl5EFcZqU71o76cH58azdW/enbno5IW9ShyRmWbsr
pTtYhk1zz0Nq/8KrgeJwRu+EYqZzpQ2Qzr2Q3P3DGyxiv+W3ThA/BUlrk8K4qvH0MFWIi9U6+jNw
Wbz+sOFDKvPh6j/DZwsXLsc28vfBfn8NXXN+ZnIdV6L1mDcTZ7GbNb0HAFEAnP2MlOCyUnt8ZJwi
vrwTx9gzPJf2zEZ5aIrfAIcoKtWiHXb4kTLcpnnE0BPR64GhhfPNLZ8yDLUxjwA/6rb78Yy/as4h
lj9Bmb9Wle3b0vH4z8tKRIooGlgyRwY7yZwaBVA7Uy4fWxkGlsolvK65BeCRuEUkkxP5q9jp3Rbu
/+8IgNJ+vCXnTpAO7oHdsTmF9RqdDOenAa1UettS5ppUrzyat34gRqvBBVnoLwbaimqvC+QooEVx
lKSxM8lw6w6w8o/puTGY+5//ADUqzxa5f3AyaBPjKrF+J5nabiOGCRre74jR0eJ8oPiL38rpGF56
xDcvZ+2m1H86+iheh/F7pej2d98EA8AdWYNFQ3HT6Ep+vmzhjArvuG1abxmpQnzd+6mtnTcxiS1d
bW7ngZBwBbJZ0rmPrmmMG7sBVAdCvBn9vnXf8DGTSqeoCgUwZXmrgAKT8vpidFjjimQGOtOs4XSH
4AbxUi+l5T5CZZ9oYZS14wvCUdJd4u0pdoDG6u0qHTrtX0tE3uLTHyWRFLn91cC7VDJRr5dsaeJm
TMm/ab+PbCvIbLDKiKy1oJHnVFGkPD1ZEEmufMzEXVO/mIB+yUKxAYqlp9cnYq8TameXMfDFwkUO
iBUJeMHOk4GQvnUmAAn/E4u/7hgcuBwzK70KiN+WiLwiRxFV+xjW2Ny5rxszdDA2ShEJMIZVlPsc
erXFTYEmMgBeADD0vsNP7rcsj1YypKxyt9hoQLn99LkenRHrP2P/DTx0rP8+qGR/wFfNW99EuylL
pTyLdyVkk8iKy6OsEDMwDfh/6Dyr1zDVY9IJ0bENlQXl5RB9v+LWf9XmM9fjzpjxd68TkNcVq1dk
Jb3oX/+VvWKW64uBdyEBSFX8flLvuE6AGERhx8ATlF299e+S+2nOark64brKJL2QvUvDeHfCN3Ll
+4hCSbJFALNfmrOWWlo1f1ymiy2AVkaZfbKvM8g1IgdZjRh3Ra0VtTNAKo81PGJv28XCYGEWoETq
DHL7DA7aMPbvQJFqN8M+mFUc6opU67wnxrxVuR+h6AUQnQDrcO3A8xrRybh5OlOemJbmxXp66wIg
eOKc0gfwEreQhQPE1zJPwIfngUxN8drqZrNKzm8Y3rG1NPy9LxvHRMA6Bccu2w7Syen2OFkIgO6/
V4u1fLEiwyl3t7g30L/NDicoiHw6i7A/Qb1r6SY/QLh3rCUAdj4foxiozxg47R/pJWMNqzXUL0kM
TplnUAhzymOXNLNCwzGRqBWpnhfN0fqiiqGlsXq+gqjKtcf2Cw6td9QpCvenuE0tIy4z1EbNtleB
hfXRhBD78Me8FJcnOCWrmd5B2DU1tF/vpjZvajyeGCtqOYbLqwXrH+aGseb7tPRyY/CiCIc+psbC
lggMoAMjin9PP/SxPmRX70WkzF/VhHlAaQCCGrkL2Ge7HVrhg4JIPQchsiGyBmlIvVbnVX3+8Sfw
mP/vxXBtOndQRR7CTr3JRBclo6hZAVAhVgEZ9xhiGQk0RXe6n/4OVIeb6s42S2COjJwe9V9RdETv
IuyYPTvaY+LBU7d5BQtM8lxX3aJ4IxUgQ3GZL64a8Ax90IigLcrri6WehYcs8hm5M7Pn1iR5gjNb
q4rvtqapOV7PjQTBk6uIwirJKLjOI54lW6Jn+/MdBcOZ0UAyk6SnGwKqNok10eXYP7YJ0sMF9rd6
zvcTNGIsAxjgA6uNuia1eOx1y2OcY2c71t5tf+Lmh+OVHVmoVlO7K078VI2Tr8EWZd+qgXQKLrb9
x6x1xNe6LfwzEbbjH3ShykMNvhwiBEqQbn3Hn9zFZsXkafQMnHBO5LqB9TDEuYmp9MrYTKwvVONx
I1e+NFOFl42T8mFkv55hfIG6nlIzMCTQCpAr8Za4v+0IieiTBnOWwlde+cNyKIJj+nV/QPIvrYBj
X98I9Kyvuxpi/d6fYINmy4qEbKZU1ecgyQQs68c1q2LmscQ7rXFHXpjtHpZwsPnGUO+Qc/+0l1bi
4YfFFYsXKM0bkGI/GON+EtaTw3XWH5wlUdDeo/ZtAYbsQr+E7x5h2Tef8cRNrW84Z4tOqruMmzdp
z45kTPS+vTt4kYaH9MrJw4wNP2EJYQJR3f/Ac5R/yqAXL9Q0ksQH+P2QkcsnJCQ7il5p6pSoixCy
hGeax48OO4+/6pdyntvfaWqr1abgKHjmhoGH1GYcqWVp7hrVUovK58Smp831IiXqVVykOtebi9Np
NjZsCzrRAbJGrCoIUX/IOQ+54PV7sRDDtNbiroOQYG5L9A0r03DRKP6MpQyB1pf0fiZDKBiiu7u2
eqnXfAFv1RiyVYjtFGqaYO5odIP4a+rHBDy9vz0Dfzxcr9z0OEOVNwEYqze8JzFP4/l0lkMfn2Pv
UmzijenS9zZbu9zlO4Jc50s0E/lul3SYSG9KunzlhwG5lwFMn51C0svxOpjVvwgw+QZif+AAtR1b
3Zmqx+c/sqKrO/2h/ZsnOEqupHRsHkFfV2IHbcbp9RY1wfkBuUnvxx/48uHt1PNajvPD9aTAwErW
udBQ+VhoA6FHtFWrjC1CS4zybNVOVOQ10i4OoF7pQMFLmorlrZh3JxAqYt115T5ClV+ip5w0+IhR
bUf171TjDcw/aRW7nm04nxYiScFejFUZJob3jSGvYeBRLzmtUq1rWEzFDHbxON6TBBxItvB3YVbT
g/4m6CIBpLAzDHSrz1nJeEmkTqBqMNTS21rZjYlqFbewfDAOCTGSCJT9p7IyaIRkNGfrWEsPDSnX
Kl7UXy1D8huUT20X0pK4THbvLv0/kVVzZ2SclnN9i6KrAFngJG7a28NPfiuyF+tRxy+L1HgEsPM3
p2ZuaB/KaIxRB8KaI2ZhIdBV4gQk5u+se7Uj+q9PEfhUzRSbczovQMK3tSurmStiT7T7At1nOs22
hcJimyJFfOT3A0APr0XBLFXf4KYuFecDVIpEHrE9bqbHr2HHmICAPQaMHQeVQrA6VKF0YDE4DAN1
DpsWfnU0s5ZUk9j7HbFuHP8rqNRPU1v4hskaziZkl1HMD+EEvlxrWpdDS+9Og6ykl5V+FztxpUTp
yUoML6qFW8sMPd42C1RYM6SPmOCxcVpFb5v4jtq339meo9vK35kEfzYi8JV/NcZYc3kRX1NSu/xp
WC0zKii3ic6SyYITzcGZCvzBMlCAq6Nyd3I4rslwrE99w7k7Oge8TYpVImPjoS52/ptPvVVjMfvV
n1vQw9At7H5OF9fe3/QVpL+6Nlvy6//dWAV87F/I74A0IjIcm6XHRiQhOZrZOI3TOAwVN5N37H/J
wP5A6e79RcO+MsElcjsqEsehj3BUQyGjay+raQWAmRF7+fEahRsJ/4PEwUV+LyRCS+0TgO5DG+78
rENUkV09DRRT0YWRYkSb7kDwvkcf7+rcCMKi7CaF5A1qDVNg7RiWqZJur/m6HFCfEjrlAV53s14r
3VnQJSJbN3nR8fdLURt4n0rhWGOQ46xzFNuNPWiDItmAvXU1zRr6Ww5XkI4KYINQ5jelDEABY0Sp
DP9nhVTBLv/nPdecRQ0EoFyAQPZDdkbaqeSjUhdAZAywld1OvrLFDlujhcnSFX53IIg2n0xG/DiX
fbWgjGICeFRqixZBkvWBTN4NYcIz5Lwf6QC6EZrORbnmV5w7MZY/oDs1L+EhTRTypBJjB6Ihk+na
XdIxf6kXP5t8q3mBzuKHrgCF0wGSz3L5O8SztCJXB0U1WFLjepR//vnYp8aZkt3Eb7Rsgu2gFsi7
mG6339RyA9Wq1RyNyEL23VbR+2R/hnre+N6GUdIhOTvmvS6HnDggdEQ4bwOru2zLXGLyKtBQko1y
a+qLzCeji2OKXsJhCNM2MHn/+9XQi9ejdTt02xdHPGJ4WHQplJqxc5lC7uhPTFcmu+Dgridam5ck
QZrpk0I9nptT8NHh50f8W0nSFjDqV2aJUkodMTANL8urwVUzd/V+OFBPAgZt98Sm/6QOzdWQ4rrW
3jHy4oMiojv7vKNmfFEgL1UAjlsoLxYU8nRs+7aTEjc4uUrhTAo1PEhe2fHkzzC3bTF3SwOaZKBt
k/zH3a3s2ugX75/XAeZqQET6PLu8+WEt8a3hmfvFod/isVKhGcwBFIgDH2oV4yiIwvVq6ccRvGDG
xJRvBOTh2LkKZsxV2Y7uQCT1OhI2oep20QwG4cB4/UdK+tCEWSMsW96USw6YhnCPLnZJ+lvwcoSo
YC3WDSVnTlZ7yUzzFc5GRzZZH1yL5afsUdLJZJSPzzDkxa5rOjywAzpcbO0lVWa2mFJ19YowrjhK
8f+ffobOOxHROWwh2/icv7kuNZpm84oqP7xmS3vYGPVUGI90Ae1B7TuYQntxwhZ/1vquiEB786YK
bzoRm9hKG8y/cdz1OhHPjlrXLkZM3NcQBroC7w/gekWwpQDgy0z0AeZt5k9qw89DKc4x+qDhoP/5
QNrQRCgXmgMp4uP6CARM8MJ+n4DKMRclAGEoa5d8HzMLpf6p9/LC99Lx/C6MTcnUkXsqSYytTV/0
TGxQcIzIu8jIVATxH+oTWQzoSNG8SGf3l3rkt4Cs/dSP4aaVU8R3Pbk0zfWpCgQvmcGhk1WdnA48
a0pftkQsTfo5x8e5eCeqBqaPXWc1Kje+D3cPoh/tdIacsNfafjl8rDqiSMnxLVp0X+bGMIh7LibL
YICIh5ciUjRnyOmhUi13uT9ZVm8s57uziULKs0O7zy7imQQVBSzo05VrLUyFduDeSrxwSfpS1rcw
DDq0yfZ2/inGl6OsOMyo2TbQ1umXXHPkrc25MRiGJmBguEWB3eYq/RRiaDIFFTm85kSzHtOi0Nb4
VfhKdLbMFtkd4mcmKNw5hvolRPbR7NOjV6aJmFdiKJHeeFjTn15Ml8rD6E57o3HP1LaWk/bUT4rY
MvIPDPypSgnHGNDoG5MTdp9IfEBmZyWFRIge9krK2j9qqogE3/smTP9007fY0HL4PVzQi6y0xkdw
Ni4G+98ZbWQxsdCuSu6zpSfwNvZ6Bxz+IwyW3GzPVr7eVAWYQ6DEKNX7R5gWzBqSfIrVDctvUMRC
L4ZEke/pDsnjeE9sghTnPcgPfTurYU51+yL6OiDoZoZAWSDp2OubTRDhn5iU7U00E/+HHFpMoCPU
EhjxYg92c/tRUzmvpmVUtvdiFCtHizcR+m9mpCd39ryerozV2tcHWObf+tMupNDE4wwBq3z79TzX
TZ/gHLf2DQn5MEwxLvSnvFhRaZV+eZsf2Q8K57M8CfFm931XyQlBFw9XKJg2f1kXrTErEaRDbqVK
rvp8+ZeZ+bmHNWb2tINxecQTkXXysQTHZFE/EjeQ13YqPChTPQCinykAzodDrEPCdJEzkd53trt+
BEAXlpnsuCr+JicjrrXzLNgCZTYsS1NqfT+jSIVh/DTglDhndPxuv8ZdJDzJgxWTZYr+Izc6hxvD
Twkyfc14xNKZ4rOLQFXXWleqFA4Y4YrN6e2apVWYYda6abqWJBsZ+CgavPSTAJRYZ8tiV5AijTyw
Cnm+bUAl09UQ6wDI84Y+YiEcyFRDBclKCtvYEnz0UdbcWaTE4exKJa5dlmk0DDCXI/vno13g2ucc
XdrsbAuJSgO8gqkmLg8RQq2V8mBoeMl4966X1k1NUsSdSc6zRG5AbkROL+HqM0GDm9lPB7v41GZd
iZfgf1btJ6Df5QamzluheEUSD58pe+9HefxezKhMVQcZPk6Q4ifWbLk86qrfuXx1LMLKB3dqB9Pm
lWkBo/TJmLV7qGkZtpe40wfvP52enkzd1mA49I5S41vShnBQdSjnv433LO/UscETe490dRmVN7FR
P7Z+G3Vwcxs/3G42uVxHZAwm3hcS8HQuO9zedl5EiqS9E91vIVzAhpoQUbjIS5N/gcNfm+4bkZih
ZQ+B7i2ipAZ+d+FlOBYA171edh6fi/KD91Yk6c12Dj9Vc1/FpqlfJgaveR3vTKzXlG1tCmHGNurI
/iRcoTfikqPI/TBBVA3Pc3W2p8oghL3wqrocpsHtuGvQDyz6OG+f1bqh2LO8uuBDRmErE54kJRK8
xAaqFGygT27lWfa4Z2pYvtngx9lKHHh3pHw0NOJ5zNBil9WonkoSB+O7Ctu4qi7LRUQraf+iSufi
jJXlPuGJxKL0YzmTa2gx3LtWiwTsZI/50G5vgLkONSBq1MeRQXJEfEg9aFpulRrNdnatB9RdB+da
m5liEGpnKWXHsGExjNmfQZWmiyGLy7A4NQk2vdYs3LUr8+ufxcmxlNKTsdDfUsmwqw1+X51yCjT6
Id3RnGSJh58L/2L9+TFFPTK21ErH9O9S69Eo37mH+kC4SlUO3dBxAOgy6aj2B7yRDpjWdg+V27wH
g2rlbZTEbrltW2k3H6JSuukPitCGGQJQBnHzGp2XZoFE2mHsf030+ib5vPSiUvyHi2R2G6CVD+zy
H86W+ojgOtqObgYPcRX7pjlBuMgox23+kcdpvJq5rXfWT1+PPOznqs+G5gl9yhJV5iXjgBCoQTCE
dXfsPrfTlO34MXneHUTiG8uev7Dh4S/svXpPg6RK5GIzeZWVkAdu/NZLZPE43V3V17ThaZFrHn5i
l41MtNazJSTZs5ShmLomLlT63+CWPuOolJSU3ikCvlSnW4j1V2A3uN4+fZdoUrAudyKug9GCVWXq
UJK3zlUUoKn2Nnqz39mf0SOAbp/NefXtUIQ/Mr7uXTPRnHG6Chffm251bqHJFeMH2yR6DqmE7nRg
qyk4HCBIHPRb/528zjldogWD+L7OTXwST7VeGciZHN5RXtt3RwzPnQ8XYUY50AcaerHFo/6VaP1C
8+lENBFQhbGzcUzGX3aYYaGF+n0u3WBzUWgDIEG8eFSJhleI5JFk5T99QNleOavgMqb8gdiFczqh
EL/Lqgk5ZquUTp7R1bJvoQWrU5HqwW6ofta+Tt2olpNj7TxwYIyPGItJjD5tH6dSEiSbMbWMw5Kd
BNhFe9/QsrqoenQFgbtHZdGtGeToMVGVY4wNMW8ZATsEJaqPqCqptkbnpd6t2p8syhHfsqDTa57y
LaTjH+aCNR/pSF6YhLO7mAhD7CMB3D7idMDKeVB2/n7NAlIskge8E0iG9t9Ijh+vrSoFNwQSTyhd
zvrfdhrshm9CsZ8lLUFs9ey+6tBNrlJonfbrvzUVCeyCz6gIR2B1UB0ifLbnPdWPASjULZKONU0C
P0mOpzayW8CiJ1GFAqx3OalFln6qT2UH/ipZYCWO8oyaCbOvhp/VAOCyw9NumZ4DH5dxGS7VyUL+
q9lbBVd3mMH4gMDE8MdF/EnMp0xRETA8RKD3nW2SvU1GypGvls3Z6hq/ZJrmGjUCBtV/UxAzKwl4
Aam551DliB5VeTHzq4sU5+NC6uVIFULu6kbprPk3h0Ncts7PEQUYyLTWtwQ+vaJx3VZmJRwcsV5R
OFoM3XzqlshjINB9adJBESACDaJvt5I2JenXajdOS/pKEA/DnAugM8K6CdiJr5NZrMpdzBH8CYKt
cjHhEBDIdObHJ2NXmh9/jrLb8ZXr1drM4CdzoExFgFqWSbbS/hgB3XOc1nvYx/Dquc8gkexl5+1I
NjHcGPhssIfA0ceTcTuGq1vDMOmiReM6eaMN+GYaPZlMBjEip+RLvTG/PSEj5uWV6RkRvWzGhBML
/N9sHhCQ6mdsLOia7TVA+5DfHGgyFBTdGdOxdPind+P9pnPQxlxdLaAaTjvtxnW7Sw8QbXLGymvb
2CzftHYsgWHN1f+AugDoegTpS1XYYTks6NaziRXKEWDMDhiFSCujtmBlYvHP1OBCrB1PEq7YLbT6
VMSgMstRNo9EgOG3XGquG1XOTB4QG0eWPagGo2iYvTc+qDImnHRN0HY5hjWOab41Sn/E3KeQbWq+
sMcROv1siEgRGk5rm7EjnJFDDOHHmPIn23k3Oj8p9LzsfOQiHDbI6oSWYC/1zfhatqsAk1B4pwxF
vMJpj0VGky/BprfmtL8aIYRoO8+sbEn/KB9gAnjJqjdI9SqtiSd56pjcgEZEkS56iq5foBMa5Qde
a+iIQSHMjZeovvEheT/Zt7pQhYfUWBsstY6F4LHqSAKnQKZbUQ9LzwW/COVq7yk2CamPYqt2cKQA
0O61MJJYUh65eQqVFbObK9c97H1kbhKYTZ6LYM5rg8OTOmWnlpjJMlHKE9eGjP8a2tC6EKnttLRP
WobeFopMkwDuPTnA5MbHlzQW5Rbtv3w9yuTTDi2KqxVvIoDvyUo9reHuKeY0d6JI/VLnrTCsZMX5
TR2MynNwwXYgoQzlx2LULMhgw9I47aCki2xXuh/zAtDNiR0YNB8UvZh7V3yXBWyAZl16bmCgBzfj
byjbCA6ub/5+B0ecl4Z+GiYuGrfnqiPtuPR4wCSO7ty5YT8dxxT7Hj3utsQqNHwkdtWWQaFyCUdO
SvEnLh/CAN7fhm3jHDIcHdtlB0nLD3Nrn0czNOBVphkZc5fTPfLGhjlAsVyOFQHb6buM19pH30sL
hnNDtkkTwfB7+siKN4dA+DQ2CZi23ARd5/o1Lm1B22zLRtS+9yuyhGaBgBnuWTO11ITmOmA1GieT
PxiST6zepNUxA6XM51Zgpyt3X8SHW971U26/hA61Oc5E0dwmtoGpu64jxDCEQ5qGhOMMowKXYaLh
5wLEr3LzGN5BO0cbSUGsL52+BcWWvsUsFIeEtAZfbNIysHT1+Umh27Zdj/QOqgzo9h8ISWqfCA7e
D8jCOkqHFxEAVvV5ziua2GHYmBsNjw2fNM10vItDot63M9IRAH908pcqWYZFwGIEwuSSY+Z+YoJ+
kGMtN/k3pmcMiKKr3p0U7AMhF0T11f8wX4H/l1+jkZ/uI9uz8SUkpdiF5QXiw1sZBNxOfc/oah6B
rHsDLgB6Mot1ceSm4208YaKdNc4Bx+Agm3oezdXSM00gk599vJ9yOcD6kNPoKnFqWjXeLkY7HX29
T4MI2sRBHsEqbSKYZ99Cx93k3KE1PmaiJg9j0Fn2qOB1PTjw2sLwXnTwPDsugQzDuV1J1BMY5RC/
0pQtateLoFRX4v9ENwWY42Y/ehFsKN9pO+avyxcPCxae41iHK9nkQjuey7duVBxEIguMm4gVwILP
p633sLdQcpE3oDo7opa0tvDDFSEusfvpK6HyvqOl0CFn9gpHgqDDOUgeBDehRroCuq/76YWoUpXi
oyqkAIozebRRieKwcKwJOZ9LCGZOXy+wvYaOu8Gg9VORLz4XGsdmYbEqXkqIkSDMdjsp1Kb9Lrwa
2aLTKlEorgZAiBX8dWMjHJlV6ZaWH2lrrK8Amcm6vrpSpjNILSCM4a5OuvBzUS/eCXE2wbVEfBup
Yzpm2L9MU7kbo0816oulC/To99eqJdI4ymmivD5v2zZvESTlAronQTrDJ+3g0KCMJc1lFt6qCmCf
7xuC3eR4bddlM9ibm0lpEzgGbGMnLgy9HwLIzJt4WJB5DznIVsA09vY0P7AUUdYXJozNsRnS2vT9
3cS2JrWvFlWyqRacC0dC/Ex837tq0MIPS+cdBjYyI27Nc8d4Xwh6rv/U4w1T9OBci09jlaXc79Um
eDUj83MQpmv0soxKAOLdOpFRWSznolnuQZi6p4CsUHH/NL9nyoNn01Lr1Mjjcf42kwh7LqzgxRdm
dkuAbzF2S+iwCHaC33QJnE5U4ejnlQpBRAtsJWXGax/hu98wl1xiEYISoPtexyY/FbJ6SCAdS3jd
SQnA2abmyYqpdm+hibvFZB6GkrErDFvWWPH3+VRcPE/RlQMIKtCXGjYJHvV15nqOsT8RjWfgJ5bi
rQcq7XbwCkgOQjUbzMQfmi38cHgGI4jwE+kYpxv4uGXgnsTlKtmpZqFo6+/UCdWKH4aPuwP5oaWw
gRTG6uGP8B65CdPmGtgYaoiY33kAZf50jiQVJ9Bql0lwD8Sd7kG76gf5vetMclLjh1jebzuOXyl8
39SkgRD7br2QeYW7059oUqV3cfY/dCSqPW4W+Va1Llsc7HGq5KP7sBvziEgv57a9nVYYEX6BqI9X
CR6yrg+YVmETprRWfCpYDo4qZwvmUYjY1WRsbHL+pSG8X4QAd0rnzAOglF5jw1jiG9NRQBVkK14w
lROQisMOKJ2MJyEKihubuBxH4Nrk4Ct6A22WCrzNMhXEOKl/W5UDC5HIQ2+qHRBBJ2T1Q8BlSCtV
+ij/KIzzIhSwIrtaTUBXHmgJ8/OPV/a/ZJ8Hvo+QWz+QI1jlYzdVzhRsrCdOAjftmJdu7SXSaRfs
rkEZiitnooo6A9YlzxOK6hfT69s1vrnGN+tfdAxPd6OMqU253vlxFNUuDw5zd/LwlAFd1irG/PYK
45uuEa0MV3RYS/8EZyaU5llcXqvG3m7MY3Zrp615rWTs0rXkimQi2yQQ4bnqc1ghVgch8D8WacwU
20q7WiIMwYJTXbEH4zyEOwBGDsrY2Gd2lj1s1K+pQwCkwwFyyGZ0Xq6oGgzLN5uqYA9VEuDFYYlh
2bvkT/DU4UXrRjDa5EMeX8IPS80aBSsSom3J/5YiE0arRnWXPOAmZKuQ0L/u6BozDkuZmmP2fo3+
NdL1a9IBZGSAVE2dSNFFy1tG/AhljCUoSaZtafSjbi3jRHbnsiySThRiqzl6giDF46d4HUXV3KAV
WavN1/5F+8ifleB15zwP4n4V1yRkKp+lsxnEXZUb0Z1e8D+KYLJd0QqBPxjlEEGf3rxRymIg5Mco
52dz7BiagkHWBlJ78nkBGqWLjZYTOFbSxNBzZJ0kIdG6l0HqXpYFlgRpq4mBNuQkE9ilaqPXNeTx
YR84QI4yDXvQ/yiAj04RY6PSjEm7YVKjrE4/IAIhYotjz/BElRKVpG8fP+93Roem9eycncP/vEDc
DnrjAGmp4ImZ4gqYFE8jGWO05JuRCD8Y/+e7yjpRfTBivWU7Ja0gsSv0zABq/oYhVEXc4h8vetwW
mdiCEAm6Ik2fSicSWJcxuz2cMkBZ2ZWKbfRMljFd4XzGEMXTi+9cj47sSg7t8jI5ae+EOjUTrLYK
IYw7OYp37xskYVl+edJx5oY9gGvmIbjkLXwe/IB0sUFpfEItnomGPirCFiMsXGBw0Ep6U5jb6Uca
ZfamZu2d+8b5YTteosyhXDJZkLAeheLqlNNIiwJer95Wi8ijgg+Kn0QJurl3hz/G2yof601AJ4iE
SvfCu2aSix2z/G2Jwlcc3WpSX1cZlPfkdk7swuHxvvvfKDMqmicOAgVnrSYOEvCmm7sZWzPsklul
vVRA/QNeVuEcCU76ht6QdD6xpYBX2Q6R1OgJVLizROUml1R/MOhKy1kXariJZrnn3oSTL6/ZUoQF
L1YHG6Soi8wEdFPu9GIX12pb/pOLh2ST4f9CCt2ZvBK0kxZnW1GeaHf356C8TICriYTzz0F01l2I
qAMdt3GcoNS/UpdnOsIdhDJZv5uVzMNsbYocrvLpDDd1LiGQSaoAfHj3u33cipp7zB2FuyIkBepC
/tx5SaFL3zMkBJMR7r76rAIQI7+2N1o/Q8pnVBCbnNtvVSm7/ZoB1umfVuhAfRvaSoDANfSLqiUq
n8jzlkZkdx79WFaVa/Ut9rq222pdHIgrY/x25asPTtYvJ3KhFT8VSmVwC+d4drAgVQszJnvMZNlc
QcP7wCm968PINZ2ZQa+fwHBC6QZ3iEAD+nrVda8BLwEDV9xf2GV/pIluTgEH8KGCI9Se2OYsy9k/
5dYavyOVHo5Uj7uwoWWVA/KwvXJd4YYPcZzmkRaktTPsA6odLdNdqNAhHlhprcjwPSus770N7VOV
ySGb5CeUSukZrkyonLuBdKIO2eP7DLm79Af8pxdGQMMRlfkJd100dMTYmTCNvtIGwLdW+35i3onT
tLeGkHPeEz24FiXeicbWQtfogOHPrvnYUNin5ZLzChXv/drS3Dbl+jhmpyXTQ6EaCOhZQ9DN+NYd
FtTdPaXrP58AFt90Z/79f6x5cP70pO7yYP3qWB42xC8Sf6eHH8t1Rqi2MEah7aPz4XHS0WhxtdQa
5pNyLCQxp9uItHyOzgaLUuS33G6mBoDNQS1yQYmKRQwGnGOHYKvOd9sCGCLIEHfCt3fOR2E8d3GV
EsM4su25eyzom4odFLww6eEU9NxW7z0ROeFQgNf0a8nMjJEN8Kx8Ujin/cWqYXrc8axpeQQ98EYd
gU6q6Hsm2otiNCFF3cAf8zNqWJ1esNpfpTwkJjFFbKkq9vE8kP1U1ZS380q8TgdyDxeEpPyj9dJq
nBAmQO6dZkBjSoB8JLksXqMbbfjJWVZgsARJG+ltA49SctHQKqx4+v7kEgzQwFhzdcUNJySUg6Tl
hvWdCHgx6N+jYl1Oc1QlwM923gj7MOLXRaE1syhIAIfgxgrVT6NrdT6yfpv/UMc4pOGsGBrjHDb5
a4gY8lBYOZuSjiytMQDVisiSwYu8NlliJ1d/L72sAh5AV1Ne/TZbPwhVdQm+8gybM+VRoEvA+qj5
a8koumDAdGKZp/Bx5yLYP1K7ghHuT0ntaJcIuaz4yzdBgjNqDKoL0Es986tf/APMf+UUB4dcP9UM
YtAkHJiZIDxFmReGW96iHyjfx4q2Rj7ufFG+YtOYarK4B55VKL1lxwRVstu1Ta1Wg/Y0v72Ghtph
GEkCfM27BpNViplS/lZPAfZDMgBjdNdOsoRFT9PBlrCAUvFTVHXHKQ0/xGTxYe3+AhJshUYFFxZa
jvUSggoUvcJaiFzSyXyfMBb+w1IAY3Wrswgtuzw1pGSNN4dlsiYr+u9BSJeWqpyCr3w0EbrJZRqb
idAAo5w6ye4Wb27u+azpbXmDBx6SZT7d3JlfsfnoKi+n3YNFAFP8Hv4eO8Az7m9DDGGXqDiY1sVj
Y4+MCWCZW9kUJmuJk8PLQnnlHj7sVHHjJX73W86zO0yK5WP9ANHNq4W2T804y42q657F1rgot9+5
1X2gGs5CVy99XMKRkY4/Fcl8EYd92Of+xsSdIt3dUnh4njTID/P9S6gsJTrUYl/IvPiqfl0pOspk
lgl1RNVRkGEp5cMNEUpP9iM3fdf8OZTikJkSg8Yyv7kxdMBfPVl+hu1isZEdyGUXE7xiloBv+NFu
rAC4L6ycVmVDWBnFNGLBN6MO5JrfZ9kI3ScENoHR6Ku/J1IGHWJb9u42C6VvO6FVhbNonojAXEZ+
2djo3eYpBt+aw8svzycsxGHxcHJGkoZWoxyLmHTm7m2Qq0bLypm0KhIwF2obiJZ9hNtRjcorhlNF
jhcJlF6nE0xdvrTVsvVVP/CN7T2ILKPSy8XtPQmzPWGOZH7F9X8Fng/Z+URE8oYnE95tp0BYcDoH
GyothnQgD1zifHTio8SH3ZcnEn2k35QpsVd0+H7ua7El/njNC44qFTvHPFrJGkzo5qE6yvjthmSD
bNiGH6ika9IJGeqkLpOybbWX1P/k0K5x2CzVkod5z4oBEEIWeMAOpUq2La/DOomF77cRmdGf8mrv
qnY1vGarxBVJ98xkPZCMeHHzS4+tIdY4WihsbJ1zr1aoX/iViQJDe6luc6T9UbDuX6a0YowlWnhb
8nIW9FBjTutUs4p767LDkjAg0/amtfJY9K5muhfLjyQ/jjnJIlO8CVzIwYirnmyQSbejIEzwv7wp
SvjAVOlVwM5E8b2N5fGOzXHqLHgb9wKOe1cNIMIXqQpZDZbWCymAaxzYkJlOs096oGrPtWFfhszB
MFJl1OH7R8is8oQWV5FnV0hhEw8dlNjORoshCCQPW8APiAFAGw3qaI+DN7ibTEnf7r1fFWjTzvF5
ScdUUbSUQCiqf+YIlsrSE88976OQer2xZ2nlLgPdHFBs3D74Ci4F/38GuRkKoblSrM2GV7fvkD+9
CDlK+dxCP3+R/8KdFf61l0SsTvW27aIwkWvw7+cwQW9LOBkvpFYl9aHpd4klR7PmAgJ0aT0g3sn+
mXRZNJgIffGRdiCO1zMxS/ZCU9DztFc1aKaUsjACnbAcNf1Y+ygKN0BQt6re9W4iZT4+wCclWu99
GIC8hY/rCbwL/oKDjRlG7ItPTuIUpz6SlhCjQCcb+mm8aG/N9EAOWEWWs7mgzU/1f6HzMR3h4jOA
V6+eQcnBNTit6xyonJ5k+0OWQV6l9/qO2iAcZcTdBqk9pufMNacVYm50LBgtn+lX4XiVnGhOJZ/q
EkI3Uic9O6V2JSBsdEAdBZsjftQEvP/x7v/h231pi42hz9UIuHjOWPiDiX04nKhjaqz7H6MFKIZr
aAiEqhHL4QSdc0iZSRXo/zjpsB7rFsuuVCwYVp/3UaTviw4foa/LYfIC3BQ4Uqv19NzMLHlnPoVr
/aWL7oJetCTxXubCmMVYj7qoljhaaTnRQNQ+imYSyp1NbwgkwAJXmF0yABB0AhroiC1SMYeoVcIr
lnUKkZr1OmTX0cpKF4EECiOeaf4d4b++1zb6cz5VG0ymme3Nl7m8C3q/38tWvJdbJm98NowEtXMm
/ZpsKRCnEoDG8fIaDxpTBKq4UHXs4n0f/UoGxaYHsmyDUSoDP730rvsOQZldlcm7e3eFpPuxrbs2
7UCsSHcILYkrkRe1CTOmlkOR7A1MEQmuRy38oZMi2yq2qbcx8jY0yRmiAV4TsCeMq7vhRVE8EsyY
LArJ8KYsWJOzazYszj7C3R1zUh8ZXqdVEPH2rKH8dTtK7M9KvO1V6PQUTTx+F7ge2RaYKFX8Xl6D
jtXmQfQEq5jytnVy65lP+tCbvrZF6hEUgyVQ1zq++1pb1cJtPsgbsOPCTcNqYZke2unAZnazlUjM
iX0KHiTk185USV+W/TA8mDCfA0wRNXTLUAqZwMfurnNOOMh1jPT+FRQpELIa2q97O8j32SX0VlC5
ajdq1ecrXKG/JfJNW9NCgdJ7GjA9wMQDqOSCTwToJGnXJXIlNI7T6bfk/FcM4hUFXpcnixci33UB
tLP6xQrvRLkBFiKoHTNCSEkO7Cl4IJrr/78BqjQ7puSXho0OuGssVxFGKNvszwOVAmF014SlMDVq
GIjjTDbaMCdyc6dpCzK/yowPzHsLjrWraHmN7pX6e/cjP+aF71WsRXNOJd7EPKdYjgRCHDKLLaQv
2InInQhsK3l035o91py2Yr9zzI+3rMZYWsCefZQGs6xqBn+TG6PV6V3QV+xQ+7Oec7vTGj74nw6T
ZX3x2yQVOKqNyak525KdYXkxMTcL7ZUlxoXSo9PHRUrAzP2PSlAMEeUA4BwqfVHjJVBK2zPvqoR9
NcAJFdyNMWv//a/Q3Ej4WTsVozc7nHaLKfwjRPufkJo7u087QUq3PXpcMGVF4cPFjkKBykvrgEI4
nFvvfOFcnBmED0eEPQMVaFIT0uiQKzHEKCD+qV0RMB/47E6TwUexCjHCj6EUa6nl58lZEOGzuRtv
PyfxEvU0uy5K1mM0/Y1ERAuNPYgTsr80D3lWHA02WSiUdbe32bObzHRZVYwD2G26P6rq84+Tto4I
AIA/GNJvEDmDT5xqPhLZQvBOEOJc33bCL6YnYF7wHRagBUR8xk74Wgeh1TAa4Vx77lSngZlx6ENm
+VwufNLowK9I2G0+lK4rxvVlCjfQEoGcVQu4eKQP8sainF16hl3IUlFNpia1S4inwnpQgI1VEdSm
OVY4WHK5I8doNN6v5/t9T1aHfdmgUxeHtInlBCwFkunzb3vCHlFwc5i5zvh8dPTQFBirhTFjr2o7
Gj3cu9BBCIZIs3ewmSEHjCq23dMkM6FjQEa/3Kv0ghMVinQ/nxA5qdR6pbA7ejUOqR33UukiHRop
3zmKnVWDe5SlxwPfsabAKNHqaGOKF0Xl2vgYUP8zSgDC9/g9R+lGP/bKvbNYO4w9qJC6C7RP5E6R
EkAR2XAstmO3sii+q2V2yy82ZEegcvu6Pyk5eRJ5JgyNn8h8yIuA5+DMN9viYM6pthPewJTog7p3
5oJvYpNiBRTH41reUOrWwbnOl2nyyH5tfr4LA8BITARMcN40LBM83bGc/sHWne1Wkv8osSV0lTq7
WQ2Aa+mxuK8JsWLxltCO7xgwi+tcfym730j/Pu7cqldvyAPKorqrxPMtQh7uDRwZozpLG4eAq7OH
5v4WlzSoaQhaMS9T3GoZ6oxzMjGN8zj0JOF0itEcNeIpCOn1o+nQFT4SkEAqWIDgYV3cJVJZp6CE
2EmW5ZF4ajHSV7PAhJ0FNXNqo/H6iKGPC/lN8FRb5rcE9/OQSXCtjZUq9BQNtleNfzzfXd4xtINv
Ki3feKRf59RFsy+AUlq8/KO7bwXgzDRFg8LYIpX1eh/my0Z7KcfO4FfgqhwBCZMMHh3KlBYp/ZrY
jEI5NmO+l4G5rVgyGCzS9Y6uB/+eRcL209LiwXVxOyyiH0x9809gqAW5uMSw0vzsTwavYyF6SSH2
eIoUpc1JGj9HhlZo1t7LKAhsIe8eQTOGm0qwBAdhc5fhUSzNLqeJvOr1jYbK/4SBpkTkWZPg4JG1
8mptAxJ67qXnlv3VlAEuZ8WFRX9Ym8fRp+p++vopWwUvyncWbjkdMVjMLwa8z09zYXb7/k/nI2ek
oRX3FmlN1SR2M8Yax2TaxTiqzLT8he9AULcPAxxsvr4ZPMIdlfAMYN9Twn5ynQ8mxIYQX7TfQWQ8
X44NPjEuiNyGVpuTgPw0xgJDsd+dELx+1yINZ1cCYUoTY4eFUet4Qetaswsv814rOYhiRtmwQZ9S
3Xt83Ggbs+a301W2ERGoYmJQ8O4bnlt5eCreU5k/U4z0beoTiDRezvssl3UgBrVZt2iHoJp5vNMl
b5kgT3ZHNqcCBKIBnkYRj6q1hycwo0ucJEPkdbQ/dka6voQ7Jrld3u305r8BaGB/v5ttSnY+k6mR
C+peRe9WyBvh8f6tjz8A9mSoMjp0/H7zHGniKw+E170LLS8/aN2q2X17uJ0Kwmev/wP5vuyCbvb7
wXljHtwC0mRPe+twv2UnXPMOQJUeKxl/XlPdJVNJzgvDZT0DAr0Q/+tkOk7LmhWuCNXMrS+TFfrM
Etn+8PFrBhQe99Z4+QFGaePaeDxIz4vnVHz1ghQb4R+b4Cz1q2syqcx27ccQQJaxFKEsYC3NSA2D
QBY/Qj+jVtS2ePPAP9eBbKJgoMA6QSPm6pJofIsMl7Tjqt6PErQ3flPHKJ/0i0RL1SQcTqUnMzz5
h3xoF373Y0yWzRcDXiNnPPvc8JMx3nMvBFHS/SK7420E2ovMudb2uMgbTMuzhQjU+ySevmZD676P
1v+knRydvx2Bz/Md3npU+IBEfr9bwBAj5fc4PrOWHd+owXtEM03gBP1XakZdb7Qa7iosFT+2HcEW
hCE3g9O+rtgHJQV7X7/8YJBoydqzM3OlMhxzVieLQ/TNfPqQedL/V0ncN0htcAY3V1p6k/BTYTFj
r2HCqzuNYRGtXruBVTcRRHRbP+i3kwNGJxRPkGo+Wdlvnf8kOz3jX6TUq9OovvgfixWg3/mpMews
B1KOJvPGW35crsVFCjV4NLRNwRHvydSlaXjbkcQFaAT4m1oRk3+jtwQSM93f0d56EWkNDr/EISQ5
y9eg/6lyqi4XrY00kNDT7zUuAmbzKFXBFLHLFVHGP7+Wvt9iunodZtkwo+m4HE/efU9OrxU+9HmU
9MYdNxKxgmygVH8cRGz4lu/EF7cgvqQvT5t6FQXxRWyo5CaNgWoupSGMSF2lbDLwrDoXPob5Iblh
YL5aoGRgZY8RfhRYhVe3HVaA2kCmnKr4amWrM8janXDHoTdZOayFDCcwf1qAwmvMwSWpYjrCK23J
yA4ruqhf4yCKyF0fdzyTKKDb49jcfgBw2bmYkS0RALLy++hMqu/7StsFYhxg2YdE08Xdq2W9kfcc
1Yz5wfwkem618+w05BTOLQDHMeYL0Nd/Ft+9YNOfrh3C0XfTeBKJSz+rOiqd8bR/7r1dJ1nWzvaH
PDTyHYFow+tFKoLVL2lbeeQ1tf7nt8y6KlIcyRgtGp8LvsWI9/oEgnBlbFoQZNvdPJzhMgeswhwJ
mKk83IW/yuB2ZqHQAQWIiZ4+cXOJIGAXzLvL7TGTnJzRNXtOaFVH3m/K4qJ8uVNMUVwP9h6uycmW
0bzgNrl4xcmxnFd0DZkIxzaXJDPAzRHOWMeTrZd0gNORjtQl6YESHqer6bQl2jgXpEFyjMPkmm9Z
eDw04xAmWqMMMLLiKf4S/wiZFWEet/g+7ki7C5NvA3O7jjbvvkRkhgt4V7Trf7WPPTYCgU71Sn13
WH3PjoUMwJynud1v2ZbN3n3zIH3m5r6CUbeyV2oZ9Y/cGVKRC1GMbrlOYVIO2RtRPoIQj4rHAz/K
lIVJ+BgkJ9JunPpTK5gi7r3oGXF2Rsinnf8Od97WM3pUdthM2RPluijhBEh5UwznkpBxYdawtmPj
nDeemtAs+Fwbz7GTWS0RmC5WFpb7Dv98mqzMiiJUvyXrs0aFa337Th7+KUKUNJVba2u0SKw/tOMx
/I8rO4IMidmzGPQBzJVLbhd9bAtdos8kWOxZdGscq5exbm9+cf3/x9RupGY1kxuGZ+IJyTt+luKI
yq5N8r0vJHs3MIzX0f8h77iY4MXf9PzLg353BE+pM4lmeiG5BnX4o5sQwmXDjf9holPdvegv4lZy
Lx+zYmoke4ypLNKKhNBB+bwipuvgY2RSs9hAGQocqBMzpBoIrk0p3D4Bew/nEWIundFEGYMvPp2C
ATvTnuhhrQU1rNpRw387kpxpTPwK2+4UW91SH1Py/XPk5SspCeTFe/ZCPn7YeOvwA1SJBD1D3Fbe
A5HE1Wflj7VEH9QEKuAQisVQ68UDOvSQ+IWU7VnQ6P768uH8YckExilAwR9qMWvnPtYj2L+ebYpU
zAqCNOtjCj69rQ5sCcNxLq500zfGavTt6PpQhpKQfQaYNKn9uBmjr072f23du9xI7fiooYqn/TUY
huJaMjRf9vn8p1A/7TNMu/Jq0O+vbV+Hh7n6/nPfON1AOTT635V5agTRYHeBJqyLXVOUklMieB0u
W8iqYjvJXXbDv9lwFZrUJZ2Joig2yPbzwPnqk3A/6qcZk1tRehQuMyTqnxpDSBBV/eIn7jPMFHJS
MDW8OSrXucpuKGVnQMs8EPSG7Wmudlw8I1a0pZ1ycRN6PKU56DfJmoy+IGQd9E/t0sERXCnyG1Aq
fCJJVvxfbt4lwUfamcb4ZUhlxWnsLr2cDx87woHNoWIyG9wisWJxtIQ4OMOUrBE8M1EkTmeADTOg
EObX2kWng8tfx2EU0bFDKSfFWmWvH/rStDe9otUfeRApXGmNd6pN/LqUbpAsxcc3Wrc2LeXs7vFo
n4TBReiTH3su3GWEOkohGFnR3vsSAR5ZDS9plQbK3mzPHP3pZO1tFHX0cSxZTYQYKi7nWFCWNtDl
+xBAkp/u8UY6LoQA205BYCqRQhCkN7/CEcc/GGy4G8FWDTLIDEjbvFJiAvVjpYm+jQXNE/iF2pwi
Snd1YSkcL4LDu9N1j3kve1Zh3gD/0nrw88Zttg7WP07axDoLHp46b7wBicXYr58Hbc/h5yMjfFys
cACM/ErWa6cYmlqL3lT0ZR6PUECXmyBQbVBHMJU9SX0Sj2q6sL1XADQKCISRgb3d7tB8tFlecrVw
KfnnUQDo4ispf+ZpaH45Metr27CiyyJuI2hpHaF9jnvdYgNsEbNibF7C/JR1Dr8WnBlN3c3qT7/V
Tux5H2dxLv2yiVXpr1J4YZWdh1FNbiIY+Q4gOKQbkkm9ezWoH6rzPiGKYvnPygc82RC0/uHkmlDY
FQxqZdoHgyWtxDVo2IaAKSVXu2srJ5/FAW6UJD389HaNI30Wkgia3iheL0+UarvbI2bd7IkG6gfS
27aDkQnnXa8rHXxwHFouCz/vMQhVXxciiET6BYgut8N8BatpqEK6PMnaeBC0kFX1p59sqxPYaeXR
juhQ8ejr1cVHT2K4CwKo3NfII2zVbkQ0b5nCjxxqH+5z9RrmO/uXS0fODGnUbBt+OYX3jBMLG3BM
nvGUPE5VY8OCuis3VeqylCiGKM4E/W7zXGlzqXzvpEdMFKkAGX4Y//yp08PRAVVe2XhPzAtT81jJ
RAR/yWFa6//uABO+AVY9UHhHGhWhrCTaBc6YcDORjg96N6/HF/gNfOThEIZivmtJuHxMwN0km4AR
wL3TUulMUDgweP6Ube5Ln2WZChPCg6dBVgcSJyCdnc04nXND4gzLX4AkDJiJjSTq/G0e5yzYH+Uj
c2hfynU7QNSOxvzww84B7cerh+mD58U9W11UBmMyVTLuVlkJWUWswcjpRFsiDouwT96URFSZiRjn
liS19ryq4wqy+7ScHPreEGLxN5bZFXhpLLH/0RCRjhQOxSro30cBmQFJy+l1FePOQSzhawba09Zw
FUxbf6jd7Mo8+S5K4T8BH4MY+bdlu2HaW3nCb41MhzZYhaQpXsxnwxKrYUn8DgMaJJzlukv17fZw
M3rN3ocpWQUOz0rnuVTqHQUSsBihCLayxh1eonm4v51vMJHcuTIpPgOz0vc87ofzju3VcIIrJOYV
9H/37Ou9VoCp7VHd+QIy/80OvoMlqoXi+XXoGxGEfkIVmpzBm3LlbfRgfvJNJXqQBTLJ/dfGeT1w
9MQKRUFd0k3Ur2OqptyH6AoQ8pJDDym1xjFPPHoStENnTeiZ5eY3ca7unKmbZRR5mi9xlybYb3+7
ghprc5rH4fCMI+Pl9tzRV0WcLcHwuOD32Yxc5Ju/7S1Sp6H4o8rC8fs8rZRWoZPllAO2BHXY53Wk
5bb2O6ujXpzJTm9wXbCuoFeQrf6oP7UWae5RLD+44CTGB7NobbV0QjuCapyx9rx2PA/N5fNe3y+l
pHiwY7trPWhAlD48+sSGdLv+yAnEF7bB4NSbvNB1nnVJu3SY4WHALbxoam0+diijXjaRc4tVHKIC
vI9VwXX5vZm/pcpDhXJVhWoLHEIi4MlprBV/mri1xMo5pvBjP1GBmFu8TKosB3slKnmvdxaZQi+g
FBJtVT9u39JSW9d33ZK2sCQpqOZ1JMX8qluxaU5hLTycs1wbLyG50L3lObcHeUNn8RexrVL0niqN
d1PdeA5yw4z0hUT0E6oAxrDnubhoQe1cuL4eMOLPnsH34gSUNccjHIp66S6mW7VlToPtzygdithq
rpqrFFqssq7IXL23IbB4iz8P0NHA+wUV5DvVoWO2hUnN/e1cohRLyxDP8ilhYYWV/dRXJcowChr2
tHe5fOL29vmWmuWI/XOfcBMX5wiovmB9NvuZGFnm2jfUkfBvcr5ml44uP0VwfuEaG9WxklTWzfIN
hppSigUEPm+BKgg93v+QpvbTLlQOFjq+zozof1Km1W4DdDxuP4TjlLLK1EnJFVyIzvXQWbH8DmE6
JUpIzfD0FiUcPM3f6t68AjCD3wNx2GBRjocRkS022opG9gkd6OC/OlNvnAv6x8ew82ycDO8QRMrq
L1jWThfUeXYerQ3HDSYA796BKpxXYJgZk2+TL8Y27ZD0o6Ftara0QbgWeKEelqq4kAFq0PwBEpWA
bdJJWD/MXBTNTWvOlhXod+ANcm8oleQ74WUQKXtvoMZL4hCKvv30Pv5LkxLVthNnDweT6LkTXCpa
jSKNTcOk6XdWr5Cb+JidIlGGbRo0xVHKUqKfkXWuhVVdAc+rx2idancTGSv+LILHI2RqzOl/O8pL
mueFsapw2nnJD6Z8EfX4a/VZMKjP0Sh8P7YMxWUEM5qld6RhPIaEckmJ/s6H8TGpFySK/M4YdOT2
euqPnf7UxSx4fr4yjki2pvQUpLmDIFaDQAS5I+/4cOm9cLlHB1IE+GRymfj+Qr69hzXTy7lQ+uLh
ztKcls+CemPDooM4noj1DLET27Pb+ZiYiTKRregRLPmdx6wDg4JfbCes6p0l+Ji/t/ZmHbj2amTQ
URiNvfCs9U+Mz2Fw4BAlzHNab+E7Nom7PJHpNErr8Y+xW6dkil8nvN3J/KA6JdochlNgaP1dMWGR
B/dOozvXFaWbCFoyCkx9VYKD+c4LuuieEhuaaA6kUclfNiVpkexHjqrSKNajaUy/MgVLFJWgJEbE
MUCFnELlT4+NhdX+StqY+5dAnwew+5bwPmfkdfyjZP4uc3Q2X8j+5q+X7yuwTi0j834cZpPYM0cc
faXEaM0v8Haf4DBrzk6lrwAdeqctU5/9vTixe/msgIv7mU9Lm5ETKKjTIoSwWleq06xpvr8tMKMe
Vwh1pqpMMLr3RXucGYFjtyM3re0lNkCx9lUtlqB1WIbBf+iFyREBdlw16MmyJmGTKXpzFZ0umzx9
AKwkxIQSo11gLJ2hE7b+uxnrcbMwXGL27g+NBVA6tGi4Pu4AMOGr0c8k+S6I+iD7IvgHRKH4fAUP
a3orVuJ6JUKuaNFQfn4rDpDvQZGQJCQD1HzeOZn0sHDAm9PYtmPnMRlltmvVPG2jnimT5poGISW+
hIXNejeFH1bpWR/rEj1PX6hInlDaV/32JlxOGDAKloZ/hU4G/MiT+MJqdduJgNtqoFV6oJZe9413
BDhCPQwTGRvB2w9/Rmu6FiDEv2ttSqiZNSr8AUMIuPgGr4y8FWZ1JkUH7IS6wn0LJeQ9Xde/rmkC
NIdRPfOUCr1L69K4kHgcMlXnzbl25Oer9YUUsk8DMojcGMrJvJZWThIt5J55wg1Pqcp/RGJRAlg/
jf5zAiH8wCyXiEUaZUIj3V+fA7havNAh3JaS2djYVLKbYonRyuhHoqKg+tIeHx5/8ATijBgc/84K
4JxPqrlsnyzek1glUHxhCZn9Ivs37tNm+1tAwhpOA0Kgo71d6GcxBt+oDV+OSbwbR6TNw4eIjQoK
f1+aA/NORbHm2h3sVwJZk6DCJCRifOZiF4uFs+dSsSHqTkdcNLC9xuFcl9fFSAVAoJm/RWVmZPqA
Hs/w/m3hFPwAuSyj8dm2R8OGlpWu5fAP1nxD6NJY76UnVwPZZFxQe0qCgX2I6pscEVbpFg/xDDnx
fGXLNgxDRPCYfq8lVWR4zchBvPPdsuHc+umsWX3ke/gPoyw/ohWaYivey6EooV//TnHoZDPDHcU9
/b5ISwEFB6D8U/SCwV7pPVfwsHMJhKZp+gzjGZs0uUkejtWeWCYi6Lq1Kqpr23h74HGbNaNuhiO3
SKirfpmGz9n5uaJnazaj4Bp8LvuiOXqCaBwWsDPJHMIvXGYRAt4Z9BjOA1RvR+qjAjAK+/0A73Vo
5TwPUGhRFNJY84ZwaAizslKcNvOBHPmu/1HCF0Zg1E8ANF+fGTiNl3UFKLuDSUVWmpOPXFv+Lx55
hnJlu/1DkvF7TwSq+yqUZCaEApDbB1epE/IQm2XPbhSeMni3HpaaSUJbeXJ8uzBeDps97LnfUBJS
oaLC5gUwnhe8XevSleWU38DcjNRS3bnt/U1GH7y3KGbJottttK0NmXI3+d55QkzqDAzxqC4sVUB/
Kk1+5ph2x98y47F5GYrFI7egcrcZhPyiit1EjVqQbJ2KYW0OxBRCN+x5mpa5SwxjyAUvnpd+08ls
NS8tLryfQdeoaOVyeKXPbO+StmQe/TVHWoWf54rHQQVfJKONWuEAHZMMU9Q04R5Tr/SD2UThIGqD
t9jghImPhZgFxOk07hFHzlO2beJgCtMF1BN6nLPi76TTztRmjyQLYmXpPsG9mGMcRUmc3U7pnh2x
u/hr2yKMNAorttUPMo10EztkOwKBDEjjvDFntmfVucs1bFGiJx3lUmLICXCXCkaND+Jc3I5zY2EC
Qp3JGT5bE+Bv48Vnzfv14cbUhcEbqfEQZKIa8plV7T0bmP6/oTZfF/+KGNg6sRIQD2TgK3qHlZ75
peluihPMxBRHXDvr7J5cg9C5IkDUFfQPtT31ki2gWTdcHjb0fjAnqaCA0CymCQGFZwpApTFg1Ecs
r7d6hGprrKBXq1LJ4h7UH7oTsZaPWvTCoWU/MFgvu0wOcQ5tfMPOQp6+hcV27os3R/wgMkQqTRel
d9gV8iFoaZ8Xqb0G814a9lvHggBmsrpWRYT/3256Uw3JzyBKb0HR45hlTY0sveoXBPBnZJAXCT5j
hdk8WM4L6zkUEttMIClumpxuxVSUNX00/qEanJQnYQZaffb0L3eClGdUKMNgu+o68H6tj7X7R6EW
oJFJOo8giL6fHFKpB9LsLN9EesX9Clp6MSPODXWEHF3gca4fX+eMY/GxXGLs+wjfE0F5ujt1+Fhu
zCVpyCkUiapWslxfiVk0wG62nKqFmZa8jTrNpMUD6FEZ+jZEEMApBo35pNmqF8oHPRq/caegYsDR
0ebds55ahEJlZmCH6rE3/+JaafI2UkMHAqSvIo/H1j1JsdFfcBPHUpiJUUQVINJLzbyOaO/6YlNT
Hdf9sAv6t58wsajpWooyRpTBvQu5OncRX9sV0IMkrDYgMqBcMS7Igo5fG7NuPA71S5BPKBZSR06t
Y/Ztlmn6KybO9sXaNqNz3ySNFHkjLp5HJN9gJJlyh5LczjGAAylY3ukRfzz5Px3DxuBrK57zm3YC
GasaGUVItj/o2v4IwCQRf6R4y7llN6m0U/S66VJaUIWqOxKv/brQQ6mWdQCVLs3B4CjPv7vl8Zm1
OIRmD06qXcCwu9c2IXCGtcbNitjgayJ0f5mxgBMSsCLOm5gu8d4COjXEn/BytsSpHSPofYtTRGGO
0IC4aGnKeGuOzJ260359bQPRJFjlLPqnKbYgHLWd3t3ZwWZlMiDjJ7BD0kOty7MQOPMuSN6SCvGd
xBfkZD2GG05NjZ3srLOVmaQdE/0+9ZTRWu0Hj5yOSnaRoo0Aw7430o3F/BJq/ejsBTbbG8uJLITE
QFVK7HEMLP6bxvqpABp5zMGRv3WHmaz+hdpSURUWtgRcVXr49DdtEJeFslWRA5PmKIlvp2OgRi9a
jV7eLvFUsYTACXOKbYc4GegwlO8C0BVdcPsg7dDWD/2ddmXkxbX9dgYi2GgU6XvJLj01xqTIll17
okW6wRyRFrXayh2MDEC37PIBKDAWAlSTIFSJ28Si+OYyVfXBA1c8L+olN5eAa3LbLRQqMz/uBA8H
LQ7RnqRjCbc8NWLypzQDkxq442EicP7i2T39yP5u+2q1rin/ybNHJp1aw9oD4sXZg+bS1rl+YuW5
P3DIYbrCyKm1Y3VtZoTcfxMpc+5IjuLdJtXH6T/TTZCy2RArBRKaOq64d/fw5HVChlA4/fkJcNCf
9FFM7BnDmYPBcgANs27ZzQpwAVZArOcOW49I5ex5yOch+KiLIf7BaozsbXXDwhKcerqa88Q/1TDB
uHI3GItFKRhiHjD0Xc8tCDRzmHISo8mqfmjqUti6LGP3h0dvqwQXqAxYwSwCW03JbAoZdhLHOE6M
qsXCed2cH4zHPW1OQOj0xtv5yM3LCA/IQPpAMkI2W/vkTQMXiJb23KmaGNVW84nII44qXCo9lp2W
9vP6uIfUCfnpTRjO+ggYfLHmD0NgHqJSVDAtXWyqqW4jOMVKg+IHe8+GSdjIT8ypAqbSCSFhXyiZ
Dfk1nl3GP9M4YICwmlYJS8CsSD2Desfj9nVoEucrbeZOU5cBXoFxZAiJoJfxyoe3gP66GR6eJlXD
l2ovYHh9lNlFup1eC5QIx+Nt0UIW4ei3TZZGI6UilvvRiO+75+kpoMuWpNy9UpalR2/uNbycHPmq
H01qSIdkszWnn8cE9+rnlHf0WpdMPY0T5hSx5oiUwrN6O1b1sO5S9NkqCOufZ3//h3Eoz8lTPOzS
smLJp1oGIVMB8OvYuviRyBTUNEmGQtXDhFf5L5zZAW8ZyLoYo7iR73n0uwUmSpz8s8DPast8LTE1
0THD1YhYs44CYBBeyIBQCG+eTmZvSKsn6rjK9w0zoNY4miidKeGc5zaF8z4HslTAsawwISFDI+CZ
tZnvK3/KJSdMHKTwv+I1IjV+OcWtgsVtZu5ZiDaBrDNmTNiGkMP/xx14b/Swic1eqkvaBXpY1ksk
2G0KJWzPaj8Fn2EVcopEhahOKCS3nK4IaNJxrKJtPLLxc5lm6c3fvyaEjMzUdJRnsh9Fj4DCiPQH
QQJWuutR/mf+HXEt6gIHoX+3qyWZ/zgoSCox1HlAlXb5IJ2TsfIMAjVC+cSchinH+wLqPW7x2EmN
Z9aS64NLlZoMwyzvUEPfZUuxqHlBVRHGkQQJ4mA6YeqALgl50NrHr4Pat5TKV8o9N0QMBEwpLAAg
+OwESOhKjdKUCuB8bIcxuVEvBx+seZZCHaIwSSlxbaKiHjeE0ndGMqy4fUUUctwZXc+Y8HU6xYvk
y56TwTbPv5/eAAxT+V2Qbz7qhfX0QOgDuJ10i5MX5uaJLkTMIzgLX8+4b5pVmGwixTY+BWL4AvpF
Xnje4NIWAMaZWR3lOEs1qt3k5Rk/ZlGHLegYvUmbxg3lI1OpZTrfvh7nau5v7EMa/MVHdjgWyGWI
tY0Jqz/vrk5zisdIej7HE7dDT8N+JyQoYbrzBIVloAZS0BVn1WEHyLVJtq36fweHK4+4azAVXijZ
Vup3Bk5kh//lk9fIsl6jXpXJrPTpT/j+XQSEUOW+V34moD1wHnd9cj1nJ7+0TB9Do4KAV03m5WBl
OhIYUiJ+uZJFl7qE3Xkqq0/BfxB7qxzZHo7ISN89YQs822RYoJ9L7hiUN6eYuRexEXJ/d/0biSRw
UM3OkGQUwsusKWZecsIOkdAkZN//4yl31WQ0B52vc2kgBfIZEqW1uYU8PNQReq9A0ImtqSh27qCY
bjhv+A4S7MWt1sbwT7RlWPxFUyknZ2ayNaD0BZOqtoHIcdnS/gVdT5LprDCd44Uyj7eb5pCnmrI0
rFh2mRMG/juB0ruv6s09JV7NDK39bg3zVlnng6JqdhhABwzLynA21Pb2jaGDyD0oAGeehOBXPgni
9EPWKADHDktXQG5wpn0kIt/HjPzl7lQFSxCccsR2nOdEszCExYvGZzNFLXJqhUzBysw3XvrD+WK/
z447z7FzJ52RTffaslafD6PZlHveJKhBlVuhzRhrxsAbUMKUm227UvctggoKDngCut+d01CC1s7D
euU4UH6+trFkLInOzY66nmBopOdEWnyJ4uKDWZOsVvaGJ6ivwKryXJcDVJMWUdglwhVtn9TQP4Wt
cXZmgY5OYx10gHySBnP2Ai5G/lRxcSwvaurHzxhnG3Pf+8QbavULQGQHrdkqE+avLTrfzF3ihtOe
bUD4TSm2gULp4TgAWZjmmMvPaQSQkG8UpASXMhMZDDmLydJ2kuBEjDzlJCXA/7x/pxjjvclUkHaD
csBMp26nqe7hcGLf/AKIGMm563g4Hukl6nAyIjskx5jKctAY/NH7ZeXcG6XBsswNQMl3LUPv7Vay
FUyx7Ie2TQ8eMyG5yDAIk8/xeb9QI/XMpi59dXKPaqn4wos8jeqK3qBnrfAbdg+TsGq5sqGEtgqK
3KqE4UqBYbl6+LNDK1b4qiMGiCgKfiorknMkhP2zYqsHb0SY2i2YLLsK7RYDg4Bh/+tZIQygpHoc
9Q1hYUrcEeh0memSIcjn5SdTyb6IZYF2MRbdUAPPms9FaI5du4xQyKr81779AVxx7QKz7kYAmViL
ccPG8HaKkM+r/o1FN+WIUD9QwWoODpTofjGTHX0nXU3AMZPgKoTAan7JWHYbfHy6Gc3icUCiOR3d
zmsMPDl9Jvfp3HwH6haTyRTSpoNqPBRb/ps9R7WPfZTBxKdvwLRn5soI8LLJ1aaqyu1vZvF0boxI
qc1qfObPA0D5lVq3Xd5kb4aq3XRp7vu5IA647AlWgo5KEA1d7l7qVlIOJ+jL5/JBpXjI7l1WnEo8
IFlS7utEZjGBhcnU7oj4yPGDClWW65Ilc/suR67iXnWI5slsGXSEQTP6g+7zMJ1FzMnb+66w8UKk
7JrFcvX3gYOgSoiGJX2X10DtDKz68NHw6z6/lrxpDReSJOPLn+y4oS+71UEf2HO363wC3QNSmvad
dxddK4DckEXhGWMjsFMJvlrACmBdiRrh/14bQnq496jV+1srNnbB/jqVIHdeZE5jsFGopYBN56ME
ou1YVZu/oc89R9NT8irPleM00ToZFnKBpknFrC9GPIQIHAdVAfGh4wdmw3jqF066bCuqYk/8+yD5
uPUz7LGSRW8WQkJI8WOsCxOnPN3UUhWiby8j2JzpOkE0+NBB2KWLyoMEbO6lOgHG3r265fwAC3QB
aDzt7EAYKB4Mp6bQY8dhlLt4ES95OYv88xFFFymUxa42xtUh0AaGZwlL2qKxTsqbm7Mzr5aQW9t7
VjLDvgYH9+aZi9w9oqo/v+Exf79CbEbNyyQLe64izXDtuW3FpiaHL+BVxz4gGu0BzKpfgk39D/Bq
WEfVWuAe086M4vqXfG3hTPKz+jWOY4Eo33ypPlqPO0tmxg8Ow08UnkCR+KPIQoNLiSlV7WszXJXI
Lm4b6zFmwL2NLE/GLp8/GCr9PVmuGMOXek1rUUv4d/FzbKqVkqtZB4ZqfaPPgs8h4rUDWEAMU/Ex
OS96FKhyesP4dUHf5QEyfoOGPTaN9zwZCvLzxhGcRuKxCYa4agFP2/q1002ZaSbEzS5LrhUBUd4B
SLWK7xwGQyHv3M18HD+/LZVBv2u8pXuki4/NQLtI7FrrX1j3YpZN4/iFhIh3vViID/9g5qeIa/wq
IwhsM0Ew2JAsg9uP5o1mZVfWRoZ0ZjcdiuEDta96u9/wnwr6uG3slsLb5UawKmd0Q9fM4zmBLROo
To26Y4d8TkV0ZNg6uOdJz+yIRWGnXy6id7qk5lnUqtAx7tgxOa+pi2BPugPAvWpYmUW6tckDrLwj
cgZu00tjzHfY9iYktcW1d95PtCkEMB9gq829aAMlS2kUaHhFbwh62VhyXxXrmN1Rz3ooZefeYIum
CK5L853o37NUlQgEuIaKRFmXGsGo56305T6TgCL2Bd4lgR2mVc9jRceQp4wgEn1MkFg3vVlpmwE8
ftPNkevb43zyKB0+U6siEWA51vQaVmB9xPRSJGUk2VeHOPC96238IciyjZNcipxNUC0zA/XyZG9a
c73iT2U8aScWwZbG7KGe7X+U8oCvAjPdKZX3rtRz9mmvEuHqXJOfH1t3OmtCPl34KELVEJJtIx+z
dEnXAaw/LE8NhxbHjsDEcBuRZ1YP9hrrfrJ1yrqyaqQtTOW4MJ3XnPfehpEl0onw+Y0kCtWG+fim
3XkmPGIGDWKbvCHIhzSiRRLQMYSQ06nS5c8L1dBFmpyObKs/zco15LEMP8XcMLu2+jLQrOkRj2t2
Ay7olDamAUbJudE603Sgmy/Trc18WWypBN873L9oArx36WNjJTAuh3cwEm5XK5RnjAn+trLt0CGj
yVjKTmhRKwcbgGJqjltLSNkXJswjSXlsCYMfiF1VRC/X1LJi0nURqNLM5aOiFH/kIi/PfI7smfsU
B/4BYmmIkwbcrWiS8V6u+KkdcoLVWOYavnNeqPHmrNKAY6NNAyvO1lpw6q6+J865JXB4mpcoF79M
3f86EWfgfFM0JUEJac2t58T2p/5RobXQaWix5rgDR9spwDllZL3zuCNWWpXgYyRGpvK+PS3l555C
e3vYTUNRCCRq2EWPP4UkCex0QN+jL/PCJ6VpIAQ+f7hop7nq9k0+zz5BkScO6mxBp5UmciGCa5+A
vedPtzV2rS4OkDd7wQPG1Th2pk22hlniaocTnohIRy3x5yIadpOVBcdWSBEqpSUKqfl6SSudf1H0
oOAa8v0yMRDh9etASGFwqM1SAVTRaAvaxj4IyCNetUD0ns7ig0SEsGflOV64rIp7M/e+mg2cqWb0
WGhRizNHmph5WIxLHePY1gBrF2pdtInMxixcmG+Tyqc+I7bACYDe33uqYh8/7YDMUI9Js5Zrbegw
PWuSE2zmydCUbIiy7JKH4yBS9YbCznTyLd/RX9TR/tvJODXeGDjkFWHN6w2glaJZwJL+D7puUVqi
zsIDPYofkKNsS1UXIa4crrtCIrT9MnKEgd21MQxEYxzX3yZqMOmswO0jTZIe6ouLPyfRBrHyx5Py
fo0/kmdBLY354ZVL4PR845YsI6kxrM59ntomLcgWpnWeezqd/VZv+rpwERWDXKtvVN7uyLeVVc+O
X8HFOOLHyPtrwJzi92njDwb8KKsSyfDwJ4aFNqPvGhZIML/szl0E0lexYJd/jOXtVrFkjWqrcjFS
Q8JU8MZ5/bRicLNkZ6+oLJm4r5s4ke7pDwa5WDzBwG84qK+oqIn+LK9yMQvZth5YLyFvTILtJW1Q
zdYOElkNl3alOgjpCUzr5lnMgoZfNtFRhXt8kVk8XOXDMXgbZvz0qDWYZO07rMjsSmxD+TXN2vGU
a9YE1R0eLls3iYdSzRL/Qv3SIUHfgOzkCiNZBo1BQPr9dw31zILT6JyopsBtf9Yz+z51DEtnm/Ou
x0OfprjBP2wUTtt2xd1aoEgF85Hru3cyq2rFqLH4W6nbjp83mn/w2f0/ypuOiCa8tmOnugIfBW1y
f86iLBaemfuocg+3hTdawk+P8ApX6O4JPaM4ihHHWDnNQCow8rE//98SRxG4PlUXrQMFG68inZOV
XBeIDIcvnQnyKJx3P0Vx2ok4UXs5PCSw8P06BLfrq9uOeKeU4uuLviux9w+r2wx7f/s9Sc4oxk2H
XHFXo4aLFxrnLSFlkCkvc8995nlCyw9dZB3gLZOcdYlB5a5WP6rgjzzUu+GwortrM5aeH6IXeaUL
+ko8KImhD2vQ0vnfYYK+XIHP/LytfFO/uPO9KyeYcbdFcklmCPeBbNRYvwZ4WEMWgaN4rvnOcN9y
hx7xWxxH/04TXArDxOl3mJ5qOicOShw2ZrJN7ysKNWsMPf6iOVqlEmB4jcByTwsNS/YxAj0dz7Op
A+wg7AWSslpb0YsveB3sd4lhntPf/fx3LvzBm2pFRTov9edIMNlrjv9rhuF8x2VKMjFg0w9AH55z
rSO1OIr7zE9EaJ+m3jW8yYKY6hpq2Dv6WaQkwih++DBYGPsGnpFiYOqmaSD8O5wHEna6U4tjHeHn
I9wDqZWsNSwsXYg7Fh6sd3SiuhYCtWpAylL/uIJcQhPPOyk75FLl0NszEXOoWQAOQ1W+tWmXsI9I
AcyUcVzvD1Fv00RgGDmq4C/QzpNpMvt8f1RsYdPFh/l+9VZD6EnaI9GsKLsaAwc48CSqu/BYEBxE
AaORtJufRjiFQeakAxS0UsCcb/dhLq7sgs/mBLJtXwmSwZMA7+1q71Tg1l1APIKc9z6TiPjNrkId
56lO2r2cD+/RXnSi0cA3QUh5YoT5GDyEIktLfBsJVKhVmUMZd1l66EXMpxf9+Xu4sys8VbEFL37Z
WicgLak/aU3UBEdTwv5qAcjnbkrTWOJ061CyQarG5f4wqG1fbmM4Z1q3BVAULEZj2RR8yzsa+jeJ
9F+HpbnCeZlVS4tJcLKahjbB7kUgRiQlOK4nimNN3zZkpod3+zT+RO/xKSTC0oa0kAG4qlQCXZju
C9TPxfPPCtVm3LhaUfn84ksWRzEI46rEFTDvdxAdhRcsC5dSlgq4QV23pjZ29sGOl7FLO/MSvupL
u4i+hYPC7yPzrFIRXDo7ZmcAiahciICm8Sem8FmOhGIxDn8TWr1e2MMkW0TP0LZHgSf4ZWgc20VR
NqNA8bWRSYNFHe/qUSAQeLPSvZYkvmRThq48Hupj2mNFOioyoHuz9AM8IUmPm5d4UJP9kUGSTkGN
GttxnuP3X4AG/gMLD1Xzb4Pjt3M0im9uxC5ZFXDpiOUyswuTrQOgH9cDCUD6oF8y+OUFzBFlvaj3
xQXqGkhIEqowlxbfgEira4UBtsZFiP/k9X6mOBkVKElGfpgoFz3KFV9Vqdib2gqE9nOmFWLBHly7
+85Xj8ZD/CFXJDzjx7E1WtZCQwSE643P1YCWPCUsS48tay3Rhqvzj9y4MV6pItNSQ9V66OYRLggl
igBOo1jcKoZHcdBKftHp2TzT782ZEKXh8LiqH6EeITW2y0Fa1wBDIoh8UY5oIylcGqO/OK3UiECI
OzzN2+2sXswkEChGpPbD6QlHnVClbGKvlcpVAUCeKBpXbOWgvXqkzwCL/Bldo8m7P644bENNAOwz
zRNhVb7U2VncMkC33PhslvPlO5Qhr0sUls7PbbwyP/pilr28fhDwgKJ7hWvxhKWRlL5Layp3b2fx
3+l/C4aR2PjKrSShFI7CiQbb6z9jUUkBkGstxUAK5M0LFibs+qIpYzw/RSEkxQH2a2TGmsR1MoNa
qWTZLobbLoLTmd3vhW1uaoIF1uceBPpE6kj8eVrF1DWdFJ5tUueRlSLXTgtxj45jzvG/FuKOkriW
zZz3vAXQc0f9YYx0EO6WhYXpTO9ujHb0IA3fpQ/rbpX5X7LzorHPeJONjCvTY2ocbj3RzfiHMzZk
h+9CoB08BQag/eRrcAZYr5/zNXx0TobCHZJjS8puSIQdf8V5OU+rhoMUteyWV2is5HryVJO0wJlM
XLdmvkrCK7utp3rCfTHGERSS49KNjCEa9D64EZbfdx8hHIlEFj7bzpYhyFLht4F/ExJ3kFHMGKg5
UGHht3d2BlKOOm5IJMoybagV8rCaeiZ5fg/UaJxWADL7mORQ0Uz8oNgx9H4hs2wWh9BPAfReHsUU
Bq9fzoEekx652H3zjH4wps+PLdDVgMwxY+cDl++zMgOsyAqkJE2EnPXSjw1ZZPC4HlauxvCAGTgk
GNjf5BqghGjYPYHPVhKbQO4oVFNGgzd1wEvlSMgO6Yg27Gug0D0iOg6iZFOgsfdHzlTaaCTCHYHx
V9PeQaIpo4pNgUJ5A4YL/39EVtObyZgGazdGKhRTLKFg4mLCImBukEG2xMv+ihudphSkfvMKCRIp
048ATbUr3jrvnxApI4Yh+UmEHcRZcR34pW3Ahe/TWfgUWOC+3vGDlXXQcgVhIo6PKzBFI5VnY+rz
fSy2tU+TBdtEX4cyJwavqPIMafui8fwo8YqjbgEV7d2hlLU3xXmSrYu3+mhVv4S4EUFSY6jUn/BC
825/Qb51GqCKn8gf51c7BibBZC9Cw5yHWHTzSK2RScuWDP5TaSrWtfbRd05h1fuRFgUCSaeqoqvK
nRdgOzZJ2ztL537yXULyfBfG2gwLz24V2Ds0WR6Xlx2do+JxcJbTMEhfLq4L6RmSPO/9BssXn7jA
fML0B23VtG1s4mTXtFlpDQqk1E30RHvrb5zz/EfsUKjebGNcIZR5b832m32XumNjJ2GlelTE8b6U
c7tzU3Ja4AzG/EAHgIAtniMqBbng2cVYXHP3zQfWW+PvWN8lyhofZd5C9eT1Pu310OnXx90zh9yW
5+e7gkdxKwYAasSDllDyYkU0dOVp/isQtGJshmeL0E2ySruDwb70Dogfh19fNxY9PuK0Z3TMmun+
PB3+O8qXtDh9uo5PT/rEmZOdGZAPN5MUcQmA2HnUlpBdm1r4iLUNUD+RFwNb+NNu1jCojK25EFT7
4uYP+iFQqmtv7shcZNlaGUR0fdMsogF5/hVxl4oOzd+lB4JryZGxkCvt1WO2ViiuWIl2hwl3X2TU
weW6gbSh8Bn1OtVhCUHMt0vX+TVodTCrqwdT+SQtSWsBNIwKpCKEiInK8zZL8U+76ZRDSWVTQ83B
AGFsKM0bxc597YvDOwYrkxYmquai/sUW+E/cKneIeclsgFSrR3niAfBF0oiBvXVoKs1KIEdaWYHK
kBvpcjuqmfl+gShnR+59acQxERs5/QNPpXtab1/49zw3WbakOf0AA8+VABuRfUG4vgYnjl8w1Trv
Ubz+XjWP3C7KU+beqMOPUbfchgyrsrSGIbPKwIC0Oiy+TfqcbhHRAbUE93fRfXZDq98w7uB1owEs
U4VeYLtOn124QPEJZY/XF10I5Cr+ULVpYDOlHq2T4xau464QoLUgCm4e2PjJVsOGvS9GeEbi2Ea9
VnsrYNLHiH863mI3+RiAlgHvdY57QB3v5T8iVoWh7zDi77WxMl68BywQ8aW5nJ2QaOEJVPp3Qq/g
EdimHoAYeF++QQZvTeiG1eDyRSeWnFXbxRSvuVuARLX0KHlHvexMerZb1bdpHNlaj38+aHxrIEWM
NQm/ps3t+86xy1kcKuRWa2IxMB60R2CenOUofRSCFml2KwUHLF44zbWXMjkqeBKn2Jkk4K3/cgGt
seI93/PojNMydsqyvrj+VrIc4E/HB14uSf1XKySILdMUJgmLKU9jYpzUjkcbOMztHa8xAfrJ6HeT
5BTRneQ9L8GW7yWdv3NfqXQr/ag8OG+dRSyixGvRuxjjP2qpivkly1Z1xLP2P9tR3RFvxk8tEsME
lpy+WFIIF2IMSMoUUIMNFYF9wVUMQB+ufFWcYEZE0nIs41PQWDVJmXPv1+roDXChy8PZK1bVQjvR
D/qV1HD8sKFeY2w4EBZU+EdNlDy43Q84RjkeDuLcnTB+927Oivq7Bo8DusBnoN0+TUlD4Ycm+vWN
nkQlmekDJZZZaJIZz6C+U92p01FMG5b4lhSRDEWZQf7TDms3EaxqZtTS6sSWmzIYCZlrm1bQixAW
qAGMAXl2AcVDBE68Tg34Z/2tfMRhksChkv9cb4AfoCFnhFiPWNCnA96lNib9MDcETHYZP/37L+wq
1w3pqNFkyUAHhyPw0VOt1zGZRxOOfCCm00taz0yeGNv3KKOBhwkraWCU5k4nCyg6IPL8QLezu5qe
rErD2DYwz3hQ5nW+r8+XuCGR4oDg6NzoyW7OCbS073OqLXOSWfE08jqCey6z2Svxp8b7HF3SqKhj
CC4uVJ+q7ZXgLIL0zAId0Npm4WPwV9afOTg14ZFFIdOTfgopw8I7lf75jKtrtm9WEtMfsPQaeVeY
ELoEic23Z7xYwoZGGcU0hpCCZESmE0jbAxMpPd2NSJCKyRWVcBWJzvpeQx/zgyX/vqmjOhgkhByT
bFwpId8npjQrXSq48EUl9Xg6+LeQK29UW47nk0bvUDW+f1ZxHXQgZBw/6w1Doi9XfQdrg5+LGkxF
7ZTuKaxPKDrTT+vMPha3vD0fzSot+VehwDg0sx3FrQZ9c8WbRw/lLzQjuDsJf5NXIhCJrXQaiPdN
JVNVQTbKX2Mk2whYUMYiF1Tzhv/qcudvODl5tIzmZvTnbk6MQh1mWyKg0J+Gu0PU0/YpVxHUxdYX
H4T2Ux6JHQhmrEGUIWDTijMw2ezIxTzW4YKQmSsZ3890ZFpjC3nZpsh0m/eL54+iT9byMp9xjA/J
xeS1f07OSfllMH837+nnz80vImf7V3kld8DTMPD5GYt7tHlMc+QF+mQqsJASU50tktSM28Wgxa/B
t3unONg8o+PsxCsyZW0A1Fa3d1v3nEnz1shzLfKUNsBg3ut/8mFYgeWAej2C38jcsnsI84x30JxF
LVfZz1cXhALDLszwuWe8UzwyvMtPuJFGR8sHvvwtZt+4Cc87VCKZ1vjeHw35P0YloyESNzES165N
O8PpNuR1SFr+tMs8SXQgwSdWixnYdKCo3P0Picvvbqi23ldY2K8EzkT4/OQ/mlFVt//QzqDmelgV
kcTMGbxsuOvUKLBlA7DMPcFoWIJVIhAUDdG4+wPQOVyJoNUXIaQUeDTSFpECrFo1tepfnG0NmQjV
8m2ntGWIbJe9dpMtty3AD54+mDpSdGQjS7Bz8hEk/0d8uD4Ac6JWBUrIaTT93QoImp7hgwhgtsC6
Xa12pkpKIAImPB7eRtGhKEiIOFw6eanXzuPPKdCrC5kVuWQZRUjpIjUX3X9tCAyEfBxZdnw7oIrW
y8HoMrk2EQC/oGM6vtCO6SOUt0oSrb2fRbXBJLqvUHeqKLatyH7EYXJoa7neQF7qfb47A7wG3fH7
wFKiCnKlZIRaVb4zdJQXXHthf0Awz2g+kwRj2ykzLz2hYXwyGOfWXImFDDwWfyghpB5RPofSRFri
bmxiGFTGnbycxWeeD/1bnB8e5xsJybryJswDap9kXuuMB1FqevBK8z9Wq2zkxsT1yrJ45v2POh/W
t5ry2zH7y7Zsr7tUxXrgumrjF/6ASmhaboYkVhh60MizU9gPg2B3Z/UlwpitsvtypewBy5qqHnn3
Vcds0XnJgS5W1Ms2AxceqlkEB9y5iMuRJ3z4vSFlBH7rJKP0SDo4yfTATNa9rjH5E/+UrWk7aMKH
fSG692TRANQdSN1SSGunyu/VnId3Fq/+fvaKimDMU8ZVvv68ezrG+bwulhRMSmu3DfUDaamHclw1
8XGkvFlxlT7qtn1sCYTaf6tp7rYb3uMqEy6owHEkzkvxlds6pZevMLJykQKoY4cEWn+/U1VJmr3m
/Re8CfD13mLL6YiO1OZ3l5+BNPVDweWCKKmBv+Q/WfMFX7l2dG/Hykoo+JwqtWrzhHryloZdK3cp
Ze4wlPSBFfJlTdJGNY5ZOXwxwdARSHiupGvuIx+HNv25d/q3oa9qig5kfj63D6U1cBl2APrySsiB
Vw4kmxs+Z99wKEBwuBGhaXzzTc4In+UbzLlEEn035DFbHk8h3a7oJxyzUOoomlJOpzIFuJ1QZE4b
Y0Ry4OktQKj0bQljCHZx4UMGsNVcpKrnXQnsHlYKJ9AoxxKUznPqq6YQcWnsltvZdedAUFqvarT7
bthqy4HSulpwnTdn2Wn6m4lze63XS9r8yVm8UeNOSOiokyW5bzuERYqCNqMYGC4BByvSSRk83v//
2ed+EniOlDh257101KYoupemgbvcLP0Mjk7D60BBTdMEKV4mRMuQb+m3JQAie2UX9G78CypUvQxk
zVfaJwKF/ACzmGvgMC7KpvzE3o0c/oWLWrYhTnAzQi6m/q9zKgvhmWx73G/EvY75RTk79kp6hPDL
TVt3pVONBhAJOBLF0Uo7CrItbMuHsvFGlftZ4dCFMVKsOyGg7srIuoCKypxGqzMyLr1Hjy8QnI54
+vozgqt0MNgLsipg16FG1j2E7MA+KMkIEA6AvRloDbglkMcVQ40YgO15buNJdWTgGPnI+qXLsVly
TEzzM/asVHgRPeLLOZ+8zHtBpxUdjs+nopW/3uOb/wE7mAh9ymARru/hGC0O4IBhiPL+i8rIACIq
ZdmnluC85aecdEXKz2am2KsBdGR2s1+aeFEnD/6NyOx5D108Aql5IbvnUhy49ROkEoQzaFEf4qr0
AOIDcTfqIgaNdsLMP0MHCYf8+sTIJ87sgBI6nzrz1lVudko2gmj6c3BMaHd1iYLnTJXb+DA9dS86
rI2Bvunle1CeBek3X+7I6AC1P1kZFw5l58ItWiORG0+bBVjtceYsiXxy+FW21IKKHdp5ZAjZXXTF
nEyl9MrwiPqa3UmMHe82SjbyHH9iwnofma586YOB8OHY9OGqatSZVzg/WjDtsgYGYiUXaSoZxLZV
GDnoRWpjExccyJH545mm0T0OTjTn0lVgvsX1NXuK+5/lzFdybi3zvOrEH6chuXR8dyWPyKiK1SWx
WMh0SKjxFm5/VjRIlWrSkqEu0bIlJSqyzYHtUhRvSefzY108WCukjF4uVVEa2sD9GXRLRDYx8FRo
oMK8QRKimgNtUOEbWNl9jLpoX2j8cwHFWwXLuGcWYC9of7jN7Sye0qGImPGDjtI/G/O2eGYmAitt
BFOYLws/iu6vqRhKdMKhTitrGWN2ZOwmzmq4fotvMaiCzDrc5U+LudBkr20hsUMf010Gk6vN3zxD
Ma/hzjYFeKtjU8wwgFmLKW/kBnf5OOPGBNlAG2cTYFpCs51lMLdsgIX/WpPIAnmpTdKDmCGI7Vum
DRB+voS28ZLkyFtC4OTkTdMR0kM/iL9pFlZRStDnwjUB7X2ibVyzLoZ1YIUxfJ08DYPlXnXRckoX
ju15UrXNXQgfNtCUwueED54MsK10bmix2yaWEOpnKXbeC4whR/dI+U+skvEsFuSSMnmTjitEl8vo
s4WSkm/tikJn5JLFv79xrSHiQP2M/Mk0BbRhaQLNc+I4akYVhtsEQraDt+T7GH8en0qNki/2oPlW
JaHzUswNzdO2WLe4YH5nG0vnjAPQdCj70adwUM3QALp4bByNDDXNfRQtR6jOfLrt7KwE4cl+AFXs
UIk+lhAyZ+HAMOH8ZnL3QOPmn0Mc46msz/WUUCzWi9Lvh3U6GOIExqULYC3QZCBT/+829tObcOe8
qm5yAAGeusJvndGiatvotn89tJDHwNGcQ2J9NyyQ56oG/JpOtnImej4vYYfqsNPcSKfZSHtzUkjo
BYz9KlVGrXiwavSc35qeJ9t+pzfhtyCnwJPDjA6vVUhznLlkoTO6EQpyWLJokCQuJ9BnJydx63HX
rCHd2GiMXbJSOGj9OaKa8oQDoPImkwF6kndD9Szg88PlyaKWlhNIt2i0VShho9iInJXM/skgpiih
XGsDKhYcz1A4qFHz83JlZ5ZWgcV3NtGnNh4ptzfbuxW9NXY4bOVZtGi54QJ+y2qGJNX/xBTqMkQK
V27u6XtloWwXeh5jfPav/7aJj61rc5f3oJV2Z7CGOgZ0GdZJY5iEt3dszzQEZCpYe5J5sgAMvpmg
m2gqqG1IWAtsDgRmNTBSVwyOZpyWu5jqKc8Q2I9+xFDY/3aANfLQ9TuHWRDODCMFmouEJ9kdVCQq
hHvz3Ii3HXuew8+BQv3grnqJc7bK+fQEWhjdlpFobVgbYJ0huROCImmlnFxEXrKObeo8l9vo1HPf
NDFtjzjfKMrkFZ26WUaGYV5Sxyk0jVffcuv7UQ1vt2MRTQz3SObJ0Lu4z+OEF8i+1a7/9SSQNlw7
yFPY5Hq2CMkWWRaRIDIWsOHdssUQGlzrWPxdHkhRxH3RujlKWuhrxokyncQvG5Deqn4ZmzIa0VuV
YTEmt7IUEnSIUBUTZ5mIzi0OrbT2xKLVAnoejeOULBMk2RQrAQthxmm9KwkcVBYav5sOdxB/oaAz
2fPgC8kfNgw4psIDWVqDroQekj5MaTL5oIIf7kyhLNnyl2siKtaWModOl7H6oeq1B2rzzlxFNGJ6
6fZFgtfcrFR0tlAqccENGtI8E7U5IvSyD8MPwWfaQwlFyrUMrXKMw5BZS2r5Kb0wly2gQA2pmeX8
xdyZ5Z9V12f7Dhogt1+JzK/YLFmosEauYaVHZaD17DJcYor35Loo0PaaAovf1az9iYuvHeMH3AYE
/sOB+ArpuG0881kHX9GFJLFQFkVq6ymi0Ot8/U/KmH/fIchkMj4Q6zuN3zEVMeKIPC999wDbp3iu
B8BuvV0iv4lHGnDswD3vE6CHuDFPue91YnLyp5gi5pPTtjPb0IxwHI8vk/vAHQ+TQRO+jbuBnLKz
nU/bffzQS9kF3PmPKWrej25G+erlBA3dKEYNmxA3GEkN7mjzepO3HTBEk2dXOmhEWurinSASbW5T
T0DipLhg6yTsGYiI4D3Grb10AJwl9Ywf68lSDd3NYNWeTzacFijEK+jvt+XxC26OVaza1KIbHoPV
c98ikCVWnDcKTTYu4r/zLlCcNLA412yAB78R+XPWyRpY+DEaV+/6sm+SaWnTg33EyQYuC0uwKM4L
FMILi384xCqDKc45mS2qwNATHPQHTFlVLjhnwMyRqStGUKD9IhHSFJFjvP2UJAIl+7GvRyOjvhpT
Wz7RCrHV6qSmWxYAaKUA4yXIo4j0lwYo0vLtRaX4YeCjCygRHEShGG+UHlo65jN/snAZ5/19QtSn
h7CQclHjKktCtZT4Ox0lFMZ5Fc6yE0C2SQ3h/BSetfgtDsVoW6Sd3jJLLdcZmxm+flx5Z3jgsGsT
BgHZ2E2GrB2xVSK1iZU7dlEM9lcv3m0rxjmmBWj0+naiD+67LTk1Sy6iEqBk7evyp9QNpExG1j+I
QKUh678MLvikD7PaBCDPY7ZgErx1l7bkPv7AYWZMoXHk1wZnpQ6YqNzYH3S7rLpiX8j1H17QYyzw
FYEThjjI0ClXH7aIkH9i59VM4p35gN+/JxNhUGfmEBd1yaOT16YFhqtN9VT8LgYTaKQEwEs/n1MJ
Wg1GO5AOK1n/5I6fgIZvQ3uADhR+qw8pulFhhr6d71Lx+YRsxGqB646UODK+bE1waWiEo32RK9IT
fvsCLgdU/fGVGRobaPEDOduIcMuFa3B1exQB5OcBwxtx+Jjkizs/mJZIoESbjOhG/ysUr+zkDg1Y
31DWwLIOk23R4nM6DgJipGRUwNNjFkRKsjnmQ0LpTrSJS7UnOCB64Tl5S40Mih38Qr03OSu+SQop
H13HawiwIAk7L5elm9VZCJNR9b3VFBeYcMVwqFN2jx1rg5rKj/klxOAbnk5i5et4W0NxK0W/5cZS
/aSnWbGEMUlbh51GldfntPK+SvRdXNSUkTkn3+gAbMRQkvfkTFdnd6BdACiz6wmVAwQt8JbY31Cv
e9dXvQ1eJg1uRJO50N9vc1RiFrdLtVO7mrX0p9U+QPBg2YFSgHxJkSaWfjuYMeOueFRtP00eMHBc
SK1TxsozDiExTmN5VWXRgxehacyLdIB5phLRRA8LY3OhmhTKNu62kJ9ldZ5YadZK1YW0V2a6S6mt
XGTp1KIYPj8jFw7T8lla2jfUbvA3PLl/ywL5wfx9nugGGv7VdakKlhOo3K2crR1J1e4TtjxPR11h
VwQ3jLMu7w9Vn/vvogzcM22pcP/zjh/dHqX+B1pmxy55CjxugYm6kOx4fg8kCZjH3el2kqTVzg4M
ECpznJ6o6RmlSq5/8pipgvW+i0H2cSx/5hMjCmobMmkogpftTckUf+IsTTxdw+qX+H09zcCV9SA0
OlauS1+wCkJAAJ33V6J/hWKv/i+p45ueSKhtg6ClQza2OIqVFO/ZiKLASRQq5vpLd+SdAHMhjPq5
zgGZ3i1bU5wM36lc5F7U09hgkLuSSiNnt1+dq03Wqf6GRZpd4mo8afrRf15ww8zsZzRfTkTQQ57O
0HeORh0r39s3cdlXmtlmtbJoeWKx3mBwevavaDuVgQqixzwYtzPJwX73OJC+/U0AhP6XFvQSo03o
RczWn5ovIHPWAj5l+/NbpP08pmwL9Xv8zeAnW/Aa/3brzFpT1kdyJD85LHZLK/YxNJ6fmh1PgsIY
VRepbsu7riOlcNILW7jQQ3hQT4fXYY+Kt8TUDzpRnk8FfXD0W6Hkg4CaAErj8bzjeh/OMfHSnCJ8
QqymK/lgUfIhUkY5ncHB+LGz/9KHjjQNozb5XMlrzcWClNI5801QsO8ZUusccfxnfQD4EdFf9tCB
ZgiW5OEvsFd81w0RI1BUfhk4uVfKWPUjsxx/AztHZDBSpNXBgpSikk0Cn5DJkDMMfiXORnmPU0g0
j4R/iWxQu2sysX5NRYxfVhNF4rgcy2Lpxk6qOLO71WX8iWUT/MVixo9TaFyo0qstyv6/h8gTrZ2g
3d9alZ8Uyl3cdcD8D7hziqMsJW3eAVd6IrRYwfZJIHSZUjkKZMimr6gF0/buMT0imdK2+5pwM8Sj
H5pKTsiESzzhCzLQdgqJneiS1J2mGg5FrLZz+rWgekIhZEuURq3BpwjsT1MDLno1apKSmJG3A0i7
APiopNioyWBgbUosTMU6WXyGQbRB9vnOp2jQS/xqWC+Hyrxey9DUhsfClQS4vzl++YmXQQ0GpWjn
+gZRrDNBgikD1YGc8XRr9sZ7DCGev/0yjq/9WRNU+SeAilhVlRXXNZSexZ+EUph5vFus1zhbpg/z
dEVkLyY9PdKscBlmxZsTo6pzhpHgpR8+7pCMdzO8EAx1VeFKPa9XPTrI7lR5qBv/NAJYy90OInRx
fXubxSCe7d8+8rpzFLG7shaybiGvW6tXQcOqigBHOdpMI78AniKYjQcRwuQlV9hY7UqdMnr0oxPt
wTVRNymNzDvnPOXN/gM6lUB3YaDV3q4wsyb7zyNWl4yyC2AVkl5YVP9BFOXGsrJawniKYy4jlooj
v5iNiWqqkWzg3ozwERei5tCBjSyb+4JgczaR2aKoDIjEylWLplJFwLg9F4LJB7R/dWG1AgiEERgQ
loV3zttJkN+WApF//dzzH6wxQZOFdRNKsgJhKwk8bvuS0ANPi8gXNF3HgF73ae3NRC0v7awmHDaV
E5UxQanVDsEM0/wWmIK87rQdfkM3BUJ7HfRIoQh/MB94zvhu9zJvQUiofe/pq5lFy2n0+mL7N74h
gcJRex3hyTtDLbX/BOVozLP/8LL5R9NqbC8hah0HNlFm5A9cR7js9rWiAIU4AWyDiADeecQcwBnA
G/aT98UzYJ8/+JzRum9bIRuYGFLC4aZ5UKp4NYqKUAVB/1R+ZavjXz0Kmo7VioQZQydMSlrbEi3I
Mpi53tvd020es3mMD/6az4UoFv3WBZMVYnn9B0KSHIiiIKjj7zDCpoJcl0tJNKY9MXbEg7NxXWhi
op+8Xgu0F7zVUja/KMJSWeJoQaeIFZQaaPigP+pPTWOb7n2PVXrel2MfI03t6Il1M/P8PzVwIvpJ
lftAJd+oyY+VVw8pPhEclW+aJ4lojmfb8LhGy9uMOvxUzMtSN4QKWxqsWb++ccqNO8zSOWIL257s
1tQbenORwKvFLiFu2ND4BBqEeGxqQXpPzzOBwhWtI1QGX0iybnWy7rfB0Iq+s/qLkZzNugckwEKD
UTL2DJt4tER7HKc2qEpGwV1pB+xkGoq0q5Y4AlTV3xfuM+kkNKjPb+D+fevqJYS2DFtr4GKw0S6A
qyuvjOl5xkJQkh8XKM8ty285sAcKG8ErFMxs2fSENSbhBUV541SJhVZUTcq1K3mZbrCyY06rWiqt
7N9JCR0t6GYXcLG+SrNIwhqlD0h1GVntdeRgA6A2dYPBDqE2g5Hzyff+e63EaB5QFY0eGVDskPMA
NgO56CciMu5+ZyofIPjinHsNQgv06EGyu6l9YER5Yuii+4/JaFU6iVoUkNWDvs8h49ojiblwSQrp
LMcHshHGMh602W+MEo9DRRy4w6W6Wr8qx/zG5qIhiokq1VymEXMS0NQZNwawikFhWZ97o3+dxUVV
XXj58iDUXHqQJI4IZWw9L+XLQrDd5pnwy/EFUBDgO084VkpXA26ATtO4sIZqzUjcNhrR/zKnM08Y
cjIOiq+FngQr9j1cEwCm7O8I4ZLhpr6h7Elhmy9T5e+fKz0j26SQMny9dZLTvO4f6zH9dem6r2z9
NdetGMuGALIs09BFdqzMA2fvAmugvhyT3rVDXpoTWNDJJupQoCvnUjeK8k7QdiWuqcuvjshLmomL
m3/Ni5Qi33TCTOhuB29uaKj50Z9jR8FtDe5MXVwNPd7kUqgw0/PkAjnErZxxGeaFvWqE4EHt+bjn
09vE+Fz0XAAPOErjGSCUiFkN/6aYMP2Z4+1kRsvhjccC9cw8Js3Y+hwpEq6iJ2QAU7oaHjuuW23N
dSQVzpFXtvmcdZCZvywsoo/dO8jtf4deO60XB4RsBKfrHz8mLcNn24rdELYBu/NC3l+Ue2UbR7um
JTd0KbzZiI+7L48BGBS0odcrT2kkM1jVWV1ggRTq+NgCyzJb6mWVNLwiNJP/ms63Cbni0/j1Akcg
5Q/DRjxUF95nPSuFcvTNlnJnEU7317MCQhw+C03EprfRYS5slZDfYJ3ps85OPGLM2diCkFPnwSBc
ReOHYowT8IbOupB5ctoR5cS1f8EXJL9yMBHf4+zOgL1x0FKpE0v/n32EQ+2J5R7s3IaMRsjkih9h
0h/o0KXVrWestzgdm91ki30v82MJP4SzoK9t5LJYbFMMkns7sRLQC+lyqCahmh7C62/tTav46H4K
r+H9nXAZyc/DMIPqg+rM+2pLOIeU5wLQmrPY7bfZK9onEY1QMLbqpFkXOAUBwKxX055T0bjWpUxo
lZ0ml7qcY7Uw28yQ9dsneupjo1T1i2j7D7DN9OW88WCOethKV4I9VYv2rPQJBjte2LzDFVxlVsT3
0DUoadeo4IzxNbVrWKMxgRJexUA5/0YkCwpJzMOjGPpMJrMW20Vb7TNqPGRtqzx+MuR3CP8xJkA1
D90FKFhzVU6+ATBQU2Lk/d1XuJ2H0IA/UxzgL+EJFe7wU/n1pcSB+N7OKSDWswOIRoUleUq2RX4q
R8c31f/W11puCI0j9bmmWZr4Nu1ShmbjxZGiK0zoHkMqYpms5aGSFv53hSlaRjDmSD7D5d/IEJFp
fSwntymlfqbY0FUC6kr3K+xwhHqU7L2Y9bsytj8Bh01YKDI+qBJqNeYVlriqZjnFq5kvKBnIDpdA
dCjpcG5PcsOq6Nf7ts3D8Jdc6KppsL5AhOU30VHdMSYmhehHrLcEy5l3QFB70g//4jPKib2JFQWX
+vpptiEpgqm28vakw//0tYP+zfwf44Rcf/xuN/ncVU+vGuMn8aZwg2OGz75p01TN7snDJ3pRSIBg
0ax67ZYMF5MGF4Le/dRUqWn1sFPNRmM2anDv5qepzj8tM4qodgRqxNW92VFRv94guVSLhibBjE7X
XEHEZTRaXff/rt21C2kZO633AUKjCkG5xzryXwEaYPV2eZeFlnDMIAcEVU01IqQPxUC+IPJZo06T
a/wzYmKK8BcBCodXPL7GSl5MZm1aXX+eW0iVifIr15outcXd0OJL/9RLdsv2w9iMkQk9HX5LoFLq
CrTYOcxSVRgnq10ecHZNe9k0GtvSmz1vqaHwEUQGc8LY0c22FlJ9Ysgz3wGQ+HMAxs8a75eA5DWJ
OH+QOV03j41VtaRJIHsj+opCiKd7U0Xl3V2Is85gkY37Bh46aoOy9r8aiFJY0//2QqmBKfIsNq+L
9+mAVfeYEPmUGy8Iwx279qiL3z3ocGCOyV+Ppzoo1caBlUGrmHV2SrT8E8qkSgjCNA74/VDtoVx9
txF93Jes1DLkd2oCEcPtDPqPdsBbfmC/HX/wF+CKjj7yO2I9esvMi1lkqFSxdwQJbsC5eivV52d1
70pXSoU2uzaiwhXqsQPYi/np+X3KY8g72me21D+OvVdMIiZnAE7JXGitlDPvXF2NuuNGYfyQQ62F
VXzxUMk5AMR670PUy43uqc/8x8ug5qWaMh+skwMY2JGHwHOAXkwi7kGVSZkYdfikd1u+5+WbO3gS
qLsXF3zFBKzP5p571Fmyrdmb/6oOLl+hXp4QNsnvaVVXJ30Qp23Qc1izkgzMM90KtFX6kGXnZVG+
7QvBpfjkaB4oGVr01knh+k3+SXaQUMcnamKFG+DGnNtk+0cfsiij0FmjikP/OPwinKLB7t4otpP4
ySg0JuvZ+1AtifTfGIoIQVR+Xz9S8A8HtI6PdxCHsFZDyJDx28z0KUaWp6BQzloq7z4jxjfJo/CN
PemMBQnhOhJS2GpeEs0WJxq+3/+RO9bLHAWaNeoLI0OBhMsnW5FdlxI8FYMbU2CVRLOihPlSfUyT
wB+4lskbtkbJc4XdQ6yYbq+B4yBF50+v6oyLGEvL5dN2SNYYTxwurbC/LP+Q31YULgshgoJ1404m
needNy8CWVQraYQQQlxgHWUIwqZS88hHvm4ddfjq6CXLMhkthY7dlRySEp85vquG/0BXULFWcGBn
rE1EJl55UEl0K4dEFyfKTIqNCEQhhE7pr61u5NW87orLpi+RiBFZBWEcJ2Ytiu4Bir/95JTQJYtt
dvML3nHIJgahFQVZeCjNSV27m2sDL/MQFVT3HBTONsGoxcxxC6BNPyM2kideSvzZLFKhS+lv+KUM
Izh1hqcJhUjJRDrxKkCFMY/sNY7zeNitTN73FnOtUaWgR7aBBcmbgpivASy9ZEQu8IDuvdQyRl48
ADO9T67+KTEZObivErdT8HWZrR1lKAMrmcTdUDrTF6FoeW+1iYlFOy3aKw3xNTTFqRtodLqjmLPb
rQumLMOH/5osT1z4JelDSTob4YdIZTImd3GV3m28SThgV0xo15sJD7K6zXtJX6XojwLGT6051fHU
H15lszWhxUsR4YqCc8i31WNOuDy8LwSP+3UkZgoHbdMY3MKjx3/lP5fOMCyvlv1/sPoVsjJOVa3j
8XGvg67v3rjibVt/R/coKU7+Swi4qvDoubeBrm7NnACQpINtByDlzpydn2yAm532EGOR9F5/zwsC
vYZIlq8l4LCtd4SJsxWCP+b0uwV4SSjG+MdYo1Y/rztM/44qi+ATfYeOs7PmENTyns/VIqb0GFbn
c1eEngxdaCP5X2rAx84HZ73fCAcpJaMtmfKkwKo1Q1sNId0+MKG8cVaqUpCShF3x/Khtb7rHNZYG
l5NglO64gl1nxB8nyf0vS5ZUP/ZooyyxAEG7HgYj6n0qPqszOgWnONXFAQC7CA7+BE0axPPtjZRg
IfWkutERsRxdgX2yaNcsVCY/bpqDddHc5GVqazcYxEjAU1GABVvCdbqqr2zTjoBtRVTocp34gCmr
TMvyCW58qlTVVzcN6wwa6tgikftUNCy6rG8SBO+RZ9KF3AHOvZNTcj332aU5I2FSqE9DDk87Clwb
NXS3Q/62Wf39BPxO/sLjA5LG79oafk4hNHBnzeyjHugmZd+YnAVS2wtRH2Xcb5tqQ1UNgb88801e
IPq8cfCi6ZXx4FC/BZmQyRa9nlVlRC1xg+rDJ7JtM7U5RpsjNmJW2T/qh9KBnL9n60bGPqx+T2FD
nrSDeQQaCRLlTWwRmWA7+XUFBFTj21qJ2pdxp27i5opJkOsl7ma2R22cCGm4Q4S+tA5Ie1Kl9iEy
sjl/B9CL7VEjp5Pe4735pCu6tGAUvVPqrHMCFUOWjoP5gfxSxy4UAVqH7o4ffHvwZe4mgRJa7Wsx
RmrVnqxSJa9IKB+NTzejxYQoHJeLpilaloBzTguk7ILUm38G7iBxyOluv6TYL9zGG4N47qEbVuGl
nXjQGiq9aWh8LLoOnvFB+UfkxbPliHet7U5R2KY3L5u5GTwDWPorQBO8wOGPUcwjUPjgfsEwgb5+
5W8y6M/ROmfAIN8j3nN74+nmFqmPNVva/hWYh9A2QNdY6PaPhf0uoSlDmE7vZbTAtFMH1JXrsPNO
F1M7Jw3Y/nF1IihY74x6PbtmAyLv/2sTXT6/tv2Gtmm9HeO2zWOJg26OS6SAqRxMo4XO/uPUczlS
HMB1vEjd9Rib6CZgMU6sJrlJwtkCVUQZzDZZlXdRMAvoZkhwDaKPU3ca4w1vXmNvAMOhrKKUBl8t
TjH+mf1aYduak/jTL1mVKev+fDQ8J1VLtWs7FmUXOBooaIFWSGOzj70mhB/V29Djtw6epk1UkFht
rKlpyDwb4/rJaoBCvRVA1wfNDt/BJOLfhYUZGGCRVZVDtaQKzVCkVUzDIv73Iz0PfEOiLwoUDAJo
Gnj5Ndmqg9oRUdLCvjKv1y9t71PSj5LdN30W4SN95Fx8uoNO6j3J/bO9b9yekb99xdHuNPaTQ43+
f40YvixP79r2Wdz0Ng+M6YTXbvGUaOJAw/Cxkebzv+xlUBxazzQ9SP4Gy8u5+bs3FGAb0wWsMLMp
xrfLvEmbAX/J0hA92Hcrp2DX0w1mFwquq3Ndh9A9oMwfx257O9jY3DZslGnfyxBErCXU3hiGf471
WQ1r/jPBS3x/WUgRmml+8ysIe4uPmc13IIIu09bOH046VpWWILri3MxKkh6I53QeJsFxoMim5xj7
B05Y2U3vsD0yF9t3BlI4n06v37o+CQ1KOuA/0V9AKwFHsCMP+9s1w9i3xeAtaCS7DsaqTIxYy5lL
FUb3TvOwBq3vWbDFbsEBV6VcJVR+nFapvWcqNdQo+X+VQokhe2tc3N8/QZGW/1c8KmnIUKTOPyla
Vkd9pqt5Bn/IbvBd4MngXilhLTwk0fhfcddDcYkwj6tvHteoWqlZE6+sTpAcKXxvVACuD1Yd4VZU
Q184POtxFjXqWfxHNOUOOhrp/f1PuJTaZik5rM+5Vzi6ux7fFgxsZneUaqJSdXm8dTMJ5cQu/5ym
g6XVNoYzr547HtqZVuswXmhx4SyUwtULLvJxMwFpTS0ZpFZ/55l4h2w2noVRzB4ESAq3ln1vL5Fh
xV7duLMCFfT8Pml+wOJ3opqg0StASnBE1BMEsQawhLt6uYtwR1aon8jvjxpB0mc3rPsF05hUI2z4
IMp7tehhhPDBT1S4r39yVyzpe27VUbXybCBsIoDHhi4Ai+uFLiYG/6+eTndWnexclQHiSXqy7nxJ
L7stLnQ2WgSMI6chIuWL2Kk81wliJduYSCO53mkpYAC1Si3fVT/MyLsszjGav4UFWjS/Ddvum+X7
C6JEQUF+g6xm+wh9gQJTix9sTu+jcCu3Vd2i8s8ZjBFA7F0dMtdz1pCgjaCA3B1hnkctK/e40xXP
o4rD0vy8SPEfXR8SsxAX5eOoO5ESiJATeIcUNd3Z1N8M8ajXIOzUmB/BWReFbtPTXwEfmjT4HJBO
ZmOXTHFmh9V+42AEctMseuSiID8B1jBIg0UY7j7NEHNWSo8TrJT0EzSp8A+4VSZ9CRTrSdOVakcj
SRL9u+uJGtYNcGowtVrbJ379XWCPWAiGKLVNm4E+Wwnd6gFoSPWYfisRUDznDYBln8uCbzJhqVUm
unqi9FCHn9xq98g+KGm7HpcJb7O+pF7dofRUT5UwCBvN5XkJvYA57Q2fQsQSdoMA0ArWwjHIWAww
2SWxHEskcFeqxuyIiUClsolbaAHsrCfEkUC83u7iR0xudU2V2UUVJJ3emuQnG3W1QGjCPZpHcPtr
d/gLovDG3drEgrCo50+LmW69ugKj9uWDKTMFPT2wxmqjE2PwmQfSGiUkq7H7zRn0KB2ceL3aPsJS
HpRbKrOFpSkbcmEnRyvff5dsUiX8PSuGIcNfDjDGVUNHpmnn8F7+smP+A4RLrzXhafWOh0gcF1xQ
rbYIfMiPxqQ+hLoBUuNTYBft80ynkw8crgi7whVepaP3VCc+LXmuq25ZgGSTkA47jipmoEYPF9r1
01rTixngThgc3ICP5OTK3Cv0oPG+E7quM9tz0HLMrWWU3mK4APCObGFmabx0ydurN5F0XjiqA+oI
/vojUZDhYX53if3ZKqGSSuuCJxV/AVHGuhjJzFajPWkO4XbEuhVYFG9cYeDCJ8TVrBOmtvHLCK81
bAgFAWA36t6ic71buhfR1rCo8h3tkSnvDAGrXMcwnmcgNWVweSjOIdnwKYjbfdU5yb6+KFRJ5hRU
KJorZ6mcs6TvCr1uomU4iO4CDuLlwhgC4syEQ0wcZZYY1HM6QhQSobq8xnwLlgPpfZaBfEddKZ3z
aNZ8IDnIfmwZfLhLnpgxMUiLS/gpA/C7oh1291LGqvukM/uFkkL2yebD2nR47nc2e8p6AYFFQaKt
oHX1sDDLq5U3RCBBU3+0SIgUw6ak4F0AOt5SlF1XQmU1oakzr3ml0i+QDUUde1dnaheandkm1Yk/
aJajMQPIbrPuOzCtEyiK0aAfyEThxUz/t1T4NsoI4wLSSPut3Mqq66Fuka1DRjvpr05M2z8KCfX7
tMMMXM18IbdvEj5nI62wTJB2B8BBcxLyu9/nYQyfiOYjCoT9iESQgMRVRlw0RJG33dVm0ngFGrb1
CxsmILlBT+2LAIwd/0Mf4y6giWhiEfZ5ET+TAg+EolEhVVadxo/nJzGvQWtk/+dmX2uqVp4P43eI
uNmdjsxdzhYyBdNSEghnGjc72zm3auWy5j9C2p4FMkIdF6FbPiD0uQGRA3bu5icynLWqoLIDvarT
XXPEcQsrq08TbrGggmWzJVeyvuFvjvn9Ow8AQK8+zzg7ki8861M6TS5XTjZms6vtg/hL4aKbj/PT
sBgTSNbwS6nsW9KZEooFzxbo0TQBfDoXobpTRPmBgqQYGVPk7rNsPejD50hk3bDx6Wd64bvSA4cR
Y/+gAT4E67INhJQFBrh9nrchXBfT/f6YwncLIlEom6ctbE4D+PH01yODIiXm6iF6TkyX9tP3m0PC
mBELhjDOjIjS4eW/DGqBUMfqGCq7rAXzQnkchqrgSW3Bfq75ovyR5c7ADEBT0R7fNxaGke1iQMls
rxzqF4TH3ThoO5hd+ZUtXriSlMa233ZPefZYZMCt05XRXrYPiQPAW5f9HqcxAzuy8hPeZIWTZbQc
c5xwmH4Hxw3w1j1CQGBjXLTLU9BRnl7xe8uOCSawQoqfj8di0eFSHZ5IiqtLyh8OBVtgpfV+SC4K
pTkINgP+8PXNkTBD5QLtYaTg7mXn3XqXcoVGiueoolHijA2UKI8dnMjjZjvrjpEqIjzoD0ILbQ9K
BsQrzEtZYrm4luO689VgnO0kiRP8tIcXpU+roipygSGR3tt90piA5jg6eBi6/q++NCOVGMcY4qUa
TKuAT/EkLR+PdebQNwe8pTJleiCorUfxxsx7FtvQALHRvYxeUEMiWM78SHlF/GHMiyWyw/gmYk0e
+P7M4cBu73zTYaUe3znPdkULpOw84mkuwl4ADY3PU1PPAfdxsTWbEnALAHSRcOw9/aJIeU175ojz
g5wefgtLn0OuBvdAXMUn3rTAj2QTxe7riPKv/nMEn3I3fFABHVxlVRGGqBMIRXg9H/WQKFsrzra5
NNAWFTQhZ0+s1KeaT38OySUx8fAmWKDY0+0KXjnGT5/6cQ0/XFO0HwWsJQPvhbeRZdxTY/jhNU1B
jEi+uJrOIMIQvDAmIs1mjFjyDULUilGK9WVcp+vtNajxsNA0mhbAj6RS/otXrGB6UkhL7T5CODml
jgmYkMfQyd3TE0MrPrP9AJUaHgCzSGVILTBuh8ZXJfwQZObpS439YKSsOUgBwFwjCnv8KxqWPnaL
oVCbnb+q73Ay2ZUlf9nhbLMWn2iR3cx00ng4+36YDTlwu9ygdecVLI9NDxUWBKMSPsX4jyM393NO
76TxzR3rlKQWEg8BI5hSYpnYinTRbPLt9MsEfKtLy1GVl6Z9w+Nw3CUPG5p6+i6d/827XrpQtONK
zNgQCbNV4Zjb4/NoF1dpTOLdlM+rlORfS3+wF2Yvn7TOu2Ss0a7OuLWyc1P2zq6fbQNA/aoErTZK
GWx8N0IORVDCCT+n4tKJ65qW7SdoJ2hFWFY6R/g+V0Xdi9Fzonm8MAsa8dsI1VYDEc9FUVPh0MrQ
/KjuSU5BORqwSnXJAsSjT2dwZXgRHkpTyztC6bi/z2sJZ4FKN0WZdle6vDI6Z2Hei1bYnHtqZc0D
c+uMPrmbPbHc6SvY82RBVCfPBkG3N6P7q26sIpFCX2P07RwT3ffPF5lHKAABDI43t+PTDpiuoZN8
e11IFxBQCbpGywe7sLumzqB8a5C3wmrv8RY2taI2NSidIC50wXMD5aENm97zJOyBkMDY+HYM7BSm
AELwaOu3vu3pYVVY3hyDBTAvd56DyMWGO+edxOmOYyL2qe65QXTA5HjcipZ1aPU6Q+c4Nmd44nBm
api5dnWybxEr9pPKqV9nwWdP6Cgh5YyD2HAj49/wucXgWorlXYHkvdqJ1g3l9Vihw4hWzk4ORg09
BUFW2lB5vbXV/P6IGlZtNSTL8OVVQKs+BaoXs5LEKOeVyQwgYs1sp9PF+wQ2/8s/TGytS4V+rKPp
fdw4Tsfoy09pKavvq5uA/q3hle4l+9ASHUIPqBWosDlTiOGI/xO3U7ew+p1JVdK5OfuAclIVyFpC
YyU+NI/N3F6BT1su8Hs4LC0mnLy4VPMIJoZeSPrLOcokrkjoEwwUTZtIn+V7+eXhr3pHEJtUA3UR
l2xCvWA03jqrNNffJNogDyLd+DDrMtOz81Wrjh+AMSZ/cHtaSldi+6AbGqhVbbzO10tWlsCZzC4D
thn0P3Y7XpwvNHs22HdGXwkWJtmfPkRfBPsV+M3lEKEz8xmUz6BQQL1Aowhz91TNQBgNpyXgkUp9
BLXZ4Du9nzYKyORKc1rnnqNMIgpoBzFNY8RrE+D/CS7PckEINvCogVX75bORjDRxAax7BckKKN4L
vf0nyTGJ5YAPsccfaRDFxGsFMItYM+cfCHFHYUrin5JmtftqRsaixXOY1bTfQ44EvdfnFhSCMMdx
hoU/YkekW5jwi4+Lm5zkIYdtvX6P+WMgKi55OHmqp3MyJSDzuWDeyReycsWacjv3Tb6pPn0YGo1m
mGxbYryRPls2sULDC8lopDBTzcV8GsGLPD7BuoDKSVqBQssSt01OTi4+jNC/fwtz/lxdmZJ10TB2
SVynlh+s3oxwUTNIGiAEQd7TCS7va3KYkzQ/QYJKa0IMZ5dn0VxbgXZ0OTanm+HvHADJ5XX3u7Yt
J1bIP6cSCytipHbaWyXO30JTZNHJ0rsVmiUqv8yOs1yt7VFuzM47r9WAlgGjgfdzn1T4jw43x7V8
LfEOjT0elX/W3QREilZF4D4Svx5yk9Xi63gHu54Xy5mi+KfCoIpufnk4gAUPVtm+nK6kPMtR97jX
83Na7+eK1LQ6kanAORKlx2TNtL/YeibceMjaZf32d4bmgdG2+X174w0iSVbdlxhXdWFfRPEmWY8J
Tj9kfDj1eBFt5YGKWY8/319UcKmSPJ2ygcQ7Q8g5km1q0oryOtw0O+xVo6qiFbFTD1Tc49K9Mijt
VvR0piF+fpzJQSLDtoQDFLLV38aupc4ZlMgU9PCkkWI6sSTZtWtycVvO+6z2VhCYy7mj5nblmv+/
UUxFb05CAjyFWXnMbPK02t/5zwX6sDDWM6/JPRz45otaWECdVhrfjxGvPBMimN11kVWBPBp8TCmk
HHeRYnE2eDC2P+dzt0zeHsDMCjLzPv1whjplDl5jU/HX27cruPbmc8GAxkVgyQswO8LPXp6bNd2D
t873gSw6JLorEdu86psDHKgrkc6+i+GKT8pYpt02HssF4pzx/+3vrP2u+Xf24/AFTUKIbWJMB9yt
KploxjZz0IqFTydJ+kfrWN8Tz5qtn+waWygkf3HwWtuizxKwovmhmuyASfUN1kB3ZtJa1BrChvh0
qmXi5gjYbNVtwhjQk5lanUePr6ICclEWSPMN65CZ2ASgUExlRzOWgo8dJzd/9FfUhaXM8aZM92zs
wb2BrMy4TK08oUhJq5oTLEpJ9RES9jqb8hfxBcfctU8/XqRypt/0M6TI+aDkOEk14LqWeEvbe1hY
+yRXOGlZ1UPFd8BtAMOeunp05iybedbPCJpZKM2kFxItzNcl8/HYjow/N/rvn+6kGWlrRrzjcf9h
Iq4VBIGuayA29xNMH0AuqAdetGVSNfRWg3r0m/ehq+xYbEUwzk/ZyW4LOoDpvy6eDWenT80J/Qbi
Kh61NhEGeW19fwYABLQyogGdvLFrR+ZwMEfuc0JJYKAMmk+8zSh0kap9Dd5LkMqXWxOda/4L6rjF
mpHEk9gW9KRCSQ2NH+1Mg17a9y46Cn19MFbavcZPlrwcDaOf0+13Q5VzJXTG13LGPYrvNINsjpBY
Pc5WARqInJtNJZsT9sr+uShBAHR+B7dp2ovJgtqy2xF2aQJoxSmqOKDy5EUQ8FqxC3Pr1BzrCRZu
R3sxe8s71YNQBk+w4MHq32xiUvV4WU2vngfXcD1Pfpd83Falc3Ge31uIwgBP9xFcrFtPAv8H4NHg
HOb1IVhi+72Njz+B56ShPxKeybRdtjFL07aakOXHaPnyOSTGjxngJ7NRrmqapDSexWX3Lay8U7hL
3BoM1TMv6+R6QaVpHDYMg4L8xbwN9m04GEv0MbtxL1q53u4llz/sNCcfVF6ndiAhOjtvn4h1Yh3Q
hOTFhimOB+pZaULsym+iXk4IgIqjy4C7/v8B3Qq+DK+kgR6c5dafVo7Z76YbIJ7yMJV3IajRNmx8
xTU/deVrJpndzpMJEPNNjPdCNM5jPT8TC4ZqJWBjCoePG7usBAtyMan+a+hkmrSqdHT4157fWNt3
OfyCgwLoPs/SLiujU2HEP/QhmSstFYMBvUWzUQY/D3M9AvwCqrcJRd6hAwqvB1Eo01AAWubpJHzJ
KHD5Hz1EUU8FjRkb8gxHEEKBoLX7Z4d4hORCzPujxKwiV1sKImdGJFJScXoFn3hTDyBMZYJlRM4H
xd7JtAXxVDLYaww6DybMuZPH5+JWle5b1sGxNi+heppRMcUVIUP/tqK6MfgYjK5gwBSIr1GJEgWh
SO/UZjaIObQgz866+00ksLiJjUPj9dVdmw1j70QUZfGaTHh+2KEHjCz0Qyv5jvOYgrHSRB5e6kv9
1IXz1yqSZTxEWyXth9nXtsFGkfOm6BW0qSwDUlLGbbhIS62CgXifSxaRmG0trPHCmBcvOTeg5ykD
p1paD95PXFQ93VaKYK0jBvTo4/KKxZI5weU2xofP+aneeaC+KbuP5VAuB8sm4HVSkoYlmSyJwJmW
CZjkEPsGhy6wgIMdmRQhdrPCvoocpXPobWUQ4wKnYYf/6GTIYasyvKXSqc+vuih6k8XhFSDgce7J
VxlyT8qkqcv6/zOJznkxaI/RvHiRmiPdHVwqjfDP6BqskSeUtFVOhF/GxdGZg/DZhA5/Pn/4gKlJ
nWzwcq14HXis2OvUluelPOCxnXFUrig7Tfh3aNOXUJUxXjYRGp95T6cal0O20cD1feUdAAmpTu8O
8nbslA9sidIqJZnczm1Z79HSzTKR0hWHxBLh87o2P3h8chCy4wU8XDtcFEZQWjz4WZW9vJkmaZug
ANM2pMCMTdR8QGk2PWW1xYRIJH1ZGwub2Nwlz2lVYg3CT3rrrF/8s1WJTpc943wGVoD4gMjWs95W
Hgpk7O2co7COrctAkYaL96QsgdTVAFDnGAk2BB/US0SzGNsUBuGxWpG3V7BuHOb516YiCeNeguqn
SgzsF/4tb81Pt0efoLSWFRCT50Iedb7MsFDb+lw3jcGcXZk3qsBER4ZS7QpLRB1tsI2kf04sUUoY
rrFpNCMHn/xlyVUbHb+z2YjvkvOUdIQ+HlK/I+r12oWIgVG1gYCjyzAZISR2DfYwrB5qbhnMuqim
NMU8NlmX1cZWr4R2vnrzZS0pQn8leO2fa8JwsdmDumOXesH62sS+1oRCwYYf8TAmiRPl/Oyonmaa
5jcVe13JUAU14CuQhwvuayutlNwA6Ze+d1mdPjcCsB5RCOe6mDSPN5AYkW7HfOgzxRsOPKAqa4eY
cNQvg7/R7wCEJbnAlwT5gxcJEX54Ok0tXsSBeHqwuxCJJNFbayHxexJAopJN9f7+J2DVv1tWO+Ra
+JLzACh7VCW+p3knY5ur1UM0selpeoZqIm2/tPHlVOFA8pstmZjgjKB3qv5igx5OUv6ofL0MOb5M
ybA2wqIHvxxfBcgJ3pKt7bi+486tXmnmV9cMMncP1C5NfuTHZK1UE/a+EcdV3xqRvy8BMDuA5xiY
yhcuH06Ttw++dD/lzdS2aEp1RG2Mk++guXCOwIq/A7JQpV4EA3lWSRA3rQ66vqniaugsllqjnF7h
Ilp8bnHsZ9m48YBWwAw3Y+nMWf3nUx/t+JKopfZG1n5iigoLm/bEKKoWObGQUC+oJtlw5fBo7JWx
rFgoL6P5wEEuX2q1FJcjX6DiT/5Kz4h242rVQhUUZN+7X0CO4D3HY2QPffa8rlyIbPKt+KZjM7Gj
y1WkT4eKnED0BhI4RhD4al89sFgOBLMGww4tK5hklIn35um4clpa0+3xXpo0sC1uxlqnkU/gFOgZ
ndnucxY5KObO5SnBXfhTNZE0UC61lgYwJWzcDdf/FUvl4abdwwW7mpY5UUf8Aj2+iTCnd3f7kdzK
y4CGuU8e7AvfRXeLnArnfH9if3Gt655ER+A303wkmmadfpdoKnkhrgmdMu66TZAwBJbPc7Hohlq/
pt/8H9ejHPdZewqY8c/fNXXHXGYbnJU8CBC7pkTSglqHX1iDmHSbV5MyHkaGWokvCMAMzeSCb7xT
w51FjvhW6V46kf++aq1v527UaYW65rKgfS9NjYA+nY3IJSMc+fUISFBrluZ3gnePlhxJD8hri4Z/
iHdr1O/VZhQCgPKsD+w36n2VW8pT7xRzK7QqzuHLe06lohzLzkeQN9PRq8iJp/5NMdMQ75YwRrP+
rw5LG9SrD3W0AlYaSZ6gCpyeFVNsu1zKrG+H5ahXv7tX0fE5QCQHcdnZqjxytmIcWouNIG/AN3Gj
xYSebnk+GAUwHkPCNApdB0DgyMb48tNx6Wg5ON3ddGTpKZOzCna+NGGlxsFTSTmsP5k6xI0BNAQw
oK+xefopG6bH7/c5/g9qWVBRaDDEWuBut9qIOT/HzOff8oqCV5J6SthitFpTj+tr1o4C2nZG/6g2
NdzhZ9ZmCx+rfHkdRr2UzkIy6EXzvqgiOfjft/BGoScwezADnYrXYT6QJF16/5ArJUQIBXpYLZDT
jCsGHQ3kKdzgnkMHTqg4e1avhRiLAGIn1txQprPn3zrwjv4rK0wPh/GvPasqsUsbutIyQ0mMjMXg
tZeH4B6966YuUHDFHUehLvLLrq560Z9ArgyNms+K3USH5hJ4zpikyDj5YBOT030Bi9uLO7sVJAJe
ow5pG3KywjcBfzr/fH7RxgyKFPG8QMFR0NJwCv7s0+m9J3Wcf3UvtEfJ4BkNl9mxTcEOoXL3ccbH
y/68i/X/2E16YZBf2Vt05WbgfZoqpuaykD9j9bi28qOHeHLLJjeIEO5TGj+OfqiCz8+k90Wjoub1
q0HxNnBG4y4QTJ/1vM4gM6DXC3DDoADEDWAd0yiKr3M82fkTLDIhcRzaDAi5t7RdvXB0f337o/r8
dAyegKs9L/8ColW5JWHDYqTFDB3x+tHMVpEz7UZZXIknuLlX7i1A5XxonvZ14x0WU/X6PCheuibB
kZaWwBC+TLJe2BeBbQmwaX/ClEwVYY3CYNlW7WxvO5maqqKYu/Z6fx6Evs23GloQfNQMPijh3yVL
AWj/1R6ZgbMrcs7yG1qRq7yeHMRVA25AI2mQSTRzBAeH4BGFuQzakCfs+Fm6B4no9aUaCUO2qljq
olDG/HNpBdJbdegJpZS0iimFCbib8qvlfHD05mPxDkxZoBnZOm6HVzXZ6sUGVvPVEh/QuHBLwrpd
q3187VyYCr/N7Q0BqzEvc3mTrGK5lNYW8ZFFdD3rSwM2qVQUoewPVM81009w4bFvzu8Tv8hMVGix
71ZFAAEuw3L+zrRrZZWasBBVTI/jjkoXfv7q583dovtG02JaQoj9CLGw+0POjgs3bHM9ZI9C9sv8
gzLzXUiKqaEpoSoNsIjMoBsZ0sE26rpoK/F4apZRM2tgqNG5NJgXbr3qNoXTJVNWAYaz0T91dUnI
4opjSi5mHvRIAw/ApisFqnvWkJztjHoXGjojzhk/of0wU6dmIHyqvTXy6of4RCp5ruY06Pdrd6pj
2hhw0Z9PXBGq4JxAM0QdW+aBZik93ukdZR2CU3rWD214MPdkJpn5U1vCB/RSsrClUNwtx1fGWXyP
rfzQBT+VZLkJAM21VXm86C009MFinLFkIpIsPmgMml5yc/kKTY/YSOL4Nzp2Qf9aPVmn75NDvrRk
Smvrybcy9BJrw1d1asiI2ACpThxubtDHdABsYf/3K+e2w+SZI+ZPS70z6p8j1FQJAouCqghYnm2k
5469oXoiUavWeWrc8+K0c9WcbnjcUzQa4kFZhMq+Na9FMdr9mWJyUCFR82fr7y5oUaiHHk5U/DD6
Ua14jLMyrT2K/F2LJHGcxaIrccPy5jjl3bq6uc8eg5XhHbTrsIIGQdP+uE7IEhaGKVzE+GWL9wf2
KRTFhNCMVOlEO4kbhkE80OCQhRdkrCRMUOLaMLdYVKjucILgMobHFRTQgICSl1kFeGv5sxX9JOmR
+zgl7YilREJXsTJSV0+Kwj07mPeGU7oRssk5nBmKRd2GiPe9WkEpiVVzNpW0V9pwSemPSyW0tbyb
34G83mYIGpwPYv7Gs62mOC30r6XMmkwTHZZMY6KwKdYLSnU+dRv79bEZTk4ii/kG5cCurCuirezC
XjgmbDQfuBNYnIRObS2YD3mVMdmfL3odBTjOtfKlYETaHpMP+pQeEfw189pUyT4LgVntMDf1qZ8r
Ql8pgH+hAgbogRsVcOoV2QGPRDDLLJXLJQ5CKo2+fzSIRNaVrrpKAbek8b/8lTeNvAWxsbTp9Jl+
HWx9bcHxICZUO5Cs4KB9+3c1AONzC6I0PaAMrsZCcaSADg5vmqYd/EA5G1gWXVhlddV54dRCT39i
0jufTalJs/w5yiWwkWXiIc2M2m22KJQ8uHrv+wGe70W2ZGPwabnc2o2hVI1adyn429W4+9SXpTfF
ADR6SEgZH0Kf0ugKb+tUZBI2L4Y8Utw5M12rdUk7h4I5bMUt7cetx4cKTKbr2spQbCsdV1puYvLP
vE59LheajoG3t65Q0e9x5n/IcubqbRWdWQh3lw7mv+5MdUSDIEYHhKMn1FMK51OritlY3Ut2eNwG
nkbmDO8yVcy+TOIsKOjAJSV01oxwuVB9IwzXXX5fs00FfRKcBzEiXnRqc0IHvGS2PzZk13E6WRZe
4nPgXd0G0FQ+cDIxmBhEmpdua8NwreYQ2jaeu6oIsfrmPXEQY2PjjFZmKKnMW2MjpptepE1GS/mz
VmmYOzi+Fm/TkE2ayvWbtCaSujb+YKzbvL2cnOHnypkTvi9AnOe78I3LOQDG5Qkhwem/ltIWNt8E
NGrroV0e+pOAiBV06snT77ir97AD/btCF88gUmKBICBNGqAXQwySJB5R7zoQa5oPfLQyD3Rd7ows
kXp3s1OsFltAupSAmMeuVSCuaL0pNz7XacRBFJAWqT29r/Pb4iB616Osg6MgHG0Cm7qK2KH4XHs5
dbA6LL7hkQDFweqfwoSKuWStE4WJrtNpqDWWoNO/EEc+dm4zsSoY+OPsCd08qywyaEWQ1ePrG1MM
+BJM3t0aunH/QCiyEb0g386PHNmZuCoj9SNZOLebz4O1mlg7ucofuRzyOF/69XM44i59Tr380ZvR
uBBAcikWoceIbc39nfZN3hwe16pYJndAINOd4Z4ZGsmRiLFooEYtf2x55KC/FwY0NGBnmn5kTATM
xwt+stWYHJP90znlo3JIsVCGhM7NP4Jt00DIRjwRNfhEtsrj3r2giBXvyg82fTfn+s8+3Ke1CvYj
TN+pLcfjtQQOuayHNurUn/TaqCf+utBjCZWcNwlaRFugY3hw99S7LR2TtXj2K4wxzF18O5JO/Drb
mm2inS+AofJUg8H5lXI0VYvYqd5VXQOzrjXFH9CKghqXtLwKoMTErtqvqcM+GmoCKTfQN7hJ1VmI
e3TFQNUSdfdFM/DjdRgT1PStF9ak5aWeqkH5c/JbMNn9d0W2SKJ3M69Nd7DvhFgM0NCuXkn5YW2h
82pdyMA94CdfTDdjQ6P+Ni7446iBLOzku02400NdTC2e1iEP0E5lqY1PkREvjZ2tqkx6YI94LTiN
MqOB2Seh0O+YD7DjfSLRrbIB4WRUD0fON3c6HB6f/FYhBbuvWWySyloGEOc3EEVeQTaSAKkaF6Iz
bUm0qSkI86TumnrOA0t3ZzixBV7m5SfFWM0ulk9gsVQtINPvKk2116viM25xMmeG9r8eST785H0K
uAjQtvPYrnZUm/D8Ngu8uiT1CbjlIIv8r05D5gjuLSCUpp7wftTtwy1YLjHMqkw1ZyvNQ31oaHXI
esrWxhHgpdPNMOIB+VwWk+bd6/G8Ob47dHpEHZClPQ+Zrm2UiVruZXcbYepLGs8NUID5+UflYt3B
dm0qWGZla5tzq9cWoMPYt7T/yZRHYAzLt0GUTemgmnV9SRokPluARYFglF+ACgxVoSdMAZBa0vcy
Oow4G+uvWoNP7fyLHWrTF4YXxJCSNrHnuWCOjoa4ymd1AVYFsSJX5G2ssXvNnYQ7PtGMD2XQNBOr
cDVbl+JQoBIz/JJ/PJDCNmazejVvnM4g/1cwF+k/BYrqNPmSGt5I/UuYJaoaRF6fSOSfpM2qoMVh
kjNhobseBxdFl0d+I+iTp19ouqG5Jok8HX7oxfWcetU9yeg6O/o+jLafKShY4mkfi+EY+4pAJqkp
pNG8efK/QwZ9FpyVEvt43wHRKViilbdyNIFbIIy5nnI3tfZ7oBJVVSWB6gvOY6ZGY+dFdwiiuWrv
0D+b27X9+0yDkobSHkaQ1MjXAGh0xX3/4gVm41jZ0w/mFE8mTdcBEZGAMjG2Tn4BbZebX60PU74j
iMbjuNnBAmiuMa5PmL/k2PQg+aPYb2b5ZJ3roi4nPFZ5ohvUArEUvqlJvwnYauc3QDEmQpFxTCah
bN/MlruXCCzc/bNj/grpdrEwUbTzsAAaC2g92snoO4TfXeYqJuFn7isMd7PDAu1E504DMXvGOBK5
cJuoav4saXU1j+eLaHudYvgCHtLneYx0ocMg7QIEPa5vVTWPTkJq/TUTA2yHGp4nCBCpNuf6DfN9
eNXzGFy7sXoORSdtS44gF1fpSd04aDs5+RCo6Dvg3BdLDiIODvUbNfYiuTVa56UUB1nzzbMm7tLY
Ebf1ZcaK10JYTbA4XXQ7t3I/YexPNt0GFJfcvj4A70akJAS8cb+WZO2nX+6AmtlGYN9xYRUrrDFQ
kEzEFLOF7hQF0dR/1K0SrayaRGFo9Bfi5V7ljFncJ81jWpGRUlETd8WL1+95KPvpP+4kLz7XUkzM
CelUhHSb/O1WDrMwmfgqniHYcbUw3q2vo3PHdKgaLxkgksww1altMeCGliyt8n/oc7YWmBkTJWzP
U012Cd809s5STMnL0sKI6BbrgBTEDG35Hj6wvbT2ZKXpJ6M65Fz0RdF+95a09BxFo8m0l9qDX0Pk
D3IsVHXLmfNRL2o9MOBUxtHDD1cBvuX1yt7lKqMgsgGGHLYl4gXG2Q2MwPvmgOvbS8TZXS38HbEz
oeL/aw+b64TltkCm/wX2Wj89BFvg2pf6Of5VsE3C27Om91JYoRoZRw95bTLT2tEgpfrUefozw/Cy
2S2yh7f6l6JI3eiUeuKL0CqEYzwOsj7Z4/4fiKRBDdC8gcbIRf2U0I0Vr8CfKvYZw16+QwZIz3SP
4SZCAVbvpjHapVKR1v9OSi+afNec1jKWXbfRgvh/OS+o8IU8tBeFPDmxkrNdv7o9r+cy/mJg07nT
IQRsS5uV8ahPrPieWchkNWGOdlJeMgAfELx1PUESpIZMyet3LzC4v3qJiCH3k4eDU2M2mzkY59WG
fAxjul8Jqqg8wiBAt2P+DNVK2uqlLnZWkNRnDlXzZyJwI3dQ8+Yep4y5EgaHDKS4gYC5WeI9Qpxd
rtyUgBT/l5eWImPCZKfEHpnr++saogBYHIFNgyr0jBiU82FZ5xlnLdXUHJl7BO/jUEWdck04ZbmG
JD2TahTiu9PMSp83DY/9sPZOQQgsQ3R9t3iWqJn5XAI7hHYMGZlV+JxoaUQvPcL+oh509LBRzuI3
GswBaboOj4a4ztKMNinusOIWgfVsSSzj1JNHTRbK2VETwzy1D4BnP17LVmLsOHkBw0PRhXqV+33f
BMZVf7aPVu327aD0I4/FQpaMMqFK2Jgaik6I8jvAJ6JcHrKx+yC2cigyyI+TSbTE9REDgdRNjzr9
ty2BLHUC/4eFwQM9hMCJUsJjyWeyMQ5lHhYFBUjgm22IsdZnF+kqoywJIz4mIplZlrWOCMykkPkN
WACRvcbULGk0EM6+taO7GBTcO1elChHc/8EMX2oAnzdLlIHTvOzpoveHpXt+BrbBvU7z9SHnU6+o
BmDYp1Td7ZGqGlwUQGccAvYzv6FfB13yl3tT6+g9LJcakiTT8WVUkEQfQ5oERqGEfAI5fWIA6vo4
TMcVPOG1tpSRTa6+W7Q4drLAXPMDiyoYLdLtW20rv1o/n/fszkfHPTQxeSO1qs3OHwx0r2clsp20
ttA1cqvieBR8cnR26fjkSC8CqIDWKYrhyaxFKBv75jM7L9QQ4V1wY36QzKjC1Nn1EXnRETj/pBdk
oUmBjKFRvs080GhqsmzD/+AkPerFfeRC1zP6sbcHQiRuNTyUZrARWT3tAHjmKWnHK/baZnwv7jNi
gXpx2wH2mXg9oNSqfkAVI7epHlNednY3yo0uq/+xsMJXylMQr9LwNbKfS00egPTl3FFBSNjqu/O+
Ey+hGCi1PGHGfIucMcmV0vrQAHZBXIHcg3ur1cDvrxSfg7Z/31XIaZGkwgBblKGJ9nsH1yviWJBb
DdHHOshfiLrxMog+AmbReo9apQDGC050tPl8ZgA3sqHeopnvSbVOSiSLDarw74d/w9zANeVkbn87
MoMPg0Dg0hu6dKfwi9yEBw3kzzplZHIx2S0IT6ZQl0pG726TeyGd/vGu7MmfJwS4Vfc9Cn6M8vem
vkIOGA8f62bGptZ5UX973Y13KEULaBMj1ytRxFy/8CvD2vbZiR3y4Px7YCbQsA0rtMwj7glVVIM5
7zFgMUY6PyAkgqOOap/JOOjsrP/lPDP+I2F6u5JYjuULFZeDUOusDi87Ng/TPOBANMj9r+dNGcES
A7Qw2Qg6xHtI/IXDDCsXisiTuEiuxXnveNLaQEcIUA09U8sK9KxJDb/96GCSgvieIA3Qv4pOUQEs
8NCeKU/JmV7MJRONRB0v1/TbwfMIkU99DwHCUeuSa/5VkG04mebXNtfl3aEVDv4/5Pr28ybMbzF5
x9HsWrw0z7fBoHKzJfX4CEX+6WvResxSyt1y0lzlx8AgrS8PZ5e6TeOUYdIBEE/XyNX+peuw5bAS
CJ0+rmUqK8xOXDFo2m9HHeXDTEl7bK6wO+u48fqZdl3s/R3g7hGaek7p/fpqi9y3+9LAU3NktTDP
FeTT2BMx/qA9635XxJh8M60FmPTRhP3M+7FiEzH+uFtDgS0OwQMjZkM9yIf2wsIZpB5AQ1bQk824
ewORmgoesGtxqSQ3XTxKfyRjSeu1Kb09L3tEKEV07b2xg2XMqibaRlhKSV35+BuK5erVDosmK8am
19cXQHPldzN+bDe7tlWak4Mz5SYOVuOfkiAmmJ+MrMabJ0T+Vj/C3yOzQ+YArWssf48/qNM+hABs
DBz3gXylP/pgI45FU0A8fPH25lhfMxhbahMdyU09AS3iekOWLkpqGSqPppSawIFcI+OKXQjDIgiH
FKnOuuo1flF4XnHEXN5O9EMCTLX7NlLO2A5/WUd4jpEOjN6+YIQLm49Uk4p6VpN/h88AWXfC0DIl
50J0cnBbS0MPWACyKIE6rRPDIv9WbUxZ5RCIASyZTwsq+l7haHXGsSGrJD+E+C1i3vS62Z4PO7iK
ZLoi7TpYTXYpNKGWcGl/jXVIC15pGwSMcXBFbWRKOI+WS8oVYwNzFCHqO9t8x+eiD1EiJP0XzVZM
3S5HrBMzyC6KLBdLdCf9O2KO+Mg/+BBJwtkPCFImte3heV1D3+h/1kxA8qaFbHke8yxVaFXJNF5w
56SSRX8C97s+Q2fLsIjadIWWzMQqQx040QFZM5HwmADWpONicXHKu02OoTrnAINrcX5xmvyIx+Mf
wZSLHAND5ktV3+BzPKdSRxDwlBEBneRDJCwx6ix6LMcD13a91aNeKrXbvBO+PDwZvNti1pWz8Z7u
KRQ3A4EEWl+Opg6V8iZmAI0BfYBzzbCf5+kZe2PNfw+5Af65RdcLlJkUycth9CRrf4TTggcVVMDo
tZ30RLu4ko/Rk9RCD9xCOU8L5+hj+txCF1hHTZXs43MxpXKAz4VLJ+7JmZMQ4pZO76rzRuPuSamj
YXimo8xTx5DZUEivhY66rJV2yH8WO7SjQnBajrAMGeibHweZhGWekbaAhujQ3ORGmaEGCO41VOiV
0g4xBtkx1ZLPxd5fF1wbzst9CMpXEi6Bm41et7gkmaT/c548Inikbzc2m02eVuk4OiwZZcR7aGT+
/HYYojtRWrYU/88lAGWpIztL3W2SrU8kIlYDQdbtykSwtGh48+Rd6BVlmWhZuaC9UDf7hmv5sI7h
YJTZZgWYk5/JOF6MyS3SSPDayAAYLSQqetAd+gnkfn6FFl+OcA9JDw6emP1mCyXTRScHX+M61wu1
B6wxF4F8S3tPtg8F6s/rRyNbYzMfSIKCm7wRb8iJbvz9d/RxLRrrepIbMYhMGRs4bcc6XS1X2sMW
YLkZS1dBbM+UltGkfwgD2GfdYzoCOAJSgeEMJfJo+78KvRn6WG8Uc78jrfdB599dK8VsSJrjqpMg
tJYQG/P4/WFZDuPApV2F13IZlwGos2Yj6uJyAFszhEVMDbbL+4tO6zentIdEvcpYD20vvgRsEWCi
krV9pU1O3iS0rQu1JWYqV764lgJNQUYn3s08F95WkGXGVDYK2057y9qTcgMNIE3Q1rImJB/D9olI
5p/KU0d1brH6Ni0OG1aeBFW6/ulb0eV5+UJqdTLzgivLLKWGgwDyXkgtQIPzCOK/4ymlZSUvCPD2
KUvRDA4TR37aBpDL0B842pyVnEKDjW+RiUkW2SRl+hf2+YWkCALQPCAM7p6Zw9+fB6EMlzN2tyS4
bbh10DuMA+WAnOdACv9lH3z4Ev2QKLIakXmRTLG2ARWTQnIlQbJEj/KTHgP4j/lpumE5ha0tf7G1
6C8YwrG4oynWk3D3/1xqjPATpbRbbTp0nHmHaYk95q+gmaj646bpS0OtSAiB5aq/6vLirfq8+Yr5
s+RbVLam+5l0+qbf01WW8y0L7EtN90x0vC8XvxLGIQ/bEd4MYeu6Pjo/zj60EN41JOg0Q4K6stMr
vcSfYo0en3mXXUwqjSKTZkPPKiEhhWzCKem2vN2HOw+Sgwowh+xclyb9n29RrCNCHg9MvD+UyLlP
u92JxR8JWDmzQo/u70PorLUFIzwo98Or0SUClTp0wmWdZV/qRcfCmQuntkfdC75DVJivcP57n17O
i9ZlOdT594d1jwVQQdbHrnSpCeJqLlqLvFg7XaB/+z8zEmvrJnNp8Pr9SCAPEH63Vi7W6UPbqvOF
bBUfTTs475Mc9ppZ+lNNWYHogTbuQ9aPRZZoNGtO5Mkhumvzj+u03HKrw+CSGCEd5N8Nn2W9ofta
xBXqnn8N5awRZzi3qiFh0f+RO0tPsO+MacmfUmt7G8DXWB57vLuf6TXI1+hx/sMlzvpEffKRNCjH
PtPz4rTm3W20V5fzIUR949R2dgBLVcwQAulXeoyn04gJT4VEkxvg+6j0R9BnjUgINN0RcaGL3M4d
Kq+ajSQOl3f8OV5sD80KN7ZAhVK+5ivr9zX8UReClEnqssGNc9bSfqyjmj73ezwfQqBHhOv7JPrg
NjUGBiL4sMGMccXYo9Mi8mOAlCGuj58NNci4LgkhdjLAUipESRD0aJnZC0yYolEFbqOBc51dPLcC
A9AIFxWmuX+Efovmz0ehsB6krNN4ud6oFtQJJ9KtE/Gy7Sa32c3QOnh4hMY6Omujdt8h39XzPX9f
V5Mp+ZDyDeIM4JH3oK+u16wS6RrRxYNLBYb2mRNF9AvtK12j7Fsai57dUJ7MJ7ZOQOLdF30oTgFr
tIs7756GDcvPXdhJsNWwsI01s/ZH6EK76ZwQ6WcIVFJCVAsa+bhe5MdaBg94TBJTw9pDwGqrHDuq
IEUW9o0PMqvOq8wBOf7JG8M2dEwEr3D9dir/wsqw4MWKDdkxC3VpAyu1Dj+4e/6Up5b1UZZ1K1PE
lG58kxDGYqE+ecQTdfyWIypdjK2xf6rqmS6E0F4auzz3OxY1pfjLNBa5ERRGSBQoj9D6DBujSOJw
yK+LxbogEVv6pxoeMgBAvgrhutCU84e5MBafcKKWlad+pANrOvwVd7e/M7orIXSNyM8DylsvuNI5
34dMSugeims0F0hwX/6ismcu/fPZQgueczvnrfvImsqePiU8sU55xbNMBrqSUVdg6buVozshXYC/
Bj5Ax29udORBXuhFAML9rouqrDBy7sNWtnCMd5mOl98uHyd8BYIGFttRu5JHBG/1S3vihsqaGH5r
Ji1ylgsFcKcpKGsw+rXHwHpF38GHQZqA3UfDB4buoMB8mgDK3ioCXo8Ow/fTX6GK+fX5Hku53bnm
wTC/O6jvpqGLIZoav45aIj7hX3zlPGV2j3oKWrcq08M4Kv+YddYPYJnuSU+VAZ4L1e8P7SIJrIjf
d3ulNA92LFQVVgAJqNVnC4sQfebd65/url6E16XWWZh+oo9xPD8vss2Hzavt1QidWXt3ILxpQk4h
cYxv7fxRHeaTxK+dozVBnK3KkjFAvbCe9w8V+EP3oZcvjCj7iFDHgWFmnMC6iZ3k7HkmEQkWYt+c
zSEsf94Plpf2efHOXz3nqo2c7mGqrZro0r6nI1NxgrdGIY615i69U+qO/GxA+ynpN2JLzJlS1yqo
bDZynclunnQqdxjh8scixiQdk5J8hArXOSkzAwK1qPiid+3yfT3iY+Uu2WPbQ36HrAX+De1NHfWO
DDTpzqEhXuKKCBA2CWzn2+Fh4Ol6K0Zq3Lm4dR0tsN827VcAg4zvYdyzHMKfX5ih9u6d9nbyUvY7
xI89olzWlbn2q075TQ2EO43klZaBNPZqLF8d9uF/HwJfhMGTYcGFbxONMwL6DV/2ErLy5DqmU0c1
BG8ubB9UJyKRUlpn+qqFBPzzNs0dGJ8ll7lAdlCwTYyeRp3hg1mATa6T1p9AT6ev0eBpjjWA6f1F
TI68dP5BvLw038/Z+5NlhwBzYNd6Oa4rFMobSY9v0iPSNlAbyzQjkCmEbqPCnpdU2JS2srBs0X1+
5N8aGnV1Znp4T7+YBHec5HLEZs2jQ62qpiti5kLPg88WfjjPhTSxzP4lqo3QslSMLeWd+XYfuy5I
+tluCf9VhkvQvLXOFQfOZXrO08Cg45pdwY9YZ6BcnupnLPc45ebOI85zoKxzy2l/QA+p3gW3D89/
FgMuO46+AcdHAbM2tpyi+pNeLGqhzYawNAvM4nkyYK0pZS4mFCChEPw6UxEdMvRjzf5eRkc6cjNs
c800lj0nuu3xl9qAySXaGnb9ZlEi1gwHACqtmAzyxxr+cpj9Ic/Fw4UIx3vGje0EZsHRCwhHd/QZ
VKS3uAY00LVKno72I51J52dIsq/szElMC4LXGLdfzW9xpJVSQ0HkbRyFmhtdpxz+5wzxlea79QlR
QBkqVFKHaNc1dLkslZJmNEEXYJHGAdGFRo7s8fxcBgWRuaR9YRUjBoem5lqWTaHLerFEXZcgDrsW
9gCEO9RGeDERsx2WXlpoHkfLL/0rdQyohXdWLbAVT9pyvGiE1G61C2JM3ZRFvDavrlj50Bu/YlNy
w9Sxy3j6EOZDHzqkiGiwhWuXsFceO5LIT26Lku9yxM6fmg4hcRybprrT7p4KufxRro0cuAceYsFf
VLQoB77RcoQb5olgy5pbAtteDQ5PoFjZj/upN3BJWo4wrlJ8SCWRxk6kMkI3bI1XLeMENAPn+hQf
Zl+8UB/dBzuP3KnO1YYH641j4aKU3cdfaz2Ud703EmuUks4dLpIlRy1QW1+n3obwVqZehQKqNUBj
vLe4ArBQ5AzVuQ4fu9nYHzbYW5DR6Uowh+gFQqOFhZI9Icuk84SyKVYtt5GnAuFEFozTWdFgNMmx
wPDSycqoiBqRjRnaJJZOHfb63Kxg/SmM3mbHuRlT5KGpo698Q1sNswLyfOQRedIJw/g2lISmxsp7
otTjto3c7bDbq59PggUjzlsR2+jU6/DEohJwnbU62gGxSH1x7c+sOz3tRC2ZlaPIBRCZbAN4SQcx
68ZpRcSCQJ1kB3LudFyswN+9rT+Nyw+aILeZat6w9gYtrCH61e3fxbX7MqnEQ072rlgV5SLquSAb
uOV1H7hzkhGDRuBFHf8Jnzg89a7m21K6JFetf53mYp0EG5MDKdO3USgBUK4GWbm1oXp6aIuLbx0K
/q3tmOlCEiTASprnCqQHQpKci+L/gwiQhO9yljdjfVd6b3UJrb6T42PHqQIdQqi8Ev9f4ujKo7nu
U1F8ABAq59B71WWWmdeLpZPTlw4AVVkexVIVsESJlDiUzBe53CD8jNDe9ZHqNln14wZDY2pdHE+V
WlzIkKf7TkT0UBEPyKCJ4IfmWXRNCHVUo4cVmHOsxUmY/FVOkDkY9Nqr7qoh9byjihz7mvGnpP5Y
M0mrtXSMxHGjz0R/zzrKJHiNqZ70k7jA3h/axJqBPHitSc7U1te80oxuBPRYERDjuJbZxzZZuEdq
cFbqENir7/LcK6xzDWsx3VNfkXoSLhYUXb1SSa5WXM7ZHmyU0H0Ug3zEsen4x2DWpGBS7K5W3CRk
YLha1LTW5X5RV+pRRpQfrcf2iohBapSZGe6mozm4eI9ga/mJIGEbW/0l2cUoxuCWWfTwgpL5ggfI
OOPY8pfHvITTkNLjDhj5tmcYzJfu6USVsa6xvVRs0EPoS6NHiQQoKWLlHkm/abNqXHtdMQmjdIx5
Lf1wHCoGqylXpxJukLNx8U/13d/MvrdyqMmIwFTd9JhxwOrsxmO32lFiYW2WTUPi4v5I37bPuZuF
zL0axxuM6kaCzUQrJkHoRGitPiH5puqWlAdmceKFwFrHuj8Npmsfh1DNUe9fFTeRolMyeo9fdTjg
8ZRVotdEc8qIbTkP1yaeq2cgeDo6S4WOVH3XMzZ4pK1j/0gf7Kb56eZAkg22LDde9cw01rAhnPHh
j8YnTWKJTYdzJyoE90sidNpjHXVndrgHB99Baxc1kUKaIM4v7j8LpaR/fYwmqmONiZlb5vXHnp9o
4nh5ZWK6d3gx8drcMYb/ga3xtMZ07w4F6zSyY63fAFz7x48Ie6YR7a8u8PU8djWbstv7FnSYWq1X
BLwNMr43WCJQtvy2NQ7b5KNFEYqZu+vPkyRYJST5a+yOHVhELXPVaZEL3fBT73RxZWWBkLa8EvW8
jZga4hsYY+yLDNYUNNQxyrHUJ4mciz4WvPvsmMGh2vFw4ducH8jUSWxS17Kg4n3JrLlEmG6xpVtu
Qp7ycIfI2I3rVihnsAExgzUe/sq7Dy8gH4RZIwDSdECUAuncGwmlFUD4A8HQbT6tUi2YMAGhF4Zo
k1yT6ee6kkf496sDdrlYt8SwhqqtV/0Yc68UXE9Cdfe/KVFASRFcNqTEbEWAnoiZNlVGrj1bTgqx
1kurVR1eJHMr7R9OXjp1qr2/GAmSLcMBdOgebqUuD/0fkMVJO2YPZUfP+VyHl0FLfH/cqva5jigE
bjT0Ze7g6wEZFzsFOvuAeS/M7RbgS0qauYUa7e89IXDBB9Vs3vDpa9M2fSe9iNA+FN9L0CcU8GNY
8F96a6RdbQlzABbmCB3gsDYXCFHv1MKaQgQDnlRqc6qXW+Isj4Nrzaffm+L5v/qBqzMCZUrOnO1a
b8ArLHkzTEerFJRKDm1GpQrqtDFiS8uPMkqXko2bvVR3mcUDvl2lLZl3ftWbzICZEUD3QmXkJrXS
5EaV51jYQlmu+cac8wmpcZW09zxOEs4ZzXiaDXlZVrbs486y2eISoGldKU8H/K6H2BTshztD3JdV
45Roy6CHpX7yRyHt8jVKgUg0K9lhS/3lNeHq7aIeRII8Q+Xw3TU7abMPoNLLuCR9msxD+9x6mw97
LAr7IRrvNZpAjOYOIfRN11KgjsCngOKHidLd0oJm3k+FPa3uSNOGWZMwO/ZaX+hdexElSzNpSK/t
9yNqh3jbiZeAFxPHDL6elfI+6cb+Lx7u8vEMf/mtRH5kPY9zkpg2O6qyEw4HmT5gXzEfdrJ8IQ8J
84FGSDS/nSgQoCPc+z3ZJckGtOrYa4ckPKYcBL6j8VKMUftYeNw3FtbUnk1aX+gyAX+TjYt2vW4x
xXk7DoREciads3DpFRO/cuS+U9AuMC7Vjr5kJ4iHWY6Cq0zkdZuyTlANj4GY3OT82D7frB2s6MXS
Clzwtfu9gpRlFSd8aw6ZMz22ZR0KcZFsbRgfyH2zNuOwYDZP1aOITRytHbJ/FYzrEKxc7BXqZe0C
CK6wJliMYCWTCtWsKbcJzzgvcYD0bh68tLn1L1vr7sOvoAQpP5VfQR9J5J3CyNa4tupRaxu1DUaX
ay1JsvLxOuWr0dpg6deuXrAhSdc7h47Dg7xm4WHky2m2zyJq1oZlBC2TY+phVqifLlcOg4EJsUt6
aeAyzON2fjTbgdsKejTwS66IFG3f46IlK0N8i3TbNWoRSnf3qP1xTC44ssvX/0ryRjn66yxN8//z
uaNpIPsIeZziQpaqMRQb1Dss045OGSLu3Uh/2QaUGJDd/7x/s+B7K0Kuo9UtD/e4pD/z5zKE0ieH
Ws3mwK3/3rTHdLDEXZIQhjI02IR3iQ7kpiC2dRhIfEBwUwWQn0ZSUAvNjYJctZurFPxtl6MfzGur
sHLgAL0/c1IYtMjjhN3Jg2UvXPqoDZvSeYERyoGG9KgMLiU4yN4Wd7B9UKcKTFGSDPbveOaBdGnJ
v2VyAUCxpW2TbsAt7FqjvSoBZ2HDzhYaXnyBokMXoZdtWNk4c1Qh0FPSTH4MRw7tbIWclcp0w3PC
Xmw6cFkmhGVt0Fat+Hx/lltG7VcLGXhVXaDd0plar7W/cHhBhHa3pFYTwKiRmIy1KUprs73naTY7
0XYvIhtqvEPO3Az3xzG6ivB/Ehs0rQusB9kb52hksoLGCYuLF3soPK0uVmx+zXEk7MbiGP5zb6fG
HqlJ2TbwBxa6W/P/DOWe3kkXLVWpV/prUsmHUMRrSpNJyq1slwnDz03toIGJ4dS7cvrbCQB8Lwrf
mcxFavmQOWgSe81pS0dDFWhIgtQ77cAkGGu+ipUpGIhfY0OSeS+XKhEcAHvlJH6M+2HkWNrUXZQ8
kXQMGEC8AeDLktiIUgpquTWrpWY8oluVzyMYkOoPjWUJi1Ead6Q9HeV3YPGl3VXE0gEGDwEF3o0U
P9k8jYAE8rhpKkdwt3lxuyznI8LF909F7aRXSQS53MP/zLmvbKhRc5E2Y+1B0M7gWDQGj6KHVM3I
TQ18tFXL8hKv3AUXL1r5+h2FxrpUvlMoXo1DuwHSaWIVg42mIKgr4SW3zWTaUVWY83XFhyx/3Nzj
eadhJDdyee5ScU5A/4IKnLjh/jioeymhYdF82Y59ggiFULdqeYmFtMSGPyiOZu0Om+W41DSy2mHP
Q4VYXTc0kr+7TAoF7CYSSJiX6riaXx7kDQYwtdTjl05vvv3JEACib0FUHxSOMKYWUNLR1OlqVL0/
tJBOtrfdvjJPAbf+DmAqk0ubtYFaE2nScnfmuWyV5Ym/RnKtZ/GxNF1Dy3OcZBZa0vcnIFg1yyEh
H5MSAX+h3W7QdKL67ZZrffOhk4UOrNptF93LAOLKYJ1SHnJou72qrqc+n7lagGud2DYTBTxIBhUL
tVqpxbVaT6tF7NHy0LuZSmn3ykDOyQ52GEDkE13ev7XmbfxFjdYkA/Adm1bGKY57gzlLYJmKQeAM
BkmK4RMMYFhJf9C9iZ/mJAlmT1mxhTB7ZoEodJBlHjQMPWd+Xxnez+7J+Ez+fb2Bb72HEgdPeRI+
LjUhhDUeV3Rpl/ijaJYV6csLl5exyYPX06FXYlDYUdNH7SG3dMWm6objzo/W79I/W2p/jvmkucop
3yfHq9+inGLWvGjRLKktRE/25xD/p7dDlsluUs8igXaB0xd70gbh2Mt8erbUBU8JKPwdhUCOMv1V
+AXWKliPUxIgBvlPdqGtgowTLU/ae+MGbord0GaE3Z9ZyVdoDte8x2EU/h1ZKhMvDvGc2xY9B0n+
BjeNXb6x4SbQEKrTcT4O/XjeuERqdWvX8+1EO4K9W+3MpE44ZuE7QLxt0BAVFuwmM6fdc+IT7PVQ
pWLqpwMFtMU+PluR5/JPjtyMxKo7tGN0Xo55yNpAjtR5R5bxqd4P7G9861igteMKNCCMRxzXUOoy
ZEO5p8BRFiyClm9S8KcNISvk5M5JcQFwJMmVShWtl5YQerJh4eHtml0ZpP4a0nyHT2aIKF+68vVL
18SarJkw8GJhwvnIeCeZax/xPW0Jr17GmDI075gc5q4pHPzSYNvCs/6Mg4iNobOFEli/+rZA/wud
RUgOnhewkD34tsqpt5qmjqinRjggjUWLLu+x0jvi+r2/HdW3DC7koHAiDq7MVveOks5g+CgcAW1k
oU0JcadzTr9lhZkQCfdDotrDJf3FuurAkT5zHeJPfhjMaVA1cAxo45YLse+G863OzEgIEASXw0Yj
zTvMwJ+cQp4eVP1uJAOo654jyjyAxSx431wXreRYyOlBOhMn2sVcLTX+8vIzSUY22KR2uqTXQ8jJ
eewsiBS0fQiRjX56AzJNAaJYheiCz53m7tYyWEI8pta95dG3xhyBXeHOc49nnNqkF64cd+Q7u3tN
JKQ3tOTUinD9YFEqe7JPXSxLfjmB5Px41N6gbcw2e+96YKohty0GTCxCADjdtPF+DWYaHAwY2+Te
fRUJCIAxorg6hW6Xzzp6qmjLsfECJSaogrn9NopINwkSR3hH+f4bfDiVe0iXdkuevxpBVigNo83E
n+vkytCEmGoXAn3kO+IY7ZchS002m2fJ4lSTDTlO9jMEbPMDOHg/y+hNEfnNyaWdvicq5sg7OITQ
lRjQFaTwRb7zLomLCqc1IPb9rEJuGCTdIcqvWUMJ+pVAVBKvUbf0juLHg3E15rFcI2QiRu/r+RJx
VyAnNuZJ2DChgnhuUklfmzW2FRoGSybWhcoNpaaizRdhWjfrVlASGgXZuki2LQlSDEJs6FOtYRLF
X4CL39l6VGQ66NxP576nI0mHJIPSsfKzMScJdVUAZufVqG4tQiUpqEm1b6o9qO26NJyGF3/+C4+D
BqFgoQxVFAM7cNKDL7HNfpM8Nn6FtvRQ/2lIb/+hSVYe6BngJe5fWWAqKImdOMWnYz8ZRpBQRSug
7DydPYVSq0uPk4QNHKs/hG9o2qmYRtb0ojYaiLb0e39qHTr9d9nqi3iRdiHxckykQcMCTRP8BlXI
6xqchkCb64dnxgV8P2gBiXJI0T5/D+1xmXnTpa2hKF4eNfcabHxa5dIm9+mU3MoD/K/l0pJkLRJk
wGNTpApNT44LmKvgBU2FRepU0Jn7On3be8xLR+w8/Y/hcffKlbHGWTv1ge2qV1Fd27b7aN1AJVuz
qHHYDh9BsRQpeKzcAdINPLvWtXmvDpYHbbGJySLCpSthdFUc785cYCp37b8b8o0/2LDqubibbTRl
WyzD4EKAlA1Kub4AUY6IQwP6yc7wnxlWIzGbRsi72VTAkVDrMiioOVM958QBTklM77E7cG4+cMgE
K0kcCWyy6A1tKSTCTZ8Q21G1Zw1lZBKY3EuoasvBkPkWmU5lacKhYL3FFEXt2FTVwch2eIfOpIWF
f3QydpR5KKv40e26uaOLbb6pkkkGsshXM57n28SwYEEqxfdBiYS08/DGlRtk9YHy/HXY5mZ3t+Ye
mBw8VeXBtSY57vy9NRsGUfWAPZxgitPsQev8iqS1yORom9HHllQZ0XQ+87HxQXKAdAKrs7uZOcPt
E40XPzvp0onBf201uWuAxR6n8iqEbJVjb4211GcUI49SviwBqvB+O9eoI1iAS49CGFbqn02Ffkwc
8GKDd4kiMN0gNO3D/aQU6HL4XDgSREAav8vcTdT3sNa8Ukb1BmWGjkvfmF8zCYWjtZ9MqAqEFX5h
miQZSD6OyvHyrvWDa4I8JF1GqAOZu6gdDoYWJ9hSlO/fCTwSdHY71g0fHjAg8uBpuSqyeb1Pz9JR
dSrakFYDTyAYsiatDO2dx0uGR7GwlNrr4th6xjSqFB2/nF/e3pHfjJKpRu9Hei4DezFoI4WMv81a
msDAITav1SOyRRoQROl6jgz/u0Po/RLSI7BMrbeUAr6ZOA3POZPQLpcsaYZREdZhnPglZtQzFv4A
X+rk8npSeQ3Xu28WXZ0D+aMjwSkco1IzCxusZF3NDIAQaDphCPHhOxAV9va5Z9J6iU7ppw6StIey
vO3EahXjj+i5uECk31lMmgjy1H5bEAte8OwWuzzkAomxy4rscgOMvgc6Vq7BDBrXzdKCXsUASWuz
HWKJbAMi87StiCpE4CrGW0QNx8XEglvNtD5gOiH9qPEbgwv9iMgq5DAdRa4zwatY+P2wWSlPXN17
I8kTsbG4/wq2MNJCXHnLrqCVkfFYQSvQtyJE85fQhTob9N1m2RRcOrfoRGlG49mZ++qEY2s5jcMf
D5TMtlKeeLs7fxUDEbsLsKWKHaEgXXTR0jwTA8JUO3EVXWGI5wHOJhr0r05Vv8LQg76S30h3p6r4
Jb6xsuNlSeXTupPUhbXOsROUL9+cvEjtw/2P27jV2lWUEMo0QlFvC2Jht7Q60cvxV8+7Nddrik/G
asMwmF+mY+E5jM+HiuGmzt6c3fOHfH0pIanzv0VYi2FKQB15jKkxkuMvylpDJueCTCkGGRfNiXVB
lOpjq9sjKYJvdvVxSmmjEuv2E0Ft/53ED4b9LgAO6/AltOSaq5jFc9WnilVXFCCubYxVs7sSl0Kk
F0gW+Y1M1fGVgkzl7YdD7NkiLhl6pkHHYWLAv9NWHOpSk1M4GpL361L0123lQbfDHgkEuJXCHhpW
CVo1/O4r3gG+TfznlCGWd3wUkqfrYsCzKWLyRMpZ9YxnlCZd5THB95BEVI7Uc19uK6nAmrnsQPl4
jGAKP8l5wWf5LNTsWrSMBU3il9k1/5rKsQIOQjcCSfmHyqXrPcjGPiFJrZDC/ys65TFbmbssCSFk
ZQbU488UvFpD/akb9rC/9AyxBgjkAv+vv2dbuH9DGLSRnXNe5AJZMLPstzuYF5lD/MmiqY1pGI7F
ZWSNBsNYZl7TV5uR4CS5itWrfv6RA3Hxxn9eONBVX/1GM0J8QIQlxnozE16/h4PAJm7dKbsW9zUG
MrgxlYHoDI+9ojbphNGkAsnL0h3wh/8inaZvXvZOnQVMD3ihaKBZSk4T4mccmvJ4Edf+HYzVj3pw
cz3Vd24c/69QBmT8g8RM9vGTbM62hbm+0537qHUfLkMEUcPH0lDcTzhY6l1Qfhfer2v7HKQwTgOl
TOVl5Ihlez2leTuh/0FINvPpwLnZO5BZFLVgodo3AIyu+vmrWEWNprpMlB9kw6EnW39vu5+he0v/
STKw3Nh+o869SsffKUJHfp+EHVZ0lNM3h9slLyJFrM8DKGm5dqHhBwI9NMdFffCDhBvRpzLzswnz
Nj+ME8eQkDWlPqbhppILgOWSj/8q/pHK56K/BzcfNUU8h8AHD0/JjOENJP07+AfwwVy+5m2uMiCA
5rmvZM1hYlCO70luQJDxDE0RjGt1dLyYrZJek8SmjzH5nzgi9B8cM9OTbvbvXIcHsqx4UgYad5up
5KV3U5EfnAJcK6veLi1up4T7wxtd53aP2kSiR/kD+auoGqaVcjo/lzxCszWtZp170Pnf56Ypstop
5aLG/Hxs2yTTsa1xiBUq4K8j8UHS19fKVufKykLL+FRxUEe2AFjTO3xMyWh5XnFOP9to210IMJ+1
eOjiY2Nu2rtQq739+yJoqzkhx/KsZy11HtFQwiQrMD04fviSyuG342dKfcvphoNdGr044zKjWz7j
SYFi9pRBoxI/XpLZ1MhFOSFT901lb4LVg1AIhfUGoCohTeGpUQe2vUADZuW8tO+oAuSWNlTCD+zo
f9t1uYoHejj72PTPoJBmSv0VrfDTVT1jNQLjnE1Wsi6Frx5teZtCAUM6cIh7oMvhU/xwQn+Mv7qg
9/ya6PhiYn0Z/DEF14+9tNyykGlRIa2iktDmVCU+pQEennlbmVydxhDC0pPVcs6KI50RvF04RrUs
2Hjw+JgxKCPC4zgln6gFkLZBlE9sRJ/sjg6Mo0smJqxS+uo2miLpxYm+j02mK8wODJC2JSVJtpfu
48Gw5h6X2kDvgdfGpnUbfPTPSLYxMeJOHxc0KO9F/OASqJQCn2bhB6pKmpbTAs/JkvmrRfZFq95x
RpoJC834qUS4EQk9tmYmNdQbYp5eVlyxfY9o1gapY3TcWHo+0/aTrqWFOZp30GrklUU6x/kDU0da
AiAOSo4azFXuX2C7ZfwLxlynCfoIh0TM2TtbggAee8+YaCgtU81MjFaJwA6rDo43uGLHdV5DSlC+
qm0uUBlFlz6aAqQQnJm8EHEyRTi8LMGe106hapachwpfQnctx81VDlw2kWzt5w0WXQ+j+ZxF7RNi
X+kpjVKHpuEvN1AZ+sWaF0j1YGTOR1rp3ZNQakJJ3VSMB9JgUPZRoPVsaCG5hdfK3PhwpbJ+84+2
kdKck789JZkouE2ELIGyFw4DMRuKoAHyCe+wuSXDmuv6hyxVltG8aSI6YsliO+GIIDeo+FsqLGr5
SctcgZCUPwAPoSGzqih4KNjEHpsmBVas6VgBjFvZw2jkxBdYet36sOxLi4WfnqMRrBT/qb+2/5IG
5uskmqKKDq5p+cr9zq8s2c6Vb+ktl/BGFfDAjfELYUBdf2DPwjAtSmG2NeTQoYsIIf/Wofx5En4d
NdEBu4jqS4TDhNPW+CaMAZxylhsOs8iwRnPJk7jHtdVzLZG/A8aKowVKS40xyQuU0/d344t+n4Mj
vFAjA59F7qS0DJkrKMTIoqKQ6Ioq+Y4CM3F8S4l7Tfo9sC3nNjnIZfiDSrRMEK+9CyvFBdvuGcVJ
U6u3g3nPmSsquZqQwc+0Xn0nRyHL2BJxDCGTcoNeqZPUiz5D+KaxMK9GqCikNy6YqUappf8OZ4LW
vnAkn/LxtFyfpInrclA7mDpAqNg4AbMg6/BeNVwbOyFTTrxscjrgEoZZOJn6hM2TelMYbR8d4EeE
mCrLrKS3LtYWq2zz1N/If0te1trepaELR9967NWXDf0zfgO/9bsle0DlOJwoeqCMKMg8Yry4zv3G
MP1B6joXVtnalwxooTohHE5jOYvcIbhAyzIi3F0we57a47d98BH/qEzI2UDJaueMQMNiLULyH/Jy
iTFNcgcyMXnJQBjWXPuF81OG2iLcU8BH/e8zxVg8b5h2rrlXJPWwU+7x98CkbxXnXjyNZWqofsTe
ctsrO2i8Wr39CKHfNl/3jgJFfqoOKF6Ug0Kj+BlQtkKPkMG/yNmH5DiCkhnGPs4ksgt6bbVH5qK5
RGAangrQeblTgb63mJ3XecjBkPLrE/Una7MGdSuRYJFduaZnX1MHbbcnB9tE2ZWfmK2H1Hxqw2XR
biJXUsv70sUkHfxmDEm278M/N5wKEpf3udb3h4Jv8d8HEFRIt2b86qU4T+NQm03f0FmDT1nJTUbo
x/Y8/MrshZZjHdyPmgq0FLXO10PZn8XIEM1Z8YClFK3UEThgDLlVrzCrHUrc2GgosCc1aYDqBZjU
L+gZcuXAynIwl0KDjfeBeekpqoWPFwFtjGx0r8yiYt2azwX5+CVgxUCXqCQ0IWouxei/FGlwI91f
USIEyTD8Yn85MLN/IFQEaL4Mjg4UX08G786bTi2axx+XFRCYYO2qIH05M+KWKFb0l9PLKOqqE3IY
FXu5iCh6+iXX3y2zcfI99xp/WNh4uMx5JRHToS23WE0OuPGJvvZCiH1XjgAt9TtCTKjD5sX9MbC5
amowZ8vq4PMJoB0I/RF02TMZ/MlQwQX1zvclqqEsVyPHCwdxRMj4rezkZn04uypGCXtYoykIIsFF
vJtxpd21I4aqVKJC7BadLwbW+65dt2WMNrPT+nl6COVXuMjRG9rW/HClMoj2gv1QaO1OHY1HEAJ6
wH5Ie9eWptnAO+nTwDzojfcdSeg5Vdyk6C+p/iKZQTT/FTME66UXX7zutHi54DwQLCp1pdyoNW5B
I6iwQ9iJKadP7yQEZGDfjX+HdMZ55ZSq1SXwX1qjdcYxAFdOi71FmxwH34hMuwDrWdHmhsc6Qdoy
uAW+T9eIudX+mP9Y9Yply1Pe+XlkyPuZtaP1KyNMcpqnYLrFSpcnDwVBu05yKukRzkfKqu8o8d1Z
6Z8f2hrbvT42b7ihnSwTTQk1fCJpL6sSbwdK9G7O6hsVGn1UEmd8CWA9VrAN8dLOsPMCRmYDlcV7
l6DeiecS7Ign9ZadpptYeqsJxVsEB1YzhxLA0aqVsspRGaIPVOoZpKzg6K9Cyj7Ez48MWYItqDXc
em0FcfTTZVwa/vdREwK76RcvUb0q9NSyiWbMPUZ2mP/rXPj7M79kBE99GmghUnm0oXcGBtqhPFRy
jBmyDBMXSmm2S4AorjayUm9oNXeptLNuMHtlpzhmiTEeROGNUwAx6QcJWkuW8p8lJhQdQwV2PNYU
gE4GSXrNAJGJ7KMhO+3v9aJ3zgom6PwrK00jE0JyC8Ql69VSFo28GUFHhW7HpVZvYus8ObPUiT/C
R7wNyMen56lIUzj5Ii4Z1G1ZVsUotJO2aV27vIXTkfczGibOWKaDwwHDCYHa+AuQmMdLba9h0+7s
sCJCYgzeq6g5Lvo+ys8txtxNHPpcPY1uvxoTQ946YIaKfG17XjZbGyY/+XkMI1TvEMKEXP/oJEJo
CCqRPlwlELVbw4naiECkRI6jHEc8sj5eOyFkN/fTtnWzMW7jgfCrMra7zgkMI/3KppNB/WxdY6FI
6H0Vr/6GCygQyX9YUXDx1FhGvsCyWvBxEtujhy5EfbaCOnFCdoF0KzjNqKp2ADuV1VQDltPYjRhb
b0rtKFM3I5oCBcElrbv35tvARtnj/wbV7m8DYdZsocG2l4FqronCR8jyXy5Ss1trkSnIfOaf8wHL
CxkqRZct6LLFUescHTfQtUKWoJbrXHCIL99aJc8qFw1SX0VytRFEx8Qib5vuQNfxTtEHLv61obMU
faeJaNFiJNh4tuBQl7JQNHPGxN0wYif0xcIYH18TLaZr5mxKs5KiU4zmVQdJMc8pc5G6TPbt8Rb5
WHmVzq9akf5VAkzRRm7imqeI0KhF/GYCimhBwDSUTzX4W9dUWpcF1fubQtJaXmtjvtB7clqqwgtY
Ih+Ro9+2I83Owof3qvzSQN5PzYYCHRdag/hdC77ij9lfgcJ1fDpFwRM3QFOudgY+Qm+tBCqU9OK9
82wBmKAoOk6JbuOR8+EM0xPpblCotcAfWDpEKMJ7XGMcEQwJrV9iuxR1kKHdYxzPRDvJE8jtjC7t
dI/2CsAnZ49MfmobZFBx4m3zfpUM6Td5Y+oiH1N9jMjKWvf4ecCkYBcfDpGSopMVoFiE9/JBqMsj
zg9iHuS88apX445b83a2K+ymPdMhS+s+/kiDAnYSnWt1/J6frXaQv/CGHcLNoMl/6pw+GHDRT+ri
GCEzYf05ueia/ojL2hwvu4iCxa6llsiuWC/tWOnHwZNzFEWOfO15qshpwhN0eX4JbS41xJNZqxFQ
GDKLjSZg/adSUiOCko4LX4FFO0k9CWflwg3wOriOYStVcWwRwe2DNz3SDLDX/I5gdzzLxX/xWT1P
aWEEN7+2VlZpgdSv8Q00o+cbu8xsdViYWyskafooQY4NLBodB1pRjbmInEY2bxUWuh/F/3xa9wQM
+DS8UN15Y+bG3JgVgJWgFzkci5Hb+mvmaTXjLIQUJdNO3J+xn5NY4s4OAvbH4p9qWiba0Afnij3i
G8k/td6wOF1aXF2rghoXws19xsg8N82ZmP+iess90y0oNVNaiYhWBbL5yAw4JyYbC+J6kVX/2THJ
lKjCpiQHTH3n9PsjKReZrTN4ciF78AiXoL12gUluwfsldB/z8vKRmKd7qDAjz+7zOzSsff1hM8Eb
5/GtaCtIa6ft1MdMJdlGWlqCzPh9QvACiqWdRY8BCAItnOOLYnAWfZmAOXJobdbzm34lIf+HN16V
FBhI8vrA1/fJVxfB3o27FGjne1/3cafNbxYsM4fVCpzttyeDW3B4zt1Sy3G32Hu1AJQGQqitE2QX
izoKn+aoryO/LERMc45yf3Nk0VF5EnOZi9kTMDf0T+LoaoLUWVoZay/YpfIovZj7EmoJDq+okt5f
qP2T6ykZepp0GNCpV+WBsgyLCX0fYUd9XYpdzMIpj3TafcvlYN6xwEyUhpjzwDCRnKlKwtMgUJJB
gPXSm8QVQynCEBkUWIt6FWDTMd5yFZHQeHkUiFlgKNqcCar8gej9u2GxiTMYh+yQ+JPCeDwKSyUC
fxGw5hUTZZCkh74Tx85w+iI07cFjCGcST6L/Z9D8cTVObzNc4yCdyWwMdFZiBlMZOKiDVA7ey41a
XzPfD8+iiixLW/4oTUiwhHpz02pP1g12k0kOaGCGUSoKumJf+gXsWLHz2bjI4YoJ7YizrLyG9+6o
1euq1reM7ar8qTFkDO3ieJw6ds4p+EeLBwTox8DIm3XJogbHlnDlCbzSibOK0Wtv6Hw9U4MdbU5p
pZr1dvmRVFMdGBGQvshutLiYAyum1LVaYyZtMy46IJvuilPfDZdCaJrEVamNvd4jONtTOQSTlsOQ
mplBDvb+gR9+AA/nMoDDxb/nrQj5Brr+p+dcB1aphcZz7Y9pVvA6Iobi8bPES3zc4D3+6arcJyDT
mNLUeGWA+Q2Z8OW50tfXB7OMV3UZ9sazOoj4sEP4yGb0+sVhWmBo5/77M8T5Ev/4jI6SjuAsrK/r
RqjYQ65P5IPRKHmLi+bJ7WDpPW7FRwC4betV9lk6mAGozvka4l7QdZTTHKlUKEb2NufJOR3zdAQz
AZ69E0VKIrF3Qd0uJFMhnfNpBjaC2Mst6kCAqyIKDh+JWY234JNoacsHCMh1PDG/gmjtCziCnlFC
fCfvmW4NoMAYWvZwQ+j7Lmx+ljQxsZhTKZp7yJ/PXwTGTRYYaVD82Kw1kDLX3XTglY3S73zThihu
XIb9MpJzWDNjF/hWWxAx8kDyEZwBqAPlspw8GUCRy0YY4V/X5QBbUR9XGc6A7bP+VJ16dYx3Uoi7
SnH7T/0hgWNSVy/mHMDuMNcjlOdAl6bDzKeVgUfToj5ZlS7TiUMVIXQz4j5H9bHhBicKCct7irAZ
8FJsfEO9+xXeQw/OH1V8i2DU9UGqYXwKlWOsHDaZzQvW8ciRufpAFJrNED0wCT3dk8nt9go3RAxe
AI6AolWAtCz33w9O0ca/CXELRXtgNlUMrbO+neBaFgnA5GN3vKcTeDdP0KYxRuDPrWN/NW6WarhD
UT5dAIq/Z5XviATA74oXwMhta84mq7ribBhctBCg8IpgHRXm5H+StxZGruOz+0ZtKKJsUjSuWC41
4iQtg7YyjixgQu8o5ro72z3kutjXOqH7UvMhdLyDX4RQcK2AlwKefgwpncq7PKwejrhwTCDgUQYN
EKIX/A+tQ7wcE4O5UNTcARcQ+q6WFBLg1I9uKEcSjzZV7DHkMwbZsK4RrIPw4Pkyx9zkgG1yeYpW
QQZgNGJ+g8UH59TV78CanWWihZzjoXaBf1Irao48QCOGNcWhcL5WeOGxrKoyWn3wSVTSDnMSFOHc
Lu25sP/6PEbVqkuZKHm8cbIG+hYRNARUjmUCy0YnFpmUebOpawJKq2tc8sNkMQevALYqBJDSuOdt
le2KShaFO3g6CwT+a7sVhqZY+0j0WPCIeKGmJwcdsJwXuCk3yWdSliQf4BmJLKee1m8dxwYIzUTd
7ZVrpvAhOBa8JDmyyswULxMLVDc2yE9Qpn/9I8qUz/RL5XC2ZrEot9XOOLcQVbd618PLB7pZ07KV
gVmbSqyu9YJzKaeDvWNnIVTAQSLmB46nl0kXxPUUGn5lC60U51mkkY4f/CpHSqJC2mFtgHMKQ7V/
o4KBqvz/j/d+QxDyjuNfsmHnnCR4WA2vKQkx1FyBrhnFnjlrNfxMJaaUlW+mouKo1pOxU7vCZC1i
GFTQpEwPiopNuETTVmtdDAhSm2IQ6A/e6MCZlAfbEHaqVms/8HpMjGrUuF9QB2cm/03/Zo5ZmObt
YKVNJZjf9R3fFhek9OIuG0w7Mmojd9GdhPwe4RnqVVThxEVavIj86bhlkKsTNfiCnv8qedwBRaeF
/6Ud8Se10NpzERMB9pbBKQm3hNC3eObU1P44ENJzWRtPwoEf5nchQh5+dGzw6pWYbB28Eb2IK0MR
rTEwchpOvYT5NKi8QYUxSVLN5aAgc3bX3XjKm0b2ayugZwZkL+dGTT6VzQlUC5X8qYcArVX/PUsk
zM5VaEaEeaL0AE5C0DJCVXqmFUHXNxDPXIDLmJclnMVA/ww4gjvV4ntKARMoELGazNFX0bOig45m
BKMICf+Xpnz+Z9PkD/D4kRCX7LSEGZ9Cw9RR2qaPGGwawAy1u/h+xcsh1grBEbDMYkDb6bP5zAJg
openfns/qMdiv2hL6D99HLVydMp8ztZGmfe2DkJviMIqUgaZLHKZP+LjnEyZxgxqWT6T6k63oDh7
fZOtrfictsyJl37Hal5Q6bf48dJL3/MR29hA6ZQ4iaxtU/foqeOTuwY5GZ0VZzAPNKxJkbevdNSy
8xqCibVwSJtZPCUM4ZMGt0rV3w/cjMlBCjMV60RJ15DTbCsUay1wzUP3gEVbbWI+dRHqw3SjQlwE
k/EJKUvmni9hsQrSk07KmAXS79b2tbgroZ4V+/2HQ4bd6Kt28dxQrkOf6wDnXGxiF2AYDkpAqjdn
XtdEJPtYtrwbcrsFJOlUw3Mkjsa6f03zJmE1izels7vGPCKXWPfCS2UIcmGsVLU6G8F9dKgWg3AL
RmI5tflaqZwYkf0E0tFu31dh4ibTKOvj+umbAcWVgKa3+a5VjvEj/ie4QT+Xnl0yQ+YwV6d+ogk2
ndi9XvpxNCLIv7tkgqVybwrj+yQMLXam6vyv21N8u0VyAx0Zf+H+NJWf/tDgTVkU42Q1q0DHIofK
eNaCi18abgDqu1RXOZ+n2tv8Fl8BvprRfKh9MmqgrgDsEZr1N8lCHEWGgfnAcen07i8UW7YN4Fii
nnM0lIoHEF8RF+JRJpMYtoWYOdblNCMCfdaOV9SaZNt1WaeFELYTG0+xjP2a3JdLd6kNSrTQSUf1
q9Rjw0GnunFthNcWPGn79Un445tfqD6tOAxqPsrbayZ4oOeP5XyXl9p7xFI3H8mZZ6bdA5qyNSoT
Sr44tvq2HOby+olsZYeGh5gPKZWQkziAz8+IDvEp7BiSgFcn6gG1c3IlJXyrVR8rYHi3OXxrta9a
Ph5wbMG8WY4jH5vVo6bXZlWrsvT5x6s8XgvV5XeXzSxy3p/frQHZw+gG9O50qipHD/1ye8f7SMVM
6Wh58HXLMME7CFn8HHU3Bpa8nGULMUzKt96s4MlT0kqDM77DqKWTXzh85iQ+e4QnOOk+q+s9+aMp
XxON9yfS5SLN9ipJ5T+Fma51BPZOFkY7K3uYsolFcAGdFXR32tWYHmN9TvpNbfIBaS0l5A+RzfpO
8er2622vaVAqJ3yNezkuN16IZ3AxjX6uEjoK+WrYkFJhhuSjPC70QEBtzfuAlvjW+//VvcDVaufv
QUIXj75dVUO+Bix/4kqkSLby/ZCdQF6ioJBmVcgDKngMGiuXJpQ6v25x1FCx0K9sUhY+GbF0W94i
8q7C5iDlrYvaYxoYkWlIzpywt4v8eGFJdWUPH6mk5N3kVnnCF/2zUldykG7IY3nqbSNvigphGIRa
tThePre23W0XF+AhmXyLPfxeNREzjcpqqVS7MpZNR74Jt+pLBJgKcyhVIDgbMJGYlxXHGZ22O7sL
CbnUYZGHCVRnSvGf38SlozmwK7mgCsTq12rEN6w6KMB21D8pwS/PXRe+ENnrZV96+FLZkj1ZQfYP
JaSc9midLKPJC3xQf/o+ldeEukZE11p/LhkBqW8ZRGlEXQGlR6Dk7iI+PvWXlHkCAXgHeicRj4Eu
TOtV2RDPUeT6jGwJUQpDIKrK5/YHOts1RFIfXtpkq9Pm6+xOrRRNjw1ZLXlyePUovyFmITHjhgUK
Ql/OWrPOPXeQlkRi04GBtCryJJC74RgNwa6U2Rsa5oe37uh2W8nvphC2QA6agplH7NBvi6z4YsiC
mD0t7LPOBsEmbd8GVVJtO+BUYzGXRWvNUO5UbvqFVBLn4tCV9+vayWzqiGUdhPpa6ELypKHDNqFr
ZOtlkoP4Od3DulpUAyhJvOfH980uQnc8Qre9KQFk0MK76RBG8vmwHooJTjSMiNipvW84asCBqAot
SZ/RmMQiJ7oMH5T+9rtp3kNLxuahLo5vOyfXPaVtdwM87Fn9Fe/w8R5g/74zIaxGruuK2LgpcUpr
7hDJ9NUcYSG/KJMVTEYIUBOVWAlefEo+S+Q7v15OAbFpg/BTDjF+c0X1+Lfxtr4+AkzFImNmisv1
LSsBmBdNPig+VfVgUw3Bxny6pdTZGSi97w4Cgdr3Vb8vLfejKUrLT5XT1opqR9d1Gw8CmMyWEqRc
ChksMKJbbXTLTXAOBlsl5S5fWOKIy31tL1Lp4+PYqhUePenjRRCcmjcMppmdPyaxXIpp9gf5QF4K
7utmOO9frsgx9ua5t32uVwpCvmSTOtREzXwFynJSel6RsCLTW0Olx4bqh5Y4stSfqRB7cBXgbth3
gMBzUC+QnOIfhWCBo3jRujy7tJSrSvv75ksrwa9JULESRfHH45mYQeZLtU9YBQjdANffNjCTzppJ
yahsZGt5KCzsimnPyCBG99h3z3W57YFaFLtdNX7OyUQKpUGUnF+mEPB9TNEHD4+ipRso2MOfeWa9
WnfpsRYw7owwEpzLrZ2QKYgNjkSr2i7jE6i32CQbJC91Jz1nhHtAYMSOdIu295DWD6i3Bwg4ktAA
NgO2jDUhADsG21202vKDPz+9Q+edbFfLSCj5y/j2U5s4nDq7yqNU+uhHlZZ3LO58N7w05kFqGyKg
bbjCUrA1ej5bcR+hmmybHQKkBQn4bVxIqNHLpTVMZuTxy2RlM/nsvrDh6GvWMm3wwmvEHymdNPx3
+277+n2QlASu+zIrLHgxZjgnNpUYVc3lmd2YjaaCwyKQdqKVYZzQcQQKpTJynCbfsf9BXuIFOmlA
DqIOig4xz3oGxDt6sOdi6BLWCutLmRk22IGUiepPfFyKHFrG4FN3ngRwmbYOFkmXgjDG/w2FMSXr
/lf88R3U3hDsSHast3L8FxAdacLpoMdH4+8s5yd1cIXY1oh4vG3FviKTEOtJ1uvlzAqwMWg8gFwT
l8S5XVsMxSFrTdcLes9rSMuE2syADqL/OLBrZSUQRMLSwF+bM4GRbQ5HNCuZvPUm26bVSJhjCHn2
H6brHlmfZ8AqetVcDSgCGPm5MA3z9kggemXYb4txjEnXKyj3tGrShNElQD955NNiB6zbfqSwsoeA
x3YFI4RSRur+UWQI2LjJunweeosZ19ibA4pRT91oL5eX7l2tRmJfRDw9D5fNERCIIQ0LGvcs7a6O
KVT8ReRNolKRjoi1g3SFFw4kenR99jOBC6gHgWgjFdhplAzSmNmIz63xzEWj3PaLvgmwX87DQBX0
FAzZpj06/PnIc3tgP3LVaRVm4p5FUIpQmia2FRGF6zYO/VNckPb45HJturzDGlq/iMicSOXL2cFP
HpiK26lVb9o4vA4KrKATkd8XbjSXPj31HNuTpm57VX+Ljhv2B8j/5t7z5D3NY3pPMNt25uZlGAZw
Jv83wvP3wHCn+AfgPRHaTwStsk7DbfztCi5HegcYEBrIqUXTL0rmX4yJVRPWo2Fo33kBiJQmAC94
q44afhpRBc+hpIGH9alCLCl2s1cpZT67H+kQ9uMznqTe236ZdGGLrtUmIVP4soRLVVfp2h8lgftJ
IqyZ6PmLtIm960P/RjnVNbJLrloXmHCyzHrACtqbNxkI0EreB4Ob8scz3UNKmspv25fAqdRLcU3B
J6Xdp4G55Mj5xXTENyIOmHZJLQyC+MyDaZRh/OfQg6+DfLJUNQ+5CDCKv6m3WGEPRR0sRKa+G+j4
Qv2lWDSTsn/dQgWuTr+8IfRHK3sI9MJKBwtPeaHIan4h1n1pqhzualg7NhDiU7KJaOuDS3X/dCt+
NZJSwmLOJ17GU5P76XSPo1ze02I+O8vJje8DTkVqJP1aG5FP99PlfSH2G3/pttxGqmMJs95Pxbx5
GgYzUWtBYgABAn1d7HPKe+AcPPgK8z1G5GakS9hS+61MQf9F30AFoGFlB8WgLGVYKNRxDf/TLSGQ
di5cw1/A7TRSrHyKarKy304V3BklLJIFWguD8dT3iCccD8lT/9GlRzF09UK7RGJ5AK7FbB+xR7ET
KHTVhfUkq6OuCdnmA43+GzNKemJ6n9K+Eowl2VAqDPSRxPKatlKfyS+mQTfSl3Al9wBFevn8mA3u
ZFle7AfbHjBTYhWO8uc9+h93FBVDTLaUiF3B3jgBvIeXN8ce+YeBt+4NoFjbk5KwAsFduI1TyXfx
mi2MNQwuD3fODBalLQOpZHk5sJ8DKchNztaH3d4fWq77uv0TkO7s1cZtlByabPHuhHgFa8hEzPd1
IanbOiugZbfYWztoelpJhNu0GytQOdCdA8uKR0QMyQl5nr//kvbrDfF0PZOEuzlLyPPVOoZoG08I
70A8RZvw/ngSkoSFP8T4hXJ+OH1h4ayOyAOVlznoCnCWvJ8KMCps/ypEdvNuNcQ4g72qk4v1xeJO
VLsRn6SxYd8sNgCzxKepGqdujL668UC5VZSK1cfCDcIXckPf1Pky+Us5uR/sTj2KG6VggWFqNknI
BkuYMy73Ul3WIqs7Yj8cYpLuKOUzV8yaIBpfBvA2agPSgxg6C1a69SaS2uhsYKtKiw1cedDdCJsi
jhlqRw0r83y5mc1TYOfBw95tkV++t7MRhIt7zG9rJtou1+bKR5ZIk8o0PmG6XMQ9PMm4GLNpkpL6
v5x5FNyUe5gEiP6VfY4yO1TC/ZEMyq/SsT8bktaeMuKwzwtEhSZJk6XH1jeMZybdGyomlEoGvZPS
z33qsyZiTYD5fKaysN7iRhHyADO53V8O8zsZgOS37X8oGjy2XxvtjKqxf6M3VKLpQzRzpE9fqGtj
6NUIDUt1oHlEkfvR+jXI0QKMYuhjEdQZ140zaBfjAILmkWqpkXJhdn0Je9uiss9x/r2YsGwxdKI3
4uyysbo0kEpx0wUYpbla/AyZlPyG7KAEo1WIokji50bmr4QWPWXAwoK0texKgzn1pSrO9PhRPPjn
+7fDNT7poBLBCOo1SMhOsQFYaRjB/nFsv6bKYdZ+Wro4eGiK5kL1VHtv1k2PARtl/IVt34aNX7VX
w5FbdSLZQSOxY8QtJUxg2hwHPyYpNUvXcjaFyRmLeQ0BVSIBcpH/DSEy6jfMUH6kjqeyFAm+HKLf
iZw/ZfdTL4fkAA/sVlMILwRjhKaFnRilm2o39NCCWGAltO91KE2TNjW3mF6OKSYAjmO+O0lomNzS
3wsbhM4KxOfQ001zAYCMjJHrH95zM4FggUTP75JwS1jj2t3Og+LeYVQtGvnB5popK1CmXmxHBOL0
q7o776YJMIfuDDSLwArTYyblhhIHSfGsaSpu77X/SfpEKCjTOstgsINXXyV8r8KF3+tStEkCkCxy
ccIxktcn12lJVZMJ8dxz4yvGlCTJcBOWi1P7+31kTB1l2iCaNISBTUMmCJjcUYd+MZIW5L4GrVbA
RqUjcx/hTLXm6iWmgxNz7rYQ6Hcwl9Eg/q2qs6ryGWfn5SVod4ix55OQAhq8br/sWcBvn7Eo+Qol
rPvjT9kFM+lt4sq64wtPnBOojSj/W1QcbPeSFtT5tjmyiypTMDIQdk2pvLa894sv0zXX/MooCjjO
l350/egOh+yAK172IQ00IwwNpAbZf/X0NoWVV6gQlSWK3oBsEDilmXOv+R8cd2Xl3x7gAHROhGrN
4zPqsKb/FjON41JQ1KEeP0LWNduhyo4VgUsfJsvyN42qNNg3N+UuvjsXycopZTmn9xlFxpDt1xzR
reoAm28OTJIY/HYFlOhIX+jut8Qvz37TBEHKjnwkcNXkwSaqIBXsnvzSaqQi07ENsP7Db/3ieiOn
wYhPt/IQNXCKaT+IkQyzJewJ7cgSlWjw90D0ktLPORXfkrYQdnnWqZ3k/nWlVhvI3JoBmN6uBfCO
3dWt9z4dtFu5K8tBfvzjng9BCPH701XYYo1c2exOOcsleRK0vCZX9r7sW3VfEWZr70lGx8WstRta
avDOhB8N0JH2xX1eA1Zb6IkKrJWvvEOCrtwN9dxdyIYpD/KKzRfxC1zqHzNSuAZqExjJ1wwo6MBk
jDA+hGSh49oTIiK5cHWxJUSa4ABg0JtNK1oOVZyg4dblKtKPNvYp6JX0duNkV3WIImbfdRInYvkp
04R1dlVEnyUjs8qHL+j6Goj/6O7tOdRIIa8TQDitU3Us6/AUbGJHQ6WluMOCb4gaBqhJxWJRxN6S
pSHqNcGskRv+vyOpfGm/UqRuRCIjUZ+Opot3ZPBCC0QVUE6/wL/CHeT5Cxz2PA5f6J5ZDqFr8it+
XmcAfRWEYJkn0h1Bj9wv8EnR4lusGjxxqpNB0dEqV5aXwa9L5o0LUP8+AhYrRVAkBFMOfxliwHI3
7wTpzlvAuFLxf/s+lY1/NEEqR/JBR8rmIUakGnXC43zvcx8lbEUcWeL6ToUMBSRqjm2TgwitjOWa
f62Mr/G9dfQ5ReBsf8y1+Qn8xfdvECGZvAWh8j0P+plWRPgoyVs9ya+DfiQKyn/NJbXBu7nsZvE+
nfB5FNAW5SYDtDmMSGxvcm8qSVUbNqyx5Uhtd56rmdzCOW595EYTL4Veb8D1ekiTh7INLv0HTJq+
bn9gx2yCa12n4sSfSi6IpAPjqsgHogmY3OdUuIlFY6/glQGBV3rPcULFgL6fvV0NSbGfwQV3b1tb
h2cAYY9hRMtxuR0jGnwU/Z9V+crCm4pUuk085uUe7RX8mP3Gw6yTWc/hViwelrpF6Prjzb0XpupR
APKSt9RPfztpvzYhsvYbRJ6/IHK0camQiqhFHVIZERHskzcUu3FgrcDdqFDjdzFyxxxLpXyIgqfq
wokHeF0kMqMuC9ISC40kox2YDab8dERiiMkj4GZIOj9lQAY4UEx0aO02u5JB8T8Yxhgj5awv+BmY
rCBoPE+1iW4VMqYateBtqdgrMpgYfeW6fJLYWbS6WXSvPmtg0WjoWibA6oCAbbdHCHdG2x7gtmtl
8cd8H2EvyBCMJqVgA0d2bfNiMH3ZpLH3VWU0ovoyDn77soj8fsKlR1ygFyTjJJRvw4DKTo03v3m9
bwUmpY96KBBTtg3ArheABXDNssKeyUQPeQO7NeqnYhOwrYaz1fWg7IenMvgn/COHcFwjEJrkZkev
VBapJ1PP15f5NKjTyFQrSfh1xUjiv4tkpo/a7EAVwJJFahPXPwnEmxTL7Tf+ukzMFKprTIp8I2RA
Z/eJqzaj6+bZ0FFlpMXNEDxX3Ju+3gNbdN9JMZq/5PGfr7vBS6vaxQIO/GBz2H+OR7vKk5T7mFSb
lHKN5wkF16mo2LAHyOatOToriQ8fpy2O+Xn+KfugKqZSyu5Zsi6eGK476BcfysfzEduHaReDPPSJ
U9ge0Vqpt3U2TOpkYJSZ9Fcqfd9apiG5ogYAQIZqY65VVEoBtEAYLhO2oQLaJarCyytifwJ4W77y
2QF2bvku6H4eW1+3BkW2djEa4kakOXOwywTAUaPzOOTOuTN2rZ7DG6vXUI4D3b42sMzAcXDzQrAU
OryfGoXAxobrc4+x8PUMzVfgjex/nNrSyK6GBtu+1VwY42m1Hzzx8OS0dSrK1/WE9n2Vhf0/KAVt
PSaFOLF09VeAvfC+EfCJFYwQG5IrecaHixIJvDRske/FQXKYYZj+TNu+vqqduq94vp03Rbj1I25r
ELBL33s/fUBDEKvalaxJkXMBKeZIeOs/qfNwRE8HnLVVkDbAAuJRU475GLyov/OJ4xZUFBjqi+Xw
d3MipCp6HaNHIFw8me0yxA/uAKIHHbvoOyAj9P1736Sbxb8EffIxBoiyJkXKICYMNHQxX9S+amUj
VuDR4Z2NH1aZQTpRqyDe6TA5nEEd32DQvlOL+AG3Y2YtthZroPs4tB5UQ2OdTgB7xtb757JJHKjH
g0lRDHFbnYrkT4zEwb763GLrzAcbCDgaoVJow1nNxdqXhiekVOByq2LvzEcLZ2J5Ysxc8bbQnOvE
O/NvkTNfUDWdstdwK40UPfvtcA7Aa9uwV06XFkCsY+YljZrt8jnmtuoCTycU9JoK6MmS88RzdV4G
kCI0jdvpqv+JquYlyecZSPbXO9UWJ08e/yt/ORGLPsdndBLpWsdYUE+74okVeP9roSNWjDnJA+cN
jj9gVs4MKpIuqb33eRpf487RZGDGWl4LsbT5JZ7jjgNGlllZPnJ6RCdqEfpzwcPjNnV1hx+3qC2f
D31oPh3pU4rNqp7kW3Z+YDqlpoO0a0Cy7+liptULk05RwiPUaAD+g4IUox57gfpsLl8qbCQ1zN1o
Aua1aB1bwgMfF18DIZRE2hM0cHya/IYhzrXDWlRfB8z9IlXZtpJqQCLuu1FeOKNYtp4+avqvOR4V
kCeIUxAYCyD9cQzXbUvdeTNzwoCigjQ2XFvsVSCUXQgoLfFnXvBZrQ/n1//xE3W+XtAG6sgykjGg
lOXws0hx+GYxsK3ft69ZLvx2na12dgtxM2w4APIngxZjAmQ2089/eUivoGZgm8WuL0O42iC9iro9
Nn/TlhaSpEzOvYH+KBoPVdXMdoNq1CGPojHUUSU65bGiZ7OqqK3QmVa+3CZmgtBf8WyKXp2CoSSq
m7ZHqn4T3cEdgxLNe5mkpEvaJYcc1mnCf2ncILX5obLa3HHcQl/y9OewLJ1vgT1PTYtCs6xLisiO
Nz7r17WDps5ypeZXLdXbkLDlsxyQKFqPtOHU9afWvJvQrCDosHoBvIsGrsNM/Pin+Jbpw7SEvFUT
8Sy5t7qz11o2FgvTkn1LODDI2ntO4tZAXVipi6tZwQhEsgTjD2AeUkBRQlpHw7hw+PNOtHbPTMDp
RJbL2OS7xVbsW77G+mI9GLNn/x9SDOOuyX6Pv2gcHavtcGG4t9DKldSHh5hBuJuDTQIo7Rt3aZeU
HzFJFB9VhRYVxsWzLo5mMXkH7TKBeQ/trS1den9v/6sFpBLVSiqE0mwlAI6SZTcjGmle4n5c+znQ
e3AwhwzDwFzuOLl/oeortOXv7CzdMi7EgXE5Rv9XNP1r1wdQJDABYAaTg+rRGnCW6TwvQ/hkMFzs
HGkVqZYHLMgLcxNgxQ0D3qqGcMTW6yk8dmNRA18YBW92u2KKi75J5vwYbW1GSjAz3nNP7iHKoTe6
0xwcHGCn18Kqc8L9U01QHmVwYh43Rh8nSOfLcqN0wtd5KRkZ0pMDKGXjBpUJR8bxsXUXuL3eE/Bq
s5RvbeJnuZdboSXr2IAG6xUIi42cJsERCLjaP9wE6q6MVqEnBE2td/kqd4HMSNWFHMX8vTWiOV4D
LVq9s+yAg3d4xekK6rwMjuFtn5XW0GmTCVToabqU28WU72YEb/SF29JiJGkjRok9j0edGDfKYcYa
lNvwxqn0aqjKvZuEBPMJu+OmRORLM1d9/Q1CJl+xHiGZSAZ6pTJJ+s3wKenm8Kq7JuD05aufc1uv
oxbMbOCHQpa877DJGf+m6gPmQ1wSh7hLW/q8MaR5taEvZpi7MmB1FhafQ7+4WPb1B5b/DQqvBBlI
xk0UTXwX1NjQGjJoykJTArsqIgDGYvdQwNE4JtGGO9R4bFti4Mc8WlK1qxZaQKu3tbpOTMEDsf+c
W95MAywKh6yxs6+/TKZViVXBV4iuWFSeu0o+JdDPe3gROZZrmr5/gwF4nwxb1UctF0UEbOAxUg2k
KMn8q1WToeDHSVCWVBNtVvNZZ+OAYz7MvT1cMMO7cmBWqHeV7Raip45jsn/O/pZCc43E2JvskOdt
Cok2tsBOTOIIH6UuBddieLQOsZZbPMW/bkSF0Fw9WQCCJ/hXCectEhy0eUQ1Ncv6N36DkMSPFxV5
eLh5BLCPib4Q+d13rBSpso4WxrHBVv8Jdx99ueOk2OTl9YiN5N/nlq/dxTtNJfLTYt0FnyDyYb3g
bvtN+VQ2IajKNeayUVTT3bPb0112CspUxwrmqH9FhutpEAodI0cd9xvYOEp4Eb10lFGkifY19T9U
thHhRNhfjjAzfi5auIDG5YoJaX/NGRntaSzclVJdrG/m9VQkZTNAMrXF9zvCdGXHjwf0mqnIjsPY
ZglxzD8WMmS/E8p9uKJ7vME8Ug6zhKHXGIcMhe/iwFJVTNU5ljdy82J/okC5Pv2M7IwLxLZ02TEF
JB+Sqth+/WyW7YHnN6Td10UV/jImop3a+lSxQW/3M0aAzdPIzJNdbHrc70z4j6TNdVjYoCJkRnaX
ky7s36a0KLVi9sWjDpo5Orvg7KqAYPk2nd0SO++an5PXCvcPm+wd+ThH9mBBydiVegrTTNUnBZ1j
ia/1AaCuyhaSX1zMW63nrZ1tV6AzDmyC/zxfkArSZZddaG7jj4S80w+pAu4yzkQPa7zmyeyKF+FP
0gTqbFuu22fl/aPlfRTaDyg0nh76F1FSD8qa0jtiCGrN0qAc/K0+AizuKgDxcdb18OQQXt+gjvEh
YnlWodbYV2XkhpEGsQe/ee7OVu8sI6yTTbWEg2Go+ymD2HtMuHYgtqsOp64EQX+K+xpNp+AkmVrO
LC6TKJM9HAiO4SdP32Rs8p+7zdKlyL8uGtzCn1HqlG6x42arHOUKPV+ps8DIddgaYpK2aDJk2oGv
v8U9m95fnoFF4IJUCwutH1rz1rjCx6OrF06iFS7Azh+tzUUpregCACr3Zn3QuSYLq98aOM4HZ/uK
4M6+AfMkq+HfzEXW2uODPzH1d0UZYoLrqDx48Tsw373T9n1HHB9Lu9RHn7ehRM20KJ2JTjDA6pI/
Wr1fIsNqXkyp0py6VTtoBjf8PeOMrByjHK5vkiBDoPrT/QkgmgtVDhKTH9mIL5HUJKxbWjcY1dIJ
ikQ5AqGLvEDSokEIRYIJSjK+Cr29aCXhlpGHyZEgvNzkoqXe+JpGcn+iVBUYdmgLsQS/LL9XFInd
Qtii2kwrW9eHG0Il3UZSIQm9pVk8SvrjTdT9+qmm6RKWlSLQ+AMRZtMAVJuxfsAeTQBm0FJBgdD2
G2EGcHemxxYSqPDVXsffpkSeRUTr/Rc/B2WaB21NYEtGJJvOZoEQFSRCppJJNeNYDyXleu6MEbDX
y/wM+iXJbOJxeGXCoyO3aQEEUYA/C5SEdNngND+LOdmUU40s2c/tn866b3cijW+5v49uI2T76oNO
QP0iH5txq2cuQUHsaRRKAjRARhHZhps2uC1E9UHQNVIIpOPdTvJHVBvK70zGibfnuMABciZEGzZI
nDLGWhcZu8SWIQs+82Efh19yT0TY2dZisur8NfVfqwi9elclRv75iYxuUomh4QVso6tHMGZfAeEP
G29eYsylQwwrmAi+zOELUXUuc6SWB4EPC47t6md5UgZZSQ2d2cxaRxtmSVvoVxnwYDp4lQ9fWT88
2fRqsTC/nsi0C89kRSzI49EUbCxgzaLVVd9/VD72qloR+z9C1w9bfSO1L2scgNAXS4GlSRjiAjyI
1vd7sIJZsbnMHl7II+fJAtq7vXAKknq6lgpzMp/vut4gvw5ITas+3Z3wv0lfuUTKrCW3R/JszW2l
iPW1IFLgUChU+GAZZG59lUPXqoW73h2BmJ7HQm6sWqQhQdtl2QWpiHJl9oNeK8MffNCLYzaezBgi
SWsgnyV9y7OmlG9drGZMYg116EAZms69UJuEEtiZ+eRA/CS/wz1Rn0gynDFAlYZRGxS1u2D+F69P
L7TwTMj6xVafMPyehOkweVnPYs3iNOWTNb/o/MRkyin3IVPMDjmXaDLpOYKgM6NCANOkQ6apWdE+
HOAEXGGVoUfC37Amlmm88e1ZwkP/Zf7ugfpjBNCAbObIUfhjNvlDdsJ8FyBDs8cSxfeku7IIcA67
BL1yu5mVrJPeEt7yuQLAti/bmOXWApzGSjkCUEeBRzP3/VVEmZ+pnkJRzKwMJUDAzoxwrMIAa3vl
eeXOf6GU2coI1mrQDHjE2c2iAihA9k2EcC2lBxCRYSHj/qxuHMP39RFUej4fIHXqChotFeHk/LxX
8q+erIP+yGjEBr30VNx1hY9fc5IPCfwWSGC2/W9AtreZyiYW7XZimvTNQZoGo6jBenUfnbLco6PP
zspO7JLoXjj6S1AX9CQ1x+zN4wVjn5jfX7ZJm5EGIJ6anglOIynM/VEkR23un9UHuGDaPlsVDKV+
+Uo0ogpnzSdRUS2+N5irV68CLBwRcO/tySGIloYK1WWNnC4OKZ+N06e2JhHqVDt4yces/Hq1H0ha
Wc36DwVGhgIQYUVUJyUnS24tv1zhAglAmuMJ03am0mf46JIsnhXWdFR+084BMDhyyxK8ERyLJrNO
cQPQ4dzOUDhiXELRGhYIWBQKtiXgcemfZNxg68ouqKiGTQsY0tuvdPXQBKC5D92U7iu++WL7vMG8
Ht/o8aOI1SNSNlFCykfG3743HJ4AmMWMnrbU16gNliHMBVcrOZ/hxb/R7HfQuCOddpQOMsY1hvdM
PE8xxmUgiKSHBZB5qgVkrTUUlgB7tV0PdiVCL7CExTnhR7EKSvmk2r4Wqq5QRfT+QfyTuSqwcbvN
rnNJWTbdISyZ7MC6E8Px0/5gJpJ+y3/NxZFk4zX6+2YNegPfSjVqZ/9wypnB0y0XdAgMKdsPnVDS
UIFbYo5eAl2I1rd86p/FbfQuaiNkeN+Msq8NSs4Z0f911LiO2CT2zevoQ+/+PmDGdB88AeVkmwDA
NgSRhNtQh1cyrYW4zX0y9U0mP3iuP1xXB1A/OInQ9ixqMrhwmk8Eb7aDVP9Ndj7QiG1NoPAAazXg
3AsN4gqxI0DLHvjNH5bguznHK55/T81X9T8jnmeXCdc0EyKjACtAf4LBcUvdwcKiuyAV5s7XVlwk
eiZ0H1UrlwEa5dunopZzYZ2HGnLO3QvD4MNXZJMpwFWbeEfCjrEp2UNfpCtLrejwkNnXxDXm8SpY
CqNylMjwO3H2b76do+uyChtCsfrAIbLqbPHWeu8+BXi0XTBf5Mz97rOETzP03YUPykmFQoB+l62g
so5fU2rAWHfrgYlISgMc4Gc/4twJJstTxlMiif9oq1i6T8QO5IHXSlxikKQcoUTiQeWZuIEraFTN
/aI2ONk7jWtcM/6QP6H00N+8O99ISsjy3cKq04OTxbvcM9GVpqe6Bk7C7NDZvof5ueV5HucwFP3l
WIlfDQ2Vtqm1gFTiT6zHcU9DyJY4EjNVkY5pe67iY0oeXTufaakehd/ymxSx/jTCUVEfElkIpR9Q
CjkmF1BF7iALpTGH4hWo0NpA6XH7j/4iLECy7q8q5ESNpN447c29VHDZPo44zxEOtZX22XtBDB51
0tUcIWbDDC1zMLh9OWtI2pfXTl519fna6kDDCtCudCwdTa/KJOGdK5jPV7HglfjW6GeTNyRRSkQB
SxHuf2tbENH7+O7fxI9qlDPsY6bsZG3Pa5HeWVrwMa8wcVsjIz1Jkz4Hw1Y7dk0N0zH52d1hU5tO
TYjnthWE/a4S9RJOYX2nXKuSeM2WV6CmoUqaGwJzi1ymcMi+muF90Gz+NX9tDEFJo1MPJLuvkstV
4iiuniKI0TyS4S6a9JgWtcwnlV6C/Wou2XFVRZe8JB4+01N7vILQ+TcBj2FjfRMxQ72OoeAEkCaj
Xv5AF9XTELKAAj1EXKi+dBhkpEOT8I58ziD5wuOqk9JjY3H3Wx2pQnk/hgAucsNwtN6t5KUkYZgs
4nEj9mwLLC0KbsgcaW2Aw6iMvq+6X8671eipyhqlOyhN9KOh0rpbnC+ILB7sVAo0BUmcAGCrGH88
9WloAfQ/Cy1H0LFLimz18Uq/1e6L0k5useB/LQPDeThKFjgBQKk03WpPe9T6rrEaF/lJkP5PoneU
5+AwIYZmqQ+4QRxzykOxdQv1FGBSIoymvzAKlzNaY9mWVPKl1TAIswwQgjod+oDtU8lQ/ldDI5wR
ahEnkMkEfV/B3e0vE1YLLzcbUGUEDsJQrk9C6/V75YuaWQaJ5awINaB1CMKyIMsdGSdH8Xe4UvpY
X2j6l3OPyT4A789j42Ebk2Ma0Qxj/MqhrluuQWtTL1GZH4X1z7BHhZ+OmX0zPRLjStcoQPTj0Dbw
FWIBzphHkAC2tSxhgKzLiZqSxuxMyB/qHYfVDiEXz8tJbiChXOXk1hlJiX8bqFK6xSWJW9kOG08u
j2JSOxdHjBzW3K5wKpRm+oEKB7+G5oToQ+uBIJQDdxa1usfka5ZtCL43CntM1o5GcPyk+2agVW11
Exs12vet6aTuVSWId3uYFvI5WvbMkjHkc8I2+wOe3ZIVb89em4WyyCkm7qJFWg4vpOzB65u9MFBB
1ZHKwC9muvfyJotOPcLUua+s/eMFCFpv8N/oq8HVpY6Yq3yrrbSrZei0SVh6mnZ42DePhbKLE7W2
LIA19JswDxsC8+jI329GB8fxm7ZkNdcVFHaJSRY/HmCdNjpgx7K0IyJLMSrc68/S8ZTUlFd82qHF
v8/JBMU5Mg7/mWbjmk/ecNz5AE5qVGmKk6sUPaAH0EyLZtHa1tAPOBAcMWsJT/t1FOd+Mw6hFQFL
ltOEMeXV6H8xc8g+l9AmaunQGfcCL/mbZe696HZJaiM3Z22Tt1GcS4op4hAj9x7iR4tqBBf6GamR
oLDauAkyZfN0CKhQ8dwNsxCvhuz8Zrx1oGnmUIZizg8p8VyJn9WE6eL4wdiX6Y+E0Gcv9vz8Xxr2
i/2AJ//ICkro7w2NjSvNaV47AKFzrkEppK8+RnMAKi1SIrATTQ2smXn+Lz0wEzIUowffvUE3L9Vw
Cm6YtfPr5vZY5Wo+/pOBGTqootIKirypyxgSMpirF/SE+ymjfaKV1o0l1Jq5/t1BtkKicf1QNAAX
MrsE7Z9FhxMEvpyID6jyFLmrXho5Lp8DL9v5QnbZV4BuyMkImA5oM3oqLAzdtHE15bdDTICInkxH
e9I2WZk+dSyVlZuj+ZwmwY17/GRIwLsZTkPoQDyzYBaKnVD87nRFApYPE9uvuytVO3YBwzZ85EAU
icY7k6saeiKxLiBoy5fwS4dhLvzkTy9Tt5s7AP6Z/G7kskReK8Hj1HKCrG50kTSqdH7bxKipraXO
xAD2CL0rvmgyGLIh6GzUykZG662tfu/6P5cPLHaJY+4HlzO9sFv1jwxP2JHegoUtly2v2z6t8ZPX
nkFaopHXiCTPO3jH/z21v67y3yJ972MqVTTwGJU+yrT+NNkk4CFviDwHEWF2QACeOcksSy/MT++Y
m09HmD+BuSNweXj1ZJamsuGMTYliQ7jL9KT61bvqUUAl7IG3Qh2jFaFTO1VGwCwzOyLVO9y6FflU
Gx6LSwjl2hlElHQj4sr6hCgstpmn3Hsl6AZcJqemj551vzf9S+IJoTwhqqUExDgC1ZrVWtRLMppx
lPwbuQ057mBwE/0mYU6Due4SUCEGq+FP6s7Fcvfx0I9VNhr9kD0cRxVndnxZFnpNZtqjCc6AMgla
/9h8iFHEf9Xrr3frg0Rk/l0Yh16lqZrb6P2kfjkwUKXZAQegke5PXLjqSFc2FnKD4RPb8O0x+jcO
u7+QQ5gLazToqWLArce3wZs4LhfskgSHEUeYztBdgnX4z+h6y8kVtlc9AdrFcYBpqQ3iV1yeFbC9
1ebVNpvzhXPHvft1/cJ8yWi3MgWjv+eQhXzF3XpaEqt2PpNcI0yM6t2lZxRiArjFflFB+P+E6evV
OOxSVEg2fIoyFkccJxH1EOH2ONyjVUIa93KZpEOGWOEAPimQhJcE3ckjmBv/o1/UV0J8uNsIh5MP
1R8pgNZoF8Dd9/3zNrcd7xgl2M7w5Jm2zoa5Vc7EB9BSzQPLWcgVIl+wXtQac0qQpJ2ZG7cGTybP
2nNN6GUIFXo9Is4PqGNl7t+JbUeddjHmqU543H4FjQwwijQ5xVPEaO02Y06NSnCV4JPvGzHP5zm1
qN4QnjK4m3Uo/KxNQIl2RvHmnCTXGtMXEErThQGrxUjiVtu2qnhBMy1jes7KX4s3ksixTjMD7cls
tUG7B7Sbk1r81XombnBV9EGqY+DyzX3+oFKSOt/0cpLUoX2/ROaai8x2uewXtyl6wkIxmgYGC/Sf
ETzYTwcdDMy84dmzFOnJQQhmzHOiU6MqZaECRjbAXKEJDn9VoUtR+1YR6H2/E97buUbWPsM4L0g+
hoqjJ4sfJUBtGaQtQe3noL17MxkDMtMJaRiYq3Kp2x0gfH4WwRUFlgXL/oSA9JUeNNMQ3b8LMOO9
0XgzVbEzQnRZ/MSP8HAcbLhCL/R6ojKWwJF0agnkIekFHohxxHEI3Oo/HZ/u5vAtQGu2umIVWtuT
nDCwkTQLNfWx8dyl60lTnxS3KzDNFZSFFkJt+2sbtdEjBkDTYPqCzdivjKiVHqBGxUT1gywn87dz
0E4J1eEjUdUmgvtKO8aX7AQWr4WDnKiWNvvpU/HI48zBkVq1U3Vkg7Feh0ZP20cHCat6XvOjE4vh
Oke1veJ2w/brWBjsbxnusiTKYDfFKU/CmkuFAT3VchjqtRMzYE4ljDRfDXhVvfevr0Pn41KNSBVf
Wm6v/s4ErWbvqAnV2OhSvqeymuCceGf8x1f5amb/iImchfG03ZXY8TuhzTZnyr8Io6t99dp5jA92
/xdmq8SXX4ucPD7gUiUGdmGJJldQg1QI88/xhc2Y+KqUm8N7fN4p28vbMbBMj7hNeTgekSV0pik7
OKAf5yPS4HC100ovK1WOk0hAHILIDj5z7swRlefk2i7A1PZGsnp1AKvBMZnmMRD1GWUyIZsLxju8
N7z8T0TZ8xmLHvbvthWQNOFduv1Qb+v8GubpkCFG0L42Hl4dsxsBpmt5l7zQiEvryVXLqUNXMlz6
cSgbupSkN2RIBNJg0/bYTbmhyUPG8DhyaPnbtNNaN8qMYCHjEhRP3bTAJXtuOZZGf/1AntKhCZa/
h5349FO8KDA0W5dctO+y9QPsZtF1iemnLf1Cn7kYlU69jqNuB+Gbnl9CLqo3ZVxVsbP53zFHWUPi
/yZL1C6WprHmYxoz9P5Re3q7MrvKkJRKvz+ZIDXgg8VxKMjOUy2LgjNQfjfQpOlhE/kI7hjNIUNK
DBYn6pzFY7valVuDryUwxhmuZeTHw3PUpy6NxPcqZ2pC8PDObMJvM4ti0uPigp8PAX98z+CAgImO
7uEOj+1QB8QRbOykVZjTG6eNRqSmq2lmUJVHzFwO/TQJrTGNXY1fydgakIDOTJjXpb2gkMQdTizq
QPT3ZGigkGL1aURtNQJ781QsFCA6pHeI2qqRUFPdbHUsRd9edotBbC1sU42SazTHJZ9eWPmjFFBk
8ZG4yP1coySNRkRorQeQlCc56cYU6e/OHcqnJW5e+Ax2/E9k+HPPeLvNfEUdQi8epJ8NovK22HQw
Nbv2jzghHT25wE03j/RQtfYph5qsGlYewL77GDL+4OVK3y3rAnwdbRtHYQJKoU0D442/6WEABiqo
as/Dl/2+LJGhg6mogBTSTPWSKt4qNlz1zhmZzLK0pRGUQ88p9TnY9CNabcqG44A8bWjwzh0ufjvf
bwC/SM9f1y48q/Om0JKjrb/79yKXxAUyzjKIv8VtCRpN4SH4U1tHXD1kqIbE36apRWplZm4WLGuK
AQMBp5eYc+y7dqsCXarIKQUyauX0M03K/yu9LsBYR5URpk3/szci+fQm7IiAeabKKfZPETALgKJP
PhL2WT8zMxBEOkB5aWEJJrouA7+KHUYhygR9tmHKwSYvuDsBWjCZweqe3FzZmeCUEVfuddfP/sps
eaC9lccAjYGgDTka2WMYDCpnPTuuhK4RN+a0cRvP1w4aRgLjgpZGfoFCOACGS/8dEqyJU1GNCOoe
2GK41zUpcaDH6brCOMvuKWwSZSTaN5FSl9sF1MSFgg38IljfxsHaPg3XvIRLxgJaRiTWwH7f3jdV
e2kc5OYwAXPV8YZpHu9/gLteL0C2Wprmjt4+5TuClfotkhoKipnph18bGwdEA16E1VyzjyEd9nhI
ChYKzwQehfHQ2DbTrzjdHUgMzg8X0+3tnZS7y08nRgzM4x1piWTqnlYm5BH4p612UCybfpiUo6FE
P+znoPM/WZAc+bdqLlM3RmWrW/b5vcP+aA/KglLOantlFa69YqTKaQGUn6dwsyO313UJmcBg5pOw
6q+qkXdAkADEv/zbDWo+XYEUoAPq58FxmIdd1KH0UOie2JZ6wutJL9r9eG/UVwjrVG6/7nioyPcI
sT48y+gmX1Bf3oPVwl/K/XS4cFzyJ4fCxwl0lWXg91tuAjw8IYCDESBBtwUIAnx/D1Psy2YZE96a
nns6mLcHsTNZqSepTS6P76NQjf730v4PJd1dAi4BeAHi2ixtL0w52BQ9pRH11BhC6DsamxzUpzvM
lGA0149fwGe8y0KF99dkxpx/zusezkD1CDilxtIuKkkzu5VfDXrsHw3yLiTKk7/86CO2bvzzAZeM
sTt7pYpzzOMSnuc62WB1cElNtzCragEtFUsrwRSRx+4OzB80oCDydhYsHQShjoaFQHQVxwXXd009
2DVZIqM2c2Y+Cu+OM9r0NQ2cA/b1VJJOQ0shOzmsZaGcQF8DeQJp1gQw2Ln4LbnRopBGBeRJG9ut
P6ve5NbfYqOGGb+R8LzKPHtkbcakgn65OMucEQrCoimMR1ZZTry+gkz8fk3LW2ye1KZUGkxwJgrP
Ey7e2fhKVjoER3XHA2wiyf28L0i69FF+tOSZU6+PrzKbYClFfVs5z7LuK7UKrQKrWfvyN/0RNLPC
+igK9dIdKHIAwb2GxDltk01beio2qk6XWqhJxztD8A9iSlOyZ/YPKdS2ul6xesby+nvvIecGVdv8
8CwNllnnNt216xV8TH3KwpORa4rs+zGJdRWhVewH0e8Yg8Xw6wOVNNK0DAHxWyaJKmvE2bKGTRGB
5/uZS3xEM7Wt50VxzN0S3CrJS1NAFPHL0znjhTrMngt19INNWxussBpuq7HhXexOiWiCkVMqElSs
jWh7yhme12Ej+IelVFUn/b375pDpQFeJbETRnUAAhyGiQHS22a3kDuE0r1e0FH9HE0Z4xGxkOSMG
iuVZvgZDrmF2zYLnuqD3LoEMZWPig17lMBSwv0mRiAoqVpD4sQDTsDt52M/wmz7OHM+UNQAJVNH/
/ZjBCNS5xE5zO3E2hdeHirRBEF4cAYL1WUHdA67E0++D2UWoKIdXguquSmgPNUXlyY+z4sgb8xvc
Voj2kTafZ5kiCHs6Ji5CIseWmBgv1KBJ6q+GbzvPfcNfTNkr5IiUrYRJPxTeMSe7bBrj75aX8MWa
38txn3r0QkNPY5qohWYva5v38vRlhz8VcKbenJlilZ7zQNoBTekj0UR26YcOaEyfKVCr4BSObwiy
SChH2AjRiX13fN97i62CDxYx7iKRcI7p37lYrUDhk2NyarYTD/jOMOUK04Vec0ItQqujUrwZz/O8
uP6F+9rHaf+Ywx3+NjLdas8U8P5OnuyNVTY5NtuVf/Z+XEU6hrcQ3C99z8QRWxUHW96we3nl6cTG
6MkFw7ApXIrA0D17lUgdvR9RewO3kijuOM+oVvBR/5ZSJLjdyILdzKQtYeeperiAjP3aWD80Q8um
P9ECuPqtYpJ5bgZ22VQRd2RNke+EW0jsqNUxC74qxyuDTejSoXdse3cM/ONNPE9MMIITbOCAlqpt
h1oagQnDAMPMhriHIeBJzSLjh9fDvYLsglagxIDU6MrwFWsWoMIGIBdi5Q/PLtPVP+XXrTbATaGi
uxuflZDmjMkX+6fmeUok/ZzzL9i/qw6Aa+/FqE2t6q9O/nJRRfTvAOEPKueS9/fuenLxek2TvEQC
HpnRaRpr9oPI4coMOBtATmss7rpL1jewoea0ykyK8d8Xz3dHYDP48gnT0NgKjDaw6od2jdk6F1Jt
7QMgV9B3x6pFfbb7oWkHsHh0eSqpO7/dlVGA/Naff2C7jgvT7DsDHUvgE0nq3L2VbEATz6q9GzF1
1oW1m4PHeJYvS+bZJJKune/pKLP1f9GEAKnW4+ilyGPj4dQgKe6jgWba1ytaP76kIBc+nk8JUC6f
qG6r04hYGZ7H7y9QXoyZZJrmG4HuN5E0UydSlc2f872Kp6Gn/DQnVadfhF7slErAAy/ZQ3Fb6CSf
711ADdjA8rnzUenPcrmDprRJ2mvbnLYmJzOfZDvOBAuHTJUpr42zYKngMBDkTxhejbJJ60N8v4N0
l7MBY53Uruhph9NccJhT3tLbrG2OZHQI8I3dcnKiXuI0jK2aTEyAY10d/PatOB12g983szXLR9E6
DAPKm/47O+prWFu2+MXuH46Yz+7oLNA6c39DmDRiKRDp7Qf/6DElBlmnnWT3sQu01xxs02b/ngvo
z9DKr1mf3oEf1di2xrPXLRNnpD8Ytce7ikQINyYlCaZ/yDE5uiutAMC36TDhUZCW9YmU/YR9XzwY
LNPZRo+74lZ8mv+YkmXE24VSfRE847/VBVmBph1lrRexdkNCb3AQFoumPf8ALSW168brKmQKz+CZ
KZLNGCdEQIzVsm8T5koenRRbm1QbCraNFc8fr0Voc0JkCxcJQMPcmUenDJTNGOP5Rg4iGwEgohvm
QTSC/8I1pRYcQOOyTm3qO3huvxDL9OQjqnN0FQX+4eLcoSzD47k3nGWo5sbIlTba4FEZVcgQWWTK
frZPg9ELdF2QkUyOKduZKLIK0pupO1ZU92H44vaEH5zDhVsGntsBzbN6EU2jcCb2LohuFo+3Zcvp
/aR5b5Q/pvuu4yhqlrxK41R8q24a/7lhlQ0TFdFbWoc+oI9prm1UsH4n6ctF4/9y/hTo7cFzRhRB
RVR1eahLCQ22GZJ9BXBzhPwzFU7WQ1jHUOkrpTKViIqdSvHBEUUjMLhEj4N0XqVAc0rQs903YZ0X
xsiQSsrp4zoAk+kNi7+DBf/0SoNIBNmomz82eXG77SjbiaU4JxMKPT9tGimME823vY8LeSGaCH2d
WiGKdqYZU8Qza9QGjgUw/xLCdaEIL626lkURfLnwAT7vZJIt8R6bQUZ5ktS/0v7yt0SqbCcib5Jb
kvpCwzAZQbu1bBI2mvsoC4rP81RYa8i2m6cK7A9sE+ZhHy1/VmpkBt78/zD5LuayOKMpig2lfkfG
K189F0Dq8AzI0DJj8lAlSv1diga48PF3LgiloHTooTSqlYEjNeHPM8vaIUGGmRpMQistGAS0LWuq
VCHqHM4r4gjQgnjHKddM5v8XQFF6EUwM5bsCBEbyOGeQV9oGJQ9H2iZf+wNs4Yv7H50e3zkFVtFx
zcz6N8Un/gD41fC0evVnAbQVVXLjRLWJ2dDyOk65RFc0GVkdaN8aAMb/uHi/TfLp6tjgGWIgq2Xb
7A9qfy72w8xZpVOkR0caBlkoxAjk7ecFqIqQOVPixQ3Ljmk2h2Jey5UCFVREgWwedYihbUMDYssM
Jaey/VJ5OgN9pL488eLZk1Xnw6mEt6GNkgTmGbcvB8dvHPhMD9MCKRD3qa1oFTpdbsGNTf94qDMx
XpBlkjusVf4ILEFHghkcRdypsApJO6LsUD0sZlJ/FkmyUy1T0MBaWZWg4kbb8e599k9UlybGLTyD
ppUX6+p8hgMO9D8CfH/FahogAPZr04HkyZUlRLIh//khjcHJ2XNpgAa0PJ1xT0QvMo3Luqg7jZxg
+nakUsBHR6/AhI9CFFTiEGEde17JyHkohlJldHwgQEKO3CRPx7uxAcdtVb28ADcrTmX9ab+BF53e
V9Wh1UVhJll9yUdfdQR2Q2bZfAUBfNQyRkebtxj9R+t4WHJmgNZs+WdRIoEPd5sGHYP6L/HweMWj
nfWodGyintqnKd4sVl62Z4u0X2Hzbrzl+7hc1utAN2UEYe5opMeABhYwr5K/oWZBGED1ZcUd3+PN
NFfuwdlrjBtIdibrday7a5bFThO+dUSx5iYaRPDuVZoS49I1W0yvOYTpfdi5rWCcASS/IVBWI93w
/UyvMOfAnp4pjXxMqUB9u2Ekji8sMhL0AbmcQk/hwG9w+R3KQItnSa/CfrTtPgltDCoxossg1f+U
1ACZcHKpEz0d+aCK9DLkeaYH65drkP1SWN9CZV5hAWIrfNWKWw5QWpw/ral6nLHsgWPmfPgnxLZL
9sxfjR7KOApVNpyZcxfoqBNoAMqoVpGhGZKeak5F+2Vi9ioioPaohD17q/IPTtcl/+PtCNkP+7ea
BBAddIMwqI7vGiff9sQD1yp1DoKP/cLfhVlmEb1r3hsQqrw/0Im+bG7agvE4ORYdpC43QOuxK5DP
K/pL/02lx/uubEwm19wuSNUHEH2R4BzYzTb6zq7PiCQmQIDEDXFPHVzPgf2bS1fk+elhc85paICx
LYVmUNL5DmerX39ZZ2p4GhW+GaZREgkB16cLYmXh0NBSMdFzSNiYBR0H4wIL5HrK2EvLlIqkf72d
Cy29Cgt9GdMq+q7A4rJI/VpCnjppDSmdiSQEpNG6OXJPQliMQUtzdFoBVatETKxytCWPitorI/2E
Cs+9rKXLXAO4T9+sI1hLQDzKd3zKtc26fRF2IrxYdHN9imaSYKzet2EZSY+meMZ/Y8UpCy7AJ+vX
wZTm3bucUwqTXDVhuYiBhsOkL2zYQaeKmRJIwn8lc+UeM16sIxCzGcV7fytpHvEHSrOrVHdUCqxn
fmWvwJIo/9zLZkQOkGqVX4HGuJIOsqGxYdtgH82yjJCj2clSRh0tmGWqjZ9VrQAu50l2c7C6FdbF
tmNceyNSg96owK0IGug4WdUJF7JNb84322pBSyRVhcfD+WduBSCYBAVLKEBK0A+u0vtivPIeE06l
OgRkssf2OeLrzl9j3qRMDKNBcT+y72OE1AJsal6jMSeq7TgFZV4x3AR8con/xwvStix2l4NizKUZ
hKKB69RS4Hmt8a2p2cdOAb+O5z+gSt5GkU6+YTM31Ca1MZAYHfmI/ad629tbZlW85WqHzaZRSC5K
atZOYw8hV8m7H6QB6pjTFeoTrPsibh1HHPcwiihDB9zFW03Bmdq46W+/GBYOCzkTTsPb6LwywSGO
EYjo7Y9LKq1L9ZA/GssQNIBVTqPB16S4Mj21kCNdG5bVSy3h/Ukp/G+cUOTVuJ28uIfpwG8f1+kL
sPsbwYIrvUcorbZuRvmD2mYsp0NyBXLal4lq6ypDsBFvwVxEv017GVt2J5TlPN3xRdrZn23tNnah
aPCWNamLcwlcuKT4gF+YGGeJYHCB5vShnGpwxliw5ocdDPV1MA/PxMCCUex/S6A2mA2N/5/muaC8
GaCtzaZugBE7NbdmatoC+GWhGseSCddOfRA5/KxZ8quJGiLe0wHXEvuOHoE/CXq/uyx+v0pCSZbC
e4XShOLIsd6GtotxNh+q29Ou5O0yMJrmCM39K7BqZ4BuURCUw0PvDtO82MkF9o9WjpugPUfjAKzO
oH8bCBUEcR8DibYNE5PATttx+7MEFL36K1DOlAbgj/2ZOEVZ9R7+obcSC/IHcTbIMPBOUHwUG/ra
/AY8DzqzNAcF66BsxcSZNgKaUO9b3EyfGStIYRydGdOxLgDZfVRRzzHLD3xx7Zl1E4GPXZD3ITJT
wzznHbfTEUaFCJ1tpMkrgOarvWpCQUssORW3IVrj8dy1yL4ubFRVF9mCIVlYLvP6YxfKKc2kfv/x
xRmFFZcdGVg1Gf6HZy7dXRyeB5JjrOLNWnqmo6ZTauJl1HVpIukdPszAw4HP+Z3vjofHAD3uoJkL
goj9yYNMV59WElg0qjLFXIuCWfDlyI1BUDCO1VyhaFfRBMwAVBWOIY0y6TKF7eChUzjTOMPv7Xvb
dbyWOOZMScGdGSpRAzQdBKDhfK61QiswZvHesYpP8RJR0Fg4s8yWSH+Jk6EMp2OHLI3GqNd7peIB
J7BDMeaE1q+A2fQr9Kf74iiFsLEhxqlHf9XCW+ukurnokitkTyYzquEOExrguTCTS4aq1J4dqQsp
3T2F/aZsn1+qBnG4YajFuZznyEqPi1AoCW8nj6KWYvUL2jPtNg1QbKuqo445hknYr3St6tZtkNXu
44ZWX/OfnL9wb1cp3ScH42ASx9+AgEISGvs/ZdCUc83it3WsQV52Cn8csp89VVCwn1nu8bc0It3K
WqVlyKGjgT0QJcZkV3nUy8EJ68trN/SvrgtYtoR2fczJCCc+FPRQRQ/a/QT4TzLDmjH3gw+K6eX7
fImEL2RL/Kg61WHt6ikKil6tovVhxGKbH58dNandF8fNNbolD5ku8jBlWp4ztiU1s43xq1cswnRS
gSqYzSVes4jRoL3qq6UxUkXYsjd7QwU15Z4owDFMWywfYABvRVr0dxOQzciaAJQSn+EOTbqH4DbZ
VFcwDnyQN1EMeS9Bidu+Ddla9b7zPq+5iPHfSMNB3e2kqM+TmUH8PcgM5ujllqIxhxSVcMaPBY6o
GN3I6+drDL1vHpKNb18r+DLgzmUZifJ5PrqroESez5/BO0gaXao2VKRMYHiFqMxcFOEd1uuHIgkI
y6C7FsfQQ30VcVU6rMbhD6py3NApQW/R2+vE1VR4PYgGHiuF5M/H7yM5P7cQ+PB17vvKBCCQJuIE
9VFaQ+w8A+sF7odqIDSqhL1CZZ5MT3pY5R8Pxd1lF+Nw062n9I09nnQPrssI68VWKkOk0Y+LiIGT
1mt/Gb2Gs0beSIq1wFEJJtgOr48nbxVWo1krQGSrtgyCJdsdwYuGbWxnqOHx4npRMRdG/VO5qWAD
C8RSt8o8uvXz49TriuNlVGkGPSxFrvAS2PMPo9Ndx9ZkJsut/PvjvZcVKmqbxSbpLn9/ura18bNU
AAxih1APF2In3We+lUTj3Xxvt0x45tepMkjditkdrY2TsizM57tQ1MGrW+dgJBvySiCUsXla9G/j
KSZ7AWrR7vU0HUfu2VAhG6tlaem1J8tuPQ5/dM6pPiRldLuimS6PY0gLMZ3C+oeNnseA0AhMgU9V
zI5gvpTNVxveHJ3+hUmqcdHoJLXMET8zrfNIHo5oNcfh0A1JK1IzS3Xc+BmUrfVpouZjBdvWr8Uc
CtxjGlJ0ER45yCKC+A2Cl9K0xsB9wh7SuFMSq1MYVazhOJNRjPEOzcCvFvczeH24OodX16rtd+3U
eorvk84bg4F0MyR8d+l/UdoCjlOxBRpELE3YNND7jRY4ciNe+ALu2Zr86K1Qy427XMQGmn4A1Y7Q
XSGYt/U0Bp2fDllGPMY3Evucz9tRXdsP/RddTsYvtredZFMYTd+krShij+cytn59na2yRm4JNlMU
RtGhLLU2NE0aONdeHhlnoJZXPU6qBucD9UxBMf5HJQ6kBbPDf1UZj3ww1hIkGIyE9C4zS3oaPi+n
FVULD3znQKUZuodOL8QAWyoOC3GGnH0OYyEgjVkO8rR+IMGCEgael/pbKjEL0sUC4gzsT1HHB2C/
ObViydvWUR7LH0SMgCskK6Snuk1cQv62sC0GrOE6UcbKdkEddrCkoAHPOA1OIPnNm1Mc4t9qtVSC
pJ9ge6NIXKEc8vLSg5Bgao/P2U2XZZ11khapavAkGMuXZuGT1P+xQCqYS7hpirBAeo20MNnYbS59
KSwuNpX1pS0wPAVdfVlhi90nYFh+7HD6HMfGCIssloo+zPmmpMuCO7H8G/2V+Kb23r9jmGG2UFKT
OZg2zWV1Ql7qVJiZ/eKS6eeZ2gTXTHTbgOQjaF98q30ey78B6zP66wb0FUN0Q1uqezANa/hpyujJ
ilfOTkqTELmF3Ut+hI5Uvm8zLQ/pr+uq9SUHsjIytgQQrqrwPtEEBCbiJ7FwW8o/6PwxjTvCrx/i
DwMu5X8FL27QIGzL3lF0cck2NS3e24Dw3tDcsKe6kmiVWFJYJgVhBoBAR8zkNzNlRA2SP7j9GYKL
qy/kLZ9UQQG1oHbUgJIpNbDnNq9UuIplCA8d6H/9aoN7rUtgqdCJgyEA/FHtgMIBbX6heninwdFZ
72GKI5vAPI3JPOdA09qnfPIvu4zoN6ekalGmE7Nf853jaEf0FPJLZJtzhTaGLE598CiTptrpKK6k
EQHW0k45Iaj5GUzqR1xtvUFacGoVmgelW1ImY+VlL6hxgSnVoNaiNXZYTuFG1fbsTqYkhURLasIm
AlkBTmEOiVNo3/BJLAXAyvOP6QUKZ3yPOewA8f263S6qOKqD9XKpT7Ua3A98AYR+LK13j8ThEw6G
7l5hzbcaj2Iu4qbdhrHRhU73dDztbJ4C0tYmri+pVdSMb5VvHYuIxXL0gOl0cYNtAGcztdX1YOHC
wiviKtLLiYXWfBP/ECOaEwYksLIjOHhxC69Myxg9r75P2u4nnoeFnfm9SMUElJoHY2eDLka0DdAu
/R1ZhVpVmL3JIBUnamcfY6UIuoFWBk7clreUY3QPMsSv954QK47mA1Gtlm4il4kqE47UoEH/xgAI
mUj1Qnl/2YFgBaKJ4F8iu06zQzWJOTkw6gWoUqyyruZtwV4PGS7o1Ubs+fAQVAz8JXuNpqL/yJBj
AV7Rn1/C0jfROJx0w5CTLAMiwmyRZESMVmgqQOMmbpPdGkFtck411TIu2V4Xjc3z1ICSXdO4mwmR
k88rF94mRqV1xMK4c/kM9ClmJKmGnP9HIXUgg/tCBmPfMCT60Tbb0sTz4oRlZzi+jT1utDBmD8HW
umsFhVpPed0xOPcPgXzOxNvLR29RnL5EkXM4n9LcD8npia5czRTB6Sszu1J/2aIV2RC81mv4/yCz
z5BhX+O1oXaJJGFc2GIFwKFzCX7s3EwO0Y9LTZSuq4T1/7vl1f3oVPaQ2i8TH49g+TlRhBmpAYyp
cBeILuYAgXgQpr8XBEUHDTb8utdM2KcqJmimgDrnvbvIPEY+GCtS7ZF+MxXZ3CoY6WBdlypoBiN/
GniFt+gk12JBT3c8cxLwuI2fIxbD3JtdVgoApB+zfYyfi9iiBVdXmRVfG1uY+veHgGJY3jTE7rCd
g215bL6mOxmTgVWyxlRFlRCkYeaNMdOVNKzwD1YzDn8pHXHIsl/TFgS7LUJoLOkWzljuTxnQ2nqq
rpAghL0jq7ZsBJTsKbOvJju/OAYIgNvYn66+flq3jwQWEhuIzEypgoApLGPKtLCmz17lau93eQ+A
vvImkedY9VFmgq2cF5p324XhwskEL2DztU5vDiT8UKQeArxY1n38zvFQn2pcdnztbj7xBdXGFymP
ffrE2SKUumYy0ZZYvyZSWiDLo6KFcG2GfvJcPuJ1W1mN5PLncXo6AM8SLdePT6IgQEs/9IL4UnvC
+wPFEPsBihJj+FOk2FjkKVAdtVBTpdkVanT4cWp1UkT8io7m2g6eggNX9iCs5HuNWdiJECWkYH48
IJPiw4OdybfnvZ728Jqanf73eRmTz7BPQETQE1koYp9/BBiyIwuP+Q06/kPRAzrLZEt7Knzj3q8Y
5fNaUs3CMVWKnC+y98um7lT8fFV7qTmrMDpiAL1LNPSpxPWQ4zy46gYs3iuRja1HeTWNqcEqwiPE
JYNmf/ag375L+hCF/Gbi9XpG08lKR3WQDn+CvvF8bLH7PoEI9fwsF73kxH3MMoidRTyiPQS02wc9
ufw9TAffL76TEnLZh9UceAA6nGTCqoA9NARpTxoc/mXza2ZuobV44Egf+nxTa79pz5XyUQlMRlTb
Qkeawh7HX0jd6c5kwmkEagNCkwmM3EBDQFmRBj2di9E42AOmAikDVDdukKgX9450Ht0iPgJuyj7G
A03nuYMIWhEhPQVW+DNzyj/QmB+LKeVwcP/HTqgFNsMfM8f+pqcX4+RLagtfHcmVllTs7QiVnSjk
ZBmfW8KQwCxhcY5/WtSFcUKabdSESHz5tS7UQpCn4ryOx7f4cV9e1YfMd0JjHJ18KvhxXBBNL5GO
wESSuVDZYUWVr9XkCtDTthmhcMR90Ghdj24EkkYus/xUsshT5fM1kiGgfoSG3WmJrtPR7i1dRiVr
ryg/Dqhh0pU7YBjadIteShuX700aQY/V4Pr8MoLJnDT1H2+ceb5jZYceXCb33m1SnEAm9TfRUWXT
xNGBU6p8Bgq00WSPdFifbqmY2Xizaftwfi2RoH8ulF0dN+q2PcepqCaBmfOLZl5j9FfiFOM6YnJa
Oa4nsuxbgB2Vx4CipEpjb5ONV+lJSL8CXDFmi63B6v/30C9Rz4WDwz7OTnpCKzVoAIzBwzmjiw0W
xsGscssDKR4NKhOX86PtxHNzJUAWPmthaiLK1r+VXrgzss8OMG+PPBAFonc4U57xb5XnioWdNnJ0
NAvbMwn3+sTvqi6xf3fp6reX4wfxj+LD+07DWzSrbQQs30A/82WC04d+kcTKdH1tNiWvixqMoRUg
NDGIFCKv+l5jple8Jdt6Tf2DVctO2SVzWubXfQnUHOY8rtxDn2KeBzPbNaZzvoJ7TSBZfOmXREZF
YcT9/4E/ZZFtIcN3GNMW3p4Jjc7B2NBDKUFsXCo3KoZkZ0oMbjXB59iu7v74RxLX6ef5NIwuKu0v
CZdAhXAfrl4e8iniu5B2Uej8aJwoxXjSgbO3aIlrZUUGFtX9len9pNCDNR1rPY6LFDJz726/rhE9
JS/PkKyNqyVJl4nL0Hu0Xi1Z7PqgrWZxlSKFMu+cqn2Nyp5vAE5iw4J03kr2FQwcpVRB8E5rsjyK
0Nst9hcIaYOuy+Kb7dzvbOXTP7CZMDYrcE+8wIQqidyTrDrN8s9g0ux7LnE8X1GBTK1w7Oj3DKHW
18W2EBAl/AGQ18rL5u/7Bp87MIlg8+1h4pUwAbugbVfUtbAoftNOGS4Q+A2vtuNbKdlYLu4dcZZ8
fTLq7v6F8Pe4PpcyiqSzaRF+XCcp6XpqRnVDVTsfRa8GLcTj9Tuma5hG8wnrtJus0FFclFPIkU3J
2IEGPKMk82fZaICzEoKRqUz1JORR8mDgXTFt/4tFv6gyZE4xOwGwZrJnaftQqPBV5PNqju/E8yGJ
/fzbi3PL5dSf+GGjQzcAQNnoWnNx1Y51X3lBeU6eqI42DeduxweBbK9wguh9Cs7agFGqxGkvA3xM
e1shVmrLyoVYAwOm3UquQeObWgYAwoxYhChQNXzHXiVWH7sepowdxxV67InAcvF+YOi+zrhXNEHn
MqxPWTKVhi962PTLihFA5fDQtC1T5fiaau5e6uYmg9eE10fvsR/NgLsi1WV253U1YUtuveqT8G9w
havBEAgzCRz/YANLSnQ2lWdXLEGN6yoODt+kfXdRmlSI3rdsDhB+he3Vzv931GMuGo7f+iMU/L0P
AwNFVVuI+Z/qcyKul9UeWDHBn/5uGtbmRIr0xjo7u1jQkTn9b9J8I7adkBfYJr6Jr5SciuIvE6OV
aGCdemrGUkoyFd7+aGQMOtzCwwtMC6gYqKtIVM5mb3EyeUDij+q9T0+9gxkplh37CtuhXzZExW+j
BZRIF8GoOrmrg+VYbrTfEJTChJEVtvSx3jj6AnMB7ZW5IpYM2xyclnox29U1ScNN2i0LBWTrPWkI
X1h1X6YQWvA8EaGpUEr+0qk4hc7VpW/XEV/cDtYm+YPIv3ZUKf0IenQXAuy4LbjnbrfALesWiyit
jjm/a5LfKggNDx5dqVAvfIcaUPAvB72iuWRIDkHIw8iU8jntWYcvGkQp47bZvL5tMoK4lCPz/I32
FaBGBRB7suwZyVuKEDJIFMzopr4MfF86MQcvKKcZEjE9HNuyKOyjumQtvx5R8k4zzdvbwP+fqZlY
Wxen41DI53sKlG9DD17TXp9e8Ogf/fFNCRNzLOMB2n+OIBGdlpY6djhFzYP8k6xIgAZaS18//0Bk
b99Qwqodms07J79aY4t9wuAeEVOd+JYp1R3j7gCRzrG/87SEENxasJxJYE5v+ONknzvC/xwG1PCX
/n4Slt4sRg2emTlqePbUfmt5Rjm7LY2TgBkdXoCFFkR09g9g7LdeYu38yVRhZsTIyyo+TxHYGNDY
AMRIM42CS5mKa0lrn8piI21bbYo9sybz0r5A0QAKZ2mzlgbMXiUp7mUqKZqCmmKEDUpza8xr3zmv
yA9LShBsJca+mD30ByrqKPSEm6DAS5oAA+rHSxZfw+TrrviZx3i+odQDl4lGDBVQnwtWSICzduIB
Jvo3v1gGB2YduGYg6i0NA8YbSw6wH0kd01HAofK/p0cnZjPF1zFWjB+KGjlxeupxyezpXlrJDwHg
Rt1BzypcyDHJspZZCt0Gp8fmVpkihdCGrzgLOnu8h/dp2lyDVL4Lv2UCijZlpIecRVDC8RRYSqPu
H4DRPMj3zhKPhId35QCWtUI3xMo5sm6TikTQ0tEubCXGnhxh/v3FM+z+8XhlaCqT55hkpzoWVHNY
4w548IK9fLbGxbhI+lTjyCTvYUQZpSIxUtbycFxiVEtVJVLfflyHrKdh7sISrQB3XtZ5l4rFBl7u
04QFPaK1/wmubtuo9a9Eut3gOqLbywgch/UhAFXaiolusODSNntyMzCaWEeGSZLjF1Am3JhHn0NR
GbQ2vTrXUKbrTX4O8xi869ELkknMqCY/+1kvQvu+Vgu47VUPFa4ageX6bVNUxP7sUdSpSr6MXI5G
FBvMpeSvA0Jt/e2Voey6tX1zbUT9Kt4K1NkWy1Btf1HkInoaeiAB7uGzJNIPqeOIlym98MwfrjsD
Nf7hSdqrFXUaytiBCA0EzvmVrDmYsw/RkrYp+HCpIPeRe98AK+I19/9wunz/OSOiU+K0Mf1HWUD6
YzLM2V+JIiMFkBS1Ul7e2OpAvykCpDR/Ued8Xo9OV0Hj2h8uQlCFDvJV+gK/9UmmTKvuegj0/d+Q
pBAFfVbmwJys+36gy8Z2sOX4Uhl5yDx2O7pToQZ3LEEa0IRL1bKtiyZ1Yft7BPnk52hs6V6e5ubY
1E4VZB9MyzwePzEF69Hgq7bg/qtjT6TywEEwJf5B4Mztc9f/u8IqX2IPMtCb763YQ4lsvs0/JRPJ
/SHzRgRheI+Z7loYyPqbjbvtNNMcUTNfFlkJdot1hgpN9pRi9uUkxpn/eRIen6OCp85zzcXDFBZK
AE4ZrTAAFU6V8NYmVFCgOAB8/9AjEjVZ/kmgNLTr1cRsIcchNMqIBuhtZ2ClI/uhntKNoJQYMg/D
6izIiqKyquLpNhEAOHYDcW7gFkZ0ZHF7Ay3NnYO/0iMDrZNIqqAC4R3n0ChiBjbOWTDJiVMbmmNK
FRMx48ze9tj28MLXdoPGrtBLHx/NF63kGeeQSjb66WeWhiN4RUePCRJ5G5zXMUVtFRJAy3eL3jMI
Cs8llCrE8/4qphZtxiawsdxVWsPzNVr+fbApv0AtFZJevLjskf/bkpDaIlfwiDYwP7FNuFqXcTD3
2O2QrK3iL5XwEfFR+EG7IJixuKjj/zAYdf0UAjNc4clVNPaTkef1KL8BaWFaUeFCEMq9y3DjCIaB
tePAFIOu5OzwBQkSs7rUrW8buLTRG2n8/4h8vc+SQQMYwCWkEFN4e5QUYsnPpeGIvRl5sQ95TowH
JqPnSO07XYbu5vOLa1w2MVg0wbySTyzlNTCPeC5EqaXnYlAz+TSX4wOr4wEBGp8n4QfLIARWyYM1
YJpSZAdEWUdAEFIg7h214SGKkbgTwQi1oknWA46c2GxGRK8AfG4z2OXz3mt7WiyRPNToxv8wS3iA
RH3iuvt4rl36ZC8vwDT7BvH6UoLyW3GDRNm7/G4y8ijuMYZgQRk+wSgEh9CRsDxq0lC1GcHDta8q
oAm3cteZZp+6Mg1c82duF4YPRHKvy4n/m0uDD6mbBBITAqkQo92SBlHQcboJrv3s6RMEJQq4NDil
Qrali7SXzpNL+HbFyYCN/dDjyGW0+8yWe/9eQijy3EyjtHuMn93YlqpDlCWP769kFI9eYuUM/C+s
6Ci5Fr+wcIlpx1+FSu/rsFw8Yj3WDp/M8EQehQEdAU411nH4pFs5fIRR/TrRRRWC2LVzGIs4vEwl
YYX45SVSC0LlYxJf+VhKccZ5CJD0AIh3ndQc6U1drvfWWW11mipwuQWGGu54Hf9ResuAoLS8cy10
n8otqL6yEH+EPFqRfG+NLDH7fBH/SqRqC45463huNcnU43RLcHd1DWCnq4ZQWbeTH3h9/94K8JYQ
ljllGOyS2CB56ZTKYXf+6kIRO70e52yY1jQD7ECdVeAfbEFIzOfxfn8XD2ZuOxIoA/9sge6//Krs
HYA2uz02mbkVpZUbB+lkhhIkULYZSWtjnM2tnN1k32GZ/N48sUVMWjkAlD+8EbjxjaYvzWjSbmGm
k3SorKXwOkhwDiXcsDUi4/almxPbLd07vYqoidlx73lsxFr1Y8seWj7wvrRm3o32xXyWgIyNXuHY
Pve7Sx17Py7hzCLlgkOo621zI4LObxOqcy+GE56O4QH/U9PSvs7WuOItVtT4PMWgjk03wR20CyIq
1NkFhq49wIY2YfMunQIMFxolVC3LHybAUrsO5niwRmnQ+Tx4AdDJCaiV3YcApyG8iUGiSH0nkY21
N7MRgRmnh8l48Wh7IF0+UvgOk9g5tBa3F+T3YazeVei6sEyaa4NKwOnBnKPkgCewfYwiNfzanzMV
T2YX5l0575yWTqh6MdlojpIP8w841QfH4XhdMWUcBtYN8cPp/8+pN4+0fLW6Cvy01wm6ztpnt+CC
NzpQV0D8M/clcKs/ORUrv6v5O/6TcRUxipdqEF3QlXqb4da+cWuFu074dRndRMwEzygwLCYX43sK
CG3l2Lte7WuDeUK4WVPzP4pqxd5fGKWb5TgMb4IU5a2Oh4jMbLL/twdcPceKMLAT9hEBaUzJFmjx
BvJxw0QdRiU/BbsmZf41QyiAOdpSWykrWltjJKndRoiTWwzyWvOfOonxvVJlhz68nplkofgkwJqZ
L1GaLk18lNA9NiPwAT64sl54Q3hKGWjqgR0A7nHeK9XVU3F11Z9wtUjsKbBwr/60YNucT3I6Wvnk
D8Z4IcUxw3++v25sOknRuzR49J8ujaMeNfYH1MlIMe6ySnYUCz+3qyS1541Ea7S4kT4t1o3m3BYL
oDxK4B8HtCCA06vdaCfxOpcoERMZDeNZcWH+Fx6++Q4pItR9mBJZAOVx+/JWo/lGmr/UIf99nH/N
wG1V/kKjVhCW2nUiFUyI1In1/eEcXbHsUdWBhjihHMDilbxTscAw4IO8PJvvBLgCW3pvQbk9FtmB
IHnrcHdX/JoWaqaYBMflyxG4t/zxO5xXwio3t7sDDHxdcE9LTNUxSKEyt8HxOAjK/3aPtcpvqDTP
dWYJnoY5vTWyTf/yfmLaWSH4QY57hc5QJq6Vn0sNZtowdMO+BpxsDqvfrCflD+pj7fUhMKoYoBrn
B5oo4vXDJo9gohZ6AkmRkfWC1X4QUVwPgnl1GqAGyVH/wAngQjdcRto+GuNhl4soFAF0tmXyLUqR
EE7Grb3HcA3vOuggHP2lrZF5noNkL1p42jvFyyENehvydUFTajolp/m8oJ3Gn875hFNbvqgc2kIY
sIyWuN671utdZz9wG1JWv7sQMBR8hgkMMTfcq1hduk4zP3DdQ/4AR8KexSK31ThzLoSTCw8yqxdP
cg81Dcf/KeNR7odrpZgdp7p0ol721gt0StiIbQGgGPPM1hMcJF49dhByJ7a+f0pYEggO9uUauhw3
g+8O4VqZIPhQPsm52qESgac+j8adRtYTSRjtcWoip7tJ2oNnqsUyoA6mr5ESCJz+OHjcwSAfPYBh
Si9AEMAB45e5K64FnwND22+pvEfhDhK6TsBOzRtzC0AvaaWF+iElWwAnbGpXEbs/6u5ZG75uimpH
JGdYhv187MMG8yXRVv1DdY6HvfsNbvhLyT8EK+bUxqLs0CYVb2GeR5uILob4oFgidE4Wr4wBuCtB
OKxO9IO6Lei54y601xW+0gaKDGo0zJaLn+iitV1twHRi3wD8x2yCo/BlBik+cXKk9PJuZL5CEIMQ
QeXuZW9tIU3v89SascqmzmclJMNvdOAOcRWHcGu2XnlyVcg6khwvFQygVJF4B9t3qJj2zP1QlsRN
DzRF/Q11PXW1gaRlZSYiSz9q3B+GUOojFFN6rHskfJ9YS1hbZBe/5ZEJC6KmKABHKXc+yanQsFEG
4xpJUB0KXR71daRyrhnb4NVHeOnm3DPVtgjjydjZs/XDDTkHVJeJPTM9RatBQYXXf5Y/J9rf//VQ
XT2iisglewzWX02FsreL0IJFevl8Pz/IIRl2FuMVqrZ4X7uPFVdhVuP3A8jEVlufiKygLid8Xuyc
vMtNeGy8+sNNJs3Hl4Dy/6pdvpd3MfjW6rtokQA/EFc64SZeGzfIjHzFUZ40KvF9lLQGFEDlxifm
kjqovGkmTe3J4GFbj6qnZqxs6RqqqYy9EIZc/6fHssOnqqezmad2vDRYZAmPqCWUV1u4Gp+fNqw8
e2nTIqi+plyEMKsE9xfR4opXOpoMvoD5xgptHxUzL/auoMXBAJlWaPIDTJPMEz+rRF1eKT/ZeOr1
KCLVGLLs8n+Hflkagh91fgmvz6D1wvIFFo99XBqUIZzJatcwsU2JaxKH0U4iVSI4M23droB5a+Kv
SUdQMcEPPIUtnOGl9nj2Ry7hZjR8TEgF6XzemSsyI+3Tlaac5CNDES51Uz1Qosp5ZdGgVQQKks1t
KbAGACvtRyfE5BPZNl9dw8/DxQQuxqBCUtoD50uM1p9ZyWpsZoYE6bbvufBcJrfKOLu63KUFhuqv
2p5FrK1dNlzpzTc0YroLZupupgP0FH+38to7BH8d1YsgSWneYuGqxh1AhR6FlOoTVYtB3tPtfXOq
ATEyxim2ovzKyOCuhvYrTsD1lRUGkqxcA8V9z5jfRm5hVLT08RtHPuadTis4vW/hxKTk/zGhdAy4
8+rq8d7Za5qeKmgydEMP7NJv8vuM+SJKb+tzPPMEx527ZEd9C3kfj4V6FoQprr1S5VFnRNMAhkzi
Suojp7s09d8tUo9wzaG8WHZoLNt3bGhXQVqIWuXLEtzLQ3zyU2Fm2roKQUb8Siqb9979ju3TRAJJ
6VDNdWCKbXsk0EvlZosUQpZPb+rVnXViy1gKogqnAWPy7dPnFy9/wXyv+Nl2BeV5VcCxdwwBfG/V
Yd4pSeTqVapdNz7FooRP7NZZrcWvTEwLAVdXlGOPoLDll/MMtfBi9MpfPrxmFaqoX2zWWZX/Ubtn
ZGRCx1oaUb17Y3DIq/ZPH6b1BjDdyOu5ufWPaxSK+AZbDNg04QVFeZK7IvCeYVMtia/Z0+I5cJhi
QgVM33YsiiHY1bmn86yv8N45N1Vvd7rMkn+Y6kIs3rnAdW5BljQq8HwJCr3+FVCQ79x78mRft9XV
Y2Twgb6tvfBYt02mAvXAvMj2un0kd7sHCyztTfCqxRMw3AZyiRyoy5r+ke5QzvPyvOz9s6TKHD5U
MqHcISl5E3xbmB2gw1vN/TFPMb8bdVuQtrk4qqNBW505og1KBbhbRIUvVIftPPGmsLCrIhCcGB0s
uKTSZLa+BSPpktCaxnzmazBfbLx9+cpAc3NM/+2SHrOB7/9VSOaNYYpo2Vt52G42EUWEsNnIMGjt
p6sxhDRIW+DJ+vLmiEEQ1VDCqDNhVKeI9zR/LZ26o98seZN+TsCdPm85b9BqFTc4ltMw2UJU6/Ve
I/xRzhpEkH0yBAj/5A1Nxx7k0LTVy672Tbzjxkm50HYgusuV5u4uaZGoJ/jZf4X60SxaC27fMGUF
OfQFiNE+VCmvdqvHoIUdhpDt7LSrn02e/91heURFEkTqFbp0JvmhPlfOQ2tPTacz8f0Yg3aVdLgs
XeJnJ2LpBxOQOLLijDrpRgLuiC670I/lfoZuxn46UqOfldD1EdY01bC87gcBnAguNqhlOfKxSxLM
e21h40r4dadwThLxPRuQ/xkXM/c5hTEKF54Tj+Hnuk4g/r8V9ajedCOZMhxyvB7yrC8K73T6ILzC
g4BdkdAqfAfQEhjo2RtVYSvCQCtt4EwpYHOzCbyBih/eFyOWzgXCiS4KH4aqF85/h4Py0G4I5Yu6
5wJVwRldLui2e/7IUbwviD+E3K9ri9ErWcJ9se7BQXz0ozBcaEdBw6G9WOXsI5GwlXsU/FnPCFF7
FXjS0mfDqkwPwQ9Zycmef0NkCm1RVbBpnS04SBqFTF9XuimopTK/jXTcf+KMQQUqihPZRLAxNjog
3cRIy3v1EXYjyw4M4htxyFb/SKzEkJIIJx1b0t+uNdRTSSxCqnz6ooWVdAe6paWrc73NKWJvHZRo
OZ4iPkpDQTxUYOSFRaygtCKpahTv/k6t2gxMMJECzWcCZCGpr9XWmiecSMOTur+1snjZqdNMkATh
Taqa5XMAyZfeOTA6XltWskxEh2aOZGCTD/EC7nXX+7dtaNbhKu+cfI31kguG2o3S3Sh8g94Ew59C
9nRsYQFMkXnIMQDGsNv6uF270iHA1OwoK03z64stY2B5CaLDus0VbulWB9nXwnvlM9CD5NnKiUGX
x1C2sv4Pcz9E6y1uSt8qT+GU7yriayo4WeWvo3t+zAzGjefP5dLxX+o2uQqnzTjrQe4Hq4pDTkQa
Gn+wknf9lt0WBmsrCKkq28iWFkofqyKUKv3ENaTyfyXxPZfGxuEYzY4KfvcgepuFhuQ98NDfCf5b
EbGz3nYbDTUd65vgvHFt0JzT00VrTWRZ9jvQCHC18JNvEvxcDNSs/3G1Lo0aZbaWVl948ObVWIgZ
tN9e1BR6IMmBR7AaaeqFj6+ft6i0Km74esDg44M+nreLg9OECQ/xi0xhFk+Zj4seKwTIPAzI7HX8
BEJDiu02k+3548d/nJ4+GuJeKoZ+XB4LZR/D9TRP9Tvv4ymud+J1vDZEpHkCNEK/SH/Ne4Fi1nNV
R3V/3j9ThvFYnKB9ie/1FbaC+NZpasRWPAQiahsIKLpYYfr6VG7jB886uSpI/KSby9QDeWWE/OPW
UnKUOCtlyloEaOS3mCxmqQ/WJwcV0A6ARGHilumZqq5utLqEKCNMLDe7SXiHqeCFgpoXVJ+KY8uc
HSmFK3WpasMCU3oF3YkyKkzFZaHugHVhSuT0xYqcONn0Cm9YwvuJQgUE3BldAvAQYMZ6LWtcyK7Z
iN0NRJuLOFZV3BVroRbdqMFtzNHr4lh9eGTlg0mm31JD9YsJN84gvv6qaC8/m3GgJq/YPJqLxj9d
jF0d+qNAPFgRvaYyb3j88bRCu6fBnURXvsG/B6i9gHdlLAJhcq8h4FTQanl8+aNr9ABAa90nH0cb
E6B6dVPtfl52wHCEtG14yg/kRxy+r39CjycdE1nwKxdsfdkwje4iZqtIE/L2PuuwllNBNUN9yCJz
PQQ2s9QoqADL6ugaQ1G9mGd/WSw/fztv0VWoLpVFp631SqnJULl6qjAOOTg114IBrhgt3ABCNRWq
hIorVsOUKKpQjsQZ3jHZYIPNwUfE03inGQOu+MQ5VhaB3YoHveyXHbcahHcFqLY23Efpw6+ULcAE
hWjBrrcht4oDfBRE1+4jieNi3JKbR++CJWEMFBnSezfBZ+EIiiQClYMW1rH8P+kn8TmuLtULKWhu
0i1sH6uCU4ADJwClhJSrpeCXvry4ohEqQtfU2kzPlzWosy2NVPMez8EZWw6lCp7WhkZyYdY79dm3
01uI7qC3NSkq14h0al2Lvup74GdB6gW6F2lGnzpOpPMOWgAmGFyB0kSm11CJdbZRQlrW6UavdmM4
Gtzxu6EjS/fBDjgVueSBVpETm1I38gQPGDwAb/vWp3sUSAXs2xUupjPervcs+HIFKLnBe81cCI8v
h2WQ6+CQDY01bQPjxMclWalDQ4FZTg5z4q2mLh/3uvKcxnWtqI+ABYefA3ZmyLSGPqag8tFgCCPa
QJs8RmolElyQfDee40Kk9W94jSEMCjiizaxkMwSDki8MhqKYmvzmradBgcfLcOp4gYHmPGKswbLA
0cgcPG+53H/qwLZYKibCYHnTUdu0z/VuUaM1ws2QQmIccY6hatVUunnAbTPe7IEi125J/KzHPEKw
8+6k/cNkoTDIO4/AehuBpVWFHSdxfqKU/VVP/hTWqsCLjj6NnjS6V13gYP4hHWCZc2x5X8GYM/pZ
dtFruoTH0YnNEo3KfLdKBXIwidiKXWi8MIZIinq3p7WdHAoG5gJJ/wyvGei2n4iRsUCdHm/xhmiO
M2T4YIExXIKw97/J7l6p+tXsige6Wwivgrd7NC78QcNvRCtp+PTtSjBgcL9kKMWpG+6coHBo1JmB
PQ4oBPUfG5O+C8LImv5TW6ORnLQE0zLAc53CL/NQuVTK+mYk2XpD8VlpHPXHDZ4z31PmL7HmJ/IJ
fgcRR6vCyaw6/V+i0tjDy7wkcb2Pj7sZKwYJCB4CXYWyOOpwuySKlw1qOko9dRXEP67O5EVqlyZp
JsmJzcwk05oyCLY/xs7IMbSkQE5I6MwedG7pfQl7B3e6s+3/U7n76ZZYUbhYxDGQsPv2qBFConSY
4hT3FT3hI+m0hrR8u17Ga8Wr6+vLSb7axwx0dCdskck5QHaSI1rmeWRc7C8nn5R5lwC7arHkM3tv
ip0hKdrGF4BGJyvnbUbtY2LJIiWj0fVEGHyE/aM7wC7+rw8PYs9gbuFFigrrSZ4fYEY3daXWlNzL
pBXP6J4YxgSvT5806svhpmyvqdlSYIW/R+Vdc4s7imtf6aW13pQ0ukpHNo6KgZkvXjiaO6rjFinR
BygibL7qVXik/NNjrC4ObNTklrikPrBbWnd/z9dN9hiDSn/71RL1jqvhgf+hgGIhj0wwuGL9+WQb
wbBhA+caRpik/6Th3wIz0b1v5A4XbcThb3BMHePS/MBOH0T+QDGKTPijNqdln/+zpvdUXy2m4W7F
eqJ3OTW3M/6bswxtG1ZWotUPZfdOTbyvmMssRj7wRFtIEg6CA3+ofIe7ztrnfwfebrFr3dhS9b7W
xmJJb+my3iF3agTEpIaHZQd6sfcysTCMAnhB3gQ/0S8aTFwvedh1HCPiYVNLGbmvhyUuavMAYBl/
OZmFNL9lK3dHwMajkypj6WCq5i6QSvMQhrss9g288cTufGV/IR3esn0pEEQOMbMKPXJyauDigQgE
8hcpEEe9ythddHOxIu58gAxk+z6apTAGx8w4VsWJIHlMonC9w7UQPb/O3ZXit/ZEYvMXFy859uHr
M2052ZBuiejMSDJvTZsItnCcQ38Fh+II3/qEODVCi2vV4OD19NXuh588pKJsbm0wzUBvG2WUMskN
wSCakNzhwXKgveVunPALmW7PvF3DueJo3Zeh5g+fRep0e1ELdyCYYwu8AkWsr8Dv8J+bUpk+YXib
06IoF7q3ngkLGPB63Siq3pjgtPt1gcJ1coq7K4tt6B5qcTr3kV3sgOTQQrYCb5Kntl/iNddY+JVT
pY5gj6AN2ONdrf8wYbDxe6L24REf8xhf0dGQjznRnLjd3VaTwC49tf/YHV8wNAP51aJJnNb/4Wmp
2H7NME9QfNezTMdU8V0VOzic08fiTIaU2p8ZiYAnbV9eWGpAcFZwDFsMIqkr7Q1n+SV9Ju9mlGc+
TtiMEWlSWI2AFvFdtaiUQmVw4wQ78iO3WmysRLxlZhh7YynOpxvVfu7HN+Jc4jGUDYMdliMIGzu4
AO+XETTPvwAbLHNQhkMc1jdWstqTGq+M326VWSM1JU0uHXiHboBtp+eMUtM4G2TMjKu9nWqikb3D
UyWuzc9nmlcdAOZxlP0GHTrS5v7sVxmhrHzkirY4+22RM55EWJgvY6GBO/4NCe/bgNzqLKi6GSNl
4VAIQ0/JfBuuHpl/4WzF3/tizTgCqoxRMaYR+aieHv4xK8Gv1sYf4TDquurozS2Q/vXoxaSC1nxP
nXa96uikUA4H7RRgE0jkS9RshSTZYhV72JBGzNrGnJngCfTImEq0co6iXQR0sncdUHg6wT1BgxZn
xXftYDH1d8ofxVLEVRhRQubLp6WmQQbypSvEQ+VaPPu1dY5BahhRCXNlrtOmE/UEVjiYUZzjsfIB
LSQGTFJAUb94YIrIdGsobiAbLyD+N3/7ik8UJKYcqVoPpjIrKEXovSZkwBeo7pd2yHPXkMhws8dm
CmVpSUljZouh6O/IHC7y6MtPtbXh4H1TZVUHVucWbVX9f6Fq46boX2sqs/W2EyLPCXdx8Lqm4OD/
HIuKSrT74EAugNFIVxLA276YhiN19voIm1qfRJwtrJRO7KsMbMkA6htSyreXVCP4FMXe1hj46g+9
eZdA0JYzJSWMcrgz0XJJ5Q2JbVkz6GgpBmc9tpMSb5QU8jBwLgZUTlK2qF+GCbxAxhzKF560i95x
7VyYRtaGqhUBdOWIwMPueaHgkTob3Fx4LZP7UGdC5qvudKSUACeZROkTKNJmrcSDrNH12+pp2Zdl
DWcouYgMatuwonP+gsnakmF9yhMqYpo1FDjKgHYhYhmmeMOqtnh61l1lo1M9QOMN4LQwl4D687qm
WN1/VDAWpaXhzTbmfcoiLJDzsCZh9+RcvwNnLh7b7xhdfoam1ep7QWnlyBE/ORL5urxufvX3QZ6N
hOMjsdRHviFqqAtmAN92wTKPRSDrb04na9JLkbawv0xXfgp+wJ92nPyJzwzAH22A/mP2xYIddJU2
3Bd7R9ZmAwNRKxJVOuV6nySQ2FWDdQyRzo8CQW3dHy+tzkYREWe4eGKiVdfyis2zjHAyYCAKwUBf
EUpVaaLXqGR/PmioJB2A/+IPF5ZDHSCTvvvfQ7HxEZOXu8JjAGutftdY69K8Vcrny/KN6v6K1VB9
AYzmmc4sVAvTNspF0J5oy8JRVIVg3hwWoOtsnOqJQFELUu/yv9PrjWZokCEl7HSYMUEnJ4X7jHyU
ItgnZ8KXpm4eOdw2db/XU+gRPwZp7Pe4Q5a00eHHcBl4cTRKT5k0ZE5j2rfEHPtg5hbnVbfJE19w
xCZZQg9s0dVtF2sSNsOtpw20lqhZJJ1R4LEh3GXkvfFkovEUEnZopj4EG2Rl9nGqA9qbZi3Ixv1b
n/JogVdSLoW0klS0wx9lshPHuehkhl+JSjz/zW0jY9+iox6loUz6r6SERdoNpkSjBrmBtaeWgJWk
vVuOUfW3yVkCguCbW7U6RnfT5UqIFrbr8lnocRIrD6BTzS+swzd0HTUuHKoKM/izrLAhxoEl8dBF
pJZSsm4xCL1eeBY7wDvGsBVVZ5A4oezBPRWxBOpLRII5E/if4YT0qutI51FxFBvau0a/I0cYxB+B
HI5jKjjfqjLM42cxi9jNSTiyAVnIPqgmn5um9AQGR1dMe/4/7xYVhID8u+iCfP2zDBfIujOa87F4
QOC7Qdx3psm+6Q0BamKM49iQN5b5ricdJ0qIcvrn06WgsiCyFYspTTEjqOIQ6r40b8q5sADaZfSD
Z5soOfD+tlKwMUZbrhcAIRAkpGg9Z66XdTZzUppPzGSDgHdyI4GTgdS3qjmWBoUthrCmZoYTQrF8
byegc+5wkdtTjSfgb3kwnwiGEcPtjEzoeTArsKMlHs5zdeXgHHCSNifRUD1qzUzkYSWUPNpXXY3Y
w9fngbzPQuoQttOi3lAIr1FKLb7e63Clb5aUCn2efqX2GHkJM9YZN/lrT27GI1qH3fS/2HMuumyP
S4rjw1j371NpwFYSyQyZhGCj36EnI9LWYVNx19INhDjUy4wuFxwezNdIfJgi8vkrh5tib2b7PJmQ
33CJ4DyCYWPpl1VsR1v4dk85lqB8OrRP+wIcRkfgHEE+x+6NYmDsoyyYB3gjp/L5+3KmO0jBgrAp
Wd/psMFESRUQlTjvQhW1RPPcC03i8MWwmzQBPwhLhK4xHAGjuzJTXFRWb7kEwAkgLVAsB+gBQUf2
yOc7UqhgO1RwuuPU7fpYqdQ43WfpdDkXdTStky8PqOB5uLfEinAmKl1DWxj9ASN9IhuDn5uIafVK
WeC2fQSjySWWmJm/O/hkpmqGoMQjePwNa+/lbr3Qg/TD+/Wyc9ZLMNVzwTDOCieOA/9la6eMkGLi
Z2lzT3Y9z4BadQaWYiK/gd9hL+3n00N46MdzSySK/WS6z6tYNt6K37cQoR6+puIuAQMf04kPcacU
Uuc4kQ3XPYV8KAr8JJsMCdoTOD3aOPsw/xItDx/sVMpEgCxeWsm17VsZ8dYlk3POe5nLsYEWS4Il
NDwszDQUoI3EBTPEBKK6QMuONN7vMqxUz48o0QkV96DDPhXF9kEBRBaMvVvNLjosMl1k7rwZzGuL
jDjzx5zzdJVJgYzGG4dv5CGL0g/0gkJUnwnxv4dki+lV4MJ17urvVT0C1mjFcQq/ghe6PcxmeFZF
AXEceAu3JIBhaRKH9wbJf7zBKfTnitp9n3DCaOFMZcqNJb4Nv38rQZkU8rZR4qmb9mzQ8PfK179y
UBS/rUnLL7feboqgfHqpN5RHxqthvJrcVy3+cOcxixof/f59FKwWFF6Pnxly5l5D3Sn5nJE6zbGy
lxWzhVJtifxl2uBfs46sBoQ2uvYbydIsDhJ8EypsHRki3r8nJehEiAj8Qc5kOt+R7c1hhYFMyRLx
HMKy1H2KW40/zFhOEDyw8xozpjKCTGrkupfi2pOVv+nh3kJlBBgdZY2d58o6TMRLrYaiHqsfU8rm
9MepvAaz5tvIfqWpF2l2Pms9b3AMTzIXuGTWi5jtVfVILuT2jnf7vt4EjjEwJ+e/eTDwDBOznota
WAbTWhzcS54U3HVJ7SHHLr6qse6w7Rs7Fx1u2rOBuBYq1//Tc3AkZcKsG25P8+24iHc+vympmRcU
uD+WkB1Eb6AV2aIRMpLqTbbSuJdIx/YXHIJhHppEDlF6pEdbLa2hIJETlcqfwj5/asbS5bngs5FT
LRBuEO6H8iU3PXvNP5W+w334x/eaiC/EG8HYjX+4vtiTXhSCeQB/oTHfXm8po3g3Al/wZBnq5Iaw
vtkeerrc3zLjDpas77j7/aUdL9wYAcn7B1TVE535f8R56uBuxk1Cy10a0ZqbfIq3eVAXYzbffHYV
g0xiYdJjNfACZbIISSgbgwUQq11gCRS+73MEs92zH8NncwqwRdfUUqquehWh6YG8ats+97ZmJkev
RucOl26wpZC2tF8nXF9CCgUEPpk4c4wRAANslMG5nAPybLxXhDqu10+EbPbWtyeqPZKVeP/2FaEr
60Act6MmzaMYmKcDWQ+4i+7e9Xwqa1zJf1fCicrDYRqMqMLXzwtHI9ZitUHUMMq0pahmI1pK4R6b
iKbAekuQPTUXt52rEdwiSNwVCcE8f/9zFCwlL2GYLuBXEvgubegx6ZsibVM+eSunPxPCGUv+NRvX
9PSbW6eZ0IDZ1hpb1orDElx8ujkamCCq1RCturo0vdz0JM1QMW5G3fZFKUWbLTopfym3cujtNYbm
/u3HTw8aGowUDc2zTwaW8lp1+f9bBA7awrSLsihwxCd9TcPWPIOMxrkSC92bJVC12+P2kFYGi7oS
UA2ubyVcmsaBI+75C07PF3pRYO+VDIGP9RHnJPhkaxTnHRWimz8J9z69iJ06SXZ/2NyamhHxNPe8
eGsXlMPK+TVGI4//ANukU5oamiotCJ7E4WWym6cPjrc0JdKnsExI7NAsr7lUk+zh+2ROnDFjn2TB
Q1tbuy5Nbs+6nME15CiXTOCVLndLZqpdZLnbei/4aEk6HfL92SYv1DNvfRnyNjqBu4JTgtgY3Qzn
CamNC7QQO3mVPsrDDJQEVS6Ks07X7KjZ2CqawhWdtLCm7CB2uqiRLkj+WPOHlimOwMgDh9UMjrGe
QN8GzlD5HfPl5XC5aZuoo1ZaYBw0HAuD0P4Q0fJaeUhRF77wbJIt59kBD9cu0/ZfFpEz63oyM0ev
Mw/bMjOFG0EtVKw35HVJifNtwQna4V9RL1aPrFEYBsNAHhjpOMwSjzIuPFIeeqYpFrRChaqykIAN
udINUq3IduysxevSELJzH/jkbk6z9qFozBiqrd5wMZtKUTS3U59KzzKnNZAogDvtbYx/WtWbLUnD
AcnoyctfbsEL+GRD+PTkdhYnXm83++EiVNthotyg0iXBJzm+hWQ3n+2V2cqk/xKX4nMCRkYyB/nL
04fWnomNgW/Lp9hBP2VCX8ZVfd2eYqEdRt+oJGxEHzO+jEBfGjidH+9gVnQCjG1R7yJnXGHMup0I
6ToTfBqsUvMJ92iVMC4IzG8gU/D50ABQGY5L/9P2ie+fkvcVJj8+XFBBSH25hQRSzXS4kAfdy5AO
zOaAZBUhvIY3cnij1oDEi8tmROqXdOqfv1cChK8RzWB7K71dBAjVnFlUUdhokaTvJlVwz0yicP0S
XFH2uveNs8gUm8Q7mNeYMb1mUw27u3/bZcq3OQRfS8rblODNNyJx4D1fHuKzKS6za6Qe2/B0CjSN
9rsoUXG9qt5wkvChkPqze+oSbiIEbItkNhDNg5otoVaz5A5GakWf7xn8TZNxroFY8TgEBN33o1qr
P+ENW0VWiNSyruyfZsgl16aMqiOksGtJ1M7j5j3oqJmB0V423ruMtx7WPAlKz3AyeRUtDPqfVG30
YlCf/vBRDyISA6feTPIUqDKFEUklh11yYy3buXMCm/yq9CP4L+r7+5psLoYM7A4I9+0YVQ3YbCCa
iHgmUkhKGBvVUYdR5pLjxjUVgn6B0XdkKtQDkpu5HRwOd97ZylIqHmoAjBmpdHo28CEA0E/HBlYL
XTTmoZSDemQTmJIsIKBnhZtdbUsE2wMAAjvxroDYqbBPINTt4XjW+Oaj1jZziuFXZ9JY7tlWKpJe
wrJFyKHi6vRJgVV2uR0YRcM3araeP1ZPH1ciZRIWTUHaC3E42o9bTDu9KoKfluL+UOb/jKTgj4cS
X9RrhZ/s5mHrNT2NZbZyJojxwwsSGnOD3GoA/DZaqMQFXJCpawEPfGnPVVXcuzpiGT5QQ83J5hYL
VnH1AZebqUXw7VLpPnB8z3OwY++KNhVSI6QApz3+bh+nC4qYCG3PkCknpDl7RTMSK9psyGkLlCgX
kUIBlKzHeNK5+PBVLbyLN4NHQFOInH92yE774Mkd+qmZSANizQJhokaJZB9+dngBxTJkFRODAfMG
96IPuDiPtvkgZv+TedtW4mqLnSWOfZcCNDXbYzbgMP0GcWzi4zRBi9BNSRfwRWWwRUB75Y/0B3eT
0Rp6nj5cGb1TlQcOi6GFg9ms/Gy/Tsc8Srnb3NuW/rCYPXE/q/GAm7ZbpeT9MKHh/uv1K+rtiEYT
zWSczmUJ9WTT0PP0/rhW1j4hxNArwU8HjHxN6wFygjefWcgGsMSQgYNk2ozlMjqR+oOGG/kWRpcW
0BGrjD1XBFOd+9Ti8dtDhe32ng/9jQSg048nZXNi0JURAduPOvwcq2cAAl7SvbxJG08I8+k+urLg
5t/gY5CDb/yCFpdJo4oyQSoI4vZc+yF9pNzDkBp5+Hy9VIQYqWu+SYEgXgb7Qi4APLSRkiw2fmv1
LSVM51DEXantaYoRu17WOaAjdpBW5BnUvCIyMkpywA3y33nf2L4jSKLMV9eIgU5rPgWntzrA4c4w
5z1/gQ/+hGBgquEOlRgre+hk6iWzYxq+/8HdbLxro2DDoxpg5fAyGoRWeBMTVKD1i5zgqVP74ubG
Bwv3k4PxYplx8ukxX7MS81q+InVEnmos8JHgbPngDQrtbgbEEW5XbSTjzW1/R0k85G7xcJDcqWlQ
FH+mFQFJFvM2FP40u7vpzIqZOXrUepTvaN1FWfWXMeLT4WrYQ5UBYN1MSoeCL4Qt2p7WWZhe75Sj
bLVbr27C6Wnasq2jP7KShGrgyZFaIKUZrwfoY5mDtPVY+xaHpBlimupPX3iCwp5xp2QyBe2MMi/u
BcZTSoQ/SsFApEDCchYnCZFPYYBT0m4Y7P1/SSyEYKl7pEMmD000+ay8SPitBmo0GI9vTpjCUkyG
LB6yKeGxJ4eNt/fSFoCrkvfpcZcJMZtz5uVp9j5or54PnReA3blFUpOfSQhRpCbrZVlax1Rm/Z8k
P5udWp/pj+gMKbFR68xF3dZ2KmgOMJ85BkjVYpVO5VrOoK/C09sRqS9rYVwn5ZL44o3j+C89m15o
nLCUsMh9P/jHaXrgWUY8z/J9aT20WyhJEdsaJkTCx1P8HmBMH1ataL5ZD1n9rftcoKSm+E59vk95
jL0Z8Gd4tG2N75XbKeIFjoiC8ed1fMD7eoWCoHqz1XAaE6xu8ahHrUjVbts1nJJvvKQMRAyYXJUi
r4IIJPxb01F3s4CcZVmCB0CBNVrWn7aq8dX9eLOaiYz7iPHbkvrOW29vR2TnNi/zMOtYp18mCVHP
qK/mnUQCy2JY+Sq44/9vEoukuMWfGug44UF5wGcM2bCREAxFqQjZsPDxnVfEtfJPB9WNYAL02EzO
078DySn5EKm/oB5BKzn3l+gma4pU8tzlPh2FYV1VPMXvtHlFzPsdTQpYAV7uPHkDop9wTgo99KSL
EtMUHxBMxEU8O/kx1eVag6saLJGz9v19wQ3sXPcYbBgjeaAySCpZYmKLNqQ5rB13bKPLPsS99yrn
jRyzdr7tT4piGHf7EafAuH/pyn5J2m23DGM6w+2tQmi2gtGMZ9GgcgJeGKTvs7ARcutUh1xzw+B6
5Fbd6ezOPAASpFSdUsf/5fFcnlGSbZREZpHTPWTuieMZDfhV+8Wn2pRwaNfqYF/hlip1ntJgUT5D
MtzNSbDF2nNJdtuaqn3rDd5XZTY6FvXVx5zUxyFsoirk7kSQ66Ig19sZooMpEL9MLdJTJ9VEOcqP
5tAdwzydeRpT5mIHu6zXoJqEldPh7GB7DcWH+Tl+g7nLUtNlhDxVrfeEz68WoXb9bQ9fa5dP8FKH
ALxzNnry/Gvh5ouNvmgacQmepylUX5E85h76hC6O/rhpz2zRLKKhvM7D9cDoz4+xYn/sZbmsnmRB
JCFGDW2YDh9UCb4yNrEsWDT3noXQRTFXvbCI2GCpiQrGqhgcTYGcSpk3HOUUP9JJJyfoGN3RBP2A
/JwnD0GmNWswnUQZNCzFBQAPWZ4hZA+Gg5fcWB3eZaP5rIviXSlXaAqdH2LAjuHKfhuE2eDw3SSB
5vVYg8ITUDFoIJFHmnotAGY50OHmzDErHNdF64iDBBy5kvPDLTo69hUFHqoYnULa3qAo/bozX490
5Sj9koZCk1Sjsm6YweIwFe5NAJkoMoa1dlW6DgG1hc7R6lGMoVU7XYXw9l2ftcHrj6TutyK4E66H
5WZZNGSEMrNT1RZWef0PNRazUV34d1byUfQjw9x/lTHbUL7HeC3lfxG7i/u7ZPu208CaZc/5+kqc
4LFKJxkXyM5TsXInk8yXKvhdc9UU6WC45rrOyq0v2RKz4EG2MfhCgI8y6V1B85g/d/PqWMS19qa1
PMuGf/R3VUoL1qCuWIIJa3vrTQRw5svsn61R5RaemfHYpZvDx8L5qOQ1x2cymWPMwYSHydFlZNKU
JhxvY2+/t+GzvX1L6VT747Pvi9yY65BTwJoH5VPaq8YiTZ3P6Gn+2QjBt+vCbpL4aOKML0E62Zho
QOHKd7RdEGhmgAAbMSDLMvGoQ4L5qH+jthNAozJ1t7NcTBceHM5YGGqTJOTSXfHYJr2LKP+W0/aK
7OtEmCyC+AffAhMqV6qbLidERoC0762BzmzVOgB+ZjmoJ5OLj8MYOWSMP50yaR81OzpmitoLiGHj
lEwazr81Ke2ZGE/2mywjKGl6VbAHW1Evw6jPNsi74U44aidy5io94KvKDumusMQCXPxVr+HZteDF
16lLsNhyVF5uKnLBhEO7mN8tMzzH80akv+HuvBDGhkuooX7pQkvlChOijmxTT5h6MO4e+LhFUPbI
vLEleLm8wy/ilugWF4aZR3onCs4h1p07NmUH9vrcWvLnxEkwFCqGid2lwDeI6CnFXVZ4bG6soZGx
8s0wBj7rARQVr1azT1OylSvq3qKAsC/Xa8PAKH+Tfusz1mAuqffsIqdcf9BBJXGaqKaTD4ZWb9Sw
P7AqtHulNVnAkh81ruHRpUdX4N0V2npCiGtr6wXDJA8ZN03yRQrIVEuXzcbjaFjM5lkRfykD3AoR
vo4T/9QxRsVdlHXSnRkOZ03fgkufJ0TSLEr/8XYhVdZo/dzyahx9pdwDpZDwC13iGeehqeAwlL1v
RpHYp7dKL2ynz02jdvgWzVNwG3pUpvNJU97at6jabrUrVEzo06yM0Z7a4d40pZxIjnqfUWVLkzIS
7uSbAQlosIcwPxH/qKjAJfntiW19eRBKtldsoseUyALJiImc9EAcUZWSuwVS9OL9o1Y041Dv8TAq
a/JuMGFsMD9AbBh5A5RU3yKU+wflkxk818KnuxLqhCchUKJCKVC6zSuMh7z14OQMbJ1i4IgZKhz+
9ShWoHNmX8FNr5qTT8y1yk3lLosDimjervbk3wJGJvdVzYXgs+OGqOCQwNlHOqDbPjYvBg+3SjYa
Xo9095xiOaNRO1WEZz/KeBibzGRHB2lTo7l7pTfok6vdx5vPfXh9qMRd6Xcs7DVAI+BLn5kLy4zN
4HbaOiutBMkXVTF+3/+5lFGK2b7cH2WjdC+XPdYa/u3Xno10MY3oYxAo4xlEoh7YYjRwwh6XnDvl
v/QkkdA3aRjADPZ7auVnKTtbzGgkm3VD79W3xILT5LiRA0NfzbFTUEaDb7s9ZXk5aGMGJKjPMM87
3cL/M9U+zqA7g6QpiWicsoF0Wojnt7hJjO/q31JZB6dBrh8I3x8BBh84SiyWTLG0vqtR6F78k25i
WZ9/JLrdLjhRaSt0SnF/XVcVZ5qS2eKUz0zsySYum5XspT8FkV9o2s8lRC14ReYXLGtNjfV1FiqI
CA1WtAjsJVDnONYqjYhvbY7u8GxPG6E0Xhxi2SHEVX5ybaAicDVAfeGcc9erVFTm56RjGS94zSDp
3zgHGo9oaWlGQZeSdMZG6DICKg7i8m33tUvv8GAe7qbuxBS8KjoyAp2SEcyckpmDMTJJd6uNyUsv
mb9oVotLAsVKdcab6E1McG/43MEVyX6arDB3ezpritJAmk8IcEaqE1tFdQ6N/UnmlKTRIhjX3wJW
FiqAWY7ZM+F2dKJFaw3YpbJpE61gXiu5Oei/Q9vLqwz57FxSfernL3FydTcxQAJ4zuF1YBts6tjY
1cVHMdne7wQivB2LViorSGUdk0F1jWLqHkiUtiAERqZJLXQERdBKmc90VCwP9MJ3C1F5sQBFMgjg
pvetJpCqK3nHn0Db6s/u4Ae8PPwnTL0qO/tKr4s+EuLCXwLoAfizok2oeWgN5xjpxZNFo8QQbvyQ
NZRsEwilnHzSDRSouP4sax2zYLZPU8P5kWUWTG8v1jmyDvP2DHQAoWy7plXo8uyyLyLzXDvHQdJD
m/3+Mw0aZ/fd8fw2GL+FpgjJzpGVEYA/ME6GRp+/yff2p0dvPqntQssorO3aAOfmnyyz3pwBrHwq
gkFpYcKLKoTiNxhHrBOP+dM9vishPG66JoBYheXoeRAPBbitQud/9xEQK9DoAKNFkwAQz0z2Y4jb
kX3N837YlDkHsq0SKO6XrbK/sIElNBE3NzURlZazxcUizgjSpwc3Lu04ReKQEWueRA/shZiSlbTr
TMkQTNJtP19VkxB/TAzo6vVkrYAOlBnhgBurtq0JJxi0sEkSV02y4K2qTuTa3ogy9biI+jeuAaFF
Iyo9y+J8UB03gfpw10PASRKGIOqTqKPQJqo1l+8UegKEPNyRMImsnCbLvubB0UziHzN7SQi325DK
ouNp+mrgI/lL5/z/HImQ9+Noo2h5nbAFbpE75yvhRuPYngDTEfD44to8ZuuPL85PDdzt9p9I39Gc
5nJCYS2B519QG0kPJDw0lRffctp76XTvZUxZ9WOwmCNRb2xVny4Pt7Y8OlGfFhU37OLhEjy8Ixjz
hp/uXZJjsqxRbIbrJ5ilSiV6UMwstsuXPkKW9eV8ghDqMGLdMmyMsONJKGkTd2wMl5zNI3pljS83
bILs9vm1EvayO83t3+KzDJSEwl94SArPFn++J4G/AVaasLhGPvEEgImSXqRLJPuRzIislinpHu32
Fug4PdCozkNV+lUwtnx2BEWZ4I8CSh/CaqD/UKccVqXylQWDzWn6fbKp1S0PxO63xs7BmCpnxqX/
S2bb2FLpK3Vv8VDU+642b1XYNSUYFQ2gSa7vrSx7OnBNgDsTo6iRKXDYdO9hIYalMyZ6EpdizJsz
RWh3QCkw6z5SXnuHZ2vIKUj2v1m7SP/BW2CmQQQnW+tCocjcJtWwoFf7PFWIGLea0W0bD4QdjU2a
VTBhI+mWPuNcnnBESzmm8oTI4GmksydOwwuANVqQCRyAsrGh2Q+1dVuytEixxr6ETSR4cZAAA4Iv
8vAh0pCicH2f6rfYSp2wjyfkd/qQL/M67femH24mQ+NgvSohnShb/EngTKav0HJMgkE6aIoXwPKK
c4gSqHGibEf8djfObwYqWe2N0qqBbrIYb6Q6k8WzPdwhG7svaJXXnAk7NR/SbifBcxiXBgNqNExg
X1/FhCTE+8K9CQEgg3h8OVduQRzAr4kRE5ls0VRUG4G/h+HwjJSjbmsOunn9jbNnO0MKdNjdNCMi
GVBJgT6upcZj0bA27XkjJGNVJsfARbtTjJu3qpVqGvpApGcQefyJmJquSIriTXzmXmBncvLjBz0F
qadGKfdKzRuPUFL3xEUmZhsZOxev6B24g2gkHSaoMX3S/6jcJvWIBBPGrXPpuSCKVSLYWuo6zAGc
make+WuL2v2DB/y955ta2ROay+Wb4ybS8QZ1FA97eWsHsD3dfND4ScQhsKvl4siNCLPh1YVQRJ5M
kZo3CsW7ATRSbg7mdAILKdLKPnNP7KE5TqEojPu5fyzUOV71fvq9+8jxVeEahxBnTnEtkuNwneqc
vHkwAutuZf63l6s05XXQ6SRwPAqK489InJrLga87qT6Qx30Cg62FdGV7EPkkY5UFy3LiFpL+HCbQ
ZXTCx+2fxNBkr4Gp+Ta10LApMtMRq0GlcYRfhgXKh73QY2SJ3V+UIZowzEbXsF+guDwl9X3RF9CT
SFkGuApoMtJM0dgza1430tN6HEfNxuUrt4dCToe7rx3pUK0N6HTLNLRtZx/zLYhrj3Qw9CmeT3sw
jv0oVdLaihnEzITKPGcd5KT+HbsYRwHIDDbVMCOZD1GoDnm79la9h+wa7/BsUlOMjD38Jn0au/dQ
gmYiiF1xbIEFP0UIx51SgkWWKCIC6FcDZGBbC0iIM2N3rX5gg3pQXBPQjk6udPI+5ZdY9SfWROBn
ZNlRHv4Wr/jJhLIgXARF9FkCjw+rBLyENbLhFL5Y/0s28dnCGRi48ZwcrJNV4GY+sdtzxrvOOmoQ
gZ8Agdvyy8IxZri11p+DtTyssbpJOSDuVaa0lvEWcgowwKpWfWvjrj2cgXvBq2H1sqx3rgiKKda/
quN95Jan4rMVy/+mxvci2kiz0pZV+36oyIlDqw7pKrsUxkvHeySVxIfsZ0Ml6PR/PEkUZX7wO7FH
ThQL5A2wouNNZ68Al2bwCMcd0of1WAZV5tGp9sIbO2tKwqnlDt0F9k6p0G6IZhCeVTIvqbflB+8O
14QpPAtC4UVfBgssuY99+sAVBxiknMIO3p/o2Nj9adKBeDmJ64RQktefOwLBN5bHy1lZArc28H8o
bU6ENL9GWD8a1oiLxRZvshgjWy7Noc3Gs80SgBWKJuk88KTzHvLKu0La6t9+YxBl+THl5AphopfC
/3k8sGbLRwQZOhItNwHP9zVsgSXX0R+EEqgkwisd6JE60ZRFRFs/ikEetTJomoub55WNI38YJTNQ
EovC/52cTYPdBEFOrcr4K36yF1Bwvs35MS44BY5xXWQviDbFP6c4KmjCDQX92qLpS4zynxCa8yMO
SuiylZVKRGZi7h8s9vkmrLZeKF+qMvl8Kq3FrsZ/qE4YMl3YS7M64gpvoFHxzgjiRAWUoSt0fkIR
4eHnP7oSF/uNxcsBTX/4L5q5oJXyf/+4dQxHYAdtP+3fQgWbdTYDUwdrBgUWcuuVFv2Y8wbdjKCO
v2u19o0Y1dmat4+l9mLTfPJ5OQpgNNBPQtM1TRVwlJhEI25p3GRb5Q+T1X1WUK88MO3QNZSvpnYj
lX121bUebV1kh7x8yWsOQhE5iuGZ321NhbhaAUfX68QjamMy6yV+mvHRubdNxtTnocqDJGwE18s2
KqoeqORkdsiO5wMWGTACqv9AzCh+V0/Stck2ctJhFx5+xHouZq8PgE5pBvptgs/iyk5GtN1E/8FA
VzRzkak9bWngaf/pnbPQ6R73/R0a8PHx/cYHEbVpRaAsd+FKfX3DD6kwx+mbIqiP4aNEHd+Q1tqi
gY49Z5mzjNng59wSbHYLvc0UFLUtVM5p8BqKpy+W53fVsNimKCdOrAueDd8VB8epvUXL6hROaFK1
iSzyQ7pX/sC/K0JVpQGeFtZpQpL5arRk/geI85JZTUMmYDd+1McGJq15rBgrr/PnDb2wqv7hv4Fo
vNefObj1KH6jWUHDsHUl53t9lh9oJpOpIH5gHddSKXzEnt2hhfxuiQ1EYcNX1UXma3wjKbIJWRAS
5mvaFD67znabHJleIeoQRUYLTIiEFEXgw7VlDg2uZpf+gHKFTVyV09/PUU2tb9XOFO6TsDtp8Vfn
H/nX63kpNaefzWypdEcThcCuVaUS4yzJ3rov8dmq1nwLyB8mepcCMocfirStmjSGfENnqaMpwV5J
Edmsp+0VDp7hvryv4rPAOGxiHcxIAMd0yKAN4FEthuY90JLO0193et8vSsARSbjQvR84ePZD1Fhs
t1ZhQkD0OmuFScROYed//J0kNq8+ow+uKgFh+RD6dJLjJ80X6xiD3MiztClM0RD7y1RCOop+NNqL
cxMl6RR9miElpdAMeVwjSBitwhPgbn8NThQnLmJT8iwa/MRG7poqvby7/RXI9zUWsJuz3Fj/rhjB
cvAicZ6KH8HxHg8yxE33ISzPMeLpcY1PCXsZJr8tEGiUd7NS36Mc26BJLlKiG3JGVzQVPJMv3aip
Q2R8YT6IuXKIat5Lcl8rvCoyP8HrgZYH4FEzwUMIgVz5z7WgcDpfVz3szH/MdwqwK62+sw2g9pJX
r9P/hUzPPgpPRLEX8FLU5/dvDq4hH9dNgEG2YXMrDryKc2oD2r1s+VkTUl4xnyYAKTUnroDax0ZH
q6VZf369QyXHYKMUUvdw4LN+rwMmwVCoxx/0sMOm/FU0MxLu99hVSrzIqHeJwSO8E3jEiAfdkAMR
b1AgPnxKIrTNME19g8tdmVrZr0FUKXdY+34LtNxDVEA3FcNX6lOtpB4oadMiQs7qrlqHnlOZ8kKC
tnvVkLSffJf0hXlfSUjOQ32UOt+nyysQYqMadyhhoEyCV+iqtsF93LOMh1pXH5Z2e/pr2LS6B+Qn
KGFiHMNPmf40pl5kkTuBCpWorAlYCwBF4UIvYuvcVBNC3PuzJm6v1RShXaVtA0bY0XCU8ZGMRpUm
pk1Fxj2PsczORGq9pQS4UwMnFovwXFj65OwZUvhsIgY0MT35X9GhwpAza5h5A0Q4SY/IK1mvKRTL
iCOTYoy603Symnzdb0PHMEykYH/7AIN8fj3fS+zjedwm5FzN6G87YGviOBkWywWmyqI2rqpqK/A7
iC+sZY90oR3yGj5UUKgEikb6DS5HwOYaPkeV9DyZdvSbX7O53w2hSqnCU6v1W/7WAkBhyLKn+fBn
fAmxKknOh+R5Yy7uLJic5eydANjJKOB6PG4yznQCoUJ4eWaroLIVZNCwVtunZvxOrGvaxKwGVwGe
73b7z/XR3RGBNCOXcZUhkg67xJTyRiM5bHdlJe9XuWXYegaon4wsZ11GSIb50tItOG1onxpbwBIn
YCnTYQYKnRmeZqVSFEIvpplsbThBWNjLUTOOvY7jAZr1FuIhRLVttR78Fie4myDck9AEx8LfRArQ
OsVBtMsfsMCcqJ2oN0R4DzaPIBkBVqnXPD2YrpH5X9FzuunxUttyebRTLJJXDZ1fcO+8yYmh0eh+
b82jz/D1CYdQ3gOJKm5cpvAazHYDv8tP3+JcndOoKxymJwCEtz/b5h6xzRF2Ace6xmP7gBc8Gu/P
A9eWmVBg+3Km+xH7UZdgWDDWpxpRQio31ZUDmtT4faumCx0Q+PidRkwAqY/0q56/Ze7sb3fVqtas
NHNNuBcNH8e4JIoFjG1TMKAEM/56eCl5+z2Xu2REh5tMsHiCOO8ks5YyvjWPsQwB4GtCSCAq8aR7
Ul0VRBwBsU8YWKCi08PrToxVOWdUxEcxHmDpWHuIHelfEc3IetD8rXjx+H2bwBBDGeY6xtfUVAZp
eRlqktFjo+BOmPQohxj4CLHZsNS77F/QBPGcbFqT/Nv8FJrA77/ZwAnwtt7Obib5T7VesPKLpmmd
ziwDyZcrlgxyMjaTPYDrldQRgorH0MZkgE9EHgH0XHntdt/QMPz0byDpvU6+zEXumyHJw676+Bpg
TZh2x4VV1yDFxXewQNa491hFvMTllkH3twFQAuJZJysYzcogl00JM8mb4a1j/KpErT6vbomOzRun
33SBhRwdTRMgBg11Yx+P8v1+kPorM2YBS8/9q8mWTVZMa5YEUh7TZA3sbLxPVlFX7sqw5rAl3gl3
AdVDAW7+JhkcrQ8F5jOgYStCZHy4BIScsJHSswpU4yJ7HZf/H5FETEMPUq4J714S5EdJv+TaDYrp
zaUN50BFAhKYJQOUsB+8FZGjLwyIuy5zBa2LQW1dz+8MB+eMVeEAVqQajanKgGTsoRLQAUPgT6cq
xpWhNQ/PVenWihyqWT/AzFEQ+atBu2O4lT06dmiA/4VChXA9JkdmMoWH6PzcOOw6HyrU6jQt7w6c
iY1rbIaWdylgOo2s483QEss0pt2bazxA4Jb12AZb6+z12LLpTOVJ6tHg/AHFFY9E9aFP30vj3jA8
x/0olhSzlyf6Cb5n3zMxXF/GUXG8IKcdm4Il0E9f7fWlKh/sKBEQp0Wq5tjqubYWehmNUJzqax67
AlRampoC0IPZgqTd2qXXI2KW7Z8xasnPdRiKR9oXc2q6S/px7c4uasNcxqlWiTgUtwL/0k67+CGC
HiTCHRx5sYJsPwsayHlZCBCA/vYxbPOAg96i0IOK4NgF/QEFp/FutK8dXLqQ1BIPoJAbh/0oc4ZQ
+vCQJpkdYo1mq1jb737I0tUFBCtb2/ooYAVx2x+bsHAmZ0e97RqjLuoiUMb/FvLpmUE3TTqNflJ3
kNOkN1f1PwZRlc42SokxqZHLitS3+wJy4X6lvwXdVvevyLI9CY3R0tyPxkNyYRIPK6O7aec5E8sA
CU/2zVtenpZn8D+oNe4HON54a4nJdnw1roBmivZHs4bNOxD+ITdRbiV6aroLPd62rJFpOVP3MBCc
mhstnoqs5UQfvnOHedPwL0UDWPbJopG7BduiDirrjUlbFS/P1H51hu0AMXjc4ba1BQbx0giihnaD
/ltS626XK0ZN1FPbh7Yu4n+Rg7P4I+lacj3p7jtrk3cLKQS3zVykS7msuE+7uFnmiQUsVX1AB4KW
F0GDpylM2z+ZocOch5w1mTatl2K4MsEgNL4l11OaYC7/kdrB42HAiOQaR1jbsSOvh9O9RhDGN9wA
q//gOlLLeCiQewOHpfH+EEp+F8FGplpconV2D2KJ0Ur3IjxGwxiAxH8VEs0t1PmPM5Sbwutk2zDw
CsENCRnGLengWYq0FkjBqwRSo4ecTaFPtJ/FNhFSiABQ7nu7n9TFkD6REYSUsKrVdUMtOyoxOsvr
jUmH0Tgumql8uJxouOIqdjbbPtu1tzUqFPPh9gGsfQsfPVKm9ssaFywsOLCbToDrZpXCNpN8Ko2j
Ureyb1KPXAkW/yH92cQ+qx6VO+ZJfk0mSztGBS0mMFVqtrt/CUv3tDICDv77wT4GY+36uyj2rmC+
FjQWLc/YerkQkcTEVeTH8tZ7i9dj10wbrD2YjTDf+iXtzvIw4jRhsIgPC38Yodkrm/cmophmDxOs
5KqxTd+fTgQu4zOSevfMgBhDdKFsGMA6X+NAMGJ3Jd8AeFBrWzy441XXLcQuC4R5/Xx6koNF3ZXE
/ZfDehwzWiwZp9162VjYysrrxVXip1pyY6Qz+HgRgMa1k/4/alHivIrundlMJZwlboevickOOA9T
CCYoCQb+HrIAffUDgoW+jJnSxXDZh+kqNpDyjonnNgmmLqe6XlbZ8DM+8EYNtyhv/Vp1aQNScLwW
H3/pxRfUXOia8+rjLyzd2aqOEX/tSCCi32zhvINv6NXjPFNoZwSMsoE/GxJGeH7zOinFytZ6e6Oh
V9xp0c1jXUU53GLn4NosbJ84yoJojSqubkNW2eO/NUT4os5rXtThdj6YrS74vL6IJSTPXLTioDM2
ULyDH3fwH3WAiDcH+ZQcE6m84sJpKqyy5FVr2H4+smvAEP8mpvjwGrY43NjhODAKb+/xyQu6CMsh
nLnxMw4XPEbjl9V0ghH+3SqWolJd5o6Ik8lcuwZIThBXgzAuamkl2+uPp4yPeD7lLnmCwY0j4rsa
cgbULyVULhsJuENbjpA7KZkRZoXa28pNzrJr8T0ew4Z7c6ZEvEEMmCaIRUDsV7+OkvSVF9k9VYz6
Xt/P/Yl8aA85/UIhjjJPw4pT3vcWPMvlxM33ZWmypXFguLsKxFvRFZotn5eP3J7uDstsevRWOLDW
Y6PonY+fBjYPgb8XMg6DHPzwZKnMd861l6SAVHNC0Zip0Nw4J8iWOPYBvKkBTE7fVj/OVX9U319U
YGX0zbhTjSaJrsJpP/B2gDbncjEQctWwJplBTHJY46k63alzKAKUZotP8aVmfcJmPkq+g40lSITM
sOrld/oibL4jV/uwuagZ7CF1Wp1ZCh9IZ0KqG7R0WkIGv5SW6FdKLRvvbUEIDGE0LtljwbiP1C2O
E14Qkl+zu0oc8lT9VzQVdMscyDaE1bCFSAhb3tTbuZgI2q6q/KfiIirDCVH5sYZYaa9euGAy/EbR
VeYgtWq76/zkZL+fX8x2Z5TsNfSuN4mFoFjlmLiDHkzZEu6SIRV/qSgFCmfxHo+aSrR/diS4Vz8u
sltLsxDVN62UbGzX7EX2JR+zcuHpHlQ8hYMiG3mVwP1GXLVtrjARU4lu3JMg8+PzYSxc8qHykaTU
0cqNCekKUHxLo380CbIUeHrpxk37fiYKQVR4DoXK1emNJzSPsnCKwvnxhclH5EsvspefhqFW+9ea
eQPjqvaNBwwEw2+AJUP5MgcmbOGrksYp6wzWLrIB6xF/JSKWr9j0MdMVAdmcM8DebO+fQDnm1HEH
eN42tCiqZUyWGABwZbP51cOi6/ea0HnJM76m62MW8gsmsAaMK6/9+SL2TL7/kDXDHLqONYeqEVlE
xCaZ8295EHngfyNM/C4E16+N+cqf8s1uidi1lJ6NtgXAAOJqSvjcBK2L2/GfE1gzXyjO4Jpw7ocJ
pUtsEcE1LA3RPekye5xpIUy9JY7zTJdSRAZQpeUCze4Ko3m1N6QK9J9SZL5UzatyfaOwoGpHf7hJ
SyF2ysA3lCS1YqWIhdmrR1EUTPpr6+kQsDWQTpIBJ8990JLrRuDpG/MgcLZ2BXBtHTXgzzAeHH3r
f5TOwiZKS1V+NRi3i32VX/pdIiC7BqEOBswM73IawucjfBqSe3V8brnw+U8cM7+0LoCq4PYcMnta
zXXpcuHphxIk5yIa4E7edADWUUVS8Y0lCc/XovAF3xiU8UhLGw2CvkqnPHSr3pGM2RILHY6AOwS3
d7/39agVY5cbSWg3N0+loAnfOJx/qybnT3wBwxisFX7sif4VK1XpX4l15ewyttRItKjnieJhWYlt
IHFzeE9EIu+/iSuOquwtrxkucv0Erkf16/9KjGTlr7+cro4FuYYzwBNkHPSdz4qhwN0zQC5CXdw9
hSG3rgPK7UT1aCmUxbFUgKK2FStoJuuASEAfWXF1Jy903gGvGCMrywjtPHO8uYM00Z1jw6oYLHtt
+I92mIuIp89PzvPVmjI2WKTAdZb/pwdPYfnhOg/WjZSCqUdHqtODbaR8IByz8xZXDv123gzT1g+K
w8uxvgw0V0/rCFTbtT17cDTI7q5O84DoyNlLYEovMi2urbWzPOVGz7ELhY6YORawv7BdYwBlkpxu
Gg6AnTrRdq4ywPJPv3MRBht9ZIMXfuPAsLa+RoRKkO3watP9aIUoSE3REuuvIs8YgdzdkoV5tfcH
HEyAFdQR9QBeUfQaXc5rH50fbQgI3rVxTp+NMfBqvNoLpSSN1bpaqQsMmQSYQh6XDV4AOPjwrQGK
1CtRcfmN4dlm/vb+3ZtA2RcHHkTO9FcCzR6Fs2OhuHpStOlEQCt0G0c/lKWavR2vsA2fHV5J40+l
t3ZH8EIH1/XliUuNFa/YRX/oiAbdnblUirmt+pgxAJRlYeGY5lVfzDxvxEaeDe7NdBw6sCpwWq93
lwp+G+Mkyxk4rM8XP+1l8unpUmkQ4TITiIv0FIq6ywAJ5+0P0tTQHAR5Tso6jA6+J7xJHvjch3Z+
7aPzrFroHKq8VQ1+mzgq5MEJjnUPc0STSoHw8HjVb8TYbNTx6clGsk0lp9SdGFpZA/QbARO1FuqO
U3yp488JLQak1TXkB76ly7U4LjnxaKW9hR/nQuGCm2EyrBaatsokqULoeJ5NSzY30WVqW/c+nOWG
dq4iM+rOznhuH0x2VmWbEut2HhOKnYPXYTZ/iMZFLGDJffzhsp85wn89m1XJUtoxyyqYanuLIAGs
4TN/H9DYiMkzphonYH24GjnEdSVvZOEbTTnv0cuvbFu32I5/EFgbbVpy22K1uuswnA0MbjMm53Ey
+/8xGKHZhmpWVrh4U9hAEuAxIrXA9xAcQp0pCagE2F26uA6TXg6xQIs+NtUff8LnW3lumuN0VrMj
EgBssDfAiZTIYglCEVLIlems1OynDNCg73CFvBynow/PeZLu8RH7GA8FuwBhpnPsqbcGMup0M6Vw
/MbTC3EQeNBOgAumCtEEeiyWzb1DmD3S4YLhAAdZjOSi0iqLXFqadkecyL1phJiaqgSpGcBoRCqK
tQ9spAb9YFD/Ftlnqtl06JWeEidurgNWJvpH5+E9NRGkCc8aqwd2Ny/O2mHEo8yBvxNV5EZJVelA
LWm+aTJC/Oc5ewF1151YmBgyyYozgLxDFvPqTmXT5CfUbtSAxh6i5RBXvfx5gufETDyZOfLFYdEI
qI2G/dm0NoEOfU3LBDKXYyOLjHdw6CC9+6bC+aWvgLZ0AbnJYk1qs2wRBnElr+JR45XWdW+aFQCb
ICq2BylAQW2MjmLZEmHMA5i1Go3Jjc9YI3thsvBCXJaLxh4IoxEPb10C6TXwkiqxgkxPQA+cLcVq
3fVp5ooyepXmqADbn64VFzwgC+W1NeVM4GyZQnwlveSHU8fUXSgv2wgPeufMHGYLWfZHk8BKioPW
kMyA/Wf3WfzrN0EnrOYZimGHMIhwGSVsiz2MDS3cXwJ6c6LfE2xqUgNqJ+U4VJPdm/OdKnm+juO8
USvT+PpvSWVX3Se2Z5kepWawnIw8li/rB/XOpfdq+tXpKr44SH6nufWsZOXR5K2Etxp1dJDbR4hG
IwAkR4c0oCsdlQ/hGN91ihh38nXc6Q37ijOz/2CSF0jTjfDOtjwPFKY22HguruYspaTJq/BaV5mk
vul5r9BtQuHOwc+WtI8u9wCxnR5lyPG5XauYc9oHQbcylEdZ1VmHB3V3ekhYUGQHFjMbl0p60ddv
L2hJhAPXR18R+bRJ8MF+S/HSftTd2g3J5c3f7hEnkUmhjtopUnL+C09HG6jdpUnbYiWIhzyCk4gy
v5ebvgZ2K4xYm3NJf+s9I9a68WFkASdIb+rD4dAwzlpze5TPbN34+rRDsZdXfegE4iyrK7rDNHUm
SHUXBuEjVJz+cgFalCmqAs68NS69KoPMS9sDWeWMK9KfmJQODDHkyUkWJsFLohd+7q5q0qbnD1vv
t1J1OQvOyi5xy/FJq4ezbhzveoqJC+1tFLQRDWI8O6Mfggpewcym63/6awLok8AlRDM89WvG/OtR
NYToxsbQmTWure+xPonXo+i78xRredoC2mEazW8u2KP7W/ZrOMeRZROvVVnwIw33oz15UpoNR3l5
xo//a5wJtCaA964zG9PKhOHWK12WwpXryTueM67c3BYLUiWCXCc7IdOXBxanmeIP5wLuLLhxeV2X
yZ4CvmSAA7hjpd0DovXpi0Iha8mDNKZwzduIu4bgEpfarJmU9LBEd3rizNcgPF6i76jfL5cpWVjA
hMTnCWhQd3Tzsl/Ja1ChNIo3JYiyJgROIcmGMpOUFcIHMD/BQ4bitKwN+jW9Y99ohQ5H2Aan3pEv
pYNkWmfxTUozClTcm08xR1K/drNVM3nk4A2Y4WuVq3zd21a4OV1mCB5PpkmuouayhMjLnR2XXTLY
QRcrfyeECvRph8+4D+ZXYgA3EKCLaYWP6ckc+zAvPK0hs7HgLva8JXqzdBMCHZ92dRjLY9LhWnBF
BI5v+qJwHfLHDvTal5qFJT8pC0Fv8wPUngOjK5P3dR9X28kZBoK10E+hCzW4OWev63LV5w40mOxi
2NJwtMsymgAUFxJHbH4zzOaguAq775mziLsMBz/7zNA5+86zUkfCIDnhMTHhm8OV2EQcr8G96JxR
JJyobeWD0eq/vb/NpryXv7W1qp/rw4P038iBeeD2GxQgmj851ugrysPBLf95Kh7t+Z63XVcTqUTX
efP0x7otSjJRnNt+19U4iQSgdaDvECz88DqYDmR5mmHz0c+ZUMnPsIQ/1ckwISdEUOhi/kcLkX7o
nH4BSpT3zOIO/lo1orHRT8XwyD5RcTf1t7fWhV/c9MsJm0rpROtQLfMHxAdlnugMmYX4HD8QL0or
YzEGeMGjdQ0IPLt1h3F8YIryMJXTcw56XYhvWHvkO/8cAXbbhCpM4Rky0wMWlqQtQtWmpTb4EV1u
sjqbiq8LNkLrEzkd7O8mu2x1X9NRhXXBDaaadZUEyVPmnGh9/Fm5y6vXs0q9ezOuahBzCx/xl9So
L8ZvMvJtSb4JfR5g5rU/BW2Pwcsenab1xZJtiOFb5BIkkxqVCpKdpTn9AiuA+Ei6bWZw2s0XuQuJ
jIUuxDhb8wgjLaFIuAMslEgX9f3akFQTlcrftAm59QV1QTPsXYxbEySJREt/Yjyx84bhRWyUkrrt
M86as1J61Dex2xqB9hzS2BnNStL5L8ja33JXRe231OutGsuRK2YYnq2KK8eOTM+gzHamDUA87+oM
rErGJh02tJH2clOwwQaTGQxjOJ1Ao0PE5oXRqQxEQ77i5jkjxekdUf/hH5FId/pZ3RwgXc1Hhv6y
8yQSF2EoHm3PNemUWqfAFw8rjp+s32tKur3dy240hDuJ8egYgiuXzstsRQnLTMhBsEZvO5NDdol7
//tAX8KbQeSOEdFQod3Qt5hj6T2oc1aWs8DD+c7rFAc2GbylJzZcgkd1w4ZFkiX+21VUz3EL83WA
DDKWGIq8DwTgZDcZyVrrNy3gHQ58WcSICXgt0Sn6uw299+Rma2TB/KPqLU/zYTZXOFypaemjy286
m3pW6XfoLTH4VLyve7y/gZSOwoOO6mKvfuiMB4rH4IghCFjz0dARTNvYHNAOwFSv9G90k5f5fUc0
AzSCdsGdSxr2oFNwPZXMgZGhcCVApxQJpXHJifrSW0sWHHqofbeM95//jk049TWdGLT2JPAcmOvl
7RznraGF3tWaXst5oasie2VwrCPEMpM3IjSqaIrMsROFTana8i4isW7jC0AmiNZ5A9qQTW+Fh+K5
ic3E0ETFLNbL/VaQQZIhgdILRn9adqsMgb88BGNQeLANPpDFvN50qQbioNstEfbcFdQLqcEckxFB
0R7L17NBB6LAOQQCOPLOHFFi9rMFClaOzEMaa/a0V4pOJVJo/2qJEEIW42to6woNYovng/PzyGVT
52C7/ILC+rUwySU4QElWhHie2cc+1tMYxfJt6MWDxitblo1SLTZSAru/grPoCRrqjBKbH0EzaGbe
rYKN5O3VH6Dc0r2pElzJnss/Yp0ceWKjsyzSgggjIRuIfj3zS82+ozQadQaLMJBe1vCszg1/Okmj
dUR3Fy6oboQB0Gu2tVG/7/DNa3Y6Dx+SSsAnO/1cAKCiUJqeMlt1CtD4pX1I8Fz4Kow2RkL1DV8S
Sxkoj7SeV7bleT/TL/9RBLp2fx95PpBUPVLFs17zymrJeLdKD31XZPB2nMTPGAH+fdfQoNuGaVPj
z+vOf7EPm6KbTELmHKGOhUi5tOETHPPMiS1q/oD3P6uxbrHCN9BNw3/bRfXKoQCOzQoK1SA1UfXr
neQnea+QuPf6yLexMx2STvvafmGMQPu4TqEMK8eK7MMOavS06i1zsrDTRdCKo7qddMPKuT5hbQVN
RvP7cY774zybVZRAqOAir5+Sbj/hUVDCXosS4yv06b1lxF9tULWU//H7gb4YdY3uI1QlF2fV/hLt
J5OQMrOmLD83OM+SZ/RVc/gcjvsrOdg3fbNVqtW16a33sU5L3y89sKt4mbURIIna9yq8TihQkuVj
ckLnCadMxvmxgnQwErHJt8ZExKMaUVCi3sZyk0scHAB9VhynSLFtGNc4ckX3nGm9r+VDT7r26xcL
3vu9hO5+DBUcur6s2MkrdrBDu4lTkf8vnu2X9eTlFnf0ZIks1Sczhi1g/xyffjp6hXx8T5b2MYk0
vsHAQPbhSlkxX+hKP3h87UcXyMngArWLGOQ5d2MaMzISKBt91iF2e4Wwzo94qg6UQ4xJVriSbs8e
lWg+0T5B8Pe84XGwE+VqO86S+0IO1KtHZAB5C+hgvg1jpzAk0h6WaI0saYX6lV2uMxX34UhiBBAN
+PbXAM5eqS/dEDgpbgBqTHd01psX4ggmgcROneo5TxjXI5l0mOtXQi7f8jFn1ukzE8sjZ4pCWwKO
dh/0nGldIyHOveCurcdo2kbOlrgLZZ7eSSYCL4IIds+GPiue5q/g7QaMo/nTo9nBZx3sketwaEaR
z2pdsHLyUtg05U6vyrJqbuJlRjKhnvVLcNBjtCujFqYJD/G8OmlhNwiJYf3wHHITLqCapTU5kQju
nbf02DOTtN8nL+jx7Y9KorEYr9U2v3aEbqoI92MpzMmVK8aUrvufdYLEpGu5eb+T3l5twI6RXzjQ
VCVw5vt3GXotwSC7IdAX+Ui5mXypS3iwVWa8HWkazvpUhRkbFBd8PGA34qsreu876f0Xkq7ftToY
2Rna7psAEgKtBGZQI4x9MNULXTbx7tOsU52rjgmp7sMAWnSnF52IXXRgWcAoIG32aov4aikxeqN+
7l/6tgvpctdeQ+jmNVyTFwCbvohWqY9GFL2gBSUuZ2rmNEDHCfoqs+GHZ0kioqPDu5xRlEbr8KMZ
QHY8mo1739b1GyphIBR1dZ0Mwz4lDlVfuQ/bOHQi9GMNqVlpP5tjwP0Td80aFPk/WNWIRjSc9SDO
3wZIKWOUdF8vWBDh2cCaDx9ywMAONtDbBEVbOi1ZLecv0zoSAjQXGpZ8XqUjrDstmxlJ+z1VIfyC
3fExPij5VQTeUKQx7c9icFEI/gkFjn2e/SldTbyRJgWihW9bw1Ilr3HL9xkdkUXKhoiMg7MNW0DD
2Tl1Ox6E7OcOLLZ0Wk1zafdl7n/MJbIFXtAz4B+4/VE1ZXNAbq09mo68gzw10figmq4vdMSWuraO
RQ+ADlR0MxccmFMzNUtWkmDUCbrEjlPCYn+D8gcOj9HdpqBys4t747NHVSM5kVamcTYah3+72xPT
V/nM3LXcaBoe8YEcnmLO1uuzHEaw1/UzLZkLofMnKS1xbPmDgUR/rJNyKrgimgQAKCx0ZZMedIA3
Do0lTFlHN//oTp/scZUtEqccTLCPyxzKcINUFp3S7FZSuAnTveg7A3lAUGGD/t/dcYg6YqjMuhAU
IJfWDQyjbkrdCUtmZxFbVeqpTcrB31UnEkGnTqUARF6Wu6a7EdoLst3Cp5Nz07ke8hB/ELol1blg
k/eIC3iAlIYUEswzuZMX1pmT/w9iFs7IS1fekYurx4KiDZEPoeC1xlYfjDQTQ+uF4AcjxSwb1kv3
hHtxnNWu5YiLZx/PZ5HsdE5Yx31z+yYgmBckRWLVafrTCbWmEcbl2VFvP2SyRd4+sVzliHM6ZGXU
33yDY7RE7H5XYgaWslrkxt7hgWtVaQ4g+R9phCCGaxy2hbbDavIxIrVMQd5UW44+tYPkZ9yhWtUW
u+a9xpfr7lHlqf3HYx4e/i3dUDITx6IYjYplIgkOG8kd1gkwxk7LQgehHOvdDPYJSO6UfIBKcvz9
aGP4U2c1hPjOaqHn8ZtftlWgPYH3onLsLq8HJShPl+A+FKaC0oHisFUTsqB8F3BSPb7azYUolTAN
r3tPHe/JbuBfLHrXl5IbDr361tj1Smtn6EELUWGic1YZW7Ic6reVkaAyz7S2lw/i2FIQvUCE/kg5
1rUEpVgYcAnFPGm2y4tixwgyYgz5hkjQqsqiPcnUXmvyPj7aI4XSwuhPvXcTfgd974V+nBtcTneD
YDqcutq3Tlz2CqTRTKbhUQWChAp90t5MXdtAdeYXBmC4yavP772tgS9fS8h2Yuf2INqYqteINgkX
noDmzLnyRxndIl3T5tUxosRrtt/RlY1okWfDdLnafBI72SaquDPslUJEWvgAxiPEooIsVuDtDOoX
sRVLkj231adMmhp4hGnMU/kMzt7B+iCIdmowdam/Y7CKTzBI7aI63xEiqZd4Oujt/rQ1YVHVjSzj
WnclNo+vr26CiOIGlKfftiEt1bi1CT84efJ/QU4hvVD+qsneEwQPdvuHW0yePlcjJPRJ7lq4Ns0s
5IWs9y62975ezbwxmzRGrCKiY8y8mu0eCrz+AEc0nFexvMRGWJA+p0qcNoRqSbRQTk1YcsiNIDDF
r2LurQHie7fsHQZdqdCw8mDNZ4fouHIL5EjPJI5gjD1jhjofNtTETOuLcRYU8Lwe2E92Y1sm/K2Z
kev7DIOK/xYLzGSIiyxkrCx83RGARCrCnPF/GhFzeYw5Kroae60MnNwqgpqer0Kd3PYbrgh1kxTU
QZn6F+TejqbzRuJRCOTzUtBCTKJ2Nvstk3PPWFLl5p6EiVwOXY6hj5KlHicED7Z1UOavllvh2NlV
CmjpxlQAKDmwijRKXqR1nue2TnPCKUmaGf4V0foVqWP0Fg1H2tCZiKgM3/gp4J1xBPQ6eJK9uYSV
dL9zhAJg5c/vhjmxa8fhgz86hiBPnZgUAQefSGjc0omkMzFGJr2KDKiv3bGGbo0XRXWQ1O7bKPdB
f/HSwqdrhtCBQxs4sUfV/F5NblEv/98i+w0kfjprha+5A5ZATyjlnKX+W9QcRbt6BVvhaIk5oLzl
nf4jNyRPoDL3ArT9rnsPiyJkQoQEtyTZr3Byu+HhmKdhVyEyM2CTjkzCShiJcL7XvEYGFgwRNDnh
rGgYoVMyMSVwDvLOphLs+Q05CRGOVqxjTq49f6Qp75bRGdYYziNexJdOFI8qKujrfb5bVY1//giK
CytQanhemiqBweXUgAwjq7typq83JWaxs1bLemH9k8gPy1/6WdMlzI2XABzWdG3Rsc6t4fTF8j5n
FqtsYMlMIxs6ie3+zf61BSaGsQiNQ8WQ9QzE/s5S1UKl86xLK+miciN63jQykotoIGAkkpgKTuin
UL3Z2XuTXpC/McV43F7vU/ZxyXNkEWGwDKBs/efFU2hTY59qNTHYSSwxYIT6upWCrQxkaHEqXPpP
7anWv9njlg+p7oXNipnK5FtdX2fGys384LDZ6xRLeGa4v0Z17p2lcSXd1+sDEuy797eFk2p17UCY
nB/F1+i8XYddFulGhh1r5QkREevtDKE50atiCYTQ3vIahiaKw6tZhyx38VXzoiVdjMQcv245RcZA
kGhXh0MOTER1TR4LyoQF7yCV7rI6ozoC4btugFnz5F8eZmDjWJq8qvmLO3IJgOkRYeHCSyCqca0i
VSWnwaskTa0KXscaF/bES9al0rf6HExVzU7OW17h1N/LTXzDakJsSVfBjRqeSXkG3fpnhiELKI3z
U/saJekI1fhCjDEfHclGzAeCPAndtUo75QNj77Gm+BUD2fQWEC0UoiDIuH2kg48QbAQx9bJlT7RR
r/r+UoHLNYF+BGk3gfVJc+5rOwQjEnubKBt8HyEIyoLYkInNyHXqf7w+e4iFtixeT7Slu6CPz5dn
ELJ+LT2846LLUBPXTHtGfkGvP07hxbgWsYgZHWViCOoTLJkmsJpo5a4uvTZpm9y0DhtLX529zltx
iirYgiciPG6gmJQxdDc62puwHon7kVZXWsibNgYMw0EUG9Rjnyli9k/oIaV/VH/VjaCC6GXglH00
DvZe4KnSL916fEdb32rIpyOvzh3cSvIHqFvd/A1V075ZYXhTQlTr8w33zpOp+ATB0hUi+IN8z8T2
sPoFY0H6eFmea2zaVg5TCiuRi4eaSl6z3AYmMxWkV2bDsXvAocZzekXzaXpA+rvQNz7mpa7QWASj
9WGtIZGL7hHwDPHLf+dR20kBOdxgNx+rmK6JD1GEoWjqPzUH3cqqC7s0MnGuoQwahHnnUJXGPdGi
AD+Mx5Lfm94Cozl4zV96IL1NmsnNtq+e9ND5+2Pp0FrMxEgww5WIoa3Pb1sbHkgR4JEFyH9N+ALf
w0bxZJQQ9S131ou5BjFsv82Ir9ANzCCk49uPCUXGhQpWqPpKHym9eIG6pYa4d8i5EOzv/oFcA8wK
cw4y5VEMvIzUmAFXNzwauSI59IZWOGCVuzkq8IkQNvztfdOj5eqlynUo4YLslrsh+Ck2Cy7pDwQO
xuecFq5ci/SsNEKK+T+lNTTHhhLataIXH3nG2uwjsndsudBHO0lan+QJTEBJDHYALobPpMzFy8wD
CpDRldzWGaFMX+eL26g5BO6gCdTIvA/VS8fdNZcaUqMmzuoe+HKUJljdWO3BiAJh11b5QA9yZMsO
03GxApUZLdIqSTpxi/AV3PZjP0nAxfppCRAiVyaGGyDDqgMHe81H0p1iZt9Vfi82eCpSizslGSZ5
8itBTm4WkR77PPGWwdJmJlrugdtQRRGjhACi/O/CvauvBf/szo+bRQPB1sZrPjzHinKmlfbdkSLB
Wk99Y3nJYwkU3qDs1aFBCSfra2auvj8VWa/tLFHvyQrNzVY00TpaEmR9pcyffFsAKJ8+MkpG3/p9
KfHN78/C2e1uQlnFm27pAtUaeuzShpGiWaax3lqaJMQRB6VP290ua47XOVUsSz4KgJYZVztv1TL4
2ESm4/n+MULXRshLrvoQJBhHneYm7IszX47qG3NkjBHRwqGRw33IAzhG4bybDDqJVnXDQ7f13rJr
ptfQKLDSJFRAklLheN1sVe7LK/tXen7+eDklPaBi21jnrmV7i9JihYoSZ3CmuwKTQSTqKYsTOMO+
wpigM6u0gPlTJtooQaioCnBCoYhED8kGEaVybkL8m99tc5/3IEkU6hQKMq3HVe7ADQJYdRX3z9x9
RQ1lFFcUYOIv30aA4ANoZM2T4eZKh5q450r2RaDzXrvIR62TosBGMtJi1Gc6whTjISoqhUdj7s7w
qUAx2Fxi1Y4eIzrNsUXiwrFNWjCOnJ2JAxJNJmAMP/XWf86jTgYCunHEDdELG9x+mDvExHNSPEX7
OQ2BDo/OKrhb5b7mIP6lWKF1naDxC5Cs6jwMLbFgfMxL5p2/66aypF/J8V1iRLyed8JSvIDWv4eW
DlVeSpHm5lMp8adM3Pm6ERMtYZeuPqAag+K0Ajmh+LyYuVlct3Ml9E9FsI2tWFJVy+DBpJZMEeGg
94WKc67attwGdUEPVJwb9t6BN2bleO7GD27+wLNJUTjDVgnSYogE8gAf20cg6Ofrd+5RAluQtnY0
TjwDNDJwRnMlvsOs73ZW0I6YwMQA6G5ajIgwpB+5aKFPslDK3sb1zsal5C086DU4gUe6wQjqFjM3
p9BwnEHPj2hFjnQrTP6NjTjRDnj76nYxtKUBDjfmBUdLUfG/xhm6DUkc7UZxI7jizakXDUbLnEKQ
zEjPtgFycdRq26ZqhrDmodWOaygMqe06n8FZderORd3PuKQsPufGhJbklOSFM+LdOZKwoGXkOIeL
Pp1MihaSNIEk+tkRt7fY8/6rKiBk9IRdN6ISoHZzH1rFB77eh1GtPwvlIIm796Ff1yPRcl5rZZpp
/zLFt4ki9Ej6GmQZ+BiqlzzbhFEPRC960kTBq9RxorkNjgOMgGeHFiIaZGBe6mB5ARlmhEHwcWKd
QDWMlA8s4y4icWE4MZtKYJ0Zd2UacA2KhPgAmh7wMMAXV18bh6O9ghPqKBsI212YKrAZOLx+uDIJ
W7W1gikl6c46q4l0zwpnxB73T+9d/Og7erXyk6ZtlMLhXqypInITWIjtbnNjxTA37MLkSO50/48q
m8SAPds+WvyNtRo1F89cPzWF/vyJarTaHoSBa8s4eCD+XjG7UxEauWOWdguNfBub5uTiR6yqLcu0
s/zMMfYxpLyY6O3OFN4CFS8ERb1p9po2vtbkTB9JzFv3NUaLzwm6AOjrDG4MxQPGK9BOiWi1n15H
n61f7DwdekfMZ5hv6XmXiNQs5eZ9Kt0jidQ6ZKxWTq/c/+Pw+Dc+GsiIt9uQZbntvhFsGhjzzSM5
q7PaOoMxIpMkey5t8GEqDjy3g9Ep6ZgTcGUyCbz70bRvPY61AhAn5R9YBvEqn6qrqF927eNfaUhe
Yw5C+m5nNLpaznzAhlgxfGFaTaV/rvwNDr6KrO+cwQ9QOpX795FME8AHcB0oy94NtewEVVlVKdxA
EcV0rpj76NEXSryaOq7CBVvLbUh7Me4ze43R0jwu2Jluf00Flg2/JBDLFIejS47kHLUeNJGUHwei
7BwSgqX+GvPnuTuJTTaes/sgLdi4Qmjrp5DFdXpHMGRqtDXZ4Hx6gIMtCp/3QXEwks6BT18QrMcS
eErAa+vpOQz9D2aJAvGDsokLLHWhljM7g/TwfYcvs4yAZRTUV6JsfBv4S0+Wwe4P4saGZhwhiPAK
Sdz0PK7SFQQrM63Jrt6g143YKoxn3hynlT5ZwT4x+Stpk886v0bUscAXdrzVWUJncCCT0xS4Kps3
waJqOjbmkoPLoFgfNDYkIoEkQR1922b1wm9VIx3FtVO9g5sjBr2TR6EuEIpmLzpIrrBC2KCciz1K
cnNmm1r5SniqC+domyrIPf0W3fhEV9XtIP455QBHEf01uwdimEDM3GRE6nlbg8w/4IvL/uRgU/Do
zJ/WlgF7sLLWeI7cbacxr61GIRcKwJ11zdjbWhKOIwwbregcApAUabHNRAxCkpbwAdzz1VOjdfSX
i7ptEdF/3Jy0e1QRuXSsXEZuOcJLPmxSBGKlhurozdCtSgwj0HuX6oiPXy++Zb1M8FxmYLg9Yi6V
nSaoyIZPcNlDLQTxzB9ZwXfWnAzx+cw0wz9QPOU7lwNix5+hiQucsNYVha0tagMtc51VRoNKiDiP
0CzSkeJXlcCQaflBAV+qU0RMVyU9KkNqMqOZROu9yM4XKYRwgMK7n91y5+cZaU1Gug/SNUmLWZep
nlbRkBzjwJ3AxhdvJGHbJa1RBZ/MHvfqnhTMlhs6ZXcgvVdwk5+qxI9wjcxlBJYeVDS1FzVmPfIq
Ik1SkgBOSG/8tYAJ/lqjAXUbMytI00SbiWIHEPdK6Rilb2YjlJ4SAHTSSU3hFFy5CUyyTg5ByvTs
CpN2opZOBA6N7GhsPEZ1sknvACYuc0z5kx5bdp7/CRmOJ28lv0aU5r6AgFc7uEQY1ZicpiWpPoov
1h+4lmtXhxQFZtAeiMVVFGHrMELYSTjD9MgFrdUaWAEzxsL51q+SItAKlkYeVv/PhVJGKoKGSkie
ZRE3dozVWbc6trX3kSZGU6wgxKEQ11x7Sa7lwWsfJsnmo1othHes6fa2wM4qccOztHiqinppn8cL
M/LOGpK/XldSlmYjm1vLsfMH4NrBXnWVWlT0leVkM2ZD/O71080ZSA16ri76294mSP2/vqVGbNcF
MXVXICvKDynXgdKhfraNi59jGdt4I6x4oyIpYMpqCkzFi3G4DStZccNO8kCnSJhsMzxSL9j2XSQT
SQPaUKVy5kEt0zfGdlIys8dm/CToQ2eOn4QoT01KbCEMdCRCHVMCFjQK2JoSZ4qfsLEFmJ6SyIJj
sX7Ql1vuBsdRPQd8OhDwr8Nu0ObMlWPw5MxJSKZEn9V2Yd1C4ftjo+B7DirNHsuz+kg/0FtWOQgy
OwCQOprfx5yJwHiuJx6F21yWk7x4M8N7zM6zBF1b9FKyjel4ZDkrs3ekXIaRraU1hCeHGhV8fObg
hJan7N59EPebHLJu0hrVLDcxIWfhxz8rtl98Z0tAuGny9agvVlE/t4IJVEze1MKHT6LalyD5i2UH
inpx9jomuupBgXN+1WK/CKDylSZzjhC0i61Zd/a/t0gCem/xGLVNHAams7moER4xIxvQFyhnEjdH
7tqQaqEiYYPuL3JQYB4AzcBw5nIi9GV6YtHoE+fzX3EOMrNkFpGT08PsTV5o4H4VW9P5DYQgfAGC
DlxUvi9+pqfcu4FKwrmvR20eutk8jYlZ2oB9/ioc6FmDDCY2Wto9auhNiT/58UztNU1vdRnDCBqA
2beiq+4q4HV362yfRJ5fLFEiQKKY/5CDFiqVjJgbBjZhfQthNgkCSIPY4lTtrHRLlqWuxten7319
60Mzto2bPZcWCe8tZrG/FbuxG3Q6HhOCGT3Ld7asAHYti2+GBIkc8qxobCXSVS/WqTD5rzIOKot5
70gJ2sdV4Lo26J3HZXCu3Y+YZRsd8/RF6jP1jr2SY0RJe1jJqgWHYiG4AJJnr7Nu6Gbe8uD791Vf
Dw/S4SfKUkY83HNno50k/J/UE1rueySeYgnxUqTuocgphDUSfkX1dAv56iyDzzes+ndHjJxrP1Kg
VWZmkJExC/UHTo0nu47XExs4OiTwxlQ9P8oNxPE4MsS6NYN9V73foAdGCi16YjPGrubMWm4wNGcY
Zr5RRbkyjZ+IvAf7kmaDpeIAJp/XwrwNbCwRwpS7D/vKd1/lQn3GMJxSzQ6tRIy9xOvHmLIO3a/X
KmTxSHBZsTKokN3+1yZpV1jEkdFIY4kkfN4j1WdRmUwx+7E/wquk0AFqGAvnJGA3rTBDmHCbjFnr
FC/f3N6JYXo7cX/nYeopjIulmVw7JWcbOlr+o9jxEAGpd/LKCqYI7QyL/bLX3tHRUoApb5ozpy27
w4g/GkN8jdk3Ck59dZ/s6NMzWdx8Xpku6cLdLXPsn2Z77sIEDRLVxMsNpD+6ykWO1BeLMgzq1uDt
Zkw6LRSwgAcQCH/e9EdibPNeNauwTuepeMCM9EOXDcCEgwrlJJFNsvs8qJYxXQWekOso8uG+BGHJ
noDJ4/4yV7r37QawqWyAfp0eb4J8pJBz2qDKxgWfD96XsFIhlMncalFox8YwoyJ8KGF6iUoJZDmk
t+ViHPtT6zQVS4+xpxRkaM9KIdiqdGXV/438Kxbr8ixNHsbgU5rPpHEaOhDUsx4bE1tWUEJ0RRh0
omarGEzGySxfWBseipGJoZSenSdkzJ7DpTLgUN21eKre8UZNVjVDidOxE0hELag6YxKkj1mimnvW
+zS6lJPP1bEiXKhcW9F1qcWg0jvDe50YgsFWZ9Ki8Fg9g305SMt7n+jseeAnevC5WI7kN0/EnCkc
9DEehVp5HLyGrvpJCfD5MaDFp68BrWqWeMvZBgKoa1KLbPuzjKrP+uz2of2jiDa4XMI2vFM5oDQE
uhO7hP4VYjgu4MPXjS7SFLCUyMoLtFD466q2rm2SbJJLH70qj+pPDei0alDbF/EBWMyLL2Frp9Z0
QiW6hFfdG8eXtjVp5pAWvVzaj6HylmTdVGCbGBIl6yWXNWYP/LJm365mvyoPNdlsfsEsyliO6UD3
moFxDHeGXSeWylWiQPpApEHbBwhhgq2/ZoxmwWOoXopv+Kwvd9s7MiyPBINIIkNwcAQ817HAlxkh
g1zpmVCsQNqA7z/9zLVoeyxAHEROjhZghpAgoYqLyxCRx5hgM99TqFQpPMxkDv+ymx/SZPv4CVw+
ZteurlzE38MjYoRPW745/TRumayXjwitHecveAcxAuGRyzr8n4Ulmn+MHcWnmyPYWjJ41wLk7k9X
LoZ9z/7DB+qDVDvGyD7n2ZlIuhEqG89mjDvb6LQBBebV1ASZu7MBSYjFVgrosrLYN0TeJGem26od
LuY7XSEVk+fHm/RjTCRf14z/IrVp8g60y6hOQTQ9WgTLpJWaYCQBFEcqS7TKJzXoXaz/8g3dpOUF
qJjCKvpzdlQ1b6y69WDxLq/fh3y/sjGcXAOuILePBhnC0cwTnnXrkcEo29T4frcTnbuw6QuYF9jJ
LW1g5V03EoyA0mLfVRhwBbBG8kehOaMzbOoQF4r45s3didHg4nP6RGz/HS/t1oPDi7dO8FVO+VkM
gCRmTuWpsM/hYP9lMuW+nmamdnMxkkDp1or97C9gdNS/mezAI/DfeGp5Yv/npasbmbEt7rmtJlwO
NHgaxtS7W035inxvQYaPntFHuLCaeLsbRR+HpwPtue3pElbaDYIfXCG1ghY0zkYZDnVxF1RUSra9
dUU/MrfMiftGbtcBftwSXOEmoGlXq7KpSF/j4lI20+zps3V+WVD4UPcOgEPXsGJ1SkOaeIUlJHPx
QJZ3wPk6qM5FZYyayv9phD9+JWe1SUHBHfBnnQyaETD2SK42GfrayKsVtxYv8dFfrBI1kfagnXUX
Ya0d0AEI6+sZ74tcxp/WLrc5mBHJ151V1c4dFGrxh3KJnNhS+WB485Yhe6CumG6NiGRMl1jet6os
CclUqQ6ORr+QcVDJwrBS481lgeYZfn9vfhP4PB6QtE9VEwGHW4TJh+5UhiUKDFDEBrVufq0vmHtE
WY1ORmBAuLyBo3P1dxM7l0tVTMy+By9TfQKt2qoFTe9bcZusdknvNcDiY3rzTi54j/+y6ZcJFBFL
t/w29kduLVQZrTm8tKHNwZoK8J5KZdntld6Nrj9E2c7hAC7dvuFIH5/KaU+on1vJgZkomEhqLlvY
6Yh3jXsN19KfEoMbAHhj9tNcH4z7OYHNqnNT1cinDGNx6GR0bncK2lB4ZlJkuxZgC4ROb/oxwVti
S2//Gg/PkM1/jWLxVaK/FHe9jPqJHauiQXzWQb+Y/d7lWHChny3SaWJpnUAVVehaDaSPM1rfLuMp
2qFylVUMWdHqs5PsP1pFH60Y6co9D8Dn5VgVhjU88a0CVH9YZkDbw807SK0Hy0OSmAbWa96Nrfb8
DHwkaArZDo63r65dwYd/rfmHzeZl0KJc0Vp2CNxvk7MyD5XdlnXFO0lRB3CrTHQdtqaT/lZiSBnr
lwY3x0/h+z/xCIlXvGj/Gi428LMbXZw3/tJj/9xmz3VF2QOOkmhhaMUoeQuCJ42JpkbAkfl1pxCW
MNFsteu15WhOm5VMUoqX8BcsJP+DqYcDmdR/8IYbPXbcHj3MYQEJTCx6xLBNygcRr7e6hmCJ2WS4
exkeqSZLuHv6wvpwiqmwJ5kZypxk8phlvDgQpR5svhl1wre7WH+VKOFyxLTL+gde7MOkNPIIihrC
6cmS8Byeh9Hwrilh/pgWoVvchSpF4c3H16k3RXhSKNFwsDw20BkjO/FMeDCCrqH+PDjZCFnojCcV
W/sjQSXojr5s3e9DIpPW3xsdSFANsedTocHo44QzZWTEIQEtgYwFSeixoSno14gRbZq1Ae0omOW2
i/5TinBl1z/TwlBgtZXkZOk6ucM5IwRpvh83bM7bAiyGckpvcQS/cZAwLGdwSTJx5/kIgpc6cFF6
fEiosKyByecweWBbCLDUxb897F9jVT+7GJcXcF3yz5sefCFytH1MgGuIYNmsAIqrG6h7+03SMcUm
ujo78xgqveAChCrzGXcVDg/tnNOfxaUZTuq8fkkcDVJg8tOps+VVF8OIrOojXSjEyqUsQ+qziSiz
aJ/rFX2AUe7xrKo25nTRxnPRpAZQLEG4sGCeIFc9G2YKYlf2dzn3fyy9cBzykASzrlY31DV0l+I0
kszZAI3GUg1kRDv+bsTI+33+bCpPmq94awzIiBRhxqsrd9x8OBZV0iYKpSq7CGprblNLYS+Lt8mM
UWQCfD/q+To+7uPrnQ6EDXmU2XIUdYVsqVLSzdzO1mLB0ombjKGVmwcLOXjsQCzs0tVED/+8snN7
ZzqcmDFmkbw56/3NgZLkz4lBKwybrh4aAISbfqJHJ3K9KmBHoE9vKzBvhAGJgWzim5Rbt2BszuxI
p/w4z2NXao4+Wx4yGUTlc8/s/Cx46i5OlR5o7onGuG9ocowCvh3t11c2hNh0kC6oK3akK2a0imkL
LLDy8qacL+4W75oiIsRSloPmS3tthwycxFijQ7WhDLZkUs5Jqp+L31Fo9UvPWcRVNjQemCTxBKxy
fgqbyf6sZisa6ynoZ6Dp4LGQvbJye/wBEvFEN1KvtPF1+kS7og7/nbc8oZu/tlBPmiVGLSFuxfZZ
A2k2HeW7WUtoPcDOq3ZC5bgD0FwE2zOo7ygvMpSvD/mzZ7ND207bf9i2CvSkSmvzNwd6A25u2IXx
mCfmLginB1FtjCEt7+WN0ELY/ILSB6TyU6qyVmxnin0l/CHh9wztNac+2qu6dcNfPwnhWMay5fQ+
2thgpq8uDjm6nBsJiaLbJq+2j0U8g+OM4xCM3Kj34nGRUfjUMgx/giCyTTLTsvjuW6TrgnK1ivce
bdgrHcsHSIucbq/z992IhUONSlTGU2Rf1xTefwc3uftR5U/CWWRQM1AnAVQS2UvIDJnFjZ6E79UJ
5Kb/MBIFyiYFwdQrUt5ntoK3WtbcFRkizQLr36qOZxuOTTQielxysS/rBG42jAef2N9iDAt9tz3n
I5+ZJQyk90uVvp2A2b2Xk0VoVjqyrbzWaV20FHDxWr5a3parR8NfPxGEI6G/EsT4m7uCk50ra09Q
DGqJHtq2LNzRRvhr6aJP3jqRQZ6GeTMxcOXwCuC2m/VS6qhHcBHVN4mf/Ns/ZayKhwCfJeGIQS2M
hvjyvuWKYnvS8HMCgUNyM7QX6VX7IVFzpJk5lmMa9u9K2cVDjMkasapsFALhVPmCG5ra1eEHiEPa
hwAQb+q8fc5z+mcmNDVjxlqsTXKGaZqQktOm3xVmZGv3YTDqqMoPPFOxK9FMJwzOGyJjTgBGof4Q
Olzm+0IIK8npZfbwdP66b2MVz+S3OP8VpOHyElHKf+DAwBxqcbPPCm3TH6FlBRJ05f2he4wj1m9G
I68CDGr7qhgNxRFhY5njSX2b1gjtTwSvqhJh2O1w2zizS/Ng7HR4T5RtQJNx2pWnKwFEyb4WHnZV
La5627FTg1O0y5sQCyPIPuBJWT5B0eY24ZPdEnDwuIgxYupkYswtuVgWWWiFcX3zp5ftn4qVHxW1
ozlVLn4ut4T/17yDd6QecNEp5Y9eBIh+aiWAvySbxLcfzVhNJ86PF8228k7bRT+Dcn4qPHN/baXG
XTG01ttHaHYj6X/vY7ewKK4QxlgNQF4Tc17l4Ce97onH/G5VvAhCSwPGjGtFDl+VFa7rD9yHNRn0
ZX0EfkVZ4Y4ibQ61GKPp1qSNprxmhrDeceQ45u0LWv7/3EnQwvHbAjp6bNNi8+9VvSPbipKgiXn4
3SS6AzalLHFgbQDV6OnFn96h/jD5JrMaft4IEqyA2pZjW00pHguMXYTC+53PYI2MeR24pi3eftye
IIJfGnw1dCdu32uLRV5+ey8Q2p95Q+grqL+ZDuZN8YU69ZpqidCsmSGYjSU/J2dr3YTSz3m5scwN
kPj1ytPo+ff39siH0JW3fjYAoufrikCmkDkSXFYGULxj+x4RJM+vBu5ozmK0p+bVhdsHHa6gDKC+
1FYvo3LQ9kRfIxr796iIQINq4cA9WI7CHOvNNK1mkXWrOYz7iWJiH9VsoXR1nV1BXntBz8f8n0rN
xCHflqPn5rve1XoZVmIK8WGWnX4J3A/5wFc79sXYq9ii8QLNTydeTk4hBYa14oaUK0AJnhXWq+LK
uDfRSh1bHQyCUV0wHUW1k0DWJObmQbTOR3tn1dDVjvkzmWy7+rTL5mjYboaay+coVFTM3ViqSDPi
ZVRsEBGrCQEj3XVRA1EGmnUF+qROEbGK+8Yu6v9QY4K0GPZKlKutp+stMXxfVq7FzP8kcXRRQfyg
lzSdppnO8lrOETZqgV83bfY86I3+j44gApmnG30L5etPvzOXZvz9j4n/fw92l5MnqguYN8Lcby7Z
dFDdf3/YoR19JJdBejV12ZsZ5Q6mne3vJZnDubGV4zdfwQPBEdSwjwmh1ip3POLCKnWLTN6LLSrv
1+yab5FAyPxw1p4FG5cvl/kA2frdztOKGRw4iGDT0NNquUlurflyYLFj4doSGreDIBYpEP9tp53a
24Nzd0npk1S4H7v+p+N8NrQPOKgUC3VCualKRzE2vdWValE3VXmMfvqk4hZ+mq2Wpwa5TAK7uQO7
zrm5Keo5TOwQSmF85wbSU87jViUDltBk61Dvd3ibJXCEufsET2JViTAU+BWaxnKVD2YKDCmP6PkV
skdm9QXQet+ifAAIgXiVgZf9IO8xNTdrui7OzWM3N7wQxGvmGCIyqEkgRfhboorEHfbwJ7euG6gy
qEyzW9sgF62zttQgX5UoH/BYrWDAjed18k/yRC3h//jjeDsQSt+ZS9dyQqmeEanERNfT943bwQZu
xAY1ToiKHI8djFmrxt/0CMX8LrGZ+NOjSDEZOfa9GL0zFYvr9U+IlBewJQYEDxrY+XpHmZ1uLm6x
BsvjEaHVBEYb8FeQD4asdeFq3IopknuzLryHzerwxPdHRebYfMy1deRUuvl6cBGw3hjQ13hS9kOp
SQmcwO5uo8h2kbUnlucn0xI2CJNG2Ki3RXzUHiDQ24r+S2OsXMLXFYaK20Abu6GtqhQ78zIB9kfY
nJsim0iVyGIfId95pHnrZPIK4P0eRvfcyw6yFI87EKPZaYTby2Gx496z1UhPYqxsVoX2ZIQjxJH0
LmH5YM8V1Gtf0ULl6gtu1ThYuHQ8e5pAVi+AXSjC/OmbQwvJUVSOhLANrMrt3XQFQjOOJvXIqejD
ssIjex1o+CxDbn3Syh9EZLOJXIJWI3O39swMsLvCNWhdE3prlE2c/1EUa8Tb9vuns8w+6gPp6RwF
EEFLkxumBeLfAApf7DBkrbpyBoTyk7h0LCTYh4Xe/APVrlLyk5GqyeUR+PsfrGdGCVFTSvPpmi89
NaNJsdFn8ZUt0BxfzgX+K/G4QeGZzARGmj4HUT58AKQWI8CP1J4s0x7h0A/kH2RMEN0p1LgkprYc
Qb7QhbpIGimepWSFrnOKmkfFhNNsSlfsbjYQmD6HOYep59XtIOh6Azan93IrZXzLPyXzkVEvJp4R
PZMi496bALjduM/OTuhbYNkO342if6+lsab7dqMOVC6NDRefeAIrFOdhrtlXkznCATeptCmMU3on
fD+S04/Q+4YfANRZ+3lWmWOizFdvwIQxghGHk2xcriuZRfSDh0VYDL7f+doprOUxuhmAFWtO2c1T
xRrd1GxrreOf8OesRWW14b1Z8/3lO7e7FHG+Mntnxg5pTGrWSiUqTALaPv39GzDhJ2hnq61MGEU8
sDR8o669+H6NYNFbbtPScS7tzXQAr0Oaj13Y+p9TmG3E0vy7jDWYbTWRBRxRdOHB5EIuk7HwozbH
J0MeJjaOa1vazKtnIy6by4zTHX1X4mbad2ZWSKK2pLGa27K04Dbg6UmT/kudxwDQD8CJZdgMUQ9W
8UJ+5EGdH1mkemxkbvcHUZRSSHc+W+9uyz4mobkVqxHzVqfG9NEZ4JXkYSHCoH5tRxhD4WAsrte3
kkIil25KaiExxv60CKBddQ8jI5yei7K3bMrcYlhVp1qRZav/48Qw7AS21XmVZNQaOvnKezYT4fLz
1Q8gqHNW44Dsi4eyh4N8BgB0tXN7I4c98+x/Q5rjzmFlXMxPS0mQGCyth6ER36IJGJ+FPpm24t63
ZXrLvRWILISVeLpnStk7AVLUC9km61ZwMJv3kThgXyeElexQ0812uZYrSc+RY71oufAwckiGwSvi
HjwVq5yHDe7eLTXv1gSz/YiDb2wpWmB5CU2Rffbf0a0HMdsM32KsioCCNW8ezYmCW22m1UAGHDh/
UkkT7x2swBCNqc2XKxh+B/sWkpOzDtupkw1UDar9f9JmWsGYgWAChf3O1GEWmMrXE419y3ckyhmj
waG7e/DRfls9IvwF6IYWrhyENC53PfDyISbF66VI1kz0UwlEloXodUfYl9xP4wg8rEcijXOeg0DF
38bBi7XxMxG/KY7OtGZnii4GqturzYgLYPqR+skwODo2cMCMUoc7usxycy1tPUKmnJzubupUHfiG
ze8OxOaa9qrHcxWoYnbxycD+m6lQP+MlZLhNJpYHfppsdmRuPHNPCwIIG1qhYmW1G1HD+jh5vyFM
ayjkL+MP3Am3IdiZNgVWc70rHEqrp3Sor1kT+lyUaCT0qfzjRbBS/tlpHWaqocKK/qG7do0t/7R6
ODKbUnqyLJf4St7KB+xf1h21jHxjU4KrLGeX7H4vxrX0lmJlhA0hOFeBxDgx1ZC6Zrl6gkNyIg4p
IdiWusATy0Q219cj6G37pzd14Q5f4pt2gwYBxnzvwvV8mtNMEdtIa6By5mN04qc41CY81t3MLWSE
zjaAqAmunTm6a8oLYHwkNykCkNhNM00GYRNfoituMHCB+5DxRUrsNg+RARX6bigEW0ikCuw2sjOM
cjEavCucBvrhAZJovG+xz7wn8xSICeO6Ki7/bv/HCDNx8zXynKPdSYL7B8SR1cbjptA2EKGHDeI1
l3svTwd9JMzQI1NIeDIG0iWCrWa+4LfvTlWsZYfhxdzTiiXqWJtQvh1WJury3k92eVoQ+DoEITeh
DsIequ/+wBudfQOQzSGldwr0WKbMkYcb/CKQeu/msG3jyurN/OggkHk4Getch+vuCMDeJ8whTi9L
O9rqCe0/V0yebru7bx5V4nA7Kg0b9uAjNnLZEnHT4ekiVaREqjfCPjKI1XFIPx+ARk+dZTjD7m8Y
2zqgejGSDV+plrwH+I9S9Rek9ij7go5AH5rkIIkkRuxmXjusVDzrXldoM+RohStDIp7VH04/ZT1M
brOBDdRxlZ+QOlp457j3w6WwwhCieUpikBaUmt1jH0pM9PoGUlNFc9CjINM7Q9CAIi3zun6iv+Tu
MIjom12oep+u++2wI7+iu0Bl8Ew/iCsWFowAa+zgziH4Y68X3IlQBoXxTm+vF+PcgrszXeD3/OE8
Qw4ezOYbZf3RtaG2KRGr6IE3bE1dt5bdCL7ihoI5tuVhf0asG09Iq2EayNj1RAxuyIpg8YXjKgim
pquH3oXGzZbHISNBRDH9HmBXLvhcpLcCLrh868CVNtNERXUcLiQI/rEebgC3F5OdUc9Sq/VnvQkY
42SR5GA3BfAmiNjR6lwJpKIjAW6bwYoFO4xRnjCokv+U46ivYFwP4Xz4r+W/KAOhnkKal9qyJ26W
wsJXl4CDyi3k7ftu0Buu/hBMjRpe1EvI5b/btwtmoBWz+XL84TLMdMQfHKrN5FwRqX9ofBUddoxE
HKiZXHjZtTtnTZwpYk6wMiXtwuH5Fc+nGrfevXNGKuqwktqNVM5jMrtY9XdO/fa2KuaWqmbvPVgI
Dt9Db7G7OEZ1n5U5hJyNa2CHpHLCN3GKZvFG3HtRMhI35C/FPJUzMtYbA9EJRLHeFH2rkbj7rg/g
V25RDIIbW7QpQrn2O3l554MO0rwdAol366ZVxH3aqTkFMLIlEyiUP8zH1TOdZmp8Ef41fzKIzlLJ
1DmLUP6j0ym9cVHsNysBun7ShaXWdmlIZD7ihM6DcrOXqheK8EFgJXO0wv70FCOf2A9KNHonhLgT
b6oxYszK+N1tKDQ9JabQRjYa35An1vtLr9W8b5EOIEnfglj6pf/lt9gpsqrUAj4mRT3cFKtnEnj8
/44hjTEPoddh6o2qN6a9yApVNUenUoLmeP9M0C8v0HhLrj7pXUoE7g8Yn+zHu+YjnaYbSeXtx8iq
UNtyqyDZrz0JZFmg8z7GL7SHEeqzL2qSeAUjTEdNvKOAAP1WDhm93+nWfYmQAbStLB1PxvYpvgl7
IqLtqtdk1k7AxJioepg+2xf3Zug8WcXhKuBHD5801uPfuplT6tfNaOuGJsZpEqVO3tsLzTY+4lp9
CJtpP8bfOoRf3+ezciWXjn202gqBxg+dx9qtd8tgh5240xA/FpwfsnVodr2DQW31RDCcBzhrLzJI
eOmXd/7rZj1xShz1q1efixx9Clplx/Apabw349UMZGAhHhRi70Kh7be8xy3eCoCpiwTrPXqoyycp
u6RhZHrpNjv8hno298AvzEprbtjYRX5CZkTEw3liDeef8/NxzMeBlr6mqU86ONaF3AQRllC47jos
4eINKJTs/45Ar2UXxO07uxMDk5NW9HBkinrzyBBj6pq4YXNF8pUrgmUpoJDcZnnenGyhQX3W0G5E
o9kmpUwJZXj/gfEbIR6H9pI8RhSUuAywKNF1pLYKB+RmqP4+rb4N3VkJSqdHITlyveT4uLF5AWN9
YEWUE4w1CiBFmjNlafHY0NDe3N+IKXWzREs51lCLgqK+8McQkdO1EzsaE0LQbh0wsNKsEK8OSk2u
H0SsBJv+gug3EJ9FikafYxVLcqgCpHZbSoTTcFYBiXTjKQm4dldl3ZwgAxl52P2A4hJj4M5cfDiF
oFPE/hlxnt9XJTIiIXgZZOkRsQu6Z4N2yjeLTHsfpWx5g1RsDfUIIYG5DXdd+ANY2/ldo7htTTkc
1G6HT2SH1vmufAjA5z+QCpRcLIQZev8K9faHin3cQ3arkUfbc46GH25TAOv2QKiOP6yQwwG2+g8p
lwt7cKW7gvO09ecuDQ8FFBDfHK95WHP7Xb0RQSwZDsAwtCmokbTzrB0sfDW7sPD/FNYdPYWkgeJn
GM8OTSP1Pwj9c+0bi71d8F67dxR/UT3V0g2KC/NGVbDu3/n8rBWbofXdPKCTumVa+z/OPOJQNOdG
I+/XVQyN/qWPeZyTy0pO2pe+mVkmD6SSbbezoG9cdhvoFf08jZj/r0Yj0ji+jnMqn7Vik3vKV6Vn
ziwq2my9Nqx3FMRRwN6pN7d4iaROzywuNrSeDT0qZxUjAO+gh6T9grvFrdg7GGbDM3oJHVyLHawi
eBzjdWNpn8AxnZYvEso1enCz2yUYH1KSrvJTz5pRR0Q7YkmAxM8AKHAVa43qDS/twNkUuUlazdXm
Azmcm4FNDgk+wEpnYVyRdUbLDYr0WdtxGoeSvog+TinUxTWG/9tA5xV42IS+k/T0r0OkXenevN4t
I33inwvlg5N6il00EWHPq19VIz0q8XBcPhYttsSCbSKtpTCghyruTpfGZcks4ftnd+IqKVusYNrs
GU324yiNO0TCSqttS3VA4dPzGfu90excMQLZjBUL3zSFK1ukB2zkuGn5yPJT08cfb3GnbCcJmGNm
zJPlT1fZOyvYqjz5f1grXGGMz3ArTsqiMY/0AkF28Awv9+xzdPOEIfi0wG5qd/IkO3jU4IxT63kY
Rn+bDaKcX9hYYiK3TYMjnTxZW+1pFlD037IQiZiNvg9Bt56kxngo8Stf/jGJ8HdDpLBNfBiACSdZ
5GPNRWkfefnE6MHrNZwAKo3T4rfFe2SCc7PLh/KDWhiV+GA/KNdPgUP6m6ZsD0m0bPpsmawhdf/L
w06NYMkqbGTDOiFqhhkTyoqzM314nWSxHoPdw9KuduiKbumk8DHLz3EwgXD8RNeGvpgRie6okRPd
EAD0cZ6f6ZE6hRwsEtpiJhruWTmtwyrnyVhnWN6sctA+QzJivk2GMPluWvedu2gbZHv+F78qHa/r
vh+cdpQBAOtJEnpiAf4OO4FXgjHlcbO+DyVWM80ZOLfU+GqBfeKVYmp0AIOPcp5FrspmdPt2xEQ5
vMSmaysg9Qt4vAP3ycHF9vCnUmaXVCI9YF+mbP0k8xqfq4XPH6laHe/si3ETptM6qa7wQRbFTKiA
+Skp3B8wG9xMyqvmxMO/SAemfdR0jsXXUaq5oU+gVdxKDXRx94qflkwhcCbO696rf5ozTj8f0pMg
Y/0jpTaYMwoRByN8mGTDIBnxuUZGCxWNW3lRhECYA2DLEV+ZmJeP7W+H+/mKlxrT6PESElp2Sq9b
wxa6Gcam6cr4yrZZMCn1Dt4Pjr9PyAKqD3pr9QMvYX4kDiXdy8I6b4i8DiASOv0trUZqeW2PmtNQ
E1YlhNF5o/ge9uox7cAUrpluYqIwDSuAWLCAzV1QCjPscdSr3wweI0IOxQy4pIDuPFfHLatFNnRX
8WCSS7WWRze6OF98ob6vJnbQwTaKpNHM0JiqIldm+B58HitQzK9gwzqoJw7UDhtUEVbYhRhCZnt2
e7clhBvgOr4tz4jC3szNGyGDz6wQzpTD5+IEfaWFlYQqWUAArsexEIxdCbmwoHuTfTHHGUg7RvCv
EEPs/5lIXC3mpULiDeqIcMHbYL334A0DNuSs3NT0VJYnspDTN/IPEdJpijQHnTpgNUMl6LHwKLaE
+0DxKQ+1mgYmCN/lU7FqnyM/LL+OFecpaQVPKj8r3udMiQIRAFJRa6y5Ixh2gurqz1898ZjACaWy
VZ1j0QDKmiC0ZRI5TmXgamvi6EGL6UxRORzn+bbZ8qWRkZE56ivECKZYyxEOIdtijW+AOSBykGhL
5UaUlvzBDcczQigi+ydcTkLw6O5Bc2rVVl65evf86jtGoPaBMsKo/ifZuTB/JMM0YPNQ5j2TgNSR
uCyy1pz9qsQrYhQGAOSWJb+IaYSAErK1hwFzH6pb4i5ph6ocqMD8LVCQCvePwTeOiHt0AzvFCI1j
4D4xe/v5Xoc/bpBmLl1XVx+fXb1M01+miUKUGvQRpIi1rsE2GWIIwVQgm12DLd3BnEJhVegUItYT
R22+370xXeA47JG4Hj0UGTdm5ITh7xrqD3Vex4rcKupBH3tHjsOdQOlGYKyUQBAkFojNBoHnQcVn
qzXaAaLg2WqQe7Y5af+8AuL7mtm2nqCZbUmSSrY0pXaw+KD9YxBMW5Ak5DY+bOSxFbuNwI/n9LVt
KshkUzWRPaKysjAmvWzuBfnNVnVA4Gy+Lb51qE6VhAR4CfVR0aJEj+wTg0L67fqWzzoihI6B5LKt
0kPIJL6wa0kurlie2lKTYSVQHN4GESSgV1kZA5IksQrAS9B73VHT2eZ/azcqQTxxfv/7hfUjO4kj
LbYlRnumcMqER1u59lqircPjAM9mnxgula6xWcBLqm8PdrgaZX2czI/3aELmkkKgJ1FvLmt/wYGA
EiAnW3IqumQQtvCzbISTzNCYC/6QnAxEyCl1OqFB2RWc7YZKBUeBULizRunORTljN/RH+aSgmsgn
LgUVJIQi30Rx8QDiX+8xZXTQKNFSH3rdNs+baEhf/O8+Ox61CKXNH3su9DLLZuiIQDDASqpCP6/o
2F8pNclKkb+JbGhspATqk8G1sJJvBkY73yIQYTtTRnYufyjHWgklkJq53Fj88qGmGfQ3v6Kiwbef
2xk9FkcPIjbjV8HYeQff30QjGAPpwbnS1NysXgNgSXrDd+wzb22YF8RB8jlZkb9ut6Cs+GzEp0m/
27pyAMrbC7Xed7A2AcPoWTfyFcTHX7F6Gn8NzS8mCltGJiFCGSiZHHA+J2iQNrQnftxcU2aLCNZ4
6PmKeDvcRolxN0rz2GbpO0cIHxlngHnM8sKrfgbScIropq9k2dH6SpGgyswOjYhpPMLGJ3jLg7+0
sz19LPftUYQwf7DfreLO4KxQH0vrpuzWRLoAgq8sNXBhKHZZ/SIw3dv4DdkrY1dR2gzE2u38EfUf
tEVgvT9bJeDLo1aCPYOEuozvbvyEaUwaYQ7XZlRywMGPHZZS45nTLEd1X8yX/6MznC6s1KPPo5xP
9x2DzWvyLxbpTWRLgczVTUBJXqMo9x0fX/95CCqPBENSf8By3kRZ2Ui5/RD162J1cslOYx90Y6V4
u+QsBcKNZNXwk09e9nVSmP8UrYQRIdH4qKIupfzHP9eFK3Km+IpiJ/EvXUoj/0PEuBPTkXnYwkyx
VSF6YXyRLcIaXnk9Dsuyje9NOdO/ggEhYmfUELmoY/5mPURCkNfhoI5IGmD/TaK/YYlpbSOcQOA3
dcc3eRP5lvo4++0POIKPpNrKeDaQy0KRsIgWgIKulYVLSyZYV4JqtHNrpS8DxdVqU8on811/UDj+
Sxyyft1nkFVFPf7Y/GYqxoRSeayqygLzx9h01x/j5I+B0rRm7/N/UQwmq9AkPdEgpa/LuRsEAVuR
TOaDjGmjPXFSCIs6v+7hufmVEd1PrKtIC/SxmLnLrHSdad5Wc3RHacdOFXLPMp+L/wAfrhQQ0ioB
QhfXYIUsYvoznWYboDMPR43nrnXW67ZhIs4adcFrNKQA3w/pQwfTJT8cQBu+heayFke1yqOYXt+y
tdvimp0ROf0BJ0Bxt+0l4Osjc598NiNqIM8TfznUnXfM3fS8hWwv/tZnirIoBCsKS3+0gOMsVWBh
TpbFq0IY3Gr4EDOGsOsmijxdApAPdUKVAOVMckXAXGcQPQQgKF/yKeuUW24cWYDcSlrbaxR8pHFw
/M5iJLW72uCqRBY8uwBRFSNoHuCerEKUCuVTlcMfgSiPK0epgRCJqvm83fgPfMGNmUvz7bsLZIKJ
RSpRC5Dsab5cmNY553qlH8LdoJpAmz04v+ft8q/CDZoTVPbAhx0yti+CsX2xFdt3741RHvWoY01t
EM8B1uQ1fWBCOQVO6wMa1kpC23SBBtpyGhJZuDIyzIqLwZjyh2yz3KQWI0eddkr2/M/vNiTtdbse
Th6vI6sMAcg7y6UrRDNS6AIkUt+4CKEVdf7wdf1cXqC9bvnV58hYhPTnk342vOtylYl7QQua98Q7
BCLWnAsJoAqEFgNIf7tO3dYrtDFWw+g6DkJC2gQcjzBUIfrDEIm8MMdzWnFAiJJlJlf5yxZu6gTz
leH5hgsm79/VUzS83BBprlADxQsPKSgziYFCZLph3kEEzSDNIW0hjpwY9FjQzFaf2Gm86foFN6en
13lpfZufJY5kYnnUQ6Yp3ZFNpVQtZOBsibHDzGj9T1MUGcal66UgcVgdMdLp7XdNhtfydzyiw+Hb
XnffUJKHKy4tbbAMmplE4RMR0f1rELGySfCEl6KAKx2KCYQrAyNIAZzmq6RDbpuvJzEEnoS6CgOH
8dbXbK5uM3o48Z0QJeFYOiPMw+sPadefuVcK7erggvnDyJKDBeVoNxEUMgD89KsxzZQbnu7oJWKn
t8Fq2DJ9FO/FCnO030qm/neO/dIoDVHQLHOXwKKLDA9jtZyoQFipS39SBUib5YFKzSuKY2jWx6DD
Ria9/o/leMNhDB/Nc7okqG4tzjE4PumtBI9zvmKeC3+o0auS99k/3PJHITMrQluKgQnXUDF+pvDt
726Z5JpVSBhsuvbc2nqs8xKFUn/z2J1hPtH9TgJznTK0IPAG1KuXJHM95hBO8zpChQtUMRKmPeW6
3v0Udi2KorVKhEr6GInegXmcCRXFMKIv+MPNOgZSPKQEarGPsZT6Yu7rUzRc6r8quHiQGzYMJ50P
aB/5ezdDfmCAHmUdtOIB9s7lnJbbY/xyCUjiEJgwpUz9MP//fUATpR0Zm3H+1EYyqTb2bfGaH1EY
VPpQQ0Y4Jgmqv+bzgbktX6FtkqQNVUXIVLwkLjYkrXkIr8Tmkjw9sj2xBKHkn5WD3CLeiaRFiIyP
IiLRz4DyiPoul8+k+4vi7hkwQGQ0b1dUUtWJRcSp3onIzge5VqUUm4RS66+XnD1txF+2Uh7d0UTL
D62VkscFWm6IWxzO4ZRREbiMi4sbOQAseOivHHdILuZmSn0Ku0l2ldDiktKYwSAn54CdlAbn9jD1
hZr2f7T/gxgtGTjM+qBIrGuXtPWmZDGhRR19E/u0DyCNcUlBtTAbI4m6fOI9dICN7k5gTakTXOdW
Xf4d9uJXHZoirQ3SCIwB/DwawbV/5QFOG05UCfyVNumAPFQNAmhPc7H8rcl0VXBUxLtnNkNpP8rV
tkzNmdQGjrAGSJbEiyBcAPNdRfnOFSzRugfwK8l8aFMGLaGynp0JuvQmWyHPCaoLSrzLvlD3l5/2
5xQpyJQVoa0yuMrkwfyuD9lZ9FAtagvmIn3lj869annFGtm/GIOkEYX6XyxaxfUQFwhIQfyEkP4o
a2ziAfRByEV1k9c3tiJprN6kQnrzPwiHSK+Hn12tfWNpd+kcC/LFTGSr05V1l8f4rxIqTI1/JZ9N
rLmwcs7NTUMD5GuhmQ+qJihebSszd0zZyUYf/i2kVrVuADHfRSou5xXllZ6EjEdgmuLJ+3q3Am34
Tp9vFnlK9FCHpGt9olnQgc6Dd28wH7Xntmn0HN2ZfHI5AofM0qbSy2NTSQTQWRnDlDEaEslFewVR
bJnabc2O02XKQQigTwvomeoDfGbYvuvM3vKktIaeLhDQQEsIH121RkVRseJWcozie8nCflo7bTc7
IsrQakTYV2rVHLwLC3yHqLg2Bl3+PIRlxEQ1md8D9DZYPizWRWaMc8vz+xN8buryCKh5jxRXWa8a
o/y5cS4ZHkyQ0FGsXDTCm4O2OlkoEduiiMbZwWKs/d/iLy8YScOy4SNDFTmHHxlrSeBXMw+v+PUh
wAQL3teR0kvD1GmeWyAfLImI/2h94ywOq/TJtnAZnElaegPOeDOmgqLu48a7HuQ5nRRIgdGtfnoB
PjjmHSsIsIqtidzzL9zWF12bSHL6lB2GZZrs8FlAC1prSPfKsuA+vjJbSBNVUUqtzdFAe6Eq5B5n
DwbuxarqGYk2IIWFLADseyejXTsAXkveMXnjtpzRuu7Ui3rUom2a4jZXr1CMJlCu9Nm8i8AovhGN
eJ8Ggyv8pninNAfFoO7IKb2UkaCWKJq3axPUw+18KS2ggQ8c8riEmbj07UwqwlKl1BVpHQR61n89
JXo2+okZfJdJRVcLXMGXrqCQjZlG1SjP04kCWcRSU0d99Ro6OzECzOb5yAQhiGbL7GhgNLpnBRez
CHj85/2TaROJUZqqUZuu9bm0Zho2zTWnF/ZEhlzLQPSX3E4Jim9q14ifLU1MkCCoC1SGPn6cC2N8
ie3kLSYu1r4ELpr/GqBBVWqa4wlAsiK5lRyMd3E8mGW2Kh6/azAh38vnW5HRck0BbVseB27XmlxM
dzNXremk0s/Wy/gaqYoGNIUZvXx+r5H4fWQxCkhgcn7lJNR/ak6XtUwAsbZzSsnx6r5GG7cIm+Bi
1JLrVNZLvPYSJ0wDPm71iGkscqFswrelbLVSo+lfhr5xOLKGl50qgBMatUZBZ2WnMR+6HMVZXyEA
nD5CbNqJvljTL/mxub7Vfe8VqLYY56NoxxF+uMEe3P8GhrH/OODZoQ0PGBAdcUrnwPDakQ0xDc0f
P4Up6ZYjoTd7uT8DVteMrbYKontB/dQ3xTXsU2EtvBYrsw5HO2iT/osA0TSvhM+r2Qk3JrW2dwlw
T46B5uOz5Qg8D9TInuPphbUmpzh3PB1C0kfwAnVkFjZ65nAle4CQmvEVNSK2TGg1+P20sqc2LYqo
NToBBKMjvOM2y551UHBwhN7FBsBy/x4Ut5xX6ls8/aJHqCzia7UBlgdhJb4ER6stcBKoqjrsdEpO
O8PlSA+yj4OdV/rtudylqhjDQ5HcFONSFlP/EQSGrMVhAGKTLiiF4GQTXZiz+aSXI/n8GCevm2NC
o1uasJMiIkOM2B42D4LPzewoHLzjujVwkb50zc5iF/fu715mQ3u/g/Pvnp2sy/fPEbGOXXEac66C
ns0HYloCYx0DuUFw8kk721CuO3ybCK+Jo0jak5elQiW8j9ldgnkio1/+xxWZhQRxJxJoFp8+g3SF
VYxzechaBQVPPG3TQplR1c3n0n2kHNqZA08c5hr/ptMcDUpVqVdywpN8faBjxlyI+uxvlTpqpx9r
sUgUxiTKb/wp23OekwnIuTxHXc3GApMj3+mj/P02lPHueJlh/90qP0CbMwldB4AINWuDzR0yxSlI
SCqDoHidKX1c1I594qw0PsUgiwJ3lL/mBd2dJkXkOL2piwKRdksOptXPr+/meDWCJLg46rILEUgz
80HXhZYrRHpTwXBlqshU1o+aU98LgZIokvu1gmrrvlYDgXvS39tpsgxYREastwVRx2ORik4pILDO
20KCUZrT7wXjy6sMnCizffmAQlPLxKkvHSvgcrklKazww4MHR1l8W6GeHyMWBMkrf7w+tspwoau7
AeLMQ8y0/T8qQ2/5XvU7OJCLHr7ZqWbbinio8IpTLTOvnEQipbaQv3pZl03Wth3AMg1/iIyXW1pR
zfdBfb8mxPy//6bOnPWeBl6nVkeSTYtfbYFjoIq3A1zoc47jS16N5jG14IQrreU7EIVWxqHHRwLN
rJbRdH75ZtBLkO+FtbSDsCW5uUq4BHKdKcDDTD/ic6ECdfNLoouYMv3k/aT4F6q0i6OjRpvbtDyg
F+t/cYT/ZZAI+YZCt2pUqKpme8UVYBOa1FkcUfivgw5OedI61Vc2OR2LCDSRTmAG3vdHWspl/jB8
Dz0Fr/+yWmkcncQhTrb8HyTgMxxqc12hoEPmrwJWFOdAIJzb2atP67ZIb/FQJJopJuOxO/bu+8pM
07Jsx9FR1y79uLomTcA9jEpLgT6nTPO/a95UekMmAAblk2bmOx6GFNT6huzbMrmpPSEo+MvHBFJF
rRqxXAuzfnnUTckMAj7VRLg+YS2jOA8MO+GpSTYKYC2+jqbFGkqPZIMXx7XdsQK/Iww7ezalzc2S
USwdnJGvquYFJ9/CpHeai0OF6YvztJLmcl1TLnSaOtG24MFAqay+dgw176wOKY9iBjpmUM5g4951
FYFRjvayG2ws8ugvOpWsbeliLicbB0nWGOaUUh3wJ+rizhwN5QV1ELB01Dch4sty/YfnTQqdgl9r
Xp2aljLxCoOmnQgzJ94gqBCwiMrMitjPoNMUu1mbreV06CA7bMfBDPV5Mdf/tgvi035trI9iUheX
OYsVTugjZKuwSU+j2tBVecAJIbRIOJAN9rVgrkXASrY7azTK8dYV3HHS4MdwjznlxTZr8qxUThUV
+joJBb6KbgsVMMJw65KntbHIyunQfowTSQvEHN8uq19XS1LmdpEmqHL0A/wg/5gwakEw5RxXMuFY
q/1lGXxqcKzBbOES5qG8RKVFx42s6Soj/Rus3zfKyHJSzSTZk1vnGuzX5Aww/n5p6Ff8V0+V5CU3
eQgL3tf9JH4Rv/i2SrH54MXnIt/ig2rluxEmQaiHcpXVJJO7FLkGUxGPQPfarSmNcKEefm39h5k0
DoLQE2IPDuCF2V1pyfW7NccY71DbL5lolKG2b4nna0TC9lumxe35HQ2Dndac5Z0fSnt3BCcdbZYq
RV8gJdWvYTv4VLEVj9FF15pF9WxsGdubr23Hlhl3pJSI81nHxfdNgVLkp/TL/z/Xx94+1OmfoqSz
0KSM1WusXaRFktUAVO+6wgwaTaGkI8OrP74KkJNlAcUHPkuIj8tUCad8MpH1r7N66bvdghorXneK
yaSjn3Jq4u70NS/X1vZiswFiJ28un/FNB0YvTcBwg/ZrMN/K+NQulgUhpTpnaRaHPycVSEAs+NXR
N9kKgIFa3KAnifcYVrlIqWqkt5L3d/8ec0zwzk281enSYmCL9rsFZJyp2nZZ/2+d0xMlUUvmSoUE
T2cHUfcrdDGP/8Z9ExQsG+kZVcK0lw+0WDpXSNagO3DDGqXFVuv0gSpa1txUUILGo7eNrb4xVQFv
jECffuubO83ESDd/XylhziIWAGnChZacxU4yz8SytziZiUcVFP9AkkCSYgCSutGC5Zu4wSbM2RI7
FjWK7iNHTHg+u7zpL6+NPIXdEaIszY0v65EYsOJdEPmxwmVBRC94VbxiN5meM5QE/V28zr4ippVD
cMqRpsqIu2T0uqwJOERsfSJ/Q0/NeW3ivEycJML/2P3DN1HqobkrTJd9H0gFa8JSiBOTgnhFHOBy
6eSfTJE3slwhJrIGdoCHUbfn1xWS5+MuzSjE/P+4lI/gPzb1lu+k5l14NbkvVgJtT4oWyjf5/gV4
u66C1ept5POlTdR7Kx4JqG6vvNDgHXE5erGaRkZbTZ9+jZANAQSZ5MTwC5XpPchb/w0+Ws+Xe0z9
XWigLgqpEGyGAEidxpL9t9ZgvZGjoGki5cbB5qFdIT7LWCbDn76tN+X3Py3qEqef5BKMQ8EmIO3k
/sDBXl5bpup38kS7BR4zrSuRBeyX92z6j1zhAHj550BDf4iM5ZyUH/Bhrt4/7hUo8BIR23D6f2UJ
LQdHtf69ESuH9/vuCEg0FFx/lWaoFMKK4FkittzWG109mHsFhDzNntGm4Uj5xInulndfP5l+0far
LLg8+wakknEtnbWajwADl0G/SPkJjeF4eOCWRXm9y34eL2yDF0sdqbQoWPvHcSxC/goYHdzhW6F0
lH+hHO6JaOroLW9y4yHzD97aAzZ+I3gpS3M2ddFtUHYcrPf9yeUe0oM2Tlgo4mEcr2c/yLgyIlf5
4xonC++49Hgnb6lz30kFltiJ1359yuKNXo4BYcDwMV+wrKup8rtgGiVxjZOeyPrKKCD6VzZ548lO
eKB2emwg3x4fC31TdFo0mr29ufLVjqYQvUht+IsEN+qW1il0FTMt+D+Wj2AhHbQT/wN7jurYgaH7
LhERDXvg5p35jkFV8fFZRu/EJC6HPzhimJLi9j1ue/iWIPUiD3cdhaN6odJ47SFITYFAT8yud25o
smPuisQ+N2gxPpQCetBEtaK8d9LnPDAv/1dCmErQLQK+FRb97Jfl/xRXRVAbcq3jBJPvMMZShnoe
H3MJz92fAlUHVC5ULqciR5YE7GjjqA7rXIazYpqnjbfOO0ivebZ7tKbm4+rkRt75KgiM2FBPWWXV
XPL65XpU8yTtajK7TGXQd74R6mKa2ERbruFaJVEVQT6NCElH1OPKqPXP0vUK3LzskbuxCW4fVHtR
VBNXFrTwthgguAwhVbk5tFInLC5DtWKyQ6DNo7m5gI0McAFW8QkA0G2Zzd5elxIVpC7eOXXO+Cxf
FIKBZv3KVNs+8xLl/k4xhB+H8rjDl+tEVr1UEDP11FQEuopdFivq4kUP4ABXut57c/TF1wBU3D2t
ErGgH8oKLQPdjNAngJzagn01ouMDnIdWONMPTuApNxlSUjXhUGqZAaJbUzFxD5QnTDMQhEvPDQtf
geB8I08jvORWfOqGItTQ31JNVl+1ydiVsdKvsMuiVAAxY4P3dWbw5XOAkJesGLvfn2BESAv/trc3
PZa7+rEj1WTw6WkhPqPprglaP4Xhe3HYrlexbmEXgxWWpuj4UMxw/+QnURUzjrJXfGf7mNRHatb4
wUJO2O48NPZ+0gh7lD+5gafMJkm0CL6EgwxxcuiXHpRPdg7ybFZqSV83pSDWl1Pp99LmKKSo5y8O
awNEwp4gC00CPpznid/mDlwb7VjOrJlyspNzTsTuAvO3vMUZ4HRMXMu7RXXve6WniK+4Kv8uRk3k
JxDh3FpkbFN4xAZ+SNB6HOJUVuLG56nSQye27LFCTlg7NgDRgpV4x5kbKV4eh6+Vl1IPyHu6ufiU
7ZiB8NK4W+UVmpqmjcB0vmL2lS5QXqA1ciK0FMXMFpQIgkOE7rfONWu/3gRfywyL9mJZGvuCoV9x
4KwoZFHBdXPz8chJIhIH1NkbLqAsx9Dy2cQpQoEQAu9ON8CVI3j0KdhsEjcheSoaZy6XDqTX+Rig
Np2wLRPcfVJ6xVpgc6qhxDONawKVvxNpkYtKFRdp1XuwNtzy3ou297Z0lAQs+kJAY0PkGj/WEJTL
bnEyt3ItzPDsTNRwl+BY+j4ZXp28vF+VLsLZ2TBqmf1PrsuAgv7/VH4i0sji3yXmXVTotJBN/W8l
e5tM6hrw8kQZHFb8nqRR+MlmcqJc/EyGJfFh+fimTjGmQj52UabCPJc2ZV7FwGRlEyv6HHa1shoJ
5pMdHVceV6Xfw8rJmL0pYzyDO5m/jujzeenfTWH31pFfFe55qaB3Do7vmA7kqcPJYSQ2pYrMPhwT
ZWqWkQHqtzVL6L+9cIRTImOqDd37BIlOsaAHJaW+gNiz2L4OK2vfK4dckCKrQ4m69ftfd/KsEiKV
BAmU+qQHkirryg7JC1s+hLzGLjCPkA7qgBAbocB51YwXmtZ6p6c0hTUjY9IP7wHA/GZ8Xl0cpc0/
IWNKsOyvFICyrutmCaxthv71Xie8udbJcbBdIWYCnd8LbaV5kYLtrVFU5msPbTjJJ5VPYhsNFpo7
wLKsWDtxzzHYcrP+qjBMNdHOSKgDeDJieazDYIfql07/OVwWwbMgaDx6PJvkB3Qgs+0DAsMyhw/R
Lmx5O/ccJi/kt9XhvXtFi/JIN2anc/tgi2XsQCC4LsoU6lsLpN/aBUPo33kBFmzDfOsvEViRwnH2
Tpek0WXkM0aIxoRVTK54KNtxDFJfQFwfX+4YoKhQe5/bCmxK4OZSCRGw6b2tHlVTS2e+GsR5Ovw1
5jJ17oUtNwnlR0FK1odCfDNJxvYJNIKcl+Vd0kEpZxhIbpNAvRqiqdEvj3vo+N4vegDnSJrb74so
ttRojEn2yAUjQgLoceWLwLNqufJedqzmG5hoMtL61U1pvK9n0yxBPV2TLcIHwKZ8+XJoEwE49LDh
FHNHxP0ard8yqC7RgEeJMYTvBcCdEU1mQBUn212t0pIv5gjkvVNUGm5Xuf6OqpAZH1BAaYtuMZyk
VM1tpE0iwmrCZU5NpzppwIC3aFyColUdtDIHjXUxe5Ad77Ff4GWMc/2xHL1nOGTt1h1jPQKAv/cH
IqlroRvYOlJFjP8qG3XGHOAj5qAFDflHgesMuZ6rNZNjhqAZegFJdrNFgsJ/hSexzmOwswkFx8Sa
+BHUXbCfIcn4Z1WUQ9uGDjfXKOKqy6T/fBi4IswkGf0QGLpVHpM9LKo8nHXQRiZ0Wr3dzBouvILM
lkmnwRo7iGjwz58UNJuNdZYTCdsV07HxizehPoqn6Futso2cfmCHWjK51lnyS8gaYaEjhLHTejxJ
gBtmZWbmePEEFLpvBA2ezjw5xxw/2BXiR2USqs3gciEkDzJGP0WTfqkzFD0F3vsE1/rdeaJDCts1
sjp5O5eBYg/RP5r6hwOpLkdTegyihSPj7+aPzWPlhwWyOtHOZlU/ZwLbPNucrKUjMSsDdJk9PoiD
b+AwcV8qYC+uTnpcB4cCxjpVKyoLtn72evlV9H6kB5i57WCJvZ/xT83OBdnKMjTG8PUxm7iHo5AE
aOvh41nLfM+Wk9qHispgymun2brqzs339dA64HBRa9Ubl5DH3mSNSnZRiwHf58JSPeAqj9cGDMpZ
voO3wMcvXsr+R3G0kZ76yRxPqM/PhRM3NMsSE0CyGUjuNRPmUeB4HzAumG/5iaP3vqdzGk0a8mv0
SXeYPWhhnIeLBotj1nJZLQhvgU8dwdAldhnA0FlCwZjX91Jf5NkfK7T5wxlbKZz/7nq4TkpaA6ft
pSvmm4whtwveLJ1P0OOcDHx9A24w06P5lDiH7S38paPWBfBcBSINBD7dGngclTK2XPag+0dqN8Rn
k+HfJsNci4pgkytHvcg71poWS7a0Ih41a4AhXYaiYAHFc7+FW1hlmhSrl7NSKj6F9F7f7qIW0Gar
xUQgxNi35EfXpG55jap/S5+GCHS8xHlWGcNXBWZMXz4RtEv+p163Gl56Puza8Q23xM3oc4mHz3+5
GzIJE6/2OFLOvlcZccMZNsrnr6eW7/XYOrN8ql2WbUGOaA1skQsw2QNnDo3+GH4urbzU4/x/Ok9Y
X/kfD3PSZaAzE5vscGhRDyqwJTLVyxNFwvXOxyGvPz+RnsXhTzDp1FBRiCznC2cKbKmsT9H+ikrz
mmIvhm+Rq86RVnDEbX/Ie/XfFSMBPcaWLFfajwByJGzBo+uScloBv7vWUY5mhf/SULqbc62cHB56
jfgRh04U2te9NnhfxH9QxPCfz4Qem2AoMPdZN/zNv8mSMKeoS5gqMFnLzom9Xh1y0dnPL5yuMVQ4
t82AYkQJzzdU9tm0rElczl3aBo7FXKhmj919YKnXsJzfxkTLDREG14cNrDpnJEbVmAZ7CCVbREyb
g8o4625S1apSZGXZ22TwZXlPS1rvd1Ww0wyKWAY++XX6EmZQ3RySBq/0t8rbRnr9uxC7EO1DapBA
ZvYeJR0fNBk2LMXQeDFCjRrVGcgTRXOAS7VMKRQz0mg3YgWzkqGF72YmsLQfRVtmHc6AeLQKKGBs
pl3O7IOGMFXNgOPqx2GZ0utL7vngisSVQTJ0UU5576d0HXfhkmi5XrxYFLj9yYe/7EGgm7ohGr3P
ddDtKXcuWyEkPgw2MOw6vgKRXvUoNAfS8Iyzbnu45TugWVI6DrVoTeJV0FR2coqOJsaEBs7kv6yR
XvV+n00Q+svSn435HflRXMv2mCQ04WbHE8wUbk6oUNjqbgCkb1oTKFzhg1A7KZgTWpSBDZByG5l8
5CkfhBs1O+tokHHX9lVYaL8o2FST3O0x28Kk2dppTpaXoGIqUiXAGon/i3ftY2UOFfzqkAOObawb
/LRIUv8r6dAzagCTXy/PbsdFxsyiRv3NZKXhxJ5qEORiS8/LD+agFQVsP5GRKILTYRnB90t/Sa3A
Yst0HdsmNBfi61u0xb7YK9TJrFJhSBGBQ+DXXZcwByAfF6vq5YyIBVUxVXYOogBT1HpPQ1vgRfoG
x9POmHniBStTdPXCq/EYXztIN+ir8vp8jkFp3CVvw2ijvw72UZniw3aSGRlqQ5N9EK2z4fIm3ycO
G+XBHSI65MTlek4/0eJ1jmoAx/MJw52g4nm+r81jbp1gSUrhcYeLrz0YhAHDwVYWd8JBOxWP/5Jd
hBPpPqlyh39w4LFqm5kxeLHkyjw6ONlJ2M0+wyxkGkfKtawoTtygR7SUW+5MYoL+rV/8jf4omO5z
vQGpvV0brImXIlnyVXEHyekA9Char99gd+6hsuGQ13x8Ir42glsX5KOkoiFcxwakIeWXfamSZgLG
93o+1RY8zfOm5c4/x5daCvNe4TuU2uyr09L65kjOP2hWjBhK+4i75vArhENMJq50TL/nMt/ocRTx
HPPfZY5m9lt+EnQn7Txtos+bWWH7ZNJ3iudjB3hCB/dbK90+GlYaQbSHgMsMle5miknXoSR0nJyu
EHkwf0qC08iUAlAZoqOpm1FDdI+gAstM5PT/SYxTOzmhMpTXe3ADuGi/m/V8OGyp9qBOW6o3tdpb
UjcB2ZM4O8iZQX+hxZdUbWJkZ0d8YjkNEvApFqAolna6Xt8CrUCT11fkn1rtWf65ROAjqHrSTUJH
FpdnhffdjkBj+Lx2jO6mfD/GfiBha0HAcpeeSLKL3N1A+jKu327Waxrh/942SabjijgvZp/wYf0c
SjKcvatDyKMN2p4SK1OmK7UShVaDx0D8+DkX1gvDLWs8q2CCLQ5kGZ0cOJC0Ks7a63+He52F+Nwb
u9TuytUixS23EhXv36YWm8LAJSVrSEIvktvbVHD8uBEOYQ+OJFjBrab/1Bgtv9dJ8UqnxH+i3Az4
D0GDIQ/ZvBrwtLQrTByatRYMWR6/2+Ey2wyO3RWKd9gucLXxliLm5wV7yXiwU2gd+XBRjWn+RNFu
sFUf6w65u0nZdYQobJsHHdl28468/lHsw0cnSsBTZTUlljdOFQ2Ww/zMmUtwL8PpVorNJiKWU6ZA
qXu6t2XUqUCebEwedaLN+OvEx08nM/N/E8oO30NmY7NmxxrC4lst8fN16HvHBloDU/jbn7KzzAIi
J+cQJ8GD9Khh22gvHLYk2jQRh4ALoFftryba75Z/8MLbtttgy5l1HjzsO/tbtXiBuUKHb+bBtNjo
KFtNRk/mAFglN2+UDkmOmIaL1IdF7LSY1bdaQ9vRNv6uBzDxubbpa1gUOHGq8w1H3viGqPrd3E8/
hJ3A89gxFOqemmbBymjFYDpowqppWNsOV0hdk5G9wHLAKBUqvx05fUQK489Qqpd2KwKfNi3XZTgy
mjXrWxVjjVFEXhrUbbQWjI7xN48p0mrwDt3LSGeYCgqJ8pzzOduWPZ3dg9XooyVBtXcMv7AEnD77
aE+MOt8YaRZClOMdD7U/s0A82ZVnGCqu5rHYMoOdfK9xY4tYosHcTrX7pz9CmhlFWSHMVhaZSsHh
OgkG1u0VCo60xONdZCKiZIkYAuTVU09jeXw12IpKhqoIEGozYR8z0FmcOOpHQADII60UmtIxDCV1
DVYSpeqiuYa6HNcYE6ek86SKCcc7KmWRMMtuv7P7+0trI6Nuy70H8LecJ7+w6Xxp+FX4asrkh1lh
85iZwJPCBkPzTy2WQnwaNSgf7O4Bhh4Mhr1T3QhOK3ejyimmVdkJuWZ4lMVgiaYTJYYR692uKMFo
h/SRDoqdoL84twVg4CRoBAb0/Fyl8do9KBIsjjyhsDAUWVpN7JF0bN7vH+9IvZlt201j3wr3K2mB
tTuaKptlRqfrx16eOytexUnI/P0lPMG/7WEqI0u+ik05GY93H+3uii0TCXIRlEhot/GuDgMxYfN0
Ci7OZ8pHNDSphuWxewD5gNFiRCNYx3X4fyUvX3rPO5AgG/Md0qE9vZN0gMOHqlD8J0ROwKAVrgvB
nqC9LpNQ3H/W595Oi3BuinZu39EX0fmV7r7jXCQ8o00nT0PVDyGBIfwNhT+9TEou9Uz8SSnzlRBa
JK1kutF5swO/z/6o1LhfUhQSUvaLF+UyfDXZzoFIKFx+K+5XKrRFBAXJsFM1rJgp7mTDY0hQw8mM
6WWsDCZabyQwmzrRTbKl1txjxie1Nf0491la1hKNtvKLWGFJJetqKLmqrv2oBu7sUGYtPCWnvt4H
Wk8K9mZ4F7Y0KJ5Ze/Z0G6uvbO869djF5C0Zwb5CvisJ/NRsB52mi/2WKZOqT+mKwiJLH5hIn8o1
otfF0pzMX8ZtTGVkU95ALldU0lGsyLNlJcnICMERPEmLirt40J3y5X2tzeTlJmE46mOhK7vL9NG0
ZNd7pN704sx5x4cdl1SniX+RiiAZQO7g7aue6kaYgwIZ2oWP6c7qIS34mwo0jEfia2ayTWfzl7ml
Al3bv59Fla16Np4GVAxA3Zq/jnXOXe0v5PTeGJL5F03DcqFOGISbP8yjp9vf1JXBGOHUBLY/aCdy
CFOLj8v9CYA+kwlmDVldi8uJtSrRLXBdzG6yDh/+FNnkD4ekwB3Q/GI3WsVhv9t72PqF7q3L2v4t
UkxiOvNXNJuZ+/Se42SGnWaX/Y5Jn6EbGD1m41+M3sfHvvZI0ehv++Ykye7ooUpMfQErBtVb7KbP
xQnlO43+dvk67h6PoYLGeV1M2BuzimIV2mt0khd1WRh9GN1Ooa4DASSG3mNnGuNPhNR4cAdLso6W
R67KOm7fadOhsX45nD9y35e6hxSgmE0DUmk/7/WWJmkdZ9QdoVLr24DnYFs3dlsFpAJzyRF9BIFe
91P6ANMIsmdXCZuEfVe49/V3BjgLaqGQI9FViRs+4/um0GNnP9qQyfztYB0WXOqLcYAfBCx3Aiqt
CZRisJoB8GhZmh/Q3wt4GocPsb3BVsELU4L+rLKjtnt+eDPSmuWpRe2KM3KeSU0qaSYj8HYoJrEM
4TtAzvj2jdO2KQnB+8f5PcR9I8PwSZfkoB0vwheG8mknSSbjOzmf3B/57gQ6ro7Di0ipQ+kf8j81
BPw56VU/qCCh2wL/xzdYwc25tTUvFxrmFd2I0BMd+crmomNWc2OfFgmFh7ghmx82VDzls9Sdzl2I
N8/roH1K+LvNpsIWD7Uo89LFKSyHh1lon+kNI81pjjclYSuu4+a4DtZV+G1WfNfn8BGr1/0U4l4p
P/Gm1D0A+44hE5OGrwzPL2D53Nat2vzlETeSYIfQnhQiy8U3Y66fQTqGCtP+i+13A1rNHqECxTC9
rz9shZh8D8evks3ic7uHvYtLDbsjz+UShFy3SaWVJ2CQnFnoz252XCUXuBepdlJvBHl00XsjTGr7
EsRJCfWY8BZ7YTOOPQxEI0Ugf+FafMlmAPW8+Fm+AeT9AKWr6MzZ5emvtP++FWtqVbaXdKYnzrUo
7ldMruNVTi91vgMgW9+2nbcGhBEZ9Zi5mF4IbefKGFUo1HrvLIKUhQKeGkmzoeVI5piRZl3kQ7/r
AmKhN3yvZsM9Lhf0pOqyuPcJhCJtkeTXlUcG1R632v+YdVjz9Y8e8kDNtD8P+9uAkO27MkgHzrBB
bJdudTPU5cwCyFtD72CEqquGJHdfpq+Kzvy25SYKh2mcwOoeb8PhsdpozbY9b2YVXxtAPbBG9E/s
B5/GEBrBquX2zPnPwlleRPm/cgdxFXM02v+wry9EObrZnLtgyMx472P10drVDm0nQEP0/gHqok7W
MlJ+lUNcNVw/dPfthO3eMTk/GNPVvYH3fYpYSuTGeYpvfeC02r/ms6vsBr1LZPyMbyH/KJNJ+Sxu
Mu3L5Y6YIm+l6fZJ79KMG7cDZQ8mipokEBTPI9WE/b8ZKIF2qjAClphe8xCGnSt6jAloFsseBKQk
8WNNdlfTwL/7kmVkZmOSg3+jKbM51B1+mPCxPgqE7ggH1HKIdCKdUP6pyU3G3FRXOVxN8UN+Det4
4XRUsZze0AYVh09jw68t2Wneef7t1QdhBpeSn3Dg4GTQlXSYb4bDSk4oQd7jZ8jAPvOilQFj5uyP
kFKsffvERSF8h4N6Os/cw/PCODkPnOJfs1xx2SXdBtk5NZqv2lgrAziWsmeaHFmVKG5hlwmAwjtz
JTq6K45CYDDc7Xy5y6FnzFF7qavcyesvrmEZAkkiV2nF+CY0zPml3j4kuwA4dzrPl+awxdR0l+k+
kXA1jcv01IZTa7Vqx217JRjswUXSgAQ7oGSC+lgw6JfpUjYcCj4wVdwOcpL9hnEO+gRRgSrS1SwW
GXE6LoKx8+DBEAU49nYr0ReoTMQbWwX78Bi7DrDYU6dFyiQdGWpWpUMN2H8TJBykKcwlLLAL7BNT
bAMRKxsucDYzAcv8NCM0/G85B7XSViPunjHEXJMqWkbi9tSpIWkiqPUmmuWdEpJvtkVzg/08lpWx
eUL6+bVl6pqfz8jAJVrZu0blRkudLa5Qxo8RdouKiAQMq7oMXzqd1FuzqJ+SIAYMR37EXC61EHBF
XwFu6NZccox1qSLn3ip57hGV+I0+f4JcNQm6qSbj3hmUIhtK6Gc7Mgzurr6HmqLgOK5mQoZMnMX/
ba7Xl15s1QjgLhp5320tChRMqjdSKF69x7SQF06cR7Au9w+PFfxMc+wrHERk+2NBp+Me6Q6rSJ6h
gxz7S+iiJiQxKQF189p0Ud1Y79rt+4fesiZd0xX6DJZQw9DE4z3nOsWKsLAWYK5xdaX+c+IRJTZ5
GMO/ZAZbnx3N3FFCFgTab0BLy6aadt5ClZyaRfl9ve9JelDUOS+0XJIfXq41YxuaMkbwuNxNaoOV
4CmdAl+8Jv3cuMBrKbyO15NMuaSa9RTYqcTmFhacMN2evKUEhNkC4dfebeFXD6VHnsVH3y5u0sHd
ovKd2ODH8Pl2I0wnKfYPumleMKhSbFHcfyNnESUhEOvJ935gWqVjaeqlLgIWyuG2XeYPEi3Nldc2
pP5Zw2Bk1D9iTujD2HIoKBhxV1AhxePqDSvUADyf8XJsM9h8rds/3ufFU4vFk0IDW1gxm0H9/6ZF
rFwggBZTnG15jGARxjXc29taz9GE043TJrb8ifewMhIe3Pbhd3vdTPsZz3A9P0wgdjygLMbMt1e/
VQQ/G8UWwnD7QmwlpNIWW+m+tpvAquFHRQraCLUgqw54JITzouC0C5YJ5WQvngGiHo9DooMrhPq/
2ZM4v1e0p6LYaK1NN7Z6P2fEAsTgRCJjkmUobUxmWtnAM4WtyF+4lI9LI2zHTE/Dl5TiKxVFuLl4
oMcDPVazmSgdleL4q9TwdECfc8qXqAB2D9poEl25JobgD3P7aa6tzOtDslXIy8bEGnZhb8msTpvX
9r7grQ5OsdvMz1rQGQjRrH678RgXsndrLy0SzD6qTFqrsIgt+ULYz/WeZo/sSy8uITZnOzgVobB6
fUIeM0NlIV4c10ZV3LAHsoqj25jNrlYRK79F+nkG6Km3WLULWT1pBXd6cZGFEJ5MOSBSUhEzwH/d
8168VtCfosFIfvfF6jCQDCc6Uh5q8qIfjh2XGrlleFZwUdfuTnCVWhsBe7lBq+F+GFIl98hK0hiF
+1CHdZbMc2nQk63u6c3KkFIs5mrDMSt9UDzSa4nCv+nE/wZB8E3JZm1/UbDXmK1FA/r/9ZAI7U5q
d/tLv0sBjoyiWb5I3rZf25lgf9VVir0j7Q74jFPfE3rQo69WYl/rNNQ7KzD6YCRzDNUy2r+jrnIh
McBhXHmx7trba3V13chE30fbwOPENF7+d9G0F03HuG4ZuIhMxEI77wi4moBVxQFHer9RYu6tfrOy
dMKLg5oUOL4ta2e50NxskhBr96hxnDP6rZLhPVTLdI+6Iv8g1ANYTXlhkUxceQOyzsVWWT6vXibq
BNe5Q+bNba9zutHd7fCG1+/wzwEkr4LufoH+cglmaeR86eWQ+EdPRlXFwsLctBWLeyGoACK10z+X
UycU4lLLKDMd3+48q45jh/TajvLcl2HL7s3WHC7538L/VGUN1S3+g81rQ91xsNbNKXBoVzcZaTrc
pxApQId5r2IXncMEtkw9c9ER8o+KLgbd00nOWTJT5e32ZSMn6p+z7Nvh60rL0e/lA0oD8Fqn5Rd6
Zs6PzhNmPozdsuko+Z0E+UkOlkR6AvCf9dzQsNN9iCy52CjHwhPfrrslYSO7/T9xAOqQeQfGfrRx
aVdc0HOihxtU1gvhPXnasj2sjDow074wtpztWs0lHX/gL/j1fvHgzSN0v7j3aRUAHAQ+3wxunRKm
BGCk7g/juDHIDHR8RtXriR9+LFHlE6K4/PtoNcI3CnD2gKHPL8CaKJoLpzwBmFmCrgUndt11FhoG
tYALyYaTjR/L0G37TMV+LrRnstA3HgU+on6IhaVFMAE2mXi6XSL8I7pCXtLoBJz4gDrReukddyPj
3mare9lRdSX6EI2dcMaNbhzIbwyso5g5zLkhYeY+aFWDiX+wcClOY8WOu8LgdClbH8X+rQTJIcEY
HDdJ3SmYjaq7rDmA6ySHhzLW+0wCZfXCfXB3enCCJ7BEk5WoNz3F7L/86NuFqChVzMrVgZDSl51b
ABiPjEiQ1919mnhNSxvtWrySvwPZFnmVWfPXKh6gn7ElUYaTP4y3GpFQfp1KUc9Wkl1gvk5oE/Jl
gRJg1QGUdaDeNhAGfD4S18wzhDQjKjqNUchymYPJtnb5cbDKmFKR1qBoe+2/3PHgsp6kxxWLgwSk
E5ZiRn9Vj2LS3NP0npPPNmO2zNjQ9XYIQjk73dfzpS6pFxPxKVn5xxUXC2GRrgwAH7gdCNORyVNp
SXDcGgBvCorIMEWa8lh3lqJgxgEo7uRlck74h65zRdaCsqjJsCq/SI34a5X164gdusQoer6/IJ6P
VHfToRRLqyXkm2CCKrCYkjHxYeRXyXsLjZPdZFkadaoT7yq4jOIa/PDdjOSBY3SxrCWAkRpwoBOM
MHeGX9VTltcV6FGyXKL4/kk6mJ85rSg7nnOMyTKE5PU9trKSw0/aUV8aj0A40cxQgiN8SQvkZa/N
uR10KZz7DiT26n03TCoPXxbDYSqsBwy8EG/a4gx6VutFCSY/gDyJBmzPiWGnTNlcZA3sJ04T0hFb
H1W7Wsia9wQJ3MpEBKRV8/0WSxSdAsdlGw1QDUW/wm7Y4dSn93KRZelfFufVcHiJcrKxhfGbCfFp
S1lmenXPTLg89I8kzLn9kE9s/chOT9lKZQ25AnjvS/fnwPfuulOzjDb+NUU47iCjw+yyb4AIJ3MI
vMwdVHWiUK0tE/zkhk6UKFbch7IMK4eoYiuNYatEaK+H1zKdmTU0AMcYq4cfTSmTWrIrAOpCt0Qo
f6PXxp66Q2N3nT9UVcSgQ1pSD0RWhRBvgCZG9aZhbYnWq2+C177/LoDsdBRS00wMRMamBG8Gpzgp
7TecCpeH+WeM5n+JX6zqto0Wa+Wi1zSCxw2bB00XHQk7EHqRwoEBcFoeFmVtf7eCEmjsk0J91XLH
hOBj4yWJfxEfOofJcWJuWKLQFM1z9pID7OW//B9bg29O3Pe8ul5hgeP8lbDy+T6kOO7X8vOWRteg
87H1FJcSHeIryhjWrr4nKWTO7Jpx43kPrS7HWsc7DeFjYZkh10HFuo7QJB1OrDMgJmhVSUkM6NXO
oQInyoXjK5vBWXfE2ynfiksxhKjxEryvos4awj5mqyeDFcGVAvnYdu/91T3shpE4xDbr/n2zYf71
9q5WDm4u4sUFkVhPD5pRqM+9MMV4J8NMXnTPoAX1CVK8Ak3AJTtG3LCFAbKseAz8BP4fUI5wF13y
d9ztl+P/iO9m884EjnehVjlemHl2UclNO1Zv5uMPD3kDZQ7qsi7z1ispQVBD1zodZFFmmj+je2/g
+r456VYAJa4l4weMUxeRIjOb+GxGwmnxKV2eTyOJ5lvAKHJeQik7kOyoH5zO4cgoGrVeTyHks31A
81lJQQQW3SvpB8x/6engMFNMrMovTvYbDzbIlfp9axjDQU1pWGlaJZveTqLL5CYYK9QHd1xLCR2x
YAZ9Gy+TsTssd0w2f8wFglPbcAiHNCdwpQK4DaV/KN9Xaz1UU6a3BcMterhmFggZlGRrVxlJjRc6
AOlU+tJgngUoR0JyHzVNvvm+6Etm1M258FxZC80ajn3Kkw0mNV8EJq2hp9TLHpFF32vGYO4+Pv8V
Yghs4/9a6ONaM8AZGpvtNYzx537lNYxvMNa4uicGsqlpSe9gU/gdDe6SMYHAr6mAd0r0vR3Y9jvZ
GDf8QMA7PwAAvdMZ5vLKf1I8vdY9F1VXJRHdl7FG4ec6QL/PlNFXV2Sd2CUWMIdYJ5MrgB1pdlDZ
Ll0+iTy3OA1FFWge+rp7mdhUk1CnUcb7st+JtKKGPhHx7vIIO0xNWaVTBhRcA1srXlGja/PPWN2K
8CCgiQUVBC6kdrcJ7ELw1FkILWjZmfiBia8Pu3AxPwlbjnIrLeMwoPx6KsM3Ew2v3iwW4nHrM4dJ
95UCtuXIgOiqamBlANZcm4/9Y5mS9gGdaCg19I9EfaNjVi9vdUEv/0FoIMUC1Y/Xme7i92Muwo1l
qPt7Pi3I2j8HJJgh+c9Pg5S7TIsvR4cJVErK8CJqudWFbalCqDtsvAW/4hIN4m43YLROSBlYytDA
ehInLy7+XPIUK5EdsWT2Mgmz7KjEAraKH1Bffrfs0gfwl27d6QPnQBnZVSRPCl/jRkzVFSYaS46s
nkuaki+ltcc7YGt98ev//IlDd9czQK+FqjGKr/cIxfZ+mCdu17b0dVnzzULNCaFZOnv/AE4peljg
h5LbSIGzqoIn8pi/ra0ozHcuW6WhwBMIfhNW/5fuSISqgrWaabUEioCBO7TFONDqX9mUAoyuduzW
KhbXl7+ycdKO2TfDJrCOHZGFqiDzG6lvdCUUSycOZRouIMDjyqCb2EBLHwJgXoIlXdP4HHUMRjW4
hJGaUhRpVsK6405WnJbROtW5fNbsTJ87heMe/Xf/oSBISUU5aDjumAmqONmIX0YdAWtZzusdTS2W
eIdTHOfUKMzf+UBD9H6BYAVAlBhKHzMkhkKnVEgJf6XWg6FviYWalEhklp8Lr6yBY0oYY/9cAcjJ
Rsln8U5KooFrj646H8GhMENC/P329An8ExWYTNJwtZsnT0mA9fMYLFR0EAEYpc22rAVMcz4esVQ1
Tff5fMFe6dGyMvhu5i49y5b9vk2RVeFSvUmOmzd8C97ZSgOjbxHkY7q0PIehd1AtxTq2wkD8kq2u
8Qo7eqWfTYqdCJdplD2VUAhffAMrOFoTu0MUApfnTGvbjET7d1lLbt4K4OSxaVq1Na87SUgwKL4R
Lgb4zcLu424OHuNq8oxK7bOrZyvw65GuazWkOJbx7Q3BulEZn/MSgvJhQPyL6gbIqcPr+h/8qFzk
J4yJMlgX5zlF3lsD+6uik0Bn2e7SJr337GbkY84vkgFpuuLAiSkUEeS+THbqQLgaFPZUEOM4LrMm
HkLF8xqEm0G3moyjAhEZbgRsmNk+919qfum7yf7TnQvh3P24L8HkzJ3LNWaxHECN0mO6kp4ZiUzX
GWw/GiZSGKpj4Qyk0ZFPqJfgpm5rN5YMPb93Ncn0nJYY5A8p1YsYdPB2zU9YUO1cfpReEWuNX56f
t8g7W6HQtOtK6raBsiIKo9Oz5jEUEynnYUzoYVLvYPUoFnnxtzGfRPLyVN9anEuFZjM5ivi4FOAl
DFunEbwWaP47vcRrkKaOVj4uTeSYjXyge858AlynewObI4VoiLHD+bwUdSX54HAuGxjjHnfb37qP
gfLQuHryeelTA789k9TINMAZRr4bT04kEZqIxYQKiZ0UGUNAIU+B+HXUXbi7xvGHnqGZ8J23zdio
lPDCWn9fuqkhidYB9L8IZgqxprPXQuwLPTKWoJBHuPYuMBJFC7eNaSmLV4A4KvsDt01wwhg1rI3l
O2Wx15jiyb7KmolnAb1o8dsY4VqT2GJbUcWSKcAJKE11uXnP0AIYgOktjwhfSULRmnHlj6ymQYGk
wyh1c8FcS5acTg2joQ7ayOyaTIq+n5aP6ZWWJ58F9Rpzi14477iwswyE2n0PMPQXQAjRoXwtGJVs
RICbQnfW84nILRyrtql9imV+xmT21sWukwXlHxdYaSiYICb/2qNx4x/okW6ragTcfnfqLcK7phP0
XA2Qi94QLli1Vs0GsZDTqMfsNbjOttedtE8ku/xCO8UIJq2jTTWB5WyIZXAjnWADjifDboMxaANu
e/9K9i7l5gKG4kH0ATZ8APT9fyfuXGcKlu4YrRrWYpvFWZYkF4aka+AkzdzO63lK7SrawrRil/q5
r+KgCT/CrwrjuVE1UTxmFsjYLmqpye/8bEQty9nV11s8vVAFV3uPxAjA/7AxWbulv2MmrQJwcQ5n
7tp08uJTAW+NXFsKpVEW1TuKbmM8sbmUEjJlz8VGCGH365++bkQ7ctYnciR5x3r4zFb+lXgmn3+E
jLG5A8Fg5cu+hg5qsoUwCjZlpvf1QX+o2PpobDaiTw3TuqaFtlPx8vG8Yac5w02IBXzSiAcaNuZ0
2w6Sonm+1w856Yv/+WU9R5SahJXm8DAsC0MOlRs91/BptJBSqhv+gwVjDNtYXTGmRsYrHBcDnQ9O
HS3LfEG4X6SOx5BkBv7HYr3ZRn1FnilnNP1C0eEqJtvb5zsguZEf6puJIOswjdYKmjb+k8c+wtZ+
EnwZVMjd6mIv9aug5XtFa6OtuTvDBFGEfGuIg0BOfN0UwJq+QyzTNZeZBGDBuWfEg6pOrJBFGNyv
JKchl/fqrTsltkMaGVFTpeHUz1gB2sQLJ93lwfLDGOkTJ0pJkkOJrH9fw13ClOimx5EL6SevdPDH
dW6bpQU83IypbepfzB0/Il6BHgBJQdrjxgitF8hlgkfVWWUdNVkwrd/LusVIiwfaZKCQRY7ZhK9l
oxn04DjJvIQ5CifaEkMsumYCgxQNcLqQaBAu2IpXlHJvQBz77cmyL3vEfsa/rtPwzlNyUiLLV3sv
hlV8Qe4vguUcuguqg7bFdRXKpJ0cRAG+SIRQyPvtuukguiQfD61nBmS16iCaypPJRLlldRTqKjEe
QzcJCaBU0ni9eu4A0/rzQPHMgzKVPZ/iGVUt0L8Frwn7+0yHaI3pO3Bc4Tq1kod5/RvFl7Wx4nxy
8tx8fuyW12MqM5jIECMZn9CieyJ8GXDI8xVViNv8RAVh/Yrfjn7gntwb9E5Czd8hJM7xwTtXrPNq
8BJIdHCXZmv+u3+QuAqz76Q7eh2jtKcewgGT5JIUnNrw5hd2btPgDZJVoOc38EeU2tx3uYduNYTz
esvn8DMchmRMIA9IeKbA8XD/hTuSMXS+qnX34l2SV41DzT4VMT/b20dAymDYAcJ+4+aWus/nsVQY
2r9DRgiclw/4F6Lj/idI/EsdN9DmarZBYahUbFRzDpe+pIt2wgg15/oNIP54OT3xKIbeI9CYJ7NS
ZIVa2n21nHiQuXf84HYBgKAb9D5Woes4+BgSL30TSe4rJHOxSL+D6NkMXgMdb5P5VVsbNdyX5OmN
NOSIAprcCyVnikP2TPoYORaxBizwzWkmPTZX323tWQVQk/aMGYjT4jWfK7hc7H0yQ07FNlf9Uddg
KdjjW3kJoUs9OiOKfkdJStrUApBfi6WUXYyICC0HR2AiKKCMh7WJo3q3h38wKgJvxoFJVRk+/8fk
MUvUOZR8aFQCxM/tHNRd6RvHIVV8OQ2TXDxhRyZPnrZZP+QMipuEcvHAksujMCEMdLxu8/NX3Xwx
bfsvXWQm1ZZFo/TEL6x3Y531IzYpOKLfvP6sTXwOzqtTq+zbxvOdkl+44rUdMhGSGz11rxL1FH6t
3Zds4PYyFqlafSaRXr5xa65QfGETqKdWfGYMwIcv12Q320W4R1LG5vgjcJ5fFTExOC68pkTswVnW
mxykmO98KWuoYZLXvv/VqBaoFkUC7rBGLAbO+o+mPd0hz6JL2frTwfhwPMeDdAc1sBrOhs4j+Q/a
yIbG/JrMuWYLJ7e2vCoUgfjvQ37nmQo8aO3NLmFYMsevGHZOAshYZjdeO3bPTKA/dgIFtuMoQPpd
bPG1zG90OJZCaY1KC1FqkG0k/RTlEFJQO64MvQvNZvnXvsmxZwiBnktF9l0u57K0NE78282BKG3c
/MISxPPLPdNJqlK70ozY5ovbxuMUJewF1uyEybNBHW9IKDJwzDh81ZsBlvfr6Gip5uLWX4dlz/Q4
v+OOPtsxjuyzvOy77cF/4S4ILQ3nLovzhLuhKnpHX3nifMQQdOOxgJJLFw//GJNztV8bdqsynbD7
jGkWevUrvi4oj9FAmTyfb6rwf8k3qRwCTzIA5ACBFCxdYjylgw8VpTapVhYNA1ucQZvKgm1MUNHU
vHUuTTMr/HuGHPsaMhUtPcDvxrCFgt9Td2mJIDwEr6uZ1IVUB+4QDCFFfj/y/ZMprV9kzfUbHeMJ
J/EdqxYMJvg8LEO6uES4JLE0ebY6V7RSsWJ0LZVdfK/nS9KQGsoUnxj6c6FTNpATTXawSs/YuWbq
OsrtCEBC/Tgjci1ymdt3tRacsKA1omQi8Jf0HCQKW/RQNWH5RFV+A/J3DXF05HVcEO4DgsOd7Xr8
CebCZbXxPNPLzyvEDwLsVU+pIQZR9S29f47nzF91ShkJ1srjB43O83tVTsWFYeV9c32G5NKDq2CG
05SNAUlKeqIj1ZcPQaHRp0mXWuGaLovIsTsCCYFXNT4LCJfxsUvRqXJfxriUs739ls0LB5HtxVxs
vraiY0jgFvzWDRiCpH1FNALjEDHwbuYdyVOAp+FU00SE1aHWyyY5AlevQsZHV57xZrjsMvojLqV4
1TU9QUs2VaLMQJyZpWwIh7GgZR1AGqUf0T1bJ7dDkc1uljQoQikCBwLh3Putf7QN7tHKJlFDmlbh
TAfz6C6wWanVgJREpsUDkf+oDrvjZxXuz3cg4fxw5mghqfR0dZZtibVwkE6ayUzRo4xBBr9PowXV
RZAiN6D3yhjsybk59AvfvIvzySOsjuHW6PZiiWUezV4gKhtC8aoM45UtxfmvL19O+GN2gjnB8rVe
hDpaKVvbmuib8hwdRAWtNYmLHZz3NkQPF7TyUxHVX0MbLsvT/GOBaexdPFA4Iz4wjQM7AJ6wTliC
U6u8EOHOvQElaww6DMMqWAn/8CNjnLzESkpn+jw5kDTr/FM9MuVRY57h+CA8Q/iMKI7dsLnfzCwp
D6qaNmUqRk+doUB3t+5j97b2OEdS81ZcUSQndHuLE1yzn/MqkjL+T+7H5UNbaHtj4+2LK9O5BHcX
wUUrp4aEUTow0RJBNqEwxubYrkMGxGp16+E1RRgZ6nDs8FGCTd1htxxu66qQ3LiiCm2+zAatuSgt
7UfrLpKhJ4gpgLZp83dGqr0fzIxka6hRT6mL0rOtYkK0F3ZGNOCX1fsCeSgeUOPQYW3mvcJ6n0QO
3PdMMhysCU+W83WNCX4hjAia1OaYOU+F1vNHoHzjVOG2jC5te/YaNNX6vFJFTUm41S48PSWwArhs
UPUxsp/da9uGUdB5GjdNu73JXx9VL8f9rzzlG6QQPaC+5HJ5UjSjehLb/8qRwstXUORa0kynlfUu
sRhYdmqWRioq8kBJiIvMl3ZSy0vcc1UjIDcudf/pBPoWQaVthJ5F13p57PPchTV61MmE0M/KOZxV
MfSd9BW3vzlsle+ZMVrC2ttIQkTmKeBExdvEw1kVuR09uAvvDqY4s2Cxql3ogOSvYJN8w9Nrqfbs
jVb5LqNM1mnYKjglP5A7nUhTdf+vf/qxyMiODCK9dXxdlowruUqzfMc+1WEmJbwBaUVclXBTguCb
8UGbt6NNf9LFbuQAh2ZlWBdXevZyhmm29ITDd4xqMxSTARnlE/U1QG/gavH/DDWMoo3DC4Io/yEZ
SUOr91JviaKiYbb3e8w2bgxGXy8kObnyiZzxOR7kkE7+z9SO/9EHSbDCHdNlIM6bl3CBq9ptRZ3s
qyz+3CEojaa6XYbgaRFTJbXwgTp13JkHAT8+fwMW6nEW6tdJg/w0/owmaKueFsQlH+NVTiJeKUp2
R7UHLcOVL55gaJIXM8ShcJGou440zWwmbbLft5fP7TbvLgdoRJkE8GWBisZPazFuFTzNXKpNjdjD
MVlMAvxltpfeFfOk5HXNEsPdBf4w1i75pzrPeLPkioZ4SLifodJgqoXpxBeI2jMKd1fnTpzjfO2L
FAz4d0Ni1jq6Q+Bek9dPfqL8Bj54Ph3P2iqLrDS9ofXc2UNXMb4oMJzfg95rn0X3O5tPcpZuwP8Y
dE1rCleWulzehczLFJ9X6RsFMqpPDwVhyUb4fN8Bb55e8u5lkGBvXX1XB+vt9/QxDvFDgIPH8wfU
gLM6ZaSPM9mWOA42s6tSxU2dwPvo4Go8xM+/NAXjPqGe2dotxTJitquadgfghZk5vKGhkyQI9BEK
+vk8bBsvtJpqnS3kgS7DG3bpKuzbaY+wMWhRkuhAvqFq6gjz1LQ5EH3rGV5fWN+kSsbENxQWxoKU
I1oPUAM7utdD8keEbOv/M+AmiaISIFD0GeBXyvThYQ4uJNjXFnUWnSQh86D4xvu+CfJ2JL6qn1+Q
P3HZzDzlM+ka55cr7bwA6tB/UyMV8OZYTL61amGgYQxK5LdoWvM+OZS59hVdGCHitJlce8VOZhUM
7sAhdMBmbABHynZVu5T9zoE/ycZGX47KSwlHzT0m1QxrYm3Z3mFtzxGOTw7/spHGAoyqtsYlnWY0
XlARgsBnPoQZixgHHWbuzQdqCC1J6azMPOQGasRjEwcz5af5kg4t0VZFSq5PUzKcarkLoVRjwepa
z8aKyUg1m4Ph9hZ0pcduF/GrwJozzHCTqtczhC85G1FmoKOuDTnEiZZ9UXz82OgVbfkIPomKZMjj
JdtyLtcWAHnFfLPsCsWMDibsFkeDE4ObeKqbQc18a8RE/tdWuNtN9674L2vGUGCXcJ6ugeWylQiY
YQFZtrhIdxAvMpE0d7xITctGCfsik/WXcuf1gpEXZcxHye4gikeVOt8tyNkX035aK0vFZ2ufmI5f
zuWuMww6dR8iZlPX92EK5itT8gpANtc0+/zR3um86VACLG/sbDp+Pdd3EiVWhU8ZNvPXSR748ceh
ZRHFTsveqmtR5GZ6uqRFpP3A6y90KtA1JLY8q4ii4CdaCbtsxXccZz1vs4I6L9sniCbgAwc5aBg4
a7rvWgqkv3cZOnCsSfSR3TpMXLBe7FA6apR8twalH8p63ei6unY9hU8RCc7r0sDg+aGgNATnYXtg
dH0PGjCI4cLfrOQaL/FcKjNmOV/glEKVR9jvqOY4lKyTE0gKGUAKL2tCR0yzztLroRcIMkUtezPA
3yyKwqT/v3PlYb53VvofCIHcFi1jskF02ja/aibqMgWsCu74GWF2S8sE5wqE97i1YQqcm82aMbei
oYT9v9UZ58LGX7aIumS1On/NH+pb3k0firycOsfmEC/soGhUrCG58ToXhLk/fqbCsEXcOxNjOgcu
v9bIzaiDreCZUnCLjh1oQ3ZaDdwA5E/I+9URawAgU2RdTEOVQBpKJzj6D8RyHIzK1e7oHpDLUcoA
y6G/pkTxUtcNVp1Eyzw9zc9AtVkIOo8Z/jE+vQrEkrz73wJbraX7USKjNF2nS7dlfEM6tDL/5wt5
90Qfy2HXdk+CjSr3pVLv7M5nMvktUcL/V82396pi0xNSdWdqwotOCpCZkLd9LZJ4qIf4vGwGkaek
HG/UyokSjNODrFTbxo45cd4bAi1KE3tmWfArPBH9OmGGuRPuMIqpsV/ebfeRE2t8M1UquMo9ekhI
Yhn5R8vQ/aTputNQ3SWWOkSn2azuzS3iTYpbO4bR1PURCj8McbjNEueZujtfRCzo5ceTNj7SkHk7
85jGXRa41bG9hr/hFUrAoAVsaFB6smHAIZFtTGVeJ0/26V8RjfvvrIzd1ThAxAVSdfckY9dZwlE5
Kh5PkRijl8vxEY08/96CB1zBoptpCM6xpSmYZ08Pht6EATfmHZUIRk+zi6UKICM4/y0bslewDl9a
f7N+nyaMyaipN326VbX/2xmHlUippRz7nPzle4fsm0YZy8HTxU9iyNlt7Hx97jOeheyDBvjGNxUe
rkSFokZIY++t6sXx/C1ekwF+9e7JpyL2KbAiUfE9O4vILjdG2DbKiZcnsB95CACzqHzrkyMqDxGm
S99pQMZ1DGqibojeZYsfIA7xoE5KFAzewBJ00pUYbwGsyIo81txFqnUmwp6oKI3QWcqdAHLsWWmJ
rAuA5ZHV1XKRvAnPLUndWmtAxz6evZvvGyfZ1brZD53kXg/q2qxM8oA0oa/6UYM6m5XR2nvG60zE
5dNosyJQ+IaOK3zrZW8JQnlIjzaCS7IH8Dtjh4opZUVk/k6FSPS7YcCRTxpQ7V0ZdfwQlZeZ1EO5
qOnTd9u3PatVykyu5ttf2PfI9Xv7Z1sH/3EkWjXjg/MQ/Wr9Y5xT7wmLbAmaJ17NIuvC3+PjymeO
mqXYNzCs95CyfMSGGeHJlMaOGf3j7gkVuFv0SPYejR91L9HWFw5lmx1T9Az8WcuSMxL1agZFgmPI
UGAfmlT0/qNqyLOdrNkFmjGF4eQ8JJOr4DotIF7QIly+KBmKY/AuycITGGC4SD65pLTSrglcsh1z
hMZa+U99YMoFsGOKUFvCc3xAZHUXps8zhKWdffbD2JBjSi6guk06djeeTOlzCuGk+DquybdJmA7N
zTXPorxj15irLIqD2SnsAN7EgE4HuKe9H33/sDzrmE4/+VjoaAqKIGYKQYa+WCJUI6PBZ41AkzqV
77YroXVcMGpoVFh0UemCVgAr0/4HZtPGEkKBeSKis63tmlAOX9CIGxtuX3oKUPIAH2oVqTJWQ/1d
kNO9qWKQbOEF14V2NbEH7oYSPKSb08TVITu2hIjfeYXWseyoUBqmbb0/wkELEy8pZStHB3f17zUp
o9RmuY1Aex5ck48+EzDeltM8LS6rcxyNcAgAQA1AT2EsTDCBR5rxTAsok5RkFktOJADwb33sg9T7
IKCof1VgrG+FE/aVIpKf0wkDkLlqdyYJqB8JXI9O/QbHQMk5y0NefO+3JMNA2KjASoeG+FijFkJQ
8xNS4EbspY85dN2lMpGYQ1wr3fKwd83LUIqkLDGBaXkpi/oSF0KFOikdweDLhl8b15EYuF/kvSN4
pQUKf6snBdvywr8AAyhnN1gI/KFTAFoQK7ZgJwb5S0JYNdqNlmANZXPsaDMzHKDs5c7k2yzuo03B
oRx7/7aByyouwtdkcYlBqZgdxAXuIB5V8mQD8KM4/qAeXdUEvIcHc39MToXm9HZ8lEAYDHxpZx9o
jCKXMFKcLY0dUyELlp2ZXCuQtq9ZAb9itZkdMYoCEMui/u2s7SPzLyJMB6w0i7JadRc1WY8Iu8/1
VDmBynbIe7N5i+Gp8QQPs7sMKSu5qAK9+MJ200fSCTY4J+Q7UWGZncV/pU174lUjNe55UWCNzLO+
QEoHe9qfH7fYh/A1t6oV17iShMI59JyeVdktbQTy9VLqPN7dDnR4vdEFleqg7lSVr4EXuilxZ/dl
SddrXWlgTPHGHFVmEQ71S+vi5tZ1SitbNaKpsstedbMEe3DgTGrrvkqIhDBueVO18sShgRsd2Q5b
A3FPpecD7PoHnm7OudcY2qBUGHDj+IAHokzKWpZ8Rw4IlV5UNHguakZ2rmhSVRaxBcSr7P6Z1bnm
sQv2yOs4wohzdyMit3qKfSy4xG+hu1tBCvQkclskRF2BCpsdQFHXadnseT3Y+qeGrYtMzpC+gsse
upf1QbkT+vzphxW1+yvmPr/VqXmyv74mm9b1pOrpQzKiB2g8SKmd6DRWaomS8ekeGh4hogjp6fFh
L17lSmaI/qYj4iZxQbjVUIW2mssiR6ixnsQhV3HGeLdxuS1kjhJ9qLL1Dj88WCBiwQ5zFvi9Kml8
cuIhjJZ90sxjIYEHfmwu+v3TXVsc6iKGh2I1Bq0Ew+2wKXXzgEx4jK0gmN2P2IBp82ngFAcFY3Rx
mOqSB+mMDghzl3rfSBz2VHar1L7IB63S99GCo5JpDWp+dQWi4RdRnFo2Zl+9V2pQseu1OiayPsWU
0ztd7ReZ8C6A4bCbIsaUfrcSUh6xlN70StM/9jZ9WBU4qpNcU95yHph2uZbP3ZtcE8HD/iUUTizy
YeIJgxz9f00bHMWajBAE7DTCEYuQiJx15zQDgz+Na5Ab0IuIEzmBjUm15GcxYZyyeYY6EinXiD6c
WxNhKM3GZjhrjS0ihWU7hH7a5wmhHeuQy9ooFqlcRzYvNJctycGCJdyD7mKSBG64Y3KTFuTj9CR2
1qX4eD9QYvcdm+3W2Dek8YXjKkpeOjxhvjAOZ9bzaeT4O9Mas15zuPLFzFeOK5yfAmbTX6Cbd+xd
wrZSW6uyPAn/XpuDJZRLGqY/gjUqWPAHeFMB4IdUN9Qt/WzcOMUXM9fS4uY6nBBj9F1Xx0e0yC9+
u/GW25Ck3WPuASkyqAQhDFjrfhza9SNzNuG0bUQmgsd0BrNWwWSnE7xvxDIombIxo4HAJW0zYJqw
iThdk4DxnjYbLlnnGsCde19kj/p10S9BA5mIzLRGKeHe4MXfaaGk1sQWJ9EtiDMopYcGhOiTLABl
BoW6gmZ6hWXVxn+rO+BuQQ8Qs6qnvveLrCBv7OQaWy8EOWVqLPcJWgVZetVk78lVtRUVW8bxCXxX
a+/fWjzfrxkt+ccxdlaslZZ4dxe4s3BMYGECxRCFp3ZFU3k880EUpNF2T3R0uJNA5ScMssYxmxAM
nqASQAe3lYYQEYTFViJXvBnSK+//iRzzMNrtgCPlWMa1QZq/D9HAdNgtbh/ehxoO5OoV3c/JsYWP
9mFSnl0resqUQ6+srH3hrBKPME7lpwfSy0r/c6W2id822gwOG8FPOt+bekyPqKuW6Y/QTTTl6KPN
WEtjzxNgqfM6UQD0TS3K/o7ylWLsLWTzLPruSHeTBvX7hkz5FWW5afuktQmxELI/UOfN0vuVInR3
UDYZp971n20WnIeHdsNrGR5Bwv2Sr+annKdmVBKTVi704iXkHuXVvnPVqEmCZ/t1cIX5L7S5aA/2
aRxIUcjhOwE9QMJMB+GUpCppXfkPfIPfnlQmfQqSQR2mAfQNu8t9/GY7AwiiNdxq4WUPzDoXNxA1
m7iGkNLMUH0xrEaZ+5MmFYLJHrfTNvLjlioHIn3oK07mfTlYiLHk51w4NW/Rhququ8HAScFdQNsk
ioF9K00PeBV+yxMs3hk6aaJ5Oi4xUsQODFmykpXjmCf9YutFdftko5EdBstncPqKolAKTvpq9XTJ
GWjBrvb51gQB0rE5ZGV4qQcBAhAZIEevqB6A7I/kuxm0oHSIvJhk0uACrVE3sReQXu4/pZUBkTOJ
aCkBdwIv4MZZRDJQWzDn5ztZj9s0NeNxOpJ27+1LwgrU5kKaXOxRAaSwfDMtCkDIhg6fIZe6Azog
R3n2h6g1pxaceyUDyHYhvnxschexodeN/NKgKxMLirhNJcrUaIqk1NWmrBY3XpVJxnFFrAhJ0HZK
pVlpo4Qw8qvjks+Gdubkli1fetK8i/xkYDZ/KyjUH0196J/scXMTRpkC0guCGGt4cLZI4Oe+FUE0
S+amfE6YZEVQktUsI2t1iRDzPCgzR46cWNLBLHbuYjd4CXP0BKt5w9yEpz77hIeegMp0yQAzO4iE
elrlczjgTvHY6sC9RgSt3fdCV42CbMbCBXxgyQNfdVIjVsMCgz67Eb5VGT50qY7iMmU44ftHcfjm
gTIBHzy4xkRdbL+xKvSv0DWt7KtoByinooNvhOgV3s3W6+d2nKWoUQ00StUkHAhsQaOF74ESjh6o
cetY33H6d+MT5+2AfCG6SobzNEYZjwES57XPqaiH15kWf6v2QYf+aeeCKm+GpT+7cX0E0TnuluxA
hQNnCfwXfDLORDnpdf6J5yUf4pvPDKgQa0WrI6Ojkkua2Toi0KKfcvknwU/wN5ehaMkQJUdcG+Y+
00nMbHEFzujNmZZVxK0Zk3aEAKj6YYJVaGxoaY6MnoAzIUVwbVkftHSPmINXxctpKAJ1vUaI0/X+
Hto/DqPU4YxkIhakX4YFwRZvzm8BSk7F9UkjSO3Fmm9jJxs9TsLiRFI5pYHsQHtTV1+y9sm9CqxP
I1oQ0yHKCAFdTHDLXc5e64rxJZhgQ4CtKkVKTUa/zFT0iPE04RH/vfXkzWR7Q+t39+Gcod0EJ4Xt
GYTkc43fFxqNrJPYwxt00FLYCg/y8AdZFthGIeeIPRUt6Ciz4ca+jhQqHVEK3Qyctd6UJGV/sUMH
SdiBcDkQM6KDMwqk9XaUwEqwQaYcSvLBYZpX1qyDHdnr5/3BST22Zgijn3Ti4SCQuPj3fNjbU2du
L+N+i2e0gOeaaEKHAmiGrEdExRYoLg8P4gsUthksyN5f/u6XjXG1HL+eE8AT8jwCpAAjJ++3RH9t
XXE1C3M3dQ97s2oEOOhn7jUq374kG71temXBgGxIT9CFhMkVl+Zhi6ZYbnSyYamme5+7sIV8xGyf
AbOBMA4eomvDFf36pt0/7sKv9PYrQYEGaO7qJQ7+sqNwyDoCcwEbxu0C52eJBiDnfKtL9Sxc4xxS
Gz4eqoxjhBa7iAn/5QYkWMfw320QhrqRPAlgrPzF4dUzu8DUfQuZQzRPgK+SfSlGJivHllcJaS7D
BrkcktIk/EcjdwAxiwx1Zx9AtXrvr62gjKZHSt7yKT4AJrSu3HC04uApO1DPWiGYTCaU97RDx7vo
7eBg6WZ7zCkRJX9a5F9RMEPC+KERDCRcIsyP//SSmVhE0VaydMuqzmQoc839QS0GOP4j2NVh9qqF
TmNUPLpYw2GB4MghBKST5iDcuE90QvUKtZvfn+UMBivuKjiASNyU8p7GQzTCqF/T6vr7OPDhfYC/
WhOtxh+A3VRwaGz1rdvyTYHUHMfwLa92ph12nqjPRfkYKIneILMwpVmTu4suW33qbohCJXjSovwR
d4GNUyzlQUGvsULXFYXOr04G/YEGU2hQqyQR+NnuQkh0pzJDPd+cWBcEnOBTmxLLX1jgqwbhsix+
rdmfG6QC2pqek/Sj9jyjzDDjmwhOPhAgYAXfNPVjyi8u14LwZiNsJ1eUHfoSn3E0tTy++hzvfqQ+
IviYYYoBXFcSod6V/bWYQ4crnegA9Dml585fs9XqB672o7QafLTIaeVYsQvmgMcnAD5vLuPEbuD8
RDigVyGK651qSoM0O7hOqtuhHQkI4WsyAaAVxygSTaiZAZ6n0AVzrXNO6C/RNCRGQwSIE655ZL99
wODAvB3ZF1WeE9lnmFXn4XIRZMIJXpv+7mE27NR3aH6+EwWX6uM9NDZPm4kcByV1f55o4y+KUUKO
emHQrEHws9JX17lMYGKCvuj5U164hSXw+euEUnE70d70+s9Lye+5sfUECY/9Ele94WOxDR5K6pog
Xp6RDnCawpD3GETIZxFpYoAryQG3GU1Tq5IVkSYPrBjNeE00YS48UpC1aZbP21uIE4t0F9ZBOu1F
v2HngYvHncJgXfklCONfirB1exDKZ2E7pdhauX6JFixuNnXJvBDk+IOp93vgJCETaYk4Iu7nxpN2
bi4XYZgVwJZrkqsABZ9z20H9ENGZ/Yu4BgIpPnhewnpZtQwZmkOxbbhc5uFvlSkvLkFPbOWDJx8f
ilZCrv3BqRoxwVN2BSYrmQK1FkhyRsUfq3+LPT3B9+zNZ8JXG9LriNK3LSrrHn+72917bxdUXZzS
G+PYqwFq1Xxg1AQnb9qpxEL67RxkHeq6xjjlyONSi6dizQ6GMwONkVP7Jj1BMqKIW8a4XYUMQbXi
Wfk+DuBZOugsDF0RLSSWqJf+nqMaIcD1MxhrQSYXUS0KQNhuo5KM8i7l1YdmFn48+LY7Bey+CdsA
NH2Wc2WhCfgb/yz+fW56ZtcN96FiO/bsKenlAlXM4LB5vR554LwYB4362pHgmoTyXRhHML/5TLSa
JplhbEB/BVBCL+pZffDimABK3omJ7quYVGU7GgHK/B6PNXn7ZDGloUAvrR9ljjaiHpbwKQT/5xea
MgRdMp/R4+5AfIhR/Csph4FVrBxGHSO3XQmx1j6AdAMvanfvWDZ6EntFmROa9m3H39PqmRIHv54Z
thl1N8qlc9H/j/WOiBxzXirKKA+GYDsPVquLi243LekILNmFTr/3zhJDWyI16iO5C1hobG82qesu
rkbL3fXdGmNBSVOCTLXFl2IMEidPD1Sfg6PIDzbYOB/dmzigQbhPIY6rQLg3NWDVwnI0px6xRdMG
K3sPvDWOSRxaqRRJEg3UxMPiSN+AMx5vPbnWcM11uWc+Yiy1B6NSmxZcrvabYeJ97+qGIQ9aAEgB
uCwZWGk+oMb1zPV+4cJk4zKWx+Mt/LVMr9LjZL4DNfWdWdqQH7+9Gg4SXj8NeHDIo8mvERkI5ahT
JHu6+QUNkn/TPAvXSPwcl3Zw6JhiaBp+uLgMIesBQzn8/rrsSzA519xcKWqyes1go845U01KnqGq
moBj3iDK8W+oC79t05TUYG9vt6N+ZLVbjzWUpLfAqinAwlAbFvxZAYMSw3yXeH7mQVLrrX2VkzIt
Qv8K2XIwMhBH8YLZUYvpPJIwvCM+v09cyhyhdGMHpUyVNa3tgEXdVopl6GHp1YSb6KLL27l4aKGF
7N4NgAgOjh5lTc0sGxH+Emjpaj2SiRyVFOBUIzlqSxW+Z2PNZ1et1wHytWXvDZRTZs2Xbmo5Rgxw
OQ6W7GiMFLR4XZNs72f5B4vLcWYEySStVjdv5hizoOM72dbyRpiUC5GzKEpjQnXsbzHu8ZebLI26
0ISl0pxDwAB7bwdTaNps2i/Rv+kFyPynOEDhNttWuO1iCqnXvYOgNRp+WmkhX0o/U0w78gxNUnDY
9FZv6n04lDfYRnxOHdr2bxqOsfvTokr/o2INsmumF1Is7p3GaYaYrj8yiGROdbpRxokTpHrFaW8y
fFm0cCyH2nORKNOVqCQ+Es9QVpz2VY4FiCgtsuJcAam4MciIZ+ABwHUbYF8/R3oynoImdbqySgeT
gLuramIcQckd4OWFKIC1jDY2Sbh1gQqCv+7O3TJeqkXBPnhx+R/gcH0tW7ji2hOq7qU8MvL30LuO
6cQDKbwvl9t+yQYC3S3gJBplHGMm97nopxb74o0prntJpBgXNqXbrrru4zKZ+d1HZcpa+W7sTTDp
dCQx/JtwHM78Mp9biKOS4UdrGIm7iUtmSIhyywRIhsSAl+ukOJh3lonOVLT9We8EEMGVnyRG2Lkk
f8aB1juQPNfiKz4e+akVHqcl8GFq59t6+XyPBH2BNI3NSmTR/N9bQ0kWgHyUZ22Qxte9tolqdQIA
DtTolz7rvuXg+o3dtwl49362VYyZyAyZ4bZk79QTe14BOHClmbEv/vMqqii0IstCDkuLj8hNihT5
vC8f+4Fy9US9Y5U/DYuCAIx8qSnrXWC1U0RWK5YhbCJZiyrb31L0qTLmJ8gTlcLEUryi+ZEPA7UN
d5/ssq87n945cNXCb4n7pHH8/l+7b81HIYLJU4Xj2Vigw76yyhQaj6HWgMHevFSkdjQXvLm8yTkO
JmQ04ySIBUIO0oyf23qLMe4iJvX4lTIr1ZR1HOurdW0mMnGWzWcysQO9MmsrB70UOsDddQCALnqs
Dmj688xTYgEvx3XzHAs7Hbif8xcoC+qxP1Ivit+d9ICUi6J0771FdE0eADeYnC272WOZmJeIjVny
rHRMlUITaGIFk1yEtSw8jNHJIg6FI9oTfNYMb+laeAuO3wUy9sUHBojQ5eMs4Di4wQ48vwBCh1Hm
57hxyS7LiPvx/X57eoppfLD5U7v34KO3o7N5UbQp0jws8zFgNCstt5OSVzVs7PhZsaECSGTSnky7
HInT9T8+7BLB59+pt4wmF1FjNvsFRsiaddPru8tMBI7RxG4SQC1EDbyAcNlKvhK4eeff/xLaUXgb
ZUxDGhdRxNdzGK2IuHhlKEoBVGqFtI5QHRJ3dcezpd3oMwpI3J/3Jlw7FO532/3QOpd18eEXAcQ2
IxBXcOt02F1siMNSD5zi5hBwyUuWmnI0V46BkozFFjya1fjzhc7pOzYpmzLKl5FLCnQBPy3TfcDY
iwZUybJi5ksasUnF8nwt1RSJ9rfwn4NFlxb0xLC6+C3XtLQGze8Ar5S747jU/vGOpnjS/IzevZCB
uovYRykSFc8Pfb1yjRdEVVG2IM8cRUI/itfbnckmGbhRVO/J9TWC5LkDOqGX3WMSkbZbqOQ1g75x
JqV4OE7xx27g3Teb4e42TJAk4runqkr29iFaIv3lKIqKiNwxftRDYJumbipKrM31FWgMBGAHlFjs
55wZA5x53kvNwzTqkZ0kh0yWfDpqHaUYbJNTNJKaMnw+tKLioz6/fti7NtmCxRnsr4R0lic7EgdP
tcVcrMZsoB6GmQzu/tXAEHuAwIGp0ykwvrjswX1EvkQZreavr68F9K25ylljYmz0hLvh6sbsRgmR
jnTHIA0/HAj3A6v226JBIVgIAS/jqz/5b2wMh77mAalzBXRtJ077cXaX7yWwbRV2gfXMqAnO9/fq
hrkRLvaI8gcQLF9vewsSmXY6nVAM4QIMEE4s4UrngTGXWHqu9I8kC6nMuuXNc9tTI3K7sUvL8Zv/
uNzSY7yPZDlyNdAFECOMNqI3+OgTKfRC9qU5vN35OrPnjxnsT/zxABZhXjiRzotmr1IgHoSruJs9
aZXZeBlhKJzePcphCOh+0EgwENDqu1QljQLlVTniYHIc+DX2gRNWebNaYmCdnfChgw+5TtNaCTRN
WBJBEOAxPLyFktPxDer2KEm2kz2hx+s0VbSaHNMgkDimD3pgB8RcOCHM4QmOD1VjnDIcgmfUkdki
amJxvUEOL6x92CfaH9SzN0uNPIIhHyleKnc3aO9/dcq+G0PpsQAE1LA2VTtA74X0ZiDdCfBX3T+o
VBpqITctpF1EnZu5xzZhRYCzm/bbMLY0GDzrCKSEr4biITG8KU+uc5lqwj4cdIo0aIiVaJWNPJl7
YZGqGqvMCpyX12eDDCWx5L7crMgP41yZlpQJO88MVxzQJf5CY57G8vHNVBURRCnaSrpZopovDN5D
qmpOPNxqcmgM9xkC9lzphfCwUrKfFHx5KPgjtn5ajv4UJGj5+1BpIhFQ145CHbrODW5lgSNvtfBp
5jG3VPp0IvKC21nyyi3cD/eNRxDP9ukF2EfPyyf19pi8tnmbYfZKbvovuCBh6W+hYUwyOGCo46nV
EnLj3AiBDLl+iP1asX+9dhl1U5oovHlyaF8R4M1lUnWgyN7D6ufkyGmRKXayLHdS7iYMSzpYPrPx
qRgSoiUfGtPRakLns5A+W/EeWP/dgqvrrifD4crKm1gyzgJIFEqsVAZOfJx2KauSA+NXOWIgLaRh
RhWRRzibgRkZix6iCJ7LPWl2Gmjq1aay7cYyyP7V2fZ4Qu/PbD8WU8E2FZHKNK9QiJzHddwGqFMz
kqUaK9/ukPDg1MpBIAboQeZVPFz0EdBmHX/K8hQKetlTxNVYtDD2sp9yqjphuSI/zuFIHQbEvvTS
OUI7mO2Q7YyH0yzPyfZoJhFD8CGeKRBhAGZyHXambIe6x3eYI+k+XjDmm2sHJNiIVq+ZuhfMUlLw
JZ80bs/ZUGIVg+TGZPbkXtoOUkkg0VM3exVKvfM902BKG+e6BlhUHPlczgQVEorAKf1Ksyo3/Va5
ZGNu6UpjLTt/hjOj6eh+TXPbYOjb1yYewa0VNDNIF4CYvp5Whw80JDuADmjUvGlZKWAUlmPTL9qv
5mcnW0BfL7U5yxK7nbW09AYaE+ChtcPuyODoNkzImoOoL+jIeF60N6UD5GEwC0WsIh6HxDHbZr6Y
zJYu5bvsPr2Ktpe9BJxdhd+0GnE38OtWeXO84q+kniW1Cooa3D289nlXUghXvuE8A9wjpVVgQCFR
ouVQz2vvztTBeZ90j6cmuTrHl7JcPxZQilvtJPwjPnkvtzJKHfqjt00rgcDBTK2Q+hUJqcEOO1r4
s9liU+LWsqHebrS7WpwX3tUI1RTD+CPHrgJUWHSMW1Kl1QC1n/wCvJKcDCqzicK3AYeWlPNXML9W
5zRupb6YERD6Pm3lmsBV/MzEJqJWZhFW6E14rPbtD1CGT9h5U9m39uYlR6VqAbsH9Pc46XykG6Ji
1TDAj1RVpMYt1h0KddufPqpcKiLmx2Ag6BpGwE7TGNa3SgvV3Z+zCjfABNH2izr5C4bdXEqOa6TL
MPoE4hwY7qWARAqxia5Tlz1si7qTgh4lkYSEJx+/V1uN2411foaD/VtqIQO8ZZnb5wSnXb+T1aEX
zMnavNj0c46Xj8WloUgLVF4w4ioNQS9WMAqhtA/zFIrilKAFVDMPcIHQMjMPPjrEqfpx4GpGKpyM
HzdsrtaQ/b+xxxT3sx34muZ11w7tqQWrjT8sqzvWcGdeY9v//xra2dSW4AuLchGZm5p0mqGn92AM
sXfDxpCUuSlBqet1uygxP4a9u+9tsZrcWdxEC8x8dXWsNRmXMIcqNa7Nv/04mCvA7PFeTni6cu0x
+wPgy3zD4DoZjNVBgb2Awne3fPPkscVzZNdRD6JV94BwQYDH5dCYAKAkta1XpRWPJgpGcUA84/Wp
O7QL99NcOkfs+oLLa2yVgcXPeEz/OU56HcuUwBja4i3dfcrHn4sYrOLqwyNz24y7SNgdcs9JRauH
Uaq4qdi1T7reAwNdSjtdqJVxfVEWjGI7IOqYKsd/pIv0AdC1rKc1hD0+HI6QyholN6bZ1FykfAls
I0QynjnI3sEGn1tz4O0zI/jnoIAxFhzlAtgOBA/CpVAFAIePnD13oaSlMrNVFTgEgVVNEwXprIcH
1z34k/0ZbOrIHGwCnH41uiHU9qTIbIm4pFt4X4vXY4j8Bi0Ho2T6ONFJymJAnb4X1uqnuINaR3pS
4gB0FP9lFz2B57Bbhpx1ONvzryqNpQJ+KrH/wLVQ1ngZDvCOVt+MgDS3n2wYnRylagAPqwacUHGU
4DpIhDGylfNuPy75ERNuRFEBjK1jcXBOqNVrcTBAfq/W7ILzuFzmRCPcDlFAnHKW12aUR9qzgixA
+5YSY7qJT/nqvZUkSTllIa2I8WR3UvBcA2hx4kDOxD6HTSTiOhF6HS9+4kWRYPad5lwM4uSXUJNt
9PzKRaSsm2kpIaVU3aJz53PRu4oEaeVam+vFkBl59j0EP8qna/EzEzupUeDaSGbPK1YQOAaEds4P
oKaypa4OaPR9hGRYe3auO/DtVO74glq3EfallE8evVBeGCpMM35/kNShJ7K4WpqOeEePci8OW+tf
PoBuTZAJgGDSKEmP34LD1SVA32ncd4YsQqjU6AtmVXmdcZr47ta15EsO5GMLpQ7dgdGZitKIB4Bu
RHT91OSjnyh1dtKcj6qMmwlLjA/pJdfBxeUyRBf5Loz/3nEsGgerRhQ5R+yg3/QsTSDBu/QuWiu4
PHY1G9S+UdCz2UB6luy96Sjn/ZS3kHQJbQMWtK7tufHA3QQ2AxoD/uWcIcazz7GpIjtNG+3+x94G
Zvr645eEX1iFmlCVPPn3NJE7LkRuAa7ujq8iHWckrKMqs1FKqt52s13b1CX6BKIevQ/zhkEbE2R8
RJ1jJJuTHNeYElFtiqpRu5WXWCbaEHIeHXX7regY2OIWZHVz6Y1xMvvbU6FqPcX5cqYTRUntBpKk
kJ6eHM2BJ1NjUjVHBWw/y7z4PDpemYL3reNPG2LdkeBkNoEZu077NYLgLOYGXT0rBwH5HWI3m3gL
wsNzfSy1ehMUaQaPBoNi6KRN004J2BNkeUAbxoRSsYxuWg02mHjf92RkRKTnX+xPZh5sMxkygKcx
GZqd9fhJALyAlioPvKgrZGRWhRnDAWcY9ZcZ4VRrdUK32EWep56ip6crNoWZcrXeJLhRLTb6ttXD
k72yggd4GCU4/sr7IxysjIJvjPxzyeTDLy/DGcnhwkxl6NSorWq9Ss91/9aF0DwkJwnntIzrCi+i
sTtZpQABBa4mg2cFIXze6hLzm7UVJGPYPe8wyptPfyaXN8CKTGWDTIG0Lr4qCntsAHozw+1SPIk2
l/GeKgpJVusp3KryvYehpZIxpAoLeNa70Ky+G0H2QXQvMr/WGnqDX6APf6raE4Renrs87F9vBpbp
gJEXksJgsCbIk7M/BP1n2vk0CBM8wleZ/dlodqI8bA+ou6nWkwRY93vltrBmHClsiaWat1eETJNP
R7gUkR62ARJh2nYtB+HgU33uf0s37P0p6jOjzVjcY94MDAJW9QePLQ/Km9/IIpncFqVsQzhIK8OC
MCbSM06NCZHJAX2eZjnVXYFuSufqQkSS0vN++51N5mNuOiVxLxYzEcCYnE5un2K0/ClLb181XdGy
ysvYyoQL05jBqO6xVfkh8Be7fmdVJd6zclFYyoj1hWuhgEQ+wzVA6ixqWxAjfw+evCOUFy48MBR7
BduHaoMnNfkYahZtvmt+u3UlqwONmeroOI7NRW6UBDLu6naGretgq5SvMhC/jNqpXnzVlpLFuFW3
/XP5Y5scODhjq6nHQuutBi5iRsBf9pgZhATB0GzWvVr25GZjAfBAYIsUJ12Fqi0+u+dfxmGhYS1J
Ydypo4HeuNmY5L9s/98pLRy6bsDMlr7eHZ0ISU/Tq2v71zfyUybo7Iqf/DLzqhITrawvzPN1FqMH
HlB0RMAy34pcu8S7CA7xOlb0AInrNa7DAKYk6PePq7KhzVP+d+lKqdAmqwdKkBO7RNDh62wjJPEp
7SEyK7NZoFhzSrMfmpQ4TmgerMo3Zd58wFDDNPNR+Xf8viW/XSJRDbgNhaMmLSu/x8OrdXoic1fb
HWszzDLfvRltQZGa7LnE0taQdvStE4q5VDR10r2xeqGPz3PKKo5mFwvkQAlJowOP9p6/k3IiBfay
qgSHnck1chm3Xy+CQIH6AhJ8hVlQ61nUTd209w+Du6ewkIBLGMDTJH0wRikUqhsuZ+iOU452jATI
wM3FnBUvtvZcEmqgFSB4v6olUw1e0BGogOYA6hXzjCriFB6BDuo+l8DB3NtQwJ6sNXPNkJsNM8JL
lF88b4Hqc7u6pWkBErtrv7FH6DhGiiWSMVpT9P567D2AqoOoQh8UV1lrTNGReteNPUb/Rs8scPlV
QMMNvRNZs4eF6EcqR+KQEubvdgjXhzgTKH211jqJKQH4LDF+XPmFnnI9JYii/tOuvwLjx7pe3JoP
2/UqIvu6+XXljer79PrQeRWjzej8LvOGjd8sFLTai1tro2qTIsiwFOHJHhlhlFVQDQG7zSpa2Lsa
sDz7biiJNt5iZL/by0LJ7OIyNx3FuB5PukbfsRktL8pCR78jTdrmjc13ea9hs2Y8MfjSTFpec7Z+
22uPJO6nHjbVwaZQe/C4x8FHtVFaNgbt0+ixPi1a0A7U4piOd3bx6kGb8803opuCTJOzzi9TI1WH
U0i6LlFvs03wh+fTBf871SPGXC/xV+4mejqYwuskSnHmY9fF1/MBUNoOEJJJJt8bOkr1oogR+utg
z9bOrVTT1h9KEZ9IISTldiFgbVRmkbK4REv/Jcl5n+HeR+fkEqqMTMEC3bnSp0rr1YjQgRjLGK8y
qf4uXcfEQ22OHzi5jL09NWKgmPyuH5T8FuOGgVLcwED792c84EynhiqQuZFg/RFZdqxCW2fCAwIU
LKz5/Nq1nU2I70VwMiun5Ed/z8tfZh51eclGC5nmiF6vimACLKbYggcXI4ePv1LvAqGkCgfwclXa
p++IQEmicFUopA9Doa5iJ4aRfxNiX2ONtJ0yy9qqbJ/jcATLBeRqOCeyR8h7xBBBbJ88gORcArNE
vdnWvP0KrMVF0I1f0D9moYF3v/zCJJyxWvLIAUid6zQ4aNRP05uDpWhIpuIxbcuOTr35tzNpXY2S
VAPeeD9hcBRd/kPNDxso+wsMYgww+6YWxpd6g9VbSwjbiNQTxYKCpmD+LuSDGGAJ4Ls9y8201mof
sjfmxmQR/yCXri1YW+9tKkJqRKr7IETSMpD5JPP2Y+U8xb5AunSPIgpKuwgAHN1dAQnuCi4mgSb/
rplpre8t0OX9vWQMl6kOAyUyTaNYBvywd2Vwz492VSf2XhYCB1AA4KpSMMJltLeAD+4ug31VfwoY
SeYSZZR2jGNFZ0ALmQvvevFlodEWL5mh6d6zovmyHtg83tLvYrRQO81/C5sx4gBsKGoEgR7ePYVp
iIPZghhMt/4hsusuPpuIEmvyP1fz4r7u+6hk837g7WnXPp1UFjYAHpsZmx1p+2+01HGxuNtqsR0z
w8pSPebInCcD2ZaMA6DKOpBMyJdD/VL+YUlBDnwH58gYhLlWeyzpYeywRiIUYm4hxXDHwUj6xj+R
PD3tnioTM6aB0n1xnvmynI+Hb8O3P2pAcNXq4WEtLvcaVhHuV1V1aDlii0O7DJ4d/C+cA8gKHBhK
YLgzyJFrtdbH6ImzQ5UbpXcTiSldqKWClT8vhm1SABZSn+GsmaxGOWlk5NWf3XuQzCzmbYOHQkKK
qocLidOxuV9z33E9LsCgGlmUVMLtuXppHQmgs+15L5PXWhUM3NZFzMS6w0zp3icg766bGSHACuXp
mfMF3TNBVEMzwnh9gFoxqSxUhvzs5Wq/yt1LU7uA/WgT6BpMWvyTfC2rNDRJem2CsDd+uY8pNSh8
TYuRfYH7ZBtAH5tI6bq+NN5o+4nbvLVzPFBVfYFPuROD7P6d2EO7Rr5R9OckGl94HrLGRUL1LfTM
LYTRVTYxvgEPb7VQLH7W4jDEu/HeTfLHIq4tWRUJwRNZL8bt1nxLmYzYT0rCED89pqfQrf1uhoN3
amTRcI7FZttLhaayma7QTMEqpHXjgRBucXamaG8ud76A8KeYCewg6yLF99ErZpebYoMjcsl915Gl
mwUjzJMvDe0ONIpgcnzGrr6QxMruH3wQtZqod8JfeLBWwbL6Khq1kTxqEBzwyP8GYqWVs/+69W8q
BdTClMCDIeAfH9vJyt00Dnt9iaeZpAE3e4NUgxVl5NEdXMTVDrqK+jRFatHFd9V9XqHGBErOXX1a
QbFhBCyjfzPw5ozte7BfNiVPAoOGuBolIGYtPiiyP9KtI6w/t7/M87Xxw8AWhVahbJL6MIqGtm1C
rgiib6WgrfpBNZV9oo0irBm9HQ39LD5RWxDpd8YDi5ggfZdIqRE3+GB+YZq0811Kmq9qLr4BRlT/
cy2k0+9zB4ffkUgsxQAthTlwt2dYC4LvDC4DHRUGB/2MIJErmA/TzguCU+qiX6wcqjZIWgOr+HPF
e0lb4D/i2JX+1CmOk93Llqgob4nISK3VowG7Fhc8MkCT+q6dkvjNax0gFuuKOGjJ9QRTL+J/kO/t
Q6Led6h91CnfEuQf7APINwR3bdW5A4FpJKVNxjzt4rdvZEjmSZBpRsvOGnAxTuROMLfGtXKoLwi6
P/MhA9uPu1EEmx7ZqI8qVY1CLvfjokBwHtD+JpDdLF3PVm5sASRlu8AVqEHuK3pZtdR7eVuw44YU
62Ti0AUSLfFsyV1hqvoUZQSnES6SW+zq7wd1mTwhLYGamfMo2O0Cdo4CozPc/+vlpcYNYP/BKA8M
EOgJnoIG/NFT/q/X3z0NNMrQmnJHKYe7vufJrsCxsNkSeXsX1VhGOqJZo+ReSgNlPcgznR3fiU0T
hbYSvju6UPOKijv/EqfGIWfaZUgubDX7wph7oKY9eMrKGtOe60VIynhqv4GVOBtHvbMwf9XVSUkG
iblOx39jm8LHCd8N8aQ0PEMEJMxduZH6DsGwfg0S9ihhQIx3w+Uap+wGPV1wXQ53QD+vgTUxZ/I4
yc7H8FfGoe64qWl2FWQkdtKz7SeljkuD87isWhEAeP4Ux3tnygXjU/CbvFnV/HK9eOK9iM5eXr+I
6+6CGebgBIWTA0rC0r1upfubWdhEWu5Xwd9BKFCT9tVg0ry+1NTaVtdz1KN+aO9oWnmRrXXm8TlO
vpxMQn7GPB3tKLWovcipAXB0c75JBpEmvWT4EdWIp60khbrlLI0pMsPb35w68CHOHx0P0Ud+Fkur
pqZpmPAKouwHuBGvlf2a8ec+3pmvTpZV2OZFgSJmwUBsCKFmwCt0DkEME7Q9OxFrYuv7Z8PmCe9j
pboLCF4vECdf3AKcUO0h0IlcGjvw70dJ/jFouRXwwuU4W34BdBnzIbySS5LuDT6PBwJigWznaxlM
euID8Eav0PGuhmUFxbKGI7OiQolTek3q5stC8m5OGdvGNpDJdsWeKNQ86SRJPsZENOKI/vAVSKL8
Ly+c33jpuyaGW/jIR5DN4q3e+ptSLrlhwya4/DMCZUFUunC7GjW4M6CqtNIrHmjKn1dZJnBYiBJm
9HOQm9V0vT3zoFZQnAb68EOs2NLN6NkhPxuV0QhENYMhYByDNsc+jBEQuI95xrNFk0feqhBXxBL9
mE+LHoNMSKdZDKQXPvvGx2b5LLeiI8NzWoj+Of//dDDyB+HbjFS22dI3uxIYA8k+wU0+juo25ITQ
tMlAykV//5L4LQU9sCeG4ytLLNGZHEFGsEQocObWBwmU5Z2iSq/BaZeZFHcn4MzzypSzY082tiN1
OIfkejWyzQOovZ3k9OoIeFFP9KZ9L4Hxp+T0bduIfr0UYiNTif632DUweJ+NHWkbk7lSgd8EVqeX
YBpbobNUUXIHfOHLjIa8Tm5CdB129G9M7mX3yqKy35drTxdiufNJEWdP60Mn+0rGN4EOgaff/fSq
xPpDqoqC3l+20jFmT1JxY9onZ8s2COGBtme8OF8pT9keTGsjEXT6Q27YMUESdWkJp1KEB6imB8bv
RG342xs5X+uJbjcwqEzvUiZbC7YIXtrumE0SszTpnE65z0NQ7JEOE4TaYqrIlwS6ODVkoeCQh2pw
6bqSoGFefWix8oZ1qVhBu38+9sXIgtqwd81fR5j7kdVnavwceMGd6vDuUe4cUJhDoVXFvDmcWUOV
/4yZgTI+3MuEv4+DRRLBEj4qrhb+b5UfiJdJLEIX9uCpfMFil/LUk+BLF3JA29SBTeijxqmAgBq6
aIZ72xB5AzvyDVwg5iisg83u7qr/YQQVTwAFHG7pGVNeenyElhtbEC0s2n58y7nNlS9jvoJ9HH2s
HLryM+PSDt/j/BZakBOZWumJ2Q9PAsTmhjIIyWkervwqW/4ILTzNUYmC51t7OMOCtc8dU68aeZOD
Ybfffz2HVCIb4V30B7dFldpA40FCIpW784CYQDNiVezc+6aGdqIqUIHvpHO5tvvuC/VSCHUBncd5
rJScCtPeYhNNipzmP+0Zua3UQo20TkyItG1i5PL5FRQ+qGGiR+A/Sgm3ecbJ+nbyQaBhahZ1MuZL
Pmd9H6HMAySJlhDx2nxjNyL3Fmf5ZRMNf56KtTnZxn59VvHbBuqfZwRjlzn9h4Y++1+Nad1poGkY
z96wL1Fx6maoYd8B5V2Tgcgn2aRfkz45wR5AtQt5Am9uuXqrW/C4R8irRSq9hlv1MePS4LX0CIK4
qxz1UgagKL+KFDbp+s67J7W2J0s0I/Ga1KFCjblNJcNzWqGKRFWqPStt8onLogl/LTvMPuJtXLu/
TUlPCTK5cTvDADJF8kV6Cgb8b7KE/irQaz63Qm6Q4/xdQwP4veIqlbtBObhSAMJ9NmE/SQwg/m+5
7Epnku1claoWh9eg+zb1ANy3ocNv25sQKE/fMQuMFrJuqh9T1F64nCccLKBgoxGb5wQmuSj5AX95
Si3ylTcezt8/RLk5/FAIJGePH3L9Mvs3DeP2kiC/Fc/Qe9kevj1nvGqhdzUE2TLGy9ereyExgUzI
e06JcgtlfbDAFB4tPyY+3zHvuvmTfSDsqKKNN8Kc//vqh8TB6pBF1Tm5hFllX9mS3Png5Vaain6z
bn/63wyBKqLtgwobdKSAu26kVfWJvsj8bNUmasjzg9UHbIMas3oT8A1gxcWFTJgL/nxUodft7ma5
ZV9xBQySQrmbOJjSN+gryrLEnk+F7w++6e/Xz11zWSJVnWRRv9s511JQqDxydXrDJfLH181KU6GJ
2LX9QRPV2WMsnhwEikSzTUhTvH0wsr+Y4XcVMUUYU48afHDm2OUkb5fj0MTcKnN5gjp6EVmspjYv
jmjoU2dnbcvbEkoLJKoOXFOJEbEzMJ5QH55W+Ab10NppMsbU/TQzC6EOXJZqUl+PdxD22tc3fDGB
yI3KY8LMHqm1ksUoD/NP7Dv7uq9+DHxQl3zZwA3HQWe4ETn9Z1EiIEM3amKYdWm9Eolu9hBmPFum
XGnaCa3JtnmmmhNbOUivNnlO2lFJXe6jLAfACM4RLdbJXvi8SPoWrTi0PTKWGMNj+u774tuSyUD2
ubOlv2mnzpZSjX5iv5B7nY/EkOlCRSQSeuJdGSxU1ho84hA/4qquOtKvjSahx2ojcHa22IfXQlU/
pVLCYOBCW654azqSoyl8qM6kUnx0TTyLdx4mxNgClC0PdUpRxGWfUp0037Xx5VghooA1p5o7ui8o
hfBqOWxf0/1EpVC92tE03d5zjDVB8w89OZYW6NUVXhocnTnk+zr/jga3/7Vxyb5wro40b/yKO/2+
COW5ya/3vfCP5CPsYd1yob//3qhfxwXktZ1UGkfUX8MkDmg4sgPyGsSPvfp6R+mb9WjgvKS3a3md
VUfx7bn6C30/YXZziAx/lWK9SiGrvF5h+ja7G4k8q+vhhZUbPkwYRb4upaQx235w2Jh4y3uLSJbT
hBB56xj5ZlL05M1E6yesqD6i4WNkPOM4ettqP01SLo7rKYwKCnQxLC5ABaJwphq+C0C8fQKVMoxe
N/FVoZVgVNdPTagO4MdbmHRmBLEI+DHZ26mTebo5j+XuMuti859uT29grcXpY0gY8UQXObAMQzQi
cvJVxTSTkZRB1aeGCgrhaOo5+jDKt+Jb+UXbUq984LVA1aTCyaZDpD0vjXx4mdotbbmOKNLLXRUI
DZAIi0yJHK/2JGHDCuBMXcI1hbfieUi7xyu/fecJH+v7a5Nk7ReH9dEo3TT/JcZC/LRYWFRBOP/7
WV2Ki1QQZqHneomIETVjAa6b7ILsBVQkHC4koJoeBK7TJTwuAkRpkNvXLd8BRmiLm3dqBGXOh38/
1rRsbsSNNghEzV+hmPqpf5Ber23M7yu/lVRINAiv9Ri+0pUm5t6nwL9Wkwm/ZfWRQkxq9PSizx4R
yAvsMdHQPrI3leTMGTiGNNEZXV4SGXCmdgtmC8gqcWYFFQDX58TZFncQ5JWtjKQEhDH5mRmixs57
db0SwC2a+XKVW0PGKUc1EK6J89JZj0/BGAuUsWfgcEBuWcFKDjZOAQ/i5IwjgohNkn7vSHvZtBXd
6Dl+e16sRFaH9FCgis2RA2SpmJChjtrk4W0/Gy9faveZsgu76LAKMMHA1wmkl9xNkge7xbg0TqfR
rk0A4cOpn2ZzopeF0X8949efyorxfTMc9qaa8uPPcc84PS0op2G5ufD26YpU7fLiBGa8eS3q3mVQ
lKxQQoAFaFoCJyeqtSeVWnXDSR+5jc+QVdMsAnmDrhcUT0LuII5ggxeCHZe1SOcNusKI6o38lN3F
g7lg3LOcNZHs1lfKyNFkRKQytA9SS29Ea6r03nqxUhJUnkDmF47+jRgqjirDH/9hHzhBEyy4tbEd
EVq+m3lS6deO/rPWfDTYS8brZjaQqfYDJEuX7WBWU2r1oNUfuSdCSWGLt+MrE7Nh4iPY7BUMItda
qHs+t4o+PvAiF/5cT4k6exPafi0arE+Vs/Y8ztWRdRPSildc9qMgn1r9kDeqyQHz7zyv+3WTDzbj
EDO8t4WzvWK6WHAc7NVcL2i5Ln2kjFj0rxHS3GeQKH10MCjiL7EOwTNl54LFHUUwR6Rg9VcI+qd0
P441iZoLlMXi9vk4KF36Cu7EvHlcBOJfV0SJwq9BVxlydW0dZhBDVWfC6WR14AvBQo7hGeyQCM+Y
v3jlPkTM0Iu4jM5czpr7mv4v+OFZaNFhV0IAJVdKJzRLSdWnBfu1k0JIRchgoUK5gsSNa2HbWe51
7AiOr55shl+e+dHhT6nPOOS8vh2ApFYNDzpXuZ6t8oKtwhP5Zd1BD9YcJtOdBd+kwGmDUTd+w4N9
PUH9iYLX9qmIYqPUVs+9zrmzbYO3vwyIdm2k1M2L80ThOhHxQeetFFFqHVbamWWjODiXP0Ap+xhz
jS1/RFnYdLDGPl80AXfyn+a81Vsja1oU2y6UKBfZ+DlFP+h258N9zIcrI+0FO8C3hCZCnY8i51uv
O0kDjmsfaJvQr1qIOSezf8He895w0gVonCAheacGKLa/yvjt1LStuUS2d6sp0Z5ZL6VCXncPQNP3
8Qw5TtZXMGWla6NqgaBJpduJJuYExVMAREfWFxdLmnYErt9IjfHMUd/l7tAx6PNsaqWEP9P7HPEA
BbvJDtjwyTtTr1JhSrB36csxxAlktCD0Km83eiky87FlPcd6FPk8MjQsInSuDKoXIL1s4bORpVsZ
0ZbMwrI73IKYj/d06YjbQ0oU7C7nmQgRXRHb2EZpbiSFedrnoEPP/y0MKfV7g5R8rRDYP5kXjE/R
OQgBYRLyvllwOiM8CritZ7016n7MkIAOBBrr3UKOULfnOgKMYUR9cSCJZaT5/PxKnLXIyErYIet7
rus65v/E3g6O+YbyoTNTSwUKqCu1V4FjJ5KXSnpn5ibknGXQ92zBklFvRsvCyWiXHrNubrSDqXE+
YCbkjSuN+cknezTN7KgxQzFBxY6sS6BwQe2enL2pmfeER0ULma+t0061GrNHAz5449+MaWUfWvNZ
6xPQh2ci1Stagnu+pCKHOfwjL4AcwfgKf9yex07XgieS3L0qnPmVV0IfIsP9X5Qn5d8rloD551rG
CpNUn4mkqAQu0Dx+nCeFKVQXhZISW7H8MmS6l5KjCPut11QybcRikGAd72GeJt29t/Mbb+mBJ02h
X7JqmZY8I56ZzEIPUQC8Zn41/TYeMopEvXY7aABSyTLvmqAxk9xbzIrJv+ETLIe/OrCo7tLY+czs
x7UtsD8Oq2b8MJ/ysRP2txBlMMA6v6SkTJe6jhJqSf2S7lbBwk2M3coaHHOjqZtls2FxV5NviArs
MsQcIA0sEcKAYkufj0jNBsDrUk/iWdIt1Dma92gzz34QHVrKV5cUIlnTlepbYg9C3xe2xMDCPNmw
/Q20US0Q3S0vPshtmhXcGynHxd0ut6SQfzpzzaIg7Zf2uEzHvOSFLcLcw982AwEWdi0MKghubG2c
2I0HIm2Ge1XVkf/Xe9wEn3WtSGiN0l5o1SIJPgSklKNQueAY1G/65qdGAXSCfKBpkjcUTXjXnhz6
o2rlQUQJQnemE5u7bwTglkn0NnbmQiEIlTRLBqpqIFqCnzTlX4/0YwEACVoYFWFkny0UNOUvRlCf
LqhpkIMX8IFl/f/IsLz+KL2PXWkRz/iiBsFQkSwrDgQfn8zL0IwxgklG29hs4f+vB47/rMIU8voV
wvBw1FKvjtSmqCzLQH5USqfdmpQCX1BAdfv4c1YaVyWwK2sLF75he1BLrZCggWPHrSHDD5CYSxIC
NbDwf1OCbcbM72/qh2rJVxainuEyg3mSfz24eEmKrhffq5OtkufaER+RrUhLTZK0z5Vn3tjtwVJh
KdcEfgk3GmejvZA6ElMvlvMBmQ4uGWJcmvi+bZ9aggzm0PKWoFJElO/Lx7hzat59M24+hS37JBQY
IJlJatV6H0JCO5qfa9Qiecx7bt33aMIs0wOQMRS1rqGQVVRv0d/qXUTeV5xU0sBC339+GP0QU5EO
CiEivJ1h4iyer8mC+YY4XGc/Vvgbg+5gj98I1o3bTLQuE1H8OuhivE+Eq4IE8PuayrL0UCIy0EW+
Kuei6jhwiItP9nQjlPTXHe4RB6QKAmPx3gNpEnOFY1lcOq3kSxK7Zee+HR4zvxmEnZfJigQmM9e6
3owVFYTZ7bo5iaoiOH/amVwkaOnlvXRucor33aiUfKpmiqc3EHsZOKNspV7l+kJCHDed0p9Ljw5n
PGvTasgLzTTEMbWUmjV2G79Zj/Oba86fruGL/0cF6ckK7m5O+zqR39EIrNelbAFpRVP0bF7rXKoq
8ywZ37sVz5HjhyyyRKoNknheEfFBOs6cQygyRPjFnFkf/OuUHmOSRw+3D4E7/duFqN1yuQw/V8ab
lHm9uld2sIiTcAX8eQs3igvJq0J2hnLzokLGD1nsdRAGUjs84wucXPU4vnaOvcF84sNkov7JOZ1E
vi6+k0xRvAfQNtaIcuUNNk2haVOGoiCzSy+4HdRWEkcqf2ObETJ57/LBwy8lcwhLuGwla4/nksM0
KHP+cYcNwJHY//Ef11DC8NyA9TgcW491e8rOTRjmjMSczjvLv45rHBGop2Ec5c+cQ8QiDm+XLm2g
t4afpz8TgW0GZ2qbuxHOnmFZ9sFrTI62nJuPp19E3BTXAWh/VbQlU2mSqhIxmP2TWXB0w5Cqgv8o
58VW2UdwM4Oc3X5STFktsGvsAleI/6fq+uMojkXoviFEv36jhoP+CnWTDS0k8o3OqRUrqBcZ5lDQ
ytZnA42tkEcp9M9waqKrbn9YRkDVXE9tfKkA+haQee4Lvc2j5glkhKz2qTpPrNuR4u6ya20N79cv
yER1x5nK50brpJKm1C9ZD3hmlKArim/v6yK09AGWpkYa5WgR3JRLN1vPNiAALYvocLoVVsat4jGu
p+oHwLoOXmJl7UGGRsoRkawrY/gf5gxSa20vCLWUiodhFqgONiNuz6wHvSvyNVWyyE1T3xF6PtCq
TesWj1M7pXSG2688x08tieRW5GLQB/KOSKkagWxTrHxMgArHwnh8mT3yg+ojtiKkr3cArwIvy28V
TYS3z5L13+SDF5K0kwaCgKAXiDgZQVdo/ScjbWzTH/PEvzXU4f66cWMZBvxKGFicu5TOXaJ2Yvtm
kMSVIk94atfM2vvcpeQfixjGTgYaQK5LPVDVr6mGS885VTy/VQ8vGTkhtWUfKpcnzEL+5Fh2i47C
jgpkxngETPdKAfsbr1xyPgVfouB4yg4HECHGkCOVwa2Xoq0Thkz0TjhzbP63gAvlDGuBoJJk52gJ
0zgzEzayhvLNhGt+zAKXTbMFrFip0GuAjbDEasBdvnY+kNIVupwg/PsUunevuN+WOFQJJe3Lhw1f
EC1ByWr4cZ8oXL4LEdwP7SL0WPAZU1KofpU/BCIQb/aNH7F+xQ0i4vV95dFhw9+1/roZhv5GhyEl
ZFQPT/hZIEEZudq7me3K2Q1+cILlmR66en3iVqZTr6cAFSaNutK5ROdL54JqiC1MoRAv+jIhNYAI
W2s//kUhoCrrDmJbq1LQcGK8Hts7ZS1Rx7MibCvE3Ywxq8J3Ml31jKy++dTAkLffEqP3enfXX68Q
Ta41b6zi8bzchT+Zhv0obdKUknJBdLfSgI/N6L+/tM1PekHOhc/eo3VPFZ23UMrZ569u2BZieYyU
8aSgrTiTlRgObgy/WP9Fk+36Q0J1Oe7ay1tF127AO0y7+YuQIfqkb5vFFCJF2SDCMY/FIcorJLVJ
Sl3gFFr4JwyPEio16cb4tOyfUeCYQW7V9QUN5ojy8jTIyAik1ILlAb0ekdZtAkDbdpeh3bgFYQJu
tMWXYHXq3gN6zyfJba26gMMpXVecACkbUqg/aMy5hxnD3a+GQZi/+V8AiPguNac2trk6IcPAWLes
5yId3ZRnY1kmc9w4QHCncrEIzEEdIovwbS3NI45kIHU3XATGECiiKX3ZE31LZEt0zYZSB7mDNpA2
4VJNlATwXxgcpIiPz3gjrNyhiAf4r2jU4Y+aGYxKIFX5nm4XOGfVO35os6aaV7zAYF1FRC3oqDmw
8nLaEbN1XzY9eDz3gGrIhUiABJN8sCHgrWUkSJx5UWtY1LL9d1mwcC2yF5UXpdGf5Y0pJVhbuIh+
ElitZZFw1N7L3kzEmGy4Mp6YOl7IkPotZelAfvXTsUmDa9S3OpFJ3PVEUPgkHzBftnVc9ZXHXLfB
j7BH2EYAYrARlzEHV9I87kDnX+gZriuI33vJdkc/2NSHSev3INqIa93bmlp5DV36YUQvXbzoVLxD
ra5R/b4aJmt9Vch6hgIrdkFp7elwudWijpjCq5b4LMHRvCdMqIvoGUk1ga4GK3ozXIRxfBzWjw1K
/yUVPJQIAzjOPOEm/eslA52wuZRYa0HU2plDZi1E9Chxa496d2KSTbME05s/6RswuIBcNgVSB74V
Avi+X6nl94nMjABFUiz6XQP3n/uvT3Dk51JtOem9ic5LTSf32BU5p/4WnP3NermNIT3ZVmOWWzR3
4bLbgb4Inu4ioUME/zBoNByMuiZPM0s6udhcRiwuJFXJB/sVBK/XyJtP44qzLVX03lqx28Pjaib6
pF8Zc4Xwdy8CVl3H/gO9EzsjekuTy69JUvTOZpk9wm7kphlQuHvyvhBgnOzpl+cyApQWXUtnIiXb
f7NM1Mni2R83qUXXXQNLRrtAkXaCU40ef2wRvE1rRUoyXZ793511YzbOTHXy2mtjFOypIB1OhKbh
0rYYcIylSEiIbTsdsi4NwDo1xeBgyUbFvYzij6d+rQicbkgYGNfZ7mDD5ofp21aLAij4snk3a3Gs
MuEJZHCNN+pcN28z7Ziy11P0oNxYPpFhe5OB0ROuKO24YifwCnWTZsTG2dQqm5p8A3+z+iY36Vfc
I449AagnXLpwaAGR9avx02pXJQbXL4QVNzM4dBN8y03oXhizVqotW41Dbnu1h+/ciBGzO524py1I
aaJ7FkMrOpBsRn67GwvuosK016HsJJF02dq+3MdydrVg1Xes4CepE3PSap8JbMggGyFe0tiI0D7v
a3mm4LjNzQfHxXanSQCqEP+Vx7QSK5fo+nKpeRLm37rqnxIkCnLCKJJ4s+keu2cSJ+B/LvxIqE1l
Z4No9xDkzhaQzG94bQhGuSOQ5Hx2iDUN0aFjoMb7GepgwTGddHKKJ9wubE4HOmy9JlqH8vFgZkxl
lvzNMnsDfWmwOm4D+o+PU2JhY++DN2yd4X6h8QiJGY8TV2P7VXvCeAb4ZjTc0fmCFfyIThEcvO4x
zjJaIxWlQ1jKl3ClQ5n46hUFgxLrvFTbldBMP6qLhcqgV7pBjHTehkQ8/VirScDEkzPtJu9hC1PK
VleFS4NwIX0RQwMu47W5q4WwBCG4eyqzbP8IZRnPhnucn9b/GB3tfStnbCEFQXBPFCu3i7T4/4gn
MW6VEaQqKSKlSVbygIRIdeOR1eFj9R+1zOZJPNw4Uap2ztHsN1DdBzlXvWRVVPSdBOkY6AtwV2lr
lVen3WqJW+XY7NHj80b9ycKtXEiNpVHutme8B9HG4rTZcaeGnnusri7T8OwHN6t0F3Nnm9hfh7Bc
BEUUY1TbXUIc4Ot/7UMLYYEYEDj/smYT/Bb0lTLfafnn6nuNYb2qGrIMMh+goEAJl9H/G6EgsLrr
MisraUkFhlfnCg/Ub3oBQl0KoYADaXHt7cVZgf9ClaHd3nhhcpqBQwFB13XiXAobvX9/j0Fi8QF7
LYgj7ek1tIDugZTJHEno5F/LAVPKNMclTl2h2RGdqoPVElxp1CpEPZ8E1uwl/bG94pBMmx0iGZOC
H8Rh/ZgHb7QXAXJT8OWWDSGnS2Xdu+HHCWU6V7jHJGJah5ZbSjrub4OyBJmRm/40HodFVBK0Uq3w
eRzTQEXLVHl8Q8yKT8MGqOpLVxxPWuCLlQIh3SbVSU26N8Mh+ZTkAPCG7IE1KobB+RnCoGZjtO5n
18gT+o5MTw4fMpJQaCaEQmlYHCFucRlqNyynhYO0sFN1LKc1s/CwMTrGAdeF5FbTzFN/kyL0iZuf
frS7nui71UgwGvm/YSZPWw1erKybBfE9zjePAaRTSd0cmHt2OJPC1jH/ykCSTGVTjVjJbNCu5a7g
UyozmplZBLXFC9wIJ4vfOcvWReIDC9fHOVn6Op/OKk+M9DD4MSX4n5rYqII3lYxDWbn18BSbeNNi
2yXWkjyw5/9T7IqXvOJZITdKomc75jIN8f73uwrDnD9947PmeJJlFQSXLFYhsjpL011UwXzFam4O
hpm8sizaTmqgz8voX/Sciml1VawjMlYYUsqQJQVH4zyDBsDAFlnCRCWomzdTfJibw2xYnnFcoItL
rSRz3F27CAgHAWgGEv4LYXU3rF75Rgza8XgbzMDVo3W7oxAXYyC3oZLGihlgSQcPm+kvd56duUfv
khItV/AJjwEUneUxU9KglAew/gtZO5Vf73Qrrzb7t4okwEZ1ONHOdhANMEP3KgwI7FXpujc/vMtU
z3QjM5xWLCuR8IdOzB9LlkKooecfeQrKAt4IGV+T5FMFVG1aXGoZ1UCvVTb3c7xpYQOOT+1mcgqh
9l23f1k7ZjDCfm0q6L45DwY8NfU+ferInBltxxPSlZamo1RXGr5TX16aNpqpdhlOXf2tFQpbAo5z
dYMZ7+qN+FIkd2bG3gJdZypQP5Lc7MyWGMIRUeW4dz//TALaIpO1JaHwPpVQ3k3iCbm7JQ/Y2fGE
9kjVmmh6vlbniT54ZQNc10po6o6CX7luZjaUpujwSblqpk+BOYmngakRXN6I1+vk0cWt2uLBSTUB
nFMdtGuxTz2QIRfOOR/qJLLwY4G+TXitt/AWcqE7iELrKPeoA7RYTQN4mm6t+UL0LrSKaMviNV/y
WW1kkHy19Gm0zJ+OljHIDXeg9Zyag8w2qjJ/febQ/9pHRGrPUjE0Qp54ZN65iyANAra4SIxSH61g
fBi8+SUUCBG0XtTj3A0R7hySZp24C7grkv4O50Qsu2Ij8TIB4Y690jcOgJ21BYOYDfKqWXrFqs9q
kbl46wS18FTZCPVZnkloXbV0IZYfLTD5MzJrMQxT+gOiXCvKBP0QkRyYTcitZ2E736NlmK/JLsHG
Z5ny01nRyHnK6nWfitYwnX/WW1Fwd0w4GLK099fo93QnV3CLjD2uUkIVaeX1IwJf5FCY1OMBIpEm
IjHTSR4kPPH97ds9/Ua0NCl+nxBb+uXmArlLbMRFZz8cIdpNfcw06ljXnilDr6t0JUtDCcpjFeVO
IXFOxowA22WsLTV6dsq0ASRTj00wlsqnmMX0vcGpAS+Uj5oipFTJRzdZB11dcJyWkFOcGDoOVuB9
zsr1INHEUeTmMEnPgOqyqf5Zm5Y8iPaxAVC2PNjHDj1bnbAToGVRRRYzrvpvTnoRH7Uyb6coXQWP
YZwgkMGgCwP++vKlF71Z3Xur1mRkbvx1rJxLP7OS0oL+B4fYwUaUfapuEtf9faikPEFBFJGkB2Ok
rwQ828lboNFkYTbYCi+mv+oxFxbZCeQRlDHKe6RpAfyVwu+JRZeSW+lSRe0O6Bf2tm2oO9aBLgEN
u8OPc0z+YmEH03cpdjnbkKfaSusXM+Lc3x2czBUVswof28+jVEer9xhI/mgYJcxxYlqrbbG+33TZ
CrS2fyXCu88rZzvoqmc2jclQoqBc5VPdmLif/Rroc/Uc3XcvMc3G/pHP4UpiHJA7C3sPojN9Fkl+
jhrl4P2kmcSUPKYtAjRf4zRS8+QW5LTnCiy0KR9JKUmAGnQ7TjzBi089pO1O0U6d7RrdX+JmFDyE
17/WOlirN+b+bXZaX8UDfdAr8v0QyjqCqD+c6cIDlS8mMFwhVXlkSq1GgkwbHzW7K5dac0C+llSK
HUTLxdYYfk8Fts8SFCgKSOolwPvFasB9DiGXGxfrO/LgkHOkzwpsBiUFRhU1oKHZNrB2eX3BBvA+
2guyltvexxtZstjP6hs5ARLtwacWv5JEoBCbeGfQiKFU0Xu4oTbAY9FkMRUegFsSRjGNsL+i68N7
MFZW31QBPio4Ba1Qazho5z3L+vXIPEBnse48SEw8mtUrT3rzn/7z0yOsQRJU4a/NLHztjEUB17hK
8d2MmDXqIYY74BAhn/3Hg6LoWSzrud4bsShpQlgb25PVhP14XbRym+SIp8VJ7kUyZ8pK4+fQ/ckF
3NdSjsVuOU3c4z9+HnPzJHwW9JjskbPpNZFz2k7/ZMot2Vl+4iXFhIxsYXMdtP3OloxrJtQh2L7D
oiJzhq0+13x4HAX72mbsXQztxz0SeJT4pTx4rAevEPuUAB2+GSfMR+P1W11RjQgtCVqxW8OOYnUy
62zg01Y3S4paT3hKoabkf0kOGjwQn7D/LXeYpQAMKkZPBPud6QqGGXb4tMgFG7nWj7GhjZKf6Hm0
KJxSV4iSzZ27RRMtZm6YTql/9+LUfhWSh8Eo8MPTyndzVJkZILyK+FkImAXtRR2Etb2LeIO5Wa7A
RHapxJyocGQvmHS+gANUmVmQNc1cWMEl9aAk7NoC9TU5/SugcArPOIEWgK4vpyL8ET60po91td9m
iTd5tlbT165aLsvT2SseRC20q2pq1/sd+kAn2SYfR4ln0fiwQ7cFrpPSHvKeJrfg4bEK+ixr3jNz
z/HtV1VcyDB9+H6NixMd1fVinTR/AF2EEXPasyO+wIC7iAcAUpqe6pMcdEVlYlN/1liGVkT8zk2N
d3Z8EjqrLb3+T+LAgCictTPG/gXk6HiKovjvCgYzcPXi4eIXxDvds3hOmOEt6I74aCZpm8I/ks3q
8LPxSkPnufTAjsDE5BjPHQLy2pBRTy8Dr/nic2c6K1A7+JmEzr4WvhPXW9bmqp4NbEtaRiMt7qQ9
iqm4X5ioS+waP+onAL9iQeAyEZ6M83l8cwau0TQWRQcPtTiOLNMXsGsMPDKLLKpoo7OZxbGFGBwS
yUh7zzbjzSTU4Nhn6EPiYBZeFnrCKMG7r+JcjkZNu0g3HfPmFFJ/FTos//5bizmEZCPWsVn4NXY1
OAtlUCErdXuJlF8MLgySuRo+sXA9+6UlKg27yrDg0wzgLeqmlTBAW+LZeq64e1fl0o2ggqbaOzYw
/suD2rui53Aq2CUgGp8YV/k+yvtx3RjUAHar7sNbQfNTO4AiyZNBvapc0EcGDoL6c60xaq5+YQhb
Gry0wm3sKYzffx3O+WlUnRyV8m7zsLuEz82tZ8MuSUeVtxBquyJ6f+pkbaPqnuJRuEwBTFULKf3N
2O0C+6J6v7WbKQOz0BZ72PR8Vv5vK2TgTrmtekzoy0xaBPoajefaH0ykPMlUUcoM54vmpwmttSmh
mO6HupZPcYW/bD46bSp1YTr6mRfwPQhsrBRkPl1aDGFU3BVYAKRImr3vQilj2mpiULEZtOoB2fYd
hoMn+6EGgAPBqXeBAJ2ptBXrBptv0wHrXiYwFojINRU2kPLK9T9FZjV4/MbDercXFmqQFPCP+pR6
MTFgT/NWyt/4NHC54R+huUHB6zV1NOEeISet4T6HVUtNH8tymk8bQiO2bhT9r2WaRjkQAZ8vDYiQ
AdacMHOZ7T7f0taCJxrwRm746B0PJf6YV1n9J0TYW95XXC4TxHQF034mrx1v44q4eKZvZPvqZd1K
OWDJ0LUYz4mJ1GrqKgC/1dms17aAEvJ6g/YHxiAdK7ZUn+sS6oG9aEeBMUFkLJ/L7QEPat5Al7PC
dixHc7iZUbLo/tfwnjhUxu3nsuLnIar4eQ4ldwIuIQ2oYa9FsQHlaBqWJLe2C9kL3ex46JnhiqQ3
ZI04VExYfy7nDoXm9yX8RalaIG3M2w9IGDutkuMZiE0P//+Palrq+inLT+uZytYmmbydvxT8TBWI
e+K31/dKP1XZ+qEH44bGIhEX402Asu0hG8tXGpjriCFHB3jJQsjvgX4FJOhOyrAMFo+abi6D0YgB
29Ts31wdWEPLsDxpA2zUN2Wnh04Y7lLIgIsh8hFrtNzBpn0LfVAQf2HvX6QOtmQSGQddQTn2WQVe
MqxYw85WaEpIq1XiyJqYvjJ0XoJMnpBvT7Gt+gMSoH312X8nSpxQqqXpBW4YTa1IPWl5xPY0xPda
N3msl9ZxESP4cO2YdDZ9xNP3g1SCiDP6LC0NVVPlLy9n+ozCpunzYmODSemTy8JTmed5GqBaae3V
bPa+Ac+jSfqyiZB2nRAM9Vf8RzFbIPsktxH5kL7LuFfC/kJyP0vTnH2Qfvugq1Jh0fEGF1VQVAPV
PdNvgTAm6TWaDE9BdsstjxFYHzzYOjasIWCrfDFh3yuoZMgZoOjDSylMfF6JAQ5HzaQCNjKKWTXJ
xzFEIBNnX5q1PKHAjq+03AtCulS6BQzzwIeErpw9AsWbQ3eastJ822HK9NGF2VMlx7cIZ0yBYZ+q
kOI/s/HXjAklzJppRCdBZc6RvWHgC6+DXg3Mrja++HX8/eVRss10yS0koUNBpjloLh4sGkmM8ufo
rk87FRBGQpBlMDlzQWtdqop60rN9I6H1E4z5XTd243Hm5td+BM4Iq9zUfK6gJ+AVYtQ9U1h9857i
qtZicMe7A1HB0+OvfGC0chAPNMaOKairF00Rk9ssLygk+0/bnipmb+RiStMmkFwzhefeaBdCIUfa
QBiVy1C+QtpNF5crfYrj3OtsUwHPNqw9Rn3TJRGAcxdCqNLhpEzlecFebmzj3Ef6JgOs1qbP6QXo
JgiM3zUYIeB0u9E6gDDglrrsb6pS+lEKdkvakSf5EKUZW1sFqtfBHZwQafZz9eDaJCgD8HKZ9ZNa
LBS5zH9iO6/AaoeBYlq3QWxbriNj2HDvS+goEGesirNnzFkIhxxXiy0Byq1eny/TLaNpgkx3wn57
Zr/bzANthEQv8Ww/BEGx9vb6ADZB/3fYcjHwdQZTh0SoZbWkmL1Cf54dsYpPEkTK3iJNr8UXeQ0S
evzPagIZ2aM37GCQ9Tr89lmLIoaodYkYojSvNLkSShdmVSBUApvtWlXdeOhrinc5VWt62zAesh/g
qauqJVExSh7y7ncmlmWxoAFYBuCOb/FmsYsa53fGcNYDHf19RYBvOlonXbIFI/QuTscnpSCqdTHh
q2SnMAW4lzmCP4rEppJ5St7vDf7vhdU0wDiWvpahYzrDLaALqLQqi4HC/L9wk3XUNGR+WNIB0hTV
cWUx2hC7jIzSsCo39ldAaC4QwOi+FrGklUs85zeRLzZ0bI5CMPzR38tI7ShOX/+pFJoPdmTGmWiR
FSO2Iu8lI6n1bj/xJNvTSv3j+QxqkQVWDPSuRsPIE+QIgFEDoxvuxBsGwC7lonqzaz75TfwvBBaC
qWfPjdZEFVpdaEVd1ywYiGQXc0T/rMgASoBOpiQObbBd1lNc8mxRcRxEOLnTAjERIGNr+KlcQy0V
alfIz+txklRphL2gAZfaJ9Cwr6CatGwTXigZbhJ1qu7B7OdDKNnzxjaL6hEwN9WUvKyMkPcWoXMh
eE0mzmOqRjXPzq4Aj1k5HHcGMqBMKiTRaKnqEENMeSxT8ATgDzg6aROLFSWjZjn/2sVlYgz9z4DJ
CIIbb98MS9QmLSqWOMTnq5EmWH+hKFT2G6LRht2wpEMbOLeXwBHoGH4zXXn9ObgWqDuX4GScPULJ
Z8uZP7bmkDxQeGJp5fxNM/74OKzr073iFRrNpiSTaZc5CkepQpkHmNqksUpKJXSTT6N/kCOzMgGq
ggeAyHJYVLqty+rtIb1ovLnkqFPBrnCPUCMidmS19vUgff2T584bxCEzqy1FFB34ZwYUw1vm/hco
qVavgSnvtpydPlstuZwvPtwQ8cgMJBAS4E4lNAaaOy1SSxrcdtbJ3Ssgd/6THQ2316mRx10NpS/Y
4IdIuhRC2DTa+E3snyC76wX3HyENgxe9kvsaZbtjRMgdPX5dxhwNan7dlQQmvRO+vXq+XX8Z79Kp
q2Yf/+8izUm6HS5lvgJ8HROtbxrk7EhkNMViH8SdW8e150zG8egfWZdFc28dG+2VaiyrYkBBZc7h
INK5zl6kw28B6/yzAST0hTEvnM2AFd64rgxzuO90Lhpa9O0nSIQa/c9Neu4N+b9HXgR4+fBZWqG4
JnzYu+4dF9DXCsicwXziKTf8coD8PRFM67p6Knvw/+7k8XaSLOGvLKt7aC6wvzeS42me/xJu8zV7
W21JGaV99F46ipmYh/oIGWU1diTSsk+czCQm5NWSO++zv5wt0NglvwppHbFB+09va1uwYFdXSe/u
WKwkmsw7uZEN8KCk9iFThcsJGrzSF7baj/VYsgXxeyjBgS/uxTVm23YbjnSwKtb+nnzKUymf2Oq+
FhuT/egryvtOZNcSaoc++0hH03fuucGq/WyKYcs8/yGYdwlm67p8Hha70ncY4UqhAV8BpdaY3eDp
AWGL4srBnczELZrgILLC25xdgbcdECOG9HEF43g6HZRQ4FR9SgCBcTFEq4VNuI7xegGbeoN299ia
+GP7g4lCGhZmehbZswG8s/yJvkuoxqHcPYUZYXOnqf9SQu1kXn3kgPr+a+MXKfvQA/CHV5hJ/vwY
G0GKmy81fDw7RInY+UzZ+UPzZtPFg0GoLbNJdH7cyLaDuY8ll5tKSMu/0k3pxb/KRZhe0W1L4Ag5
2a8SzNmg+NqSVSCNeKktzSMmD5UGwGUZd1pPzheQuvy0KhskhOrsRVu9VkEqQ4/GRMRkik9DbhoE
vx26B7E4aDfDcYShT7zhiOnJ/vHgOuVzaX5mnr79hrWuPuQVP5ZO6ixYBwoeNe1TzgYWRSNMWp+b
J9thPpnGe5KfYRNqCX1JgGTLG4hr1x2Wg/nNX1r4nugP/CG0FtKN7GzKJWX8HLBV+soJcc4fQhpk
NQzE5IsFKZXgU5PFvkKJE0Il28+BN0+vuES8jBClc9Enai3QpN5ZqMwW7CgAKhKc/ycTX81uwv2q
jkQYEPkywvsP3Y2DTgFxRYkrx76ajPPfMcseiV8/q2tKuHnqmCU0fin+1NaNHF76KHgYHG4DS+0E
54lQRxpIctL7Rmck65NFdFtk/vS2QuQ5L75EYlQfRT36DDVGLW+B5dlyPS4SdwuPN44UH6eWStaX
NwR0JVWgs8t8bOXKhdo1Kaf7y8yL7IWrDROn4UEKQzLfGevK6JvP8RoXnD0iyGjBWBR8rF/BSAwJ
GpbfBm7AEeL4zZW/iZUHndbdJxE+h0y1Nl7ixQ2/gD4pckzP7fObXHOp4aodD1LquY4Ggudk0Ad4
u4zlAHbfQQbar+LdA4UXdb/zWPOMk3+eFsRA5VsoAzSwindMzrVFKwMu45b5EDr+0IBf0e476PNW
2uaIGfbh6IrTytvHThMb530bJ2081EzNInch1sI4I22d2QVpsSLKrg4sSm0y3CbG+ac5pySf84SI
9PrEDx1946qh+rrI0CcNwwtOlAQ7AbE/xV6DyIrA98l8z7f0jnpFaTW1v+DsAXCjUvsfIr1GvPyJ
z1NKia/LqnLVrb7l9UrNCYlvZ7NytukUgvS48u9lIcu2x2iLnl2tG1IT2sSCg34HfNcJoiRrAzuB
eyQEy/y5PbzYcZ4mplR0wDs1PNoV4KbrP7YaRAFyGGO3DcL92vni3xpQx3HR1Xk+Gzpr71jzratX
WowrEKUpHrEU8w3kTAmKmt51MdMosgcKxePf8/lXKHSNvL3nBv0b2/cqsGTQDlVtLV9VAoHXz7HA
JVI8dlwul+TpKH9ELO/UiKHh9ZK0giLiDzgRDHu+gfb8OHXGmn3w3ge0ipDnX7gOuNQEA2AIw1Tn
3s8a2/CyAtomvGiOLEPtvxzfX9preioB9nMNKlcQ04k1NFMBplmyLl0q85DLpyG18PqsQ/aF90Ja
i9c6MJGt6MAYBuW7cgLTz3r0BVvV1GU0gSpsRnphnn9EFoudIQVcPhYUsaaCxE98IZbGLMKFWVoT
k9JEcP+D1cLigliLW2CaeV9bsMeOaMcZgFpIEjj1CtZMbDImVK0ySZY+GDXpqPorI+BQO0dFKbVk
GLa9eFPQs2ptdSvrkqy+v+TxqJS0NsqfNIfQFiDmTsdklSFY6rrKCnP/DoSMLpeVWB1ONpBjmukG
lh75MHMHipHMqQQFNVDN6Oc2hNxOvnxDiYsk7aGVfIR8CBRXRVW+m1Lvy63MvC6h7sbDreffgKYx
lMFs6MdSa6hbWS+cMLx087IZbQSupwsYc0Z+uyaVq1NxJcxAN4oP0Efc0RVnNN2tnWG/q8da7hiO
R9ok95rKsZ+bAxMn/NM9aPn8F9L8E23s+ix1n1Z/1jKtIX2NBtQMl3JIWqCdDFEdbwKLjvpZnrYL
GlvK59xMeV89/yfAFgEfHPILU5wWqAfUaCv3KnZZ9vr+mY7YvT2ciC3ldzQhMXtB2blpGjIc07fy
qRoX1Tj0l0cJ8QLch/inbsIvmYr4HCizoErKMtC613EYMmzHQ0e5say9k8+Uwd8vPWYdhh9OtYHa
2GYg0ER51+qkC+CVOcGFsLInSrQ8TYoiT9jFD4XYSaXVqv4LkEmLTyqbU5LX2ovzuLu4osDQEvmH
1ZIQRLwGcFOfIb1zSwIUMuznrLgLDsWW1pKPgscRo8dvJbGgDwe+NpvSLjZHVB2ZqvXpS/mUG4hw
sxSKydieTCt0V+18B9gKHd82x/rP/AkU+ny/zmEYOhzBxqJ8L1KRS37zlrXJexv3B89neoxB6YRp
skBRHFZ/dKC4TSfnpBD9yMyRV4eM6jxGWdcuLd0qD8zKwCKfHGuAP7z1kC8WP2/QofkxWNk+C+E0
fwdgrIXMI73qjwldFbf2FqMuIx3t7ZLKhyMd5HP8issX3d09qQ3WzienGyQ3xjqPg76zYKez2+kA
grittYQZideYsNgxM1vRJDbLsWhx4Vz0bRqILlrQTuEjmGTEVAbkrGJ/jbeR3ijw2aCIf/M8kSvi
n8aqYexM6nISGRdiFZtfkw4/RjgCfWg1Y04Y/WaLn5iMIMwckXu6djVcMltipkSij/wl3dba2UHz
j5daudl5vzKlCTaeIWbAEfCU03MzAQrX56njXUq2Zn4sfGgMamGeIyHtAA67zWvxL8EhRkaoI3KL
NMfrHEvGBxfHA/UWogEb3zTt1c+taJPDREsHIIEtYjD2gwdRdKyVmP+qC4l85+iXxUzYcFbFL//B
eefhhLld0bC4mZ+pPrt4c9+Ivy7jBtxjlWtZ97AwStB7Np1Zs8T1vhJSduFQw+tWEXLMZKX2s5jJ
P/vQ3VvTZahBayAYOXWn2FiP2rmqS/5b00s/TsS0SwtIKTJzo73PCxg7W5Sz1h8GNwWJNVJ7a2wm
2s6iBQ7lk4mzk6ARC5ukx7oK+pkdq9+LfNIxOI/dtgPJtI+yOECx1JU44bipBFz4vjNrz20ySdVM
4G/aDTX+r1xrmSeYVo0XLNIufnIL6cWYqB71zMiQKp5o4zmvXu/RjVor8dFIhvU4ZAXVuzLwu0y4
jdfkfCyEhJ8vabwISjammwvvhx3UpnYjaXyS67p+oBUuycUVvvg/5cTGWh9KQee447axPqG49pY2
u0jStmbC/O4r+dExcd4xldgi30ghw33pH2nEgdiQQCWbv4KFIP99fBIHAiRUJy8yHP6B8709+Rgi
ZwCYDD+VB/gWQIeO/Q167KgdVT9W+LmpZQL4kLZbLxMfr6MLxg3p9EcOQVq+fH21CIPaCHDJLi/U
JdfXE2a148q0r6o22R9XP6MGy9oPup5kYkQBw5OdEQoWqXgxe64eFkY04Nrrk/vfOH+mtoEb+A+I
wdl7Q7TnaFMKAvDjI6SnT/nXQYBPeeY/z7+jt47YgvR0THINlRpWzrIzLT4RNaAEK4QHCLaCZqkU
6aqPpOdX3h+TdaC7w7UoQwQprP/fSTMdC1BnVQBuHtQtdaEchm7O/Jnlvj24LA56MZJm+CXUIt0i
yjymhuC1nsNC5IXDgxB4pwvgK3JE0TjKQH70yC6Xp4dsJ53N9GiNesip2ILp7jd5nhP2PHeS+U2E
jGCulv48zFqWNcdkgpdNK02w0pGLDmdnhAPYB6ww3dxdIii3yOSVyEZavGodYcPYDWDQ5fhnVtND
PnE3OKgwXSGFQ/o6hIWGIS2YYvgqTUVRwV6cEvykIo47ZgP0r06ttxkePzBh9Y/Tewp4Sg3LM0wE
dJUOZQXBdUAD/XUmOeNU8zP4hLEeQ+tFlSZyhspvOwtdrBTJ9eFI/CN5lG5IAwkXr3ynR4j2Kgns
sM7+aChFqO7txTR1cp1kbFPJp9h1VaR6p//BNsJJ36tLGDZ7fojani8OaRATIVpRPJxNVXh+5OvW
bPEw7HtH6oLkw0HcespQjdowFpS3kfyjhMX7JwIlBqY12aLgypiKs+ETW822CYoQqBbLXJglXPoF
DvyQss7eCpt4zJ/CoYKHVHjAxWZvIVfzDNM1Cn0nKXGA+hDFK2tVzxIWQ77wQoT24LbMIqLn+CcM
Tdvy/gFbOUKdpv8VdymbAIvNbq5oF0OGhwBC3Ra1JJS+e7rGv6mAOpwrarL+d3qOFyabI5O16fWK
hmq7WR293L6d3VVVrq2D3J0USDekfFaUqruCnxBGnmEdlJgYvUDwDW8FA6sxJPizv5tVSRUi+1yz
2kmFvPnXFzVeJxOIRvpt98Pu8JPlztsgDmHVJ7mkKgsIhI/of+deZIUCd8EcvHKwt3L2N3SfC1FB
f97gczITodIoJfeWiIM7hlrGi0ispvVyK2VFsExIXZ36itrquHSW5NoOspvX+ihIUx8WGyWPzBtY
OBzsXUhdyERguuiNTtrPTPKHVYeis7dOE0PBG7w3cKBXMffmtKaBCZYTEccWldZKuC3IgkX9huHP
cjMfOtjnD6WsBPng7f4k3fwm2Y2fMOee1K6XO2BWSBIF3SqergnwUg8EhGeqWTfnhpenYbHTe9U/
8hiQOIJLK++vl5oI5CztqlNPPR3HfA82XDBKe+nwvSnkVXveSMgFyEFHaMeYpAivQbf8RBBhJsaz
9t7dkcwweerunIFAhRbbTTzfKcGYOFzj7lU7szIWO7fNooYiu6G+qNs8YENbHgRlfQON4eZYaGU/
ak0nvSZzmwH9XoEHMyeFPtAvVCGku8kWcRHQ5gQsmcbFXW5wkMyWytAnU38Y4IQdfqMcLnqK3tv9
WOHGAcK7Sfa0KWCxocjmoZfyGtjP00UWAVk5DqtHwY4XSX6uM0vBg6+VrChE5Fk/t/Ovnj0MEoCl
zkpKJbUtJ9euny2QoH0ySfgzbQlLA4Ifn15X7oMNxocFpbgzQ1vCYKxItCQHh91kP+jnRhK4wz0z
ANMXzmJrd64Z2IX9PF+5wJkwbu5WUP9lGg2Of0vl4IqKkz3glm639XQ7Np4fYP9R0GC8LU8Al04D
Cl8jkIx5Dd6DXhMiZmylpgPws+DlWT9xUhvoWWEjB9EKtwEVwbmENwTQtD835FLDCel/KVmawFlH
9Fq6PmpVlRrfdu3oa0R3nHKIlifQUUK++Gfi5DgOwDq5+Hw+KYPuK27e/Xz46cYN7LjuQge/Irvd
loyr2+kxFEM0ySmGjauNZuJrCVkyB9yhp8I4PCCM7l5rRoYpOS+mAAf491Q2CdTI00toI0x6eWYu
oq6gh0PJwhLgYZrmEdoEvlEGRmOCu1k/LvqlPC/50uwiXxw18g1jG4oHdvRxW+4gU8kpVqumcsJW
cEWtJKshPnriPT3aRL6xY0EQ6B/jLN4i42nC6rf38MfqVmkXpWK7qW9H2aUskyNqUABZ0PRFoqDZ
6PL7luQBCkZcprW17wjA97liKMEoD6WtD+Iy7Q+UjVTv1xuRFG8/pySq2IzG6+DDudI8uDeKX5TT
XY5hDzeErjyQvm6AM9Ml3M/eiaQaDtNNcHvJiVFJQXTN4rYXqM4fJZm+THHdgewI/iRzCE72hGZ8
n6eEgr/4eeVHD4KwMHJ2v+orZbDGaV0RTYcTP76Wdad8REKxQM2N/C8VE8iofeCwUcswMxXouE9t
2/SshrQxFAqp/PSDs8jAKk1xmkogStzyoGl+QMU6mQ3CM6ooDNbWgMnP/Y3l1bmZ+o3yWcvrFdRh
vARsphqdK++vIo/+qPNh3d+PGixwNugYzgaS7Qoyy2OAxvcsa/Azzv/KxPIOypaG3Z09vOaiIYI0
yJKQ80uDdhoQ/lXhZlihpUbf0egRm7speN3pdSsjGG1x52jhjosGAvQWGn0XlP7icGrcerL54uOs
VrpdQlgjvclOo1nx/04hLybSkXMD2jtlbE1MRgozoGBs8j4l4Zvpf/NqaTX6b9XCdbtz/haNor2M
z4lw9DEf74M07wkVM4yCLRkjBS6Jxcot/aZ/jXaCHjSuSTg5pzyB289Mp8qq92u2jfVflUQ/OVmA
EfomCgV4LHkYBHbP822gHuAAhCfDBoSW+zI25kWIupT4gP2Bl6+NPNlyug/GeU3HjwzN5mVZhrUP
lskRa6Sa15YVHEi+0hw/cwF0Y9R06WM1i7qF2uCt08/wURsLHjLE1/0aB3Gi2EQZ5+omprarX8i1
0Ak+JfVwmY5yrsPSiG2teN27a4/du4H5GIvjj5NQkbGw7yRYFLY5UIojko5W/wJhPa7tLaIT7zGD
OAJQIfo2cZWE47nOMgDq2E2os0scoJhwZDe92DMaICnW6lYFS2AknE/IXILxXR2rK7B8TnAeW270
O1eESKB+tDHeQf5gym10W8X1rtV6YwMnKJZuIS4wmhi4RB+PvP6SofhYDcNO0nJmwZnRo/tcD8fj
5rqRrcaJ3fwdZeFgr4xmYbZgUxgsXZhaYzjtpfDtiuMMODMjVJCdKQ/t716A9j+rKk7rE9gTlB1e
mVtMwGT9xDNtPoPel5qMQY6+sSIZtBv/xzObTJyayrLPUu6sVkeov/pr1gi+ONEK2vN++aO6JW5u
DJhI3NQpZqyRzauyuog6hf9Dmqvrp2CjuBds7bV7CUj/CUs6i2hx5EmBmTvvwadKDLPjJHtdoJwI
WkqT3psiee4Gyz7Ok38SMiWNjdbFQFRWaCT3TLfjnMMGTkFeMKa4kC/aB5UYfs7sHCdsTWcCzC95
c3y+qq9Z8z5fe82jV/myWtjVnsRzZZiL/O/Z/Nicr/9ueiXlkRJyZzIJEBKdSD24kloqURa/ANka
n2/DE3VO+5yoDGUtNHWEDlgkIfwgC9bh1fcWSltOYWZDdjlnknJUgpmJautOwK5/h0yEy17IJFpf
dwVfCWbQdLhK7FIzurcaH+LiXDjGdRHALtAh9lCRtaRHlvWCVXFHKBUPRCfyyFnRY0rEKZpapDhf
IcpzzAKlwr6eBvysHskx5WJJBZAkUddjXd/w3qAihHbvRkEntLYNjlovgoVkz2TH0WoPqujTQxBI
03Mi5DuPYALh6rWDwlc+4YdpWkKMr2px4136emGUcpp5uYg4W5z8je/JA/bBHRENXG3wy5UyA3W+
dDKaCm5yN2ANZFpiFT5/Zk4CADR91Ncgpnagb+at21Z3Y0pXUEt8GzFPeUkgdDVfwKQG3K4agr0F
D85tpWyz1HnyrYkegNFh3rY6TbyVeR0iQFOX9jma8M13bRVEcIiFznpPYk07RJP2jfM13GcOJXsx
cbCVM3EWvQb/A3wsWewXAlZ/Q+AahfeWz/6NzIRWV34MYfxPFYtDzsgHpHgBg3sK0T/HpZgg0pNN
VvuYOuhcomhJvB7/iTwdA7gJqPZA1XGeXYPOoKZrctdpaiC59BgyA+C0GuQGQAoQMrHZnPeNrjgI
CmOpjd/UJ6AVSVRUpCYZkiYjxUN+jFpGuAt++mcln5rd2j8JzCthcZOCWZjmxSGWTkwBjjfa+waB
OhWF2WWTAkKJyNDN0ASmCiZDe7cVU57xAo/VYEbN4neThOMbExkvsv/rB2LiWeLlB2xjFFuF0wQM
7V2+dyasmUEtrNmsGK4GXAkf6UEqH4F2hsHDMGoMW/NPsNMrFqJMLPyztgRuXrTkqJHHGyLcGuv2
xiS6y+ZE97ZPJb+9Qhzgkn9foV9AQB61NJljOAZHy+9Pk3KEPOwsNDfEtuzPxGQSkncrp7U2TE6x
2E8RLV4L2w4xIBzDtIlPisIG1uQwEDoezpit6bkjqc0S0tlShufpAstQq3OGZo+v+dlBkBRS/8/c
QuGCEXHIkHj+PcnHGubkt2CLkFzGD2M4DhSApLTipAn9Ki0B2o1Qu1DTjJb9JUQJ2zRZAI5uJOdu
VV8EVxcceVc7iWZL0iYMgwrCpwR/Rb2GyqbW5ObyPW9idfRbkQLnAsBfdAoukbXJt5Cj6LSY7EtM
rmdXMT+TwpLeJPgyLVl3XOzy+dRklZ/I0eNTPDGzFlGcxROWxo9CwymwPI9yRVWowUSAy/7tezXm
k2A6aAg6inU4SKz6HnymQvoeKHup32Al00YQKt41PRPRz8F0gzMBOvtnIiLCGPzr3g8MnT3WdOsj
9cpG88apH3ID59eoSj/1tY5tufJdLaOZNQIcheZFwD5O2bOnO1K7TPXaapi/KCrLcDSKztxv0aCo
rYX1NFEumIq5UbTzIfCYRzHsDUjPTwx6D4HxY8Z6D+/3PZwee8zSJXM2Tqt9+Ju8HDTfHlTJu4hf
nJXwByeHQuWIDaPP/WP5TgriiFUthJJvLOMtZE70R4jGX8TNL/WcxFcZmyN1zVIKjQhra6u7Bzs/
K7FNXpPs/BqOW/RXc/awPoO733+16ACGjGNy5o8TjvigMNZIbrzpyYPaCQ0fpcYoTIuVlhPajLL+
T/w1NTC253CNbl+yK32ehyOwSiostnlG3H+bqqRZJfYrcQbxKatyO4mLLdUHfkmcUFCSGKNpVroj
MfC/cv8OXXLqeHf/X6KukYBDV8UqS0SWqYmksU2uQtL5mHidkfLa3+wKU1tlLRukQKARCmdrN9LZ
GmL2eB2y+Zd/THoGr7zUP1z9XVGLDmZTUMBir5IDHKNdzqMudTcIWvbyE+IputGZ4MxM7RGfhgEu
bOD5yM6Nu5J48c4X/UFweAjbb5KrpUdHo7+L8dbqqITTi84CceSvkGW9OuO0Q7zvwB2pVOL3b0+L
XLcB6wSSIm95jv3NpwgeFKTKobSmj9knBAzylN1VCQ8QXPQiAe4YZAcRV6mmm7yW6ejFl4qgO46U
p8hzc1fIWU8lTDuRwJTW8CCAUO5m166IAcKAuDXZ3SY9kpUY01yqk9fU05wcQNbJlRGvZiH8MWjU
1do+Db4vly46eKppMjkIMw5pxdkpTUbP+dvxCacmdcU8OvGwxAO68F9miT/lRcNAqLkHpz61hUBb
tfON3yHeYe1TNAH6nQDYAWPabhAxCkXY+kqqcvxOAGNt5a1tHKWY872ZV5ffnxd6MTwAXKUo1Nrl
2ZaKsS3aWwB5EeLz0QAYxGzBeC34kz7Kr/rnyj+uV5YhEA3LpMf/wDY8h5+Pk5hNNsJkyTM1d/Ud
vMFXjTMO5qmNsF5t3hWvD6qK3S1VKC6XOl2fWNq2RAAQ+OOEyzElOvbtPiORovlcM95fjHThHZwQ
zi3knrgSMNPpcHz73FM6bhmX/J99HydtNClixRl71Z1+k+pcS3G5YC5gutLZ/t6q852MoKdXMBDe
RUjxqN1zX6wUz0El7CFodLSswnN3k73FdhM1jfriTQV8FbxhU9VxCh6MoroozxoQd3yW7FPF9Xjm
rBG0+JkNEX/lGEA2qBJQTXm20LUK+U72w9ZDeF2F62Ykwwf+UIlyzpmdjAw0hWZam8zgLa35gp3a
SZMpzAnV5TG4vlroXyGK98EOozMadEJTQCxLFvPYdz52axagXCLYxxQg2KdF34pW3N3iKZm9oyCW
hmRXOsbxD97n+U7GD2/FfCSmzho2UXyaxoCh4Nh6mkscxzgiJZsGT0PzZ8n5gZBdk+KQmpQJ+hvC
KZnU8mNQLMKEj94inUj12tsFVXUDMrTpZpmyC3w2cnb3OfZDHwPmffqLmYPtAXxwQD9WVtnfFh2p
63F1Uaok0odcJBtj36watiudchS3LF6n8AYRmtB0K7u3u+KdDYYhxLjzn/oUOzVEhznIpFj3Js9u
fawJrrM/Lmg716ztn6y1M366e1r+38enpqeWXNan4fd/MBWVPErkXrL5YrIvZBQB3tY4oDUtdKth
g7yfDU64XR1jmlkZlaOke5MMdiHdmU5+YysbIAMg3qFWJ+FO9KLJL13r2OrUygqHgZEJSzBYZ8xE
n6Z8XTDCpXDGJzM6wdXvHOsGFpkXBB8XkIkFDHT269ZLB4sPwCx7H3BdzxRuA6iEF/oV9K8srkLR
d5WuKVqah41Gnc13vfAEKrPehjlIti5bepuCpP+tBZysThUwGikAupk0st+owIG3+1yGhCLAxixn
UyqAJQjZL10jwDftg1lounDXpvi610sjKp0vkblEr6E793BaaUCyVQoB9rTH05oS9muq/aFEx4+y
4dNfHghnt8mLIVAtvkVxsloEZsCW2tX8d7KA61nyKaWysS3qbRaBCMf6iZyfeednkH3W7q1VxSxn
mi17N9bTL/VLRJneTekMOzS/M0sktB7bQ3YcxrKMNuQnyZ6XQi2B63j+rfL1JVXpcQIWmNIQgg8p
5mqTmJA+/th0V2dII1FSNw0k87zOatLdgSkpKS1ms/LU7T1E6u1SbEIodXv1j5YzhxXXZaaWMvdx
JWrP4npRERtOG5uPnc9xvVak20twPs6w4iO0MII67TBImlsQDf7FgU0Gl9h7I93WTZvKI8O8zkJd
66i2h3BL7QC1YC8311/huRel0oWviUf50+HLnNPWOiiPsmtB4dj8yzNXB4xhXEoEa6AVkJtgFWkK
srhf25VRJgT3jwQONQQXpyizY2JaOHg32Bgdn5J3oHWtEQBx6IyYXif2+luih8m/tyxA59PJpF68
Tr59lVCyx/jh0bxZvIbN9xdKv2Nubp0S04xpKWSwm2EK8hirAO2qmcCD+aOYloOcp1K2BLLUYjXj
LHETXnqIfjNUTDutet0fit82yYJpQLnOAd0K4xM/mGfmzMd3l/30701yVKB5kORwbsIhH+xf1Wpv
DiJ/OdurRI1ZlWdswXDH/iJJXdAizQ2qHmsboDVER4HF/ItpAB9pBIVDvvSq12Eo90WcFLDY9oQ8
kV4A2Vx+BJdDhOzQfuKTjwofLZBMmihHxoTXSK2xS4dKjdfAFYfXAWTMu14F0CN80LhIM8B+su8A
LWlRaUbRIm5EdDVjy95dpsNmpCV9fJjXvUYFxZMzClXpyZK1X9kEpi8W0y3xxT+ntCfAxfbpFM4v
41WbL724e7pTTCzWRuqY/nRYEENQbWKb9exiAukcOpmvNUMt2jkDYaU/MbqHjQ8Kt++f29cPNYBm
ZpLPCPk86LKSlqwVfkzRsYFAF/BtYw8eULQHfJE0fGW5IS09snkrUO3felMFhHeaOBwRIAeYVqFx
JjBs8OA8/YLwGJW5wEvMi4NmGl26D7VILBJjH2lj62iOLf3bls27/jT/04SaVH/u6nZMpmqt4Hr0
t+8FVs0ifnEHJ7ThriZMOzEod7XIb9Eh1k/Qfls6fMzXbsSe8lS/lUAUac8tKCkATCMUah/pbaEF
xy9tqKZ35Fmrs1hvFFSoqyLw3qmXb1JanGBRJanGLnJzFcLW2rceiVLyEh2M8VfCedEzbL6vw50s
7AgAn1fkEl12l2+6dbN826TYpvjZOXCyEOQQB+rOFNw4hwHuGniGWKccFQ3UTB5Wa3O58lRl30Gc
8KfBZwhrNPzNKR/CX/597DyMzjYf8WjeNi+wrgK2+Bc9q/hBb5f26x7vwzmo56mynFF5NlSvrTZO
/aWI8tzlkEq1vH49cl7sz1opPf6KvWdYqV8ZiDqcoxF2WTUCyqujI17pmMw3LTtBTtE/tmEOC9v4
io6AfHUTwZH783e40hCaypVE0bUNRcDuB1SQpeSKQABR7DibbiBGa2oEZLx1elpTSrcYx0MZwSAL
tFs3uRTWqDrW9d34Efpi8u0JoqmP3pYiLjz6M423rtYNf7JfXHkppLt07vm7qGXpm8iFGKjbSP9f
weENWwt22PkT17QXiwv9R2xaOD5w05r7ebUQSwoGHw4Uxv9COIpWwB+F122DBRG9Pyi6P3KeHZdZ
AebGuz0HXv0++BHEGQ6Au78CMAyHvpAcb5xN67Cy57Sn/6pSZ6YlP6J+sUFi320xF/qu6dzII6lj
BKdDzUEg5tzd1CL7P2sgWPKgI+NEhGQ2BOcu7ztN6vSsI8pKbv62xmujUGKrX4zd2JP0EjjWpSTC
cpAItipOZ+p3jDMyEOFRkevL0CamArkDwqpVwgJ9H0jKhCeADWZCLG4hZshebGcoa3d09BfKRMvg
xb1Uf250iGAme6Cy6rzb1RGgFeaxEiRxAhdEKxGwocc3rj57iBqhmRp2k8Y6EbCAyCMdAw2KJZiU
GdFhIscIl6xCm9EjMExEGyVPFDGddOnEcyCY2stcuk+AaDDFqL3s1l9Oea0Cf2K9ushbyVuIFNB6
rjDddlOE5bzkqEAXARJNRxRmjmmk42IDDecifBp70Woq1O8Tf05CI/bm8EOeL/PsF4BIFn0YVsp7
g09mDkpESS0nrotYi8t4u30Z+HO8VzQaD6Z910aSIFujkXKIVpomOCDmNLMjVPW7fnGwUieTdHXU
vOG1kddyafEUb1XsMiNd1gj1xFA58JFUmRav2Wv0LsgVkclB7xnfTBgq+SAjIXxH4pZAe+W3z9qX
gYw7rrJuIL67uHHO4/ppb+ncihRjwf+5e5vwNR4kHm3feT3pIbQSzBEuF2t7GlNoMnXCOVH9HOeY
pOT1MaQrlwRtmZ+1MB6QisrrPeQogHWmVpvsbMYWWu593BV4D4hBZG316BFSxHBPewKJRmTavWjE
BvBUM5SPHXXLyktwoxlMQ14e9FDK3KC6wDgHQprRFzjIsZ2K6vZrNX4lcJsQvy1OtXRKUrbSiZMt
Qxka8kKFinVBAqQ7K0LAHn5v/OxMnIJjmZfgwBOOD5wwmzjmtUEZHb6mWyIPsIjpIYRxQ40ZDhwH
79LadIczoF3ro6RPw+ZkpldlACTescilxNtON8UAHtMZ+lnYXuqWeImZ2wjOuehnJIKZZmGKjYMN
ijueCU9ZbgyctZMtejoFONb1/oju56TkpmeV1s/HlCX5tzWLF4eyptrOk+pCODfO+2JnFA+KRFrB
B8a7SBi3j1qKcr/GPV+oALJd9CP+j26FLw0bphD80U60JVxJ1lgtIWIMhHiKqRVfLuKYtaSfdKQZ
fc6FOJgKN8MK9hIBsI8tPdwDp/ckYUG/9koUqyxE9FjSFOZUP8ooQhzaUtaQMfK8h69CwAQLT/gC
GDjCvog50cboJusqY31uh33W9LeelznXqBbt58YY1A4z9ZqshpDCkeNGfe0o7zGGs8v5p8Jf+DN1
Vqez53agIpBTP5u3OruIHUv5ErDpRcYj3N0Ge2GmRmca4Yj6gUaS5HG5+TizEM2abRoNoJh4n5Dp
ocsQNGC4TVRHpcvfd5HWswrnT8aGAs6XDPXL06BgFtomqII5YbB04wszhKOGBssAo6+3Sapxdj6+
7WnfWSp/UMXqP6xLxZZc9bWY4gACDGkDvMV2DsFU7Sxi8eYIZxBBJ0jX0W/5HoCKYIv4NQ4P9JEA
4y6uFqfYO4CSs4ntlDVcOr55qGRCDTGj+eZ6T6H8sgG34q73UzyYHstBrm5s6HYwjKAUwhuwF5jn
V6NkQI18fumy31j3Qnv5T3tW2Be2xF9wxt781ra1qB/M3e8+1Ct8J6/pKOMqfr6lpqUT7Gdf8PRP
qAHcMFNs0joN5OmXd6MyXVNjoi6r5g8sL/yopLBZsbjNgDdK3aCO4HD2ThB7+X6UXqFeV4QztSq0
VAWb2M1Z7Ya9+9JOo2gNPCuMPOtQRSoiX5xRkw9uEU/romRnp/2VEsTyQLUwu33YTzSCEEO2Pj41
ozruiNIALllOF9+7CXtjN72Ropxv+w0oswxER4/stSMr4zigIePUw64SCcrtaNSCDeFQuG/TDU1z
mefpkzzIq60UR/fbDv6LmCmGlnTqkbmof6TVohRWjlGgKmnqUOiVJhTtrpQiCXFQcAsd/Xv0XCLh
qdHH1Hm0SaGWf5OxusERjj3QA7lMhFpSJy1TY53deIgTxStTaA02Qb5tABdjnV55gQmcF5ixQzDI
TTAn85oVA6uP4lfVsTRPK3UpjyArgh7C44q9CYk+w3+1cb/sbXjpDgbXy+LIq4ZJUfIdMXOOgGCV
Ocr2C0r0a0USKlE+VzU6nQp2hdEpNcvMU0QTgsSSd03gz1PcgrjVna1pVDlLS5SumLO867QnygF9
fbhzTcVpXWmfsSy7DHi+kLRdqExUfxZEMdBD9ogkP76DABkHtyadHb6a9c6gHc21SXQIhTr/SR0J
d/djj5r3Mc1fhJzOQHBLWGbNUEIBQGnNGDlk1elHabPlipvHGY5FbBt7lido2Xyxp9zNV2ZqE+/F
AvKKmeN1dS2CNKOyhw/BB/jgG8qZ5NEYBS6qEjAS3YThoDyLdgep87FfFXsAx9uKEVzr1Cyst6yR
mhHWRVrxtB07Vk9r6Os8q8jNm/DkNxVovUknruyI+393cKgxdKCn1Rbk/uflR39eSrIWrwhaTDZo
Bg3mgEN1/nNmJPYYswKU0a5MzDZnuhv3WfUuB6+Pg8rNMXKBOyJzzsSS/VMyUp0+VZ/vVoeveTaZ
obN4pJdc3SvXZ46eXpb37R9GTOocM5GmXigrbGSZr8cF8pIiRH2vZFuSoaHrKM0hhgFN6WouYxuP
n8Ivo5DvFZZuecP+znxZNp2RgC0KpiG0TBwrI0GSWS2wcA8URXGALfLQQ7bRqRnFDGc0YvBrRQjw
TnV6GYdubOyLWlq3QVm6P+/W23F3zoJOgBEoRW3eQhEDfMAfB2bkG3j4N0ndtPFs1vpDqWc83afJ
7p+xu6mLdLDFVsB+do8OHXeUssFJKIvTkT5oAem1dQhtYUMHPXEPoAWS9C1bpbq480MeWYdGxsI3
yBVzvNQAAw+YdHxrLGsmWAriP9A+YrmjrQfnCvo9dz44JtGRdellq+C01dXHsCQToyvpSOuG0lfT
IUPYpwcBsqTi3Lh/PzU1rzImtTZ3WTi1BLvH8u4zuboI9ZgoLNdnO0XzGRrvFvBFz8pl/RDGIYhn
EVUFzGVELxGAzAPl5Ont1GTy9ecxP+mlKQFZ0AaF2jU64QU7IgYjQiD/yRQ8W51IAWsr8MATUJcE
vflHPWnm7E+814WdRWrCqqRs1p7sL2kodz/ugaUQn1gijZweJbvO2cx0/aiFVYLWqRxKldiE0Vit
EEiUW4F2s5dlt0kr/4hwXRa7tHInykW9Wu2VRnOF8RgHKC/ywponFg9wrlpjWDMUnAm9AXr2uQBw
u/qA/kB+JNqmQQ5Iz5YqUgUmCmCcXLBTKEXAH/UvpsG41OzbiiEnBqQqn8sXIg98cwmED+TsOVYe
h+lf3KstoDKrwBsECX0Uk8szrMzpd0hRIbj0bZdxLVcNd9j/l+9Q6pe3r68rOUHXeB57ZVzPyszK
edhrcMRCxBCfkCcoeBVqjDp3CwxEacSno4kdcwvARV6E2TXbjKnflujz5V3mTnumYpDTy+2hro1/
797+FXpYO4AdPdna/eB9+cK1VqWina7h3TPjeTJ+mETJ80CFUJoP0UPTR91/GzCLGcQNKltZ+iir
gz2AE4LZoVnkanGPiGzhniyWIJx4Uycwz1swucnYKcH3EpD7e2QaorR/O5GLZedzm+Ajw3voYwgs
VVQNvKxJFf+UD9tHOgKwCrPFFrVVB48Tf2TXwFTiSH4q7+3cesuPA5QRirMR+ZQRRzK/nPmI+v39
BCd/xdZkIFu39QcckwexbEfGdEh83Cw5tvN99dnpj5/xnV4LciRBuMZdNYkpKPbMMntchNUfck5w
A8VTKwaTEToTsE1B1A4KkxQgYYEIUvUtQN27WunJOtBmzuOJexBTqen0s5AMJSa9GzihywdERyYY
Dd96Y6PQWM0w0jcCGwIbYGB5vMpI4OTyusk4RuouY81FIKRDf5ZOV0cOkyszxfn4OAw+n0sQJ6jK
R4gBmybfKu/vLVwa8f9XDU/LV3X0HVZqfuB8IXsQa91D+HWbHyG9hYRB3X56JnL+SDL8pFvSjGMJ
MiY+9aWZkgtMZ5Kg9006aN4PjSkNPEaadw5dTqhwuESa7e4lE/f/RfLYyzmJ1QCjL37Sv8n6R8E7
6EMYBKJNfg24CIH2P0Q+vWmHzvm+HUVd9vNMYBLeQu60FqFiTVrNAVq2vtK7YWTUz7W3IePb8dsF
XmcYskcan6WSdXjYLFtsNiVCDuUasMl9kcpBjQYMqUA7X5s1NN7O2NKhpy8dwndPwBqTzekbC/Ix
loNwOw6jSTp/ZHIsrLQXcrEyx8mGBpWB2fxtmeqW2cKEQJhRLGRIFmw2LJdztJcP6N1Mtbmc3nnn
w+UptsUyRpxn4CJP5lbBZFGTP8lLrUFPnGTODtnRWiDFNU2+2yyy5Mh3Bcs9q73al07MevVB0kw7
hdALXu+sq5xkgFjLX4z6+80e2BjXZtPq3+xR9NLhRcFBvTxPRnjCWGLKXlRWsnW3mWrxlqjFY47Z
j6usX7Dq7tU+uIZp/Zox/uCTclo2vzKEG8V7bz/dgPCSmOt1DFjLdYtTS/LP4MJVAj8S4r4+K/WV
beAuyIBt/ZXsHrT0WgLkmau3TlozFzbMGM7x+S/8jfmr5RLx2L47/SwF8zrAkI/yVysjiSKj+DIu
VcTVTAivcnmMXitAnvgR/vUbWpg5eXl0VCe8nlxmrWWymbBzng0ghtSDsLZqh1jJIiN5CT2S1fKH
rXr5aTym88FC1eqAhLB1v6yvq0J+jjv1pQ/sMAAJAmuZ2Y1AEXxfk2pXMHdUS35nGGZ3RumLGYmR
VEq1oo15GayfmJ2BoJEnRGlWuEpo7PoYJEFKOQXMYCSimVheE0yK5cCrdEGLAB6Mnh80c7IhF+Xp
QCqlQhLHneUl8PVN5ohK7UKlvwoql0crQCp7U12brYP2Xge4/3//PJBtPbDAinWwc+2Sfi0ipB62
oKL2AKCeQZz51VlVTd0x2Oc6mFQWxY5V4Sm3jIpcSaqXanJAfcKOTEeFaentzWMF7xf1Jq/O+eEu
pSe3vtAZfrH+smU6Yv6Webd4brpXWkYAqC6c7WpPzMqvNQgU/HST4OzJJf0p12Vwy9lzo+GNvLOG
dK+OyHl5AEI33VxIvW1JEismukIuq8d+jcKVkHzGu5rHzhdeAdDCv9z4c59V3YX1d2h7c91TVpZE
2EGbPixEdbg5d5slH9bUFsUJY+RSXy0gAygvBZWFSTwkMAZ2sqsZ6NH4CtpkMfsPPXpz93TtAi6u
4xqfFMEOERmhuQiwH1WAQpt7p5KWAHkApFjCL2Gji35utMvhLjn5QO0OK0eeAdTDWxlWmBJCt3Ec
xUpQArsi69ypbwPZymuOsjpwWmyXR/qBCXDm5JJ9NdWzmOUcMVsW/gfQynBeFyQWpvlqyRDSgSf0
vyVHOvn81dV925qXKXa2qSaIYa4ZwhtN5P8+ZgG40n4otwDTAHoHMVB2TVZCWt3s9WwvCPi/4vLO
zkNhCF+MPZrdkFvhyXdaMqHs8k4XgXkm/BQjMM/GM1YIPkCrKRpUd/cUIjir634T0oXIbMk5co4e
LxJDIXc7K9XVxkIwuZGMN3h2+bWqnJIwCcgDSEm5xYTdp7EwB+qe4HZddm7MCpsny2NuI0Ez98Ca
ZHV6Zt6b6STRFMLUbNsLTLSagE5lOL3IVEy/6rN15VoIE+YXHDZNVR+j42q363d7r+2sK89E71nE
JLZkttYL07h76SsvYBewdg1LEDsL53+XTgFv3HSHfdxBSAUr9XVuDw9RMCiR21803bW33trFkeSm
TrXbRO61mYRBFPGaanaE+4i87bzrOGn80/bQqXdqCvslBQHEo4wUQcGkkmbSC6f47aodzrEdZ3IO
daTOfUz1aujBbMwu5GSeO2+xrD5w0gC8Jyb2DYqDW0dGWMK3IhOWHBV8ZX0zoEJCh7hnEjnzhLvo
bsOSnqjRCpz2BieuzHU33MBrp2w2/Qd5/o58oI6QhCx5yxpJJ+MWwV4yPwathdBWCVKFbxN9Mdx7
WdPZaOXBD3cDsqNCWy3EKbQs0PIpGZv4clv2GaHq91BbeoP07On3cjQLvirWkZpnMfjGn2sPRStL
G0Ymhpku3UiyKJ7dcbmEH8mcZvjYkabgqNWKFCkx4VjzQZXNSOJOF49vM9UmhMk1PR6KsyaV1qQo
59cyHIdx0Z72PIXEnGbIGak0yxI3Dd7Iig0Yg3WlyfiSYaKlwZ2SMDUq8t974NzOTDlU0xWHdnTH
ahw4qZCDHtcFGAroaJPCrJ4z6ThGh8zd4LekAFsMrVKE5xVwF9Gzl52pGm2AE+2in/YoypnStqZl
OMW+60lTkZ4C8OkeZuEhEJdL6V95VlP6u3rKg9d6pKJdKS/zIBXt8eLbcRAD/mujMLQfbpVn648g
M0w7lET6tI/+wgYkSsDExyDjUW5B0BZzuhVawVLvyC18u3cqZNRQTwGXOicxdBPFe8qnBiKfqBVh
R9T21TaE8V4NYkpvoanqxdzVYRQ/OhLY6M7k2jpcuXMl+Hqg6D4Qkguu294eImxdWDOkVSUV/U6i
p2l822xgVFlRr0bPem/GWSPiPkZRuW1gKc0PxDNIt0yb6MM6o/tlUdDilSEV/biWU5mab2kcpfaj
xaL2flnr/A14ujMu9liek7taW8O6sjPUdUu7Ty+KwlLT6SUjzjEjkH5WMaTwwlVzu22QubpSRbFx
QFtF1FJNsSRYONlWPbeE/nI8NEUK5TITkL6yaFyROihSxnL45jaq0WDF7MvPABYzvcgTvQ7NMeIA
uuHnRNwqkjMgxqxcr857TFb+iwi6ELZDwVz1VoX7N0XmlrmqIhf1WJxai1CDZUHG9tUAOGWZXceL
A7o8bKhxiI6d34fhlcHiy4HjfyqzA6Zwbbj4ngI8Cdc98C2e+2pbUEdaOAMs2m4mAtbH/yV3yGPg
p4qG9wu5Rsxe8yEUgU9UBry1h+px0YjLpqgjSlH7aZIwSr+JoeWxl4oUI/wY5PGa0pwGWQrI7epg
7v7niSk0LkNYmYZes5ImtjmA0ZJKGeffHKhBHv4s1gqVYQD1YsuV3wWwYvFoNaPRjNLa9I5VpEFR
uBBPh7zvXlMBOHmDV12l34ty5mpyulrddp5nFMVx0Vqy2vpDwYBf6KOFnfWrzt0ES2KzoWE+lOmk
l309yxRJl3U35TN7rDXlEa6toZ5pQvdqLSFWva5x4vhGLeaFutjS0U/TL3PUHX9TdY99H93USbZQ
/texdEvWngdeoN8lr37hwRmmpt6ejfy4IPmlRh4rAMUEVjAUE1y/tQJI0oI8x5sjMlyXevzGdUtk
GDcYfeb3ypHMw6Zo5G/NZCQle/1ywHJoLzB82jmJmjPNehciGWEIPKgymdkWkPSf9qwrPDp0jn77
btGGo1+W7C3LYoz4b0drekGwsuIA1fpMj41FSLxM4113MAMfdeZ418zRs183C7F1h7/fmvikp9BI
cL1bz2jJMU1qwplwy2JW4Zv8o+JSfF82ZpmA/qZJyWnZGpk+9pDjkn7lOfMSkYAhbfIha5T42i4A
/m/RA3HS7ZW+UkmCRDoj0w0C6OsIyJu8hrKex/DlICFb9+4ZmNxKhZA2LK3Uy6MJ/ijMC/HaJSCt
GCc4/mhal1k6R0GWIV0f6Fyr8DvOAoRoZkgGsVB5KCn9b9e0k59d9tgA2XE+/BviJH5pvWlvG30h
xX/hvOnV7zgy05XaOji8EH0/iqLB+4Qf9P914a9xH8BIO2wkKVX2EJ1t8CaMUaEAH/e86tr2WFqp
6BK0VQCGV/thXGdh96Rc7B13jws6ujY/b3naS73/lWjHmaFU3q2RjAhPadXu9x5X+r10tbcj/SJT
6ADFqitCgjLmPJOILQX3gCBMud5bwdc4+tY3lVh36PVfYq4RAGbD08OmopgsrdroOph2xXnu4jtU
HNEmkrjMOXj+s2PysP45BQ8X+uEB3sazaYsssCM+5zGypQ3CjOuyvHiD8nRHwLO+7tcKkTYUqUCA
fMxB77ncgiPQMH9PdMR8tKQquYeG9e052OIhyg0b7EEM0VM3bSrjUipctyXjzX0zPlJMvfJW3PgW
7ntkKOU7qgqbAX5XQ7YvoX4hFKWWPOPxtbZeNKeHjFD8Q5go+M/NWosWzTJ243rPKE+C2NMxAPje
v5+vDyjJNY69LTbK3UENO0qxSTUMs948oqGpLPky4amGlqoYLNkyQpOFGaoHtLOzXoMIglVWHWf4
WZJrdSFUvbjKn9CqTp/bmWS6j8ipo2yCBlvzl/iBlYCOcBcvIDnNwG9qGhkLJlUNV3DRUC8PwnfK
DBbND+BYNMInBZ7nDgc0wBmHBeJzBbCi85g9JuDDC2DuAvIOBdGv01Y+OQjYzUw2zCXNoDAkulfn
fyN286RsXR9lMTVFfBo9S7xlvdAMkQj8MxZx3JJyvR152m+GVSIOF/6rI1iGBFawJzsNhjb+CYx2
Qszy4MCnYe1S/Je+PBhpuPfDwdYquASWE5YHeAulYc1yyKksSj/hRPJqQN4CK93J5rx7LDcDtuEE
ZxP8AtmOQaWRfsKifyWedD02g80IQlvawyXP4mYNYA2FNB/vu/3WJHgzy06ty9QDwRAS2A31KOIf
cx1xjwlofFM6/cN6B2fy9UY6o6+K4wIK3fhHR9YAQtrejsZavb372hIAQDUvAPZvC6FxOV5lQnlV
GtA7l6eGKj9dIfvhLdaJK8Ry4qFLXrgiL3rAKHfRP6kPOkDiCCOypMK1FLXOQXlbZf9BHAJFjY6y
ye74eNOcBY+HLfyqQpBtxszaqu+MUUI4VV+xTlZcaA2T1ztL0Zm3hO2iQyCNK8eY1jh6B8DmEdOw
SvA9Hq7cckEOP1pE8PY//vDdB9wJQWJRxQ7f5rgrLllR1UIxgU0+o3cuEABAHK5dI46POu0+TY/m
d6EC6RrOJ3pxyrp65pYdYmRJuZ184EkvETN8sPXTxHeUPgiMgf9t9zG8QZzNG4MTYg3bWa2E+DFt
t3O0Q8IY/mW1CPgg+hUeY3uVGBrad9mko3zQ7jkeVxYwrPr6GasyzaaqK1fL6NDCJpBf9d+eDi1x
dep/LF1CPTWmi8JoCwSqsj6lH86ocL7Lo2zLTt1D1BiPCZ5kzn2QNxnTA5N5/dJaAe4yQanPzkM2
7aiabeIWRNH0/5O91OuHhMRxQ6aCKVoaBQK2IXWYjNXLW68qo/gjDU00zv1h9I+cLrS38+izRp/d
SCaNamh5e5zAcIN1unWt0M0D9PI3vfslcLFFZKCGA4vYeWG0U0ONJYnkXv/GhYKPnnqycU5dXOjk
eCXNKP7lW+uZJFl2WyBVZSdb4P1F2rs4WqZ2NpQBOUA7GWsxWvEiHBzlRGZydS2FLtUG30Ady9BB
P7dLiByQOQ2FgY7320wSfyHwVRr8fS/eIt5k0GBk2XN0wMgX/tC+XzGfsdhOb+ds9wY6EkVmvoaa
7pFXWEEM8IiDTU7y8/aRKexxtUt4k0+Yeo0x1LK7rQuItXOMpL3jBTjCXoJ5PsrHHVbU37uyf44s
0sLpUgRr8XVPIQaxPGl8Wl0iRJlncsHuNu3fqgDad3u51ZlOM4koNpMYJjs/n/Qn4fUOz0I6D2cn
3wXvdyswjzOIyAGpIJrXSSLJGQb7i3xexx1mQFj68Sv9iQM0nvsy2QLGBvyS8HoL8SZcRLX+1xOs
xTMaiPeBASyr/OiMhRRJb7gc/qbR9U2mfXqU5FXHy6iB+GLnm0Wqo+5eDZdWYCSPDSumuA1FyX0T
XNQRb95qAtlrJeAUqphrwXGlHtP2QcJkA/JqgUyy7wWCy27t2O44ZG6rY0XLB8+L66eDXTCSMkPf
W+TU7LdrXFEjkQPEnGkTjM1iKJ3tI2YcVE3QwsBSFI9ROMFpBGA5EIJmp2oJzqCEhrHCZ4k8mKI2
K0IRGjmTwMvKQB+wfNRy9iG0iS4qmcZXR7oUmPp7s5mg/5ar8BgqQTnPBZVO1cQLEI+813ch+zwh
W536WH+HRawi3exTkg0lWst1LPlfQRBzHnUTbAqk1VLqHhVKWjAwbtRxNKlia9dUlmC3HX4k5TsA
ERyQBX3VhZqOliW42QwCzVH5jSBfTZM7lRJgCLG8Hyyheu7OMnCPikpCaM61yxmXSeRuSy7/5zV4
Wx8a5f4wAfpR1MN6hHKLDA6pcWHifY96ac35D/1i3ErZdhKuyua0ZZ7biz5CC6pNnTu3duD9zV4Y
hRtlalQU3B+n8TMm+5ENDxBRzW4zLerVg339Hp7ETwSNtUj3jgvhUutaOE7rWl9zTTvQ/cVXZGN/
0e6LyyHVW0jPJSjgA/T7YJNyulGD/mWHi1Lmx1NSYXfXSp+k5BzAwl5TxC/FjFLeGVPgvqOfqlr8
8ux6RCkpUye8aCx3CNin7w63lW0U4S11frP6v0rY2FYg2xZFkfHqomg9wQAkcpqbWfx7b0kc+H/K
ZZVxJiQIzKtd/qYRxrrOV12wYG8XmtVDhC8N/9iNKNZmIiXaTMXhi/rhHFN728KyRdx4Fk2cPHYu
IFT8Ml+gAaiPMdjOfguKEcTpo96fL6MQGKwvZUO7yk7qKVPZIIlAXkYfHN6/k/y7EcGRRGTvv9ou
9rj8LI7ypZ9Ma0IPZUM4crkYYCQqX4nMa0NTEZiHwaZejg2O6YklSpyT7w/uPk5pM+TZ90YxIadJ
ie/ZSsFzMYsHYkzICbOkSlR4Ra78M1kxJ7f3pMwh+fTG0d/etsr4qNaDtHcXS1vgM/MIDMUdY9a1
ZXzNqld2bdxQWiBH1gfI9pHePrq/w21TlGvSQ5kCM1fqBqQdT+dRSNNPU44ChwRpvUs7R4ZDgXLC
R2YJcPmQ0GYjTjKvq+zNC8lsKophABzDkYKOMkckGdpFE7V31qJYKUp4XqlYPZNflvqtoAzu9slE
huUHV84SiHiEOxkk+rsp7cfjKYdj1YHsAwQXSbga/8KC6ExRV/9quMpdEZu4Wx+Xt6KcrEuG6kJC
mxFveE8eO+XckOwtQRUP3ispV0H1LeHVf84DxZ91d3f7GY+7dsKGsVXf0Dl7gFsxtXUB0hxpjn7l
S97dv+dRLWEQTcBhfGei0PiachTpYWCmC2FC1UcQWMddDMZM0H9vCmA+qk7O/ARjEhbh3HOjj8df
+NtJYpb0oVZOCQfwb5D5jivbc7ZBJAtGQ4am5tK1zUtZOe01vdpqCu4fPxN9ol1v64R1jH5qdM08
LhW5om/0J9J+CHOK0WZ3mvIaZQWuWxO3NfdwS1y8l1NoYQP9yX/NcK5zVIJ5boxY2o5rpHLjg0x5
Dc5WR90kP6Ohao0EhxQx6dSxdoMgLA59+NzOoAayYLbUiE8WgpYhCqPeq7U24JTvJlUOnnEsvf5d
fGzZWI9kDboTqGbiW5F6uRwzkkrH0oMOBVxjB13UCcVa+lsgCdCfs55ulrfXzHOmU5y7QF0KP+U8
U7Od2BJa/SEmbEuWuZSjXdXei7+mKqQUqdPaxUuCP5d6OjBEVZU8gBVG681Q8CarsrBm/9kUZf88
AnS8X2ORWaMkvXQEiB+2TAXO8RYNre3IMagc1PJJmAA+LcdMJUWtwee3sNuINWCcg2aW+fqUMc4U
CCQOH0ocstJzn7KSZ2V3YTckftCjw7wwEq7wUD7OihlStGEWGzFwWLovPH+btUcO3v9WtlHJP+hH
DqlR6SvrPmkOPzxEHrClhCCohbOQc9qaP5nPP8MV7I+gez05nFoqjyzqJU/YdzObGspGdW9wX3Hm
R1xK1HVumWrz8567GN7GiMQ8GtmvYbp2lJE+/wq4Y8VMPygWe929E6yQBxljyzvKNbGmibeGU3UV
sAuKTtoZCtAI4yFrzh+3GHfY0HnBSiX4tBnGdWNl3N+BFHbI6pBeIO9A5MovG6XgZoj7k0F0UhmG
6bIt4QbcuyZ/O41OmZhsT33Q33CRpRW/1DnnpFgs7aDK6QlxaSfpWJ/YTRXf3lK5f+TGLDmisDC2
dutjC7MBOKbccZQZfFdtegRWoi0KO/7NIO3KwYRZ2CfE6napAhavhgU/NOGhpPdKxATf+X9oN4Gw
QWWJh3XVoHudQL1fMfy1dOv9Xep5K8HZvnYnoSPDjJ9qwCnywJOkA5weHykBFz8M1vZ31kG+W826
V9T3ACJfeL6lHLtT1SWCSleD2KnUZPPgEmkM/z8+pej4IDZWNgtp2G9SB5p07XvcwUaB/NX8D5yN
xPI5OXGo/9ix/UZ2AYHZJ+7SKrp0BqHhU4SZaHO/j/fAyDkfwcwzo4meDlHdQ+s//V+k3zvPKxHi
rqd4P0OKf2WDs3Ll7S1Rcxhfo/yXyRPDgclkjPZGr5DtpWfWYJ7PH+n01x1+5b92teJMS4N9ci4Y
F/WAffLraHO57uFsfulCgh8TJcIdqVhu2byJjGkUiL1iMPX+dTlfrm7AQ/SEtYnvmTPgRyD7D+7n
e3wk8cwE7AAVahVwWz7TrWz4ratlSBqrLxWsTlLztMrDV7dZwK/r82+f8Q/aJE6sq5vs75yR9LP7
w98RP9PQUzR9bMrVkJLVBtU5eUwzrJoOljxbhM/R/X7HQTadx9MeqQzf3MCrHdtcnC1hp3NQSaoV
0fWI6kwbCajXroOVlWPTRFKJjJPiECnqIw5Wxh9G8OZQ+rLjnjHzHRVwLsPoh2rF9szISo4XbTTH
FUJbflEwFeyO4InuxZ8V5UL/mtATEoRRIFPYa5RaqnOuDriyDfNh863UgC5bM4wLzk/yQKFe1z5J
8z6cy9w6CRSKMoSUUxGYNsAiQkMB0HSMUGrkeBYdb0F0tpFyKD9YtMf1gRTYPUYRZ5A2IP6TyCwi
hn9JPO2P/NEZlmp3GAhauV2ba6AlfBQO1PAO/7viAcFGpGlXc8eyBFgEnrxKp66ZLHOOlAfSQBu8
uxOjW2hcLzSKyDHapL2R8ndid8Ui+aPacZNH1QsdUAPETC7d0RIPI96e5gn0UZHIy3qKW7HUJH9B
7H6BNiOJckZb8aFTSQ3ELDbfFa4vyPOPUnw/VRgI4T+0XRSoTexFT8RzHci4lZ8SRTDTWNj378p5
7y6iFc/9fim4W2P2eaaeMF1fZpIGhhmBMlCXtvbC5EVHin+c7cVFre4B6JFqgCc0Fyx99mEha/WS
m2gDDYhuClEvyVILGShjgXftfW4SPW8Bea8cLhtj331RSOYNBGMj3mit1hxHcLXZ+SblQsBd3FlF
uLiD6WFTGGiRogs66AolgM2G5EN59cl2VRz8Q7i2TrGCF26bS/0YZ4aSOIw+rfgiaXEFTcqEKA/j
x1MxI+o5WP6MFLJ5DnS/nWtKr3v97Ss1WmfE2SQ+ImSZZDDo4In/Wj9PZf6Bfr9XxE2BdoGDiqeZ
dQRIIgeIrZzQ6O8Vn8EKJQjAy00CBOu0EWxGE3DJo0pXj32aW57fLDqwFAAJssbubt+jXKVz8Y+P
5hYAJuryjtkQDSr2Z1gQMiPo18GwTUt4QtC+9sGnJLuarMDroBMxUlFqF1GivUS7J7cLcFJ1lLO+
XhxiUjLmbb4v3V+HwONgA86klMOFDh5arzQ9x6q54tLtfGfuo7iBMBLTgfPr2SsnmEPAG1XNd/9w
aLwkgbV8VPsQAf/Ude+oOISV73AIyRQ5xNiuvP98sU2pTwC/C54g9/qKRZ3QfpiwnwrwMMYhX8lu
Vhp/DPMSgmy9isJc6CXbtmAvf9wM4Bbq0mZetx6TCStW1VBda0byycWkxq7ddl0Km3JBVJPaq4hE
wD4W+QlpkIDYn/SARstoBD8gK3xXmItAjKA9LWSLRI7sjKQ5HBFjAyxI/Rn0NXPvOvI0x4UtA04o
sq5xm4ckk5z9dxEoyy8c6ZkF6G4olVWhnzeAYNz+bQG9m23Id/aGqkY17L31/vqXTi6oGnTdLJQM
ZB7EVrSjwkZQcK4Ndp6oW0cJkAM3Aper7vS7nIkP0Nfo3ZUywGLoF5Vip8TCaWUT0mDzX+hfn4VG
qwm4enAdjkae0bosBqp1WQ4Hmdk7QYuILqPcB81LpmmB3u5gq3z3nKLeWsMwcNZ4GxtSkTlrKtTL
KtbzwtgJQ9MntKS/seBJ8NJRc6+X2Wl+b8I336DLP4beW8zWXSJMyPJS2EYqZa0/9x62J9Wb9oNl
6bhKWrCtIUBPyPYjhlP/w06VWHXemhHt228MhAKrf380MdWq0Lh0FfYNega0yQrSgRr5Axd9uKjh
8Nr9EZW2Sn8tuxKWoJGqw9YD6kD3+qZJhUZsAYag1bYuTn8SQkV0xQmb7OrQ+YpSO9TBuHMfw7p9
kg312XkiTq3CNjK+uN6v6dzfYd/V5vphaA6G1a8pSq1HCqdY/74k7HSDsKaDkwl8wyw7OTj02d5D
nDhSoB76y1I+I0XARfP1Zd6vhJK/r9BtzAceR91FlzZETMMX/HiXEhBToo1jgIcbvJXc11sLiz0v
Q/Le/C0O7sZCRyde304mnnPtCebhvX8Smm/UZwEtKbuJn9Jw8npYm2UXGFRy4bjSLQiRdJjxLoX0
JJgdM1oVxTDe32kpLyphPqVu4w8wQuwBvKxM1CGOb7qilQSCB5PIT/8Lujw+6Z+3uSWfzTVz22Bn
Cd5xBsKMy38LLhcRJ70psfBZQldglCTmFqIzQvOE7Zm7Lz4ScJwrBKdhAw7+rTakRJISmT8JdpEw
XEhJbKc8+67DpsyyMYA3nEbY2tYeKmUQbW6CDOZdQfkUu/TxcJ8zDV5gdb2AZMciUm7r+slVRxIh
ZCQGEF2M//38rxBZanErL4dNTId58uQZKtq2loY3oAbfXP3sG9Ea0SEJU8i2lyskBodlkJR5hY7b
ma5KnppMJzXKxFihhv08C52eHAM/Qd2GltN+NZMAbw+bAeg0mpprC34SGW2e06Sm8BsS1izegVRl
7FxYhVYZcAjSscd42oGrpK005TENMZCsBwn/DXKrU+LL9ARAggjeXKfWuSmQe+tpM7c3mGhyV4fB
feyNkPT4t+pT4g4nN3JGeTOvpRYJWtr1GqCo4t6blJOZCcwCxY8lczKVKfXEuoY7f5QL99aTd1D1
qWFEJCRT2iyWvPcLNU41a+YZZKvOjLI5sWdpwXiqjBrBLmBwoc2jQboGtGlgRrUMQ30el0xM65Dp
uvj3/aksXWYB80yLDVXC2CEom8pZi9S7VGC64gmZOqL4fXVr+h9Qovf0yz8+s7dkROAKPG7OEUwq
/0tq8FPdHvL3nOeNkFMeihrnQycBPBmOW4npMtY9J2+UreJbFung+MX00NTmITtXiANC09QmD4t6
uNILJK/sKE6aKShdo7I++G0VTxMXD4bM7JXJGnFW7nDmL54o02iTsyWKC+A2SdOOtO/CPfHZaj2m
kXcEss40wVZN3GfUIoE/1NgEUoYz6Af/ecyPCEzvN5xaN6tYcmgZ4ph2gdssGJe20Anl2vwBPKNS
6ddBXG1q7Xu2fU2MvshWfwq4xJYfPoy0ONxRr37zh+Zr+LP6rSfLwCO0xMmtW74w98DKu22h/IEk
s64I2yt78eQcRFfwKhbO/HRNcULkX2V6hfBUNJFQDzSiNDekGZkLkpYPouY1GlmrKOhmKJtCwER3
0y9E8h3ZFmXfTlbuC3lxKf+5S64VCq8dyUmFw8pLUfAYMQLNa/gaOYGR4TiGKmupLcAcriXYe6dE
lTGMNJn6RwNxEN5reVDWWFCm2q4bRJAQf6MFEJfFH58Yo1PFy/1H2GDMFTfQwMaZTo5XiAExzhN7
HUrZTTalBorWiNL2Q4Enxw02k2n2mrPB+CY5BIRep5KyLJrD0XqkzwphsGn00ic7WTdmqbn1yOmY
lGH44ZZCr4VO2e5D0XWJx+Bn9u7uDkfEAC6W8ITxa4SbUcI0lTfaPEzB6l1GH/aMWjYGDxhyNqnQ
AG3ESoV5gLQvcwXOXrqfjwDK/N3qR4Uw0q79HfoKE7mmnOXQI6DN8JjqXoggN1nCpNFyj1AQLiJz
vwjZyAApx0vKKn/hqUCVckbbtgyC5zUMkHyM1ujmiqDiXhMNbBwb09xWQOHBVvy/H4juAMmpJolh
rVPcXC836/Lgtj3/4vXIAQsEKSsVzitcMWfWmtCMkt4JYcyiVGzLQ9IwGU1namSOF3tfT7p9rVdz
mu1Nx0QpBYPXc4WF3WyOLjtiRz36NW7/vxa9ZzMOuYE4Q8fYXCsmIewZJBByOF4UBiMwmxlnOvVc
RlafYhM34yXh1z5rt7Vex/Kk+llsmDJrN4hgKgZJy77HnKrDhxImmIXUdC7t2X4tq+vVoyiJOIe+
cnKYzBFLz/XB3xco48Tt86c6JH1lDwUxyHBUP+fJrb8ygeoB1KlBJajtOVq6sIQht/6wLJhmG96W
LuXojVUY7Ja4LYe3W2Ag9cI0h0zSPbDKS+jpeEFuMq+I6ApXJcT0B9wk/zs1i+YSh8XOLJNSWEnv
qHw6whdjlxLZJl11iz7f8dEffXPZIblnjz9ptLardwRgnRxkgo0fnTnixOsb+Z1Gj0wplpE74LdG
1OCrTS5WP5YOBbLN/bZg21XKBnD63xNUfEs0q0bGty2Hkv01caN2xnBuEPwtqAZSN22Meqn66FNX
j9kaipmdUh0DxExhcuVYP7RL1AWY4F79KaaDU1dmyvpDYYUKSsxI14pL3RUtnTLDwgWnhuQbIakn
ZVW6R6oyCdGKZ3QToyOqnU/8QuBfwOsjwYVwFzD8H1cgBAqiKsUhRzynP3jU3BkTsJxZ4Fea+Efq
/g32gwYwiTGvfAqdTg1HUXe0zm19C1WvZ6Nlt8tVc0sPcW2uayha/5m/jDl/CQ5BFE8Ta5xfIExF
yvGd1T9LtTPR/tL6Fqfw3r9j7qbJXSU+t0xtSIZTrGH/8ihB/yK+LbPgBXk6QrcabcQbugeJ/jjX
Z1QhX+leuPnAoFJ+CskGhWoCKvRyDTuB1jC9+6WNEr9tvUv+KodU9kN57InfUwKtgkgYuaNkc/YL
CRrthpm/QUhQItel1yWvfM2M6X+JnJcIMbgp87+71L80Gfs9JM877PtzWAoGxneUAvhltoIvjFrL
eM39g3f92L2gjlsxYJNOcZSFsMuCFLkrSEkgjo66CzV6noJpTgoOluQsOdXodajUnSWChOHmBLsT
rYcT4FYnv6tjAY+AdFLjGc2zP+Y5zLjsexfrky6wZVLpfrtXEGLK+rmSzCotmXRIDOJMnELdOvuB
ZexIOBvYiBEXKXGhl0G94Ijk9GH+Gg0qTN60BQvYTMyI01P6/QYQ4OHayPG8PeNSknUmIDh3VsQ2
qfT4y/1O+Pl+nqjW9rd2ByKXja1xJfRKR/FnOsxX7oIdziZdPiHH2kakft1G+xvDiBCBSB26JgLZ
rf/H0GDnYrosucgkLQe4w5kQ+WaVSuBnOUWQEI3fWI0/RhYpIWnPnAnQx4tVvt3szy3GyzTGEs50
UMPJsYRUJp1vNPAQyf18yuQl2PYHz/Fd0GzfmFomkLr39AXFsbfHIbQSGFxM1RHkrIov59/JZIpP
bzz6n+AxKfWvvppQiZ+CM8WzKpg9aPSeHFZkA2g6s9TIlzj0NARz/0Z1PUZ9aCnjH83F5FovyppF
bkqVDFwd8CIpwE1pfMlGNmdaa8VWkZI+zk3JnDZkybl6U8to2wunTj0pLh5R5jYM+vjR+v8idOAF
bR9U6RGeesRVv+VqXkPRP8erE7cuJaA6WJnDm7m+SVgiA4tnPO3ofCLja3YT8inmW+g3PoX2wSpU
K6aDtF1hJLl3dptD4Y4O0ZLolHBLI7bKvkTPaW7MiONKRgysz1lBEZtHE9N5/8/H9QRABga33GSW
iaRkiUSmRQIgOBEOSbPXwbTO3LAVegzdZd9uPo168n4hgNK3koYATWLByVV8yB2VBzjr5cw/Sg1s
Ct/U5d1pcMj0ac12ZdrLm9TVxQEKn4a+op7DjIKTQWfFAXwvIYRujDRUG1JsZC3aVtU7twXu63iA
K5alOV5S0ZQH/J0MrHUDWp0w0KVj7LSqjkd+R5fiard2aQqZc4VZuUs5pFEgDXnEu4DxY1W1rG+j
k7anXiNZSWmRQCGXS/qmiCkQX8ZV1/2swyoJkRpfgntJ2rU3G1VYxMrA4C9rvIZ/nQIq4qtYPp4F
1ujwSHp+fX9vv25opOQAPZjnaYXPzLDP+iS1CDO3lqWDcqwjEq4OoFsSfhn4aiWHA5A5QB93BHlg
GKRP6MWi6Ka/i5zAfDahzsbqO5O45JjqaE58D+xNJztCCWvQSf0SXQu+9t6qEMicxe+JHP3etFiz
hefdNJyT1fS3cWQJAd3wF/MgcT3VFl+kx/Tj2SV70dpYf46/KNBeuLIWnbB83jaxhazq99UA3Y3R
KrZwbAU8UoT0IGBlix7ZdeVdyOdtGDVj9FVGA7qQ5yrCurogEraYMVVcatWbFfAyqxd2/GpWjCHD
cODYYuj8189pR2k1+pQJiaGRTeFDJqVQwlQtsSYtqiXn7rt/N9ECid+N6X4F2qRtW2eJi9OV/vKb
g8Wy+4JqNxF615cDi+QpdCgqKYUA6QKj466QvYiMbc9/WHsJt/etZQtCLmgbzO4NPDDHFZsM962x
33bfa5qXkjkiJzjOMlqrG0HkcyIl/t0uhn3+Lg93K/QZtIEdgbpIbR6Gq4LkLwyARlmUFg2oCssd
9tBw8yYdc1m9/vjXLTXeShqmHpTlD3ACG8uy3iKYeLSWLhb5NEC9YD6rkYGIWHlqMTkb5riRFneq
oS8DPKE/IpIudRDBwK657kK03Pehc0RNJ/MlsbcSm7XDXcB2hFfQoam+K78Hz2wkIrNkcalKLyDw
dj4DWXhrjRM9C0vYYPR0CXQw8NcJVEtXOXQEfgx3slSFEP8LXsgoxmmg81xGQAXNxcnCMg7CUPy1
4CffICXF+SQrPXMiepxIFCbSeQnxzgjWWx/4LDIKaepN+eF7RsZw9KirY0kNjxXMffAAgaRJ+/0y
szZED1oX2UXSWz0FQRV6UUXeZqd3Tp9hGgmqizFmti1nLhjAXxAkAWAK4bUQia9UL5BRd5fZOJqi
5Myz/ygDcjc+ylvbbp3dOgGOaWXrY5OSVe8kK+iI1UlP0Vs5t5XQhkFwXwbRA7EO82tCrTl2POoj
zSeDIoaKY3fS/9LznthzuOy7JzLQucnJSrTPeHDTJB0wgTnulzXrr/3WOLsmY5RHcOQxX34gP+UP
7D2A3Oo4cf+KAT1Kb8o5n+5SOZ80pGTh+grmiRmdLz4XgmQI/mv4S9oXr66Mx6CxGw6P1E7W3oei
N81sE+DRPcyPJo7WoPDrrNKuv3kL3fPBHMVBNLTrgVoT3B35hHj78L1rOUOQ6/l/bWfdF6flqlFe
P15FEfc+s6r0Byahq3Y2YcscSeGyiULtBshEkfpYRwIB/eFpwsSed952HRQbObZAbxBiRrM/oV2t
vimqBCp0Gig30D6Eq2LUEePKzLPi3Cu+TehPz1xIj+5dKU2KcEZ2IlCVCoRabtZfzb0fRyKst/Ix
ClAwYrwvYZKslLfv2RV7L+rksg+01FvwBgmjr9Ahuj67zd01A9WH7MIRQ5JvUs53n+/iN3kQJOIk
JybcqNiFfrFUGTITahWJ0Roe8sw+ETy0nWn0SCn7x1Isew9rCFlpWOOTF/OP746QCSD0eOJ6riNL
IOnMQORpGOchaccafq1OLdYAPvpBFqstpzA6ZyeJ9kgLgmcjVFAO3uADHRJIUU+wreChvJ3KFmNu
s3JxTm5fryllIMwPQvpjOWg7ikPIdrXS7QY4O6y4NCRzubGLeeusT0zr/jjFCETcW9xJLLqKMB/n
wjDd+HBw9j7El5zROInL2ANdlofcxIrqs7hjT+/uUPZcYZDySBCexUbawL7lgbuFlYU73nH3QUri
PKsezkoEb02rjKDL/RFMWY6gheXxnVNw0tVK4H5vwULHOGMfu+yTgjk0f9RWi79EiD4aQf+St83r
E1ZzS7aPGsLZ2mnJP4CToa6KSG3x7aCX8ld4CY55agetYFOofhkToaY74C8wixBWihy3xdpH11RV
pde5lc8oBRvohNOKj6qekAD/zRm0LZhUw/OdZPbTQ35phO61PmME9wKpHFieiDmyDAVltHp9lpPK
cSSpNr8MaLAcMos1VrrhhvknejXEhq7qS1uN9FyH0GM/fKoSagonGSNA+LbefzQUFk9HS8Js5DR+
6aPZKk5ys3sd1XRVDLw+sanSvkYIMab+tpnSzZgMqlSYK6FEtwa2MVGUT03Xcc+UjPCj6X8We7tI
rZP2iupQ6TP4UbRSxusaEYu1gCOb6OPI8aYPbYb7zFdIrMdCsAal143QLlM5hljVvq7MB1zm7Lcd
AKDGdD9nUc5DpAI3GKS1Z3M39tvUyzYaH3VJR45XwLwnGJ0ynlQ0mQ9uxyms/yQ7Idmr5aMYTsjQ
KeayhcLVK0jZGYaRQow2c7p/IYuc0Dih5QtAyHg0b6jBRWck1C8je05OTNfsATYEMRlesrkfg0ON
icQIwWkJPCCTX4CN9dfzc8MbbUyIsUXxNlB5U7QYt5uXxqQT9RDtqbkzbEQTB9Ne/i41fTI2w1c8
870v7rktwIJ4OHvWLDrOSv6a4IAx/FTgA194nDFIHHTAH/FUxeKTiOq8xavxvhnJ7F+BtCOC2r9Q
doXV5Yx94MWbZi85L9aTgiPupqNhSa+T2qYp7sPBpWVsJ+yMloXC4yVY5C7aMGZy1rRIRsDgUKhZ
YTLqKM4COlg34FJEvtBcIDqI837qBAsLOF6bN/s8IeUguksZIVFnh6J25rvt3zSrcfMyCPK2U+Nz
3iKIKUwaoSDW1Fw5ldUEAUoS6h8Hoyp1L+6zaetzI6BR5T+aj8hrZgHJF3Y8s1pANKqkWrgKJ2ab
yAki8dM5M9x+vHw6Aab2zLw22D5Xs7YGEfvsiTBQzwyUhFz/u/qfaGj4EJL88UK4wWKY2NGnkbCr
zm+RL+MT9AZtHjB3d3Hf2Tc/d0sRnJE/wd1pKB/l72a6qY5XPmlNNaBlF52NXAKOVyGsLtF1SiUs
hHll6K4sswmmJc1gCF7mJu0/Gtt2qmS7LyhQK8dc8QjoudnNoN0m2gop+XMTzfflbNpGXvJEd6iJ
wG6V/kyZmisXwojOMV26bi6D/hLZxIIwORWvrfu/7o6u6JF5+sMlx0TL/jD/JB2khNNC5CpE6jvk
AtCtBvUlXg7UO26D9D08cQSxbfqEr+MScVZAxHmMeiBobPGEchafOF7oz5Q8oKwq3rWZh1RxQ9XH
2EEmw+Ms+xFQ07DTvq5bqvgqAe5sW42Mr812UPlOdmjWiNJ+jw2PE7DJU3C11/jQy6y28eYG5zMS
LGAGwmGiecgcqPzPxp3n9LFVUVgStDE3noJCB0oSqah9HBrjdAV/8ZqrwPp/jB5BlP/6KO31Evv3
reNhjBlae0DpAu/AUnAnGzNKqmSjG4wuSln0kvHmHi4HZVvSRscLfFqecDMYsy8x/lZbhGHu0LVC
jAzW5A1SD6soXXEgZsqLIP00Ltau5RH4DaljlOvAdRMvNRcBunXj8nRNEy4H6WtbVppmy18qjIG2
zcM+XCDWPXYwaG1bulasnbcw+GJL5rAcruT4Th1uPCTKiJKVDpjlm0QqBpjQp51/A9nYFubkbK0y
RpS6fvsx2pJzko2x5ec3R6TLM+3IOHpQIwo7uO1dVCzlQjETANQxZABYpRRmQnwqj/aIYeRMq9ir
FXOdWI5nw89ttD58cuJV3YiThmi+Wk7OGSrF5UBlvt2yaMW7N5FJIdfAISAcvkUzzooJoHrCBvO5
ccOr5hUydkJA2KtBYvnkpuYxWTqTnEaDx7qbd+66uahB9yVi9YxqG22FwEhZWxaSnObfWbIODKsD
CulURy5fAnD7XpkPXI3pjNn2OIJhcno2PxwhMYz2CkeO6e5QZ0ej8N5uqsbLkVLn8gE+1X2CPYQA
rAXg468Tz44qJam4sbeq1D7pZOD0a4cYzGusV48ANThCYQOxb71fDL8sSHQrgI+WNPF3AI48yih8
P1NqoKQJetWdSLPwzrVOw/KbCHv1zTnf+QYGYbn9EXuxBdB28RgLuAdMWb9pR/2uv/4NGonhGP7Y
ExE+roB11gf5bZH65l5UUjTXzjA+vzSo2VDQ5ZDHVorpDo88ypEblgaBxGLGISBm5dbZZ03d0Vf3
p2hakWxlTc94UQlN6FekANIe5l5EBm3Z2M3CYYrrem1SXJPH9K8SK+0a9oUcpZVDRz9Xc8tfMWXO
MY95JG6DSTVTViEA1Y0ywLX4WU6r9HAseRy1XZM6gQb0hEv/CUEUbb9j/IJDXkG6uKj0LMzWy3Iv
1dYUMl9yIADAR4C/cDOZ9C7yPXvU5dPuzazgunstzwZCKzU35Zpb88BJXC2brzsh3Sl3XfB71EqJ
5bP6xnyEGLulDGnLZ90WScZI6M5K8g7Pw8H305DBbG1+Aa6IETiWg6R4fppRBauL+5RJRZr392di
Ha65QT4wRM/q86QDMKUlF1jkJY8/AqxtR/q4Q0ue5s3ESH3OYlKoPPp2mxlxXZP7XftMsM/+gcwp
+6WK+ZHmX1DvYv6AZYZ8wKn4YzxeooZqRQ4OloqheKbsx/p0sn7J5ih9WjUvVxAl1NY1ncOLSkcH
t93F+Zn0/LY6+bhx24IRJEYrxLPafxf5xTpiLsfKNiwJ3CLKixCqubRMb1qIP1DHR2vbXlH6NY70
pSakBDuQu4OjjoNEJLHhYBdPiA1VyKJyzBX+6XODfSahf2WG4VLtN6FyHYacOOksnJw5/PO69A14
BEcgfdYxVdc3lmCXQscvQdldngdagebG7UX1wOF/PeSU4omEO2tOWZnMRGaLBmn711sCkrJM6Yex
MSG+tdxxAJ2KDc2jwMU5eVrfka3Pj79E74gKvzIhB3ogfcd5MS/ORJTa6/P8uT/kZgI8YJdzIwKR
iisEp0JUagSN1oRU3jSwtdbiMWfJoxMjrmf2ZP+TkC2OqUwKXvCGtxIeRG33ZfzvvvOHXzytfW0r
SXrVZTYUXfqvTEuBGyVtMJUv2O1CpDAg2/EiO3wlDxEuPoqZz3aihwMuhmQ6aps8ihdgkQE4c/9K
blXMlgY4Ciu8hYuWVFmQLCPNlN5R5hTres+8GQkNZ05sXi4rFUlPl1MDUQdSm+n3iqpZVVqoNLoS
PZ/pTV4AVs+U4H5BQI41b4ClOwQ5SXnhayMSqEXQSFu1qb9DDYlpd5xn2FWhxCH01PaMZwmidWYY
h8UXo4cpaVjRAjZ8UJZ7gTNjRICPfEd+noixyYglLwgMipNbkrhf8qUwzVtYiL63na4pEg+JodCV
fPq9rjcVbaXJzmaU0UzNQMy4rYfaIWjhcOzOUo6bFRNaKlPjMHV15Aeb/cePW4AOOJo6TB4XiWgy
p94wIJ59WT9rGPV98Sn/4CE0G/lK4ivmlQbOXz2VT6/WizjcZEkebRmqtSM9b9bfCaGB3KHwL+TN
UkzdKADdorcK/k4Mn/ZyBPG4JGNRpds+BqFF/iOhxYXTQCIdb2P0jLKz9X1mlN3JJLIfgJJxKNOE
3/iMXVpRAg+wTM7gamtBuxkMvbfVzNXNj5RcKMcEgHCMmv79pBtuGNsSPddgEtcpBJyCjzDHzuh7
DlM+RrhkRBWTLZupbTiooONR/jFSwfKSXHqcaFxmVaEYA8EIbNreLBlNUf9W0SqYq+VkM6dOCWsK
//XAL/IqCGW2m3zKZ9orDyRoNzSVmVNaDOV77+frvOLJz+7qANTnxJ91iXOImpe2CPiU+re2a9wX
JmQGYcpZo6IMixrKJk2qMO7CE010rAIpesLHtQ8CwsjWc7uTzbRNoNMiEXQdO3kSCF7a9+ch1kXe
vepqBGBHBNORp/3mTyjIzUshuGg2r2nSq/wHKY1Ezr7hxrWRS+cC9IOOsu/KOlfyGha+760IIcdc
jVRuL7Bdr0bBrSIKbhDxP1r4ch0Eu53iuywcQCvIUhpJU87B4J4r/eSIOuUsFfpdl54WT5L02sCi
o0BdTM6KcjIbtf/hqZJMy/UHONWSBR1nwdqoxs2806IPyzPs5ow8uEHpgtuU2+3npOHVY8Vat/yJ
jpPX/PHHeGc5CMeyZ9U9jNBy7N+J+ray4cf9UNfvU4NxTp3LfVXwBFZcDajxWKwtIIlnxt9exgHU
t7VN6Ik0cVnXCS+eSomNKW2lJjMrJFii/A3ADFv8N7k8jghP3e6ZtoFVkgWVq0WQZ+5oLlmftP18
wxXph9Mof+1Cm1Fa9h7M8AOA1LOJGha3KYnu6IbVsiESpHz9YATOULqDn0ftP1tgVpOKBo0pCnDH
juhbUlS6aNRhQ7LzQOsAQ43/sAcf4dr8FqbmGRd1dtouBGFe5PNupyLAKgd4Nqs8N7uy2T2a7GDB
qYsiyMjsFH6dDDXMdwb+0x+sNhcuWLkbEMqmmi7lUlHGBYQC72AKvtfd5A1FiHkYhMlYsNqL+ppV
W8qkrtA+DuP4/jxkfxS2IMUiGfhzsCTXr933gMUT3W5gLVEWSu0q2Q/yxmmumlnhYD04IVj6h8Tt
FpwMH38y3Z3wvbSvUoLz2dnEwXXc0FVJZbugxN91MV9vhYwBB5JyH6Bf0/ZEdeYXKeMJb2F+VLYP
bogEoMh6HKYyt8oQNQb1JVqzZVCiKkK4T+LRDDs9TvVsdvpIiuf3ktJu6h9zSuoLLHxvkRj8KwwI
VgrxqMcAIgd+/RLUnFs8PWDQf1oqrzaho9rO3oIccurvX11ssqkBirk3tEKWvNNa1VfVbZxZp+HC
vLspTYKjoca05Wpmjem24Aek9vcQWri7Tu8WSxu+skhp6KkJ50QYDzsBXXUnREFqMoc90TC0ufqp
ifAVJsVLppHD8I0SILyyF6yCRv3CRIWKM4sINA3JT5FNZqLPLFG30GXBEPQB9uK9NUbNFYcEiMWB
WjjdxCeQZpkeKYSXM5wntX8NkCApgRIQYGPr2I1g+YuDYxrG/4ppU9tjttBJd+crbW7gFMb2v1oZ
1nhA45WxDxnSMN7jiEYx+ckx3int7mfbgNGx6jvY3GZ37gU0ILCT6N1xG1nkNJlLa9sU4RtynVlc
qM7/RTg/hznylcOY0HvG8UqVpFyHsS4IiLDF19P4WM6zVzG5qFlThXAuQUmXOOEbdLweKr6NLgVG
MbEBcQAvIlQK3GmtFj3J/ZA4spyOAdVXplCqm2euImBoaWRv9Q53oCBwtYwXidzJ4BifIGevIYwe
e8hNMvwWyIezVgevdzH/UDt+wCKdR94bfZLc16aHqaXssD4EOBm8pl/JW5ogtqnkc7ZYgi1UnBtO
Q5/GBmTsXYCN4GHsY/HMemOxrrzDWk/V/WkkFrndAD0+0Vyrcy+5i6OiUBlezRT4u9dPPqpPKiKS
5aGy6Bf3fSiH+GBGrgpCzInusleG4Jcrk+xJ6iRJDb5NkA+4jKJg2MFd09KGttfnIfzNJHYtEVoG
P/9S1J5UgkXHgmFQPYVZW2jUC/8YVoSxuZKfNtFsy7E0exMXLZ7SVfu8XTl+/xP8kfp2Eq5HtUWl
qBuJ7OrK/0G6UeOA1t6KEMgDliVwPpHOy8JzJEwO3T5czZb3AlqqO53x/jBUZXC5g585JFmCaK1/
OfyskmKHq3mcSy/XHKz/KrTeAQW4JPZH6ItZUZTw7vVItWato6agekXdmjP9y8LS63syBYcDrgCf
IvO1chNu/hL8YfyZl1lzQ7ezxBk4V0sZ6w1OYJNWAefTBH1EPOe2LrQsA0UZTrqoVeIO0OJ259S5
fbG/dPtXcUto6v6cQ5TSB7seqpw6LX2mpkExt7uzPtPGcz/FAgmyV1rMyPDAMCGatUrQCJSIfDBH
em6gTfY/WH20Md6tzS5pMkeIgG6taR8bKZGaTbzeuWqRqh7gFKhLQJB7idnml7K/GDePGnkOZ8XR
Bv1iJbh8rZkAH/Q0N3hByMq13iFLGDLjv8HZik39FA/WcPcPW/sAmVXSC3VFCWJ6suiiu2XU+aoS
RKeKTs8yNyrmwCXmIjKp7gxCrewtloac+tisRou+TaovM6GjVDw3D8VXYN7yU22lPnAbA2B3ITqW
C0wQaDy8nuo3YuvVSZ+lO3NeVwWhfHovmMSXJSVO25N4OJLRQdqow5G68PKM4ksLiblHQ1EUmYVO
N7ZMl+4vZKkATQ18G7/wE7G+6gUqICigHsV5g5fd1hFbTEKNQKIv68oUKCJ/ONdFzNguFT0d2LYw
haVr4L+7KbruTUkF0Pj35PPkpClkFcHgxvJwuHUS2/IuJpNxPssMkHH/bxf7ZOSYPAhmLMAz9ivq
C2NfePd5IeTrjtMtp0TbgkK7w5Uq+rPLnZx/Rvz3g+NsMtrfoR/86zfZIurkcGrYJh3e529K7/Pe
ZgjMmWicg7y4+w2+WOiUY7AwIHNonNfWB23CRaGQ8inXmAsaXr4cNzq6K9bGui3gT2NR4nFpwLAv
/66MVt1K+5b95KkVNz7V6B14v7vg5ZAKOZm0QIpv5lI6meZcR6jm878Kv2SSe09c+JujBfI5d9qw
69M8NwmIZfP5SwRywLrQ4N/h/IUi8MNG/ab4BcDVyXVI14kMNuyDxUSBZ/My+sStgpS50s3rUaJj
xORn9uuY2yhY0IMVfa/L43mYAz7uvQav2NH6qPsSQ1aYFF5jOUwUXNPGjEH3I1YdPvvALx6Uk+4/
hVlMfk5pS88Eyu1SmkL3IxNgabGs4Ml7ZBYJxHIAQJrMMM+wjGw8dTCQSyEsVyYf8qbKrA3V53cD
hLCXSP01Epru9JRniZgAyUnKEkScnjE9JOuNnvFuryl+S3brf+iKGevmv4M+DP6ZG/ba7VDbut74
QUtfRtTMvInbp58zx1K48qaLo8CUqZvOGvdcAIF2m4YPRgkQv8DdOuTT8VaQE33/1uUGsGPDY20a
rdITU7zPwIq1ukcPiVgZtWjMyou2VDxRNR1NYNxLfRQmW6F/Gc0onlU5oVYkPQhZXlX4v28XkiIR
W2KeiJss3/exGY8uOiApaXeKvOFs4RQhS7ffdFA4eGXZDYKQe8BTB0tKxX3aNDs+y3Eqvi49uQd+
rA4AzWuqOli4gyluZK1/8I4ru9RlQyJFaRKX3T0MaRkUpJPS6L+jQrwImv1mBuUHwOTGduNE6Q1A
Wvfj/QuQoLrc6hnYaaAThLaWz75/FLcXWdnbtBdxpdpIWUm6J2bi+Xx0YrrXfzRypFGaiBUxMbYj
fha8tQnBmitgSbg4xvCCT3KpKHUE+biLlMg+w6u8naydrxvLhWyzKviOokm+wH0uY7G+FFeUhJnr
WcdFDuKXXzDCxQ7mFaaYPjZABIz7hhOr9FFgXpJTi/03buXgupk8qkhiFJbyt/SbpaPpVVeHQn4A
feWeN8nE9T+yyVtEyqjeoguWPCMHRr9vvZFvekelFzNFLMq0NM8hBOiH035JuLWCx+Y8TLpZ5aqp
E2j8VKC5Zo7Dy5XulL+09czdm63DFlsZZhp8iknUW9KOwfct1+Gg5S7+K4bj0ROI0+0I+WB3C/cH
xs48ccZG2PRBZzW1x6h5pQ5u6zc4h+VBvsynR8VisOyXQMP+23WwqTedDD45LyEiJjqIA7tL6Naa
KeG1ktUluwvXvsvTjamIT/oJ3bho+XZYmF8ET1mivZGzUdOPYKFAQqqEERmgh8YM0Rxqbt472evR
JOrW1b7JU45VDyMTMbnICJUbB5Qccs2kkxyL/CCptUYrgP68r4iPAuAq0U8XUorj9kH3XyGYXDBk
v/WS3x7XD4ykeX8LS3K6ZGVzznH1YaAtMpY8uNiGGFJNjrKzUi561ze29OaPZXpRhgP30X6Ju0aN
b7s1LKzVjumWxoMasgvsykd+oqELwVoVU00Na6/DfRVwIYI+lE3ugF0yBcKLyAAFsmCIKdWuzUIQ
wguR83bAGdNavF5qgIDQ3rKyxthDD3tc25YyvzG60gGAnMAPqExPNR7/G0niI59N1gBeSwRdBLgf
IG6W3liGxw+bnHwi9tRXJ3PdTJiys7OvwT7Cy6o8x6lWOlQJ+f478E76DPREqFY0lfkEQgavW567
ujBZFXVuGCuGCPjkJOF7zzxyWi9CyL7K4lT/IICpBChsoOvjxHcR5htGVGUZhgnt0UjfuR1MzLV3
0+ySp79AbRb7YW4N0LAC0Ny5cLZGUhSbaVq545Wy0FEVv2GyR7I58sczWeBvNa1oomOZvRsqRyql
6OH6tjvdGh7aAltUfn0cSERdvqo4gFZKGay+/BxVTtu9KL1jBijOM1ASVtQabFaGGbWPD9KlH3vF
B38srHstpM/EAZl8jqQY0QHtUT7zokt9CfzwNcR1Wr5WEuGMK98p9bY7xXLspBVIWZdLxg5wcha3
5IzMxicXr0u0gP0HTNvQ5VUBmPCq2qwB0i1lsxZ6vtihTGbtx/YXAmiGID9ueNs7vm7jQuWKKzu+
XEkPYPXfCWIgUz0SqY6wVmX0TiHVLPWUlKACwauYylW2F3Zj131xGBxps8VJYI0BhXOy09V3WR49
BbBCYu4xnGUhkR3X3jQmDL5ncQQvWHoP2c8hg/ijz02p6EZjZL/EqKDQaSi7rSaXf6+JvJkGjT7Q
9FLy7kuWJV6/Kq1TvIs669xawNHT96mz4bb2nE+bGdbAhGsOAC8OxiNNsmiqMpDIXbPCZ728nGMb
mVm2VHJvPfFSPzzMYXaTdjGDlUCzGBzWm2HC4TGfMcj+L/DX7SbOwDxhHwbsfbaF16nWzG5t+qGQ
ucovgFvP96C/6eJ4+Q4c0d9Fq3Oys1c8SYASQaGCCJ3PWGHZE5aGwv5/d8y7jd+xEjmH/eKdHWQT
5U+s9+dNqUWF4IbLF0KiQKaBQdy2d0dywhltni5rhl3oooYohNwZGw251NaF28tEOMUOq+ZKz8r/
9YszTcBl6dms6vEsYxUMjHdr9YdP5W5ds1dGQegWPkeoNrXZ5RVSkb+2/Me33T4NShs554dsmxPR
QRJDlm7Ph+vVCB2ZbEa2WyuVCrRrlh10dqfWgh1qvQlgHzcXsS4q8+/nEQ/3bp1Se/xI5DaB++ZU
0D9JKIjLXj6vcvIEmTWGhz24T8ZuxWX6X/eYvbYIgeq2+YLyJYF3utZQvQ2XwBz7KD2IC+0aZz14
SpKXqa7iu6R+PHSdtYS8gJ+JbV5UuRcsb37+QCvkMDFP/m0IIj/CChaDTN0T5BKKVKXcOQZmTqd/
3zV73eLoVOT7X8a+F74O169fzQdcr46FH6vRsYtUVtFqOPp9wpIjp4waeaEz/U/o+WjT3z0TNLzU
AP3wwdeyVUc1hmcC46k1zR897o0gJFKrrX5UQr/If2GADQmKcEatcjqH0iYj0eE22E2HTTuP67Dm
a6KpOw2ZMDyYDamO4zkIZG1LYCHd/A7/PlSnz4ixunGLzXqlBGngE7Jk45MuTMyLkxPSxYI1V6/c
NKAtGge5Lbvsvb1rQ6eiHMmGumhRT8WSJIwCUmRsq8Iw/Mp0C03kZMi1xSgpLW+saYt0gnkyTJ2i
vTM/GaDEG4NH6M7gBH/efIKynhv5cA8KsgY7hd+Zdwjn5vEFKkNP24vtS1Jqlk2SkS1l7rP8n5D2
6ghHBQ4xBLPWA+SNJMy2KEMvKAQgbT6IALcWn+tw1BZUJAiHFcFK8X9RiU3ioWI4tYm5l+nQ+VQT
EmCJ/PAiU7oKy9nQbNrXMm1Aac7Ua39bN0YXDldO9ZKpzyi4AWDZ29v273dMRmQPLI+kd//aRwlO
Wim7HFvboou10uYWqzZzQtLpcAEkf9FYumtBK4AlE7WYl9/f2FocVjQaOey9jeolUK8gr7Rj6YRT
3wFpbeHtMSjP58U2kf9+zrmeNWZiGPvZlb0P2bM0NjJ2RX2H8A5dwbBUT7KXd+ZUQk2MYMxSzykS
EI+HL3AAs4FliDDeyjf2T2GJdXbw8/kaPdQhv6bAXDImSSOTNvTDSt+rh/UnW/AZqd4gXmVJ5ecj
MuT0RmsICWLfFFk0Q1JSvY8N2lXbPReflhL0JRcKddvGZOloCsr031L7EaPypKErbcQBjL87P6T0
wcPzP3D0II+gHx/0GBJf/zTCSKfs950G/oGEXvI/4Z+iqMI+CPTbzD2MiIbNQS4L8NvzCL9/dbo9
BmJepDTtJxDpLsWsms4w5DqS5aDaPzXj1kMVSyNbpw8WGbJrpgNz9p+jbDGAn0efMP5fkozQ8OVV
rX80QhOk56js1nqbE9jcOR2Sop0tnURYgZSOZ3Sn1oxTDfjpAsCyh1arbYGQFq3XkR20PW0v5ZDe
NUYcJK+Wj+LRcNF/q/7sw/A8V3dRlqDbX+42EwbVDcVx9dYTthagY7xuT838ihb2YPEMLqGJKQC2
CKMppV6yrpGANqjm2N652gEfsjIsjLrX2p5VNx1AgN6g/KwaEsm5XJ8cCNMWJ/F1nFVKX1qwXrS1
wrcgRRlg1fiE7QQJRthdcKe1aQZAmj8Esq48ohxMyoi11zlZOqA6G3kNN4m60NNZZzCQVBLM9srV
IBZpZt9ao/Qg3z5QDlagm3mCTT82j7iV87Lv+u3cWJZZbfugiq9CX6qdsc7oAydLPzQxMeiTMJnQ
iIMaXttDcplpfOPe4A/5G3i+031kMuJjJ0rAtRVHX0Hj2BsDNCcqtNodsTYZtVD0VnUoScSqAJFN
Yvc61GDsaSeIEVSCMLvXT9lNYb2tud55xQI7qmoqJ7xPGqozMxDj5dYUAh4F4CZWfciYkiokPQap
aU+8B0lynmmgLa4rFOFf28P2oVaV8m6jSO2eTG1bJlmakGIFw5I2uyVo7vRFLdBkrMx99WhR8TfG
GjXhAyRo1CSyK5bxSuItqZJ9t3PU6yvhbDyP0soFUzb+6XH1pGZS2hosM6jgVhAIxIIvFKroj8NY
J6s85s4ybGGqs1D0ImI5LikZ1ddeb47DdH0gPITm/S535OR+ttqFKhCSLa8vw26Nc3z6k5NatGPP
MpZy5wsui8RYKCCEUcCFrUU4MaGOkxsO4DlXvlW3s/zcY7sZY6fzWJFz+nx+/3eKmYWzEpRm9tK/
dzZxDVp+ltsmSt+E0bcaCuhHWO+P6OKxJ0LMZl2oztVnVmxbYXMkORU54Y8VQxD8qHfsW2PhJ+EB
9nquM9k6fGxUOvJLQO3NohPJ3l3G4HT5itB19ZZuD2R80/1sMYA1ra7TgZfDzTbSzAKUkSXUCWLL
83pyAZkrcRubIMsdL8hA6v3VvYvXrFxZzpIejwJi/2aYQ94VSydpV23N91MfCgkr5VhzRjbGdEbw
UcwrDJcRRwNIeq48WNOE5c83g+Dfs8XAok5cJ2O1Azg1Emxft1Cs5NPc8cMZAAnG/mIni1pY3Mmc
knHPgj0/Fi+SeYAhRr4bRb1HfwHV/i53p2Ow/BaQzwYWqLS4iOEfb0Fs79FYdC8E/+TZpYueWV9H
LK9f1BBSUQ5xvD6Z+NX593lmFovCnEGADHfY5CLtLpBRYjXnIVn+EYHpF4dKZrVTrFcmd+zUSZbY
23DPbwVPivbwXk30UwAH1cbUNoMFm1CYPzYtJsRwsiEbx1uqysPQ7UjMquKNzvgME6eu+he/hYWf
Id6hc4d9GCAmcPmxqj6gzSfrcfzqJGo2SkUPzubRmlwij8BgMOCgIEyh21weNViiTHi44sJ5fjX1
ptfYd5H3GNBve9Ys9OHjE/K4w58oJ+Gfv+sFDgtTk3Y+/6em7QEB0MxPqagiRltFmCXvOXJHQzGa
DAF+BZLs99fCu1pLAjHWTguROhgDwzCwqAeuuHLTqxWLt6PTlVASJo4VZoX0gaLE5vNL9I4Uzqs7
mSzBRZA7fYLTTy5/mBzundnfOSUwybVpAEJzOIGnZcf8Zt4R/NwVk+hyb4hQlRvX7kITn4XxeNXT
0uZZoBOsl1hfxWW+jjyW+XYRiDlo3kMi8AMVpGfsHR5rQwRlJjp3EcC9G6lbM3X8xJpfdIN7YQJE
V8nh2US7/SfcqETi1p+6dDmLXBiwYOBGlQeRSyLQgWiqfOxMRT9UsI2lHpfXfkF1mdk5LoSc9zja
Zj9HUJCNP3X3eejf1jUs/5Adx7AsqC7nSJTGGwT46BwA7h1cNwihoE9+JYnIW+ctk7MX5LMDxf11
xfAlQV12zz9EyaTA870O44qVpC069D52Xz4QREOZ9MHwBy9UP2mcUYZ6dpuFukAdg8PPi0kLs/SG
wFdGrMym2AR9RDoaLy9FmCscZ3qNkWc7mEqZ8tE9VNGPoFOBdHll8I0yS//UKW4hwZvitXllImQT
EzbX44Ac2iFk7kw2pIADK0D0zbDvfOc9Cv1wobw4haOdXrRZBoermiC6uA+tMbJoU370QASFdPSI
6/lf72V1XL3zR2UJrqInPni9AaZ6Z0geYxMxwqNZv0McfmloqdGtGjKINw9qnUL7+X2ZuhLiCShQ
aVOLmfGdWWWT+oc2oLTbD8FVCPlhtXYJ8dJVz23tiA4rlWqXG0j17dkkOhEb2ovsTjd6Q8sUXYAz
kxYzaqOwbH5DQWxOPN12c6Hl8ejnY4q6Ait4lcX67XQmeEUXK5jBECnbvT5veB8sxpyej/WoEzdf
VuYvFSJ5WZDnaqsDw6VXFdZoX+0uJ57nGGwmtVpUl7m/mEsL2vYQqnDVvzbl13KsrZh344GKpCPX
/daR2FxgTkxb0gtGZhv2zdL9oQptQGwUg1hcfPhDks+qWyUpC+zTuSb5sY3ddE9TXgE0M/fwvMcv
djCEOS39X7ENU2X8kd/Fq+93OJTPnWp+CanVi9jdYXa9f73e50BDaDABWW55uB7zzxnysKIaAkjH
7U6oimsqBAtJoWCdGqAXXz4OHhyvMHt4W0LEwuT4U0TbnRHQ7owzDWuf5xWq01bcxO6sjnZQA5iW
z7LkmkjTIjQsyD3ore188Ejaaoim3DdOFG2lRPFLg6DKPvyvWu9tm8GQiEhcvxQ/fnXdr3WIyoIE
qXq4DblZxbeDfCQmDiSwuNFWBGaQWcgot8ksNtlukU94x+F1NSoHmCGRhxO6ekE0fH9Lc8lEsiNn
Oyo5jGYdZHV27poLijgEsAABwch5rJePC7dZfz/QecMuuca7VgVYuF99uyunJmUemdZ44PeiVstT
+UcH6fY8e+SjGw4RohChWYD0sRicTtrTQDMUek1sI07kvhIB38gg61V5F9wCxAp0ir0SNc033JoN
hJHXHy31baBIYX5Osmz20YKkc4EECkggiN08Ghpim09hwMx8n33DoKxUMRzBFxlen2R/V9JVs16I
KB7Tv+jiNYhJK4XuKqi3L8d12SUhkcfHLeh10z9GPCjsR/Fvgj2XjtrF+QZcbz6Gealnlxw7SNON
7RnqGCmVokSPcCgbkNkTejzYeCeMyMVoZ0IOVXld0KMfPIuUVoYiqTNrakp7CTc1Ftt/0BrVZrxd
fedU7vmI22MqKR85LIF4RqbthgkWwfP9rbXcwSu3+saxzmuZ86MY0w5w2rSZnIGGH41MPLg9QMnX
kAxuVYoqr4ntRHsIc8UIDkshjrzdwKLyhrXgvThdQRm5wE/LjWNcAtbZ3bI+0XcpeqMzEJtRM8IN
5RkCDNj6RJs5bhq8AVillgI5RDwFep1nv+ufBnz8pByNTLt/MOYHBcofoxUzCe5woBxRDCbwIvJf
g9G3FYknwm1k1puyUA8Bn4gGuYufSWt/w4eXrvIKS46MaYL3NqVOIMBEgsTiL1Ycwzl0kuD4ykTh
g7w1Voy4/wf1STFMwrhTyf683J+Q1nPzCZ8teKFE6GAiJo0sprY4h01YWboxUX29pHTvzAfIDnBP
u49Xf2E7AqAF4cIJY3kh6/EA0N8DYv3FmPZV1CGaPU656zpABW6UJklkfWAhOjOQfRrNsOPAwBia
7LVvjlPO9mZ6P/GOmPjIR+lH2Eb+xMvxhpHws/6UURZCIwclzJwbTN5ZkK2AUAfXqSgojfbR1pt+
m68koOJT2xc7kaVbThpK7qocqgNdi56L9ipSuPk9RbY5ixgENpznhTVTK4LwzcEE6apoU33AUM4P
Iw8iO9mChU7shTijaAaR3gX50rvBMr7l01hnArUsAmkn5nOkyCIGQZXaUaTa+wH+tW0zdIK8frML
rR3PmX6rtAapYCOGJvMm2yus1omOfl/wXll3N2tub35mlquRWSOez8nz70p3IK2onsmEgva7qMe0
QHeqavlf8SPd/MsRZ385GYhuGJP7Av2rFO5iVlDdIrNuxVCNX/xPeM/CsV+wTZLcCaA+OdGmP002
KeV7kgccGa9yFxL8zcfrfC8nq9bQaai1l8nZg6tig+ClXi9Z4cVHth5lmk0sxlNQVhDRIILcswoB
PdDOvASpoioWMcECvKJTpsuo26FGHMIhmm0xME8uOtaGeh4SXF36o/aAfKaWkF5dMyCsvPKjVCkG
BOlKG3Uy9dKQgZf2t50KASrISc+a53FCLzFhXTxHxdnO4LwxQ0oa2A2lv8+b4Fv9ohyDnrIsDBoC
2giLTomwKTnyRzU2Bd3yM1VQ8lijhVyVzmTd/Cn5xDbM+e20GbpNCq2SFB0jk+C+vHGQHOgQbkSo
HoXSovzqCQysOure9rC7/jJeaOPipfllvFoRD8DM3JWbRtnZ6s4lDA5oJ/ftnrA00RZeXfWsYfap
lixe21hTS3+n/7AdbR6jLzD+om3zbKpBCAo9Yjy5TvJzl5gUocJrqLoJcMUy4uFtbfdYO5Yof2sr
6JLAJXyaO3MLJRY0ZqrAAX3nhwy8Fzo3Q9jL11j8iLC1neNnIzNb7GnQxS9R01rMu14p8/fOqa6l
Uv6S5/sOg9S4O0CTTuHO+lbJ45koQtJnaiNWTvc6HUMkeAgti+mjZGLosExnz0rwYMIKrDyqoNzy
yuddSACjCd/qKnYF7UvxLm0D8/CO2VENwrVaiIl8gvd1tNyRTe8/AEguTnqsOk8N4nKNcIKmhVvb
6bDvE863g1FX9WDrC6eqQllX1P7GSblbZuug/hLkO6Q9Vx24SqmI5+U1/Yma/SWmOic2fdon6KIZ
uAjUJEgeA07sfNA/t7PBDMAhQc5uY2dPwy2tJG8aPI2WL5ls38awg/KVy2WHzJAz8UqE8RbZ24iB
jLnwoF6hQ+pglE8vu5FADq3H18YORjjxJwbd2pnyc8rcbsMryURSM05iQw2rx/VFjWGsqLf7BwVU
l/W5knjphzeVIo+Mmv3DEyBWZ4UiVHGhtoNLOoFFPgXr4ppOjOh7WVJNJ+2tWBjokoGuFRnj1jtE
LIhlmKAK6+1R7QlW0J8wtOaPWrC3O0G89OOsQPRPVWmwwAkWIHiV28hfV9tmlvLW6i53Y2sOwp2i
0qlsJhZVxRgPuTr0IcDOpB5+og/7OrQ6f/cafh8C29umgwoyU9Hxe4quauJdsXCaFK3G8oBg0pQj
4moQJaZXx96ZWI7aGcIacJ3D+PkJBy8wH3GhtFvKySmjc5TLdZMZ/DUWnhLDzJpaYFZ/V6f4Yn8T
sdanzV2iMFHigt+FOJphsBOVB+jQI+OfCHOJjpwA/GyvI79801f/96qOIED6W/W5OFYXNyvrdlM0
SQRuIJ7Sb9OIHaDXwm8Rj+kcQWYwTtgLGgZx1htzusewhltUV/VfnLybBjbXaAQYcb/v0+5jTPyb
mt9iVFbBmlkc3eQqR0EwoAD48yFZXufSy7/q/CyvxHAWajPEmKsuDZvAcaFXI09G7ocjRpy4MJj5
G4zk4FrAfciJ6VutPgTnIfTcyi4sfwlcpo8BMK7LXNvxiiOERuiPKtRAqJcM1KqKjiWfC2cppGYs
wo+29CeiVIw1Z02nIGpL+MoQAn2aIi2S1BqIOHW6Lheiirtm/KPxd/uNi6UCB/hS92nxaRdGMJ6v
DHBpMnRMvQJ6LQFpNj2n2aL0kjkw4s/Tw8ZPcrvS8mCDfodUB1DO+ImhlVpj4JKdpTs/aR1aFY9w
B5Iu14A0x2rWjKrvqpdPK69uO8BlJynjiM8vVlLBiQc0lCM35bT7NsDCM7oNEWskTJV2UAn8coee
fyfKGJO9WErfcN3L605etCCd+MoLR54VElbEDBnQeXwAgmtNnO92yo+tnLS1dxbszWiwReD1PlAZ
Xk3/TIvwN5TA9mO8de0YqFvc7fyB9ixItP32YabTs0NxjCV6bwfdr6prNYdc2vtgbgEa0Msq84cB
2si7PRi9Q35azmNc19Na+Z1hu74cLnBHa2bXDhzIzPoO45YI8ES8tr4zsW+/qtuS0b5YmkmxpU1Y
Lvq17FejCLPgILMybqsJCyIPI6ENaYtp9PlBarsCMvpEAUcl88VB4NkHQ4yOKUOLzpFVbGwELIY4
JpmCY/jA+Z3QJGZ+BRl2XJ97UtAN5yks0hb0wiXPVnf9zAQAgEufJAhpdZAqDNkCWrLwFpt7MSV0
6+CNl1DEd/RSct5JDh+4m+rQo09ew6fEoO56wOv0g/gUt7vF990MlgF/RbhWg5sIIyMq2XnRtFfK
XqsN2Iu7amLKTO9bGsnLY/s94hBVO3BoUcxcH6mnB3rensNd4P0kp6cVZmXuSZOfv3n1+QfpEBVX
ug3dU1q+QeyAB6xT765dOEgvwd153Sz5VWyojU80SWtkNaIC1+gpuxdVj1zcCjySh2ufRK/LGBZF
LaRczS6n+9BAiHDYNzvrWyNo14kSSwz1+PhsLP5nZVCLmIEwtR1Io58kfb6rqx4HVIezwLePLZVn
5taXnkVP1zk9uyluLph1BPkbK4TH4QxBMIFxMV/Vz4HlztDQXYj3RnsJ5cqFW5Q1vh4LRRopTFQX
6K4X9Dpgqu1dvzWPFYZ8+T3YYzpifkan671l6iSBMwrpwE0FA+yVEuzIuMlhvFhc1xZ80xLimBxa
ivB/yP/Sv5Drb7UOIeshK7nDovQPQ0Po+xjnZaYQMXN4/stDGxGoSAfLqZxwNOhOPXu/mk5w3A8l
cbZVir3q4hBYNSRXQ+Xd8mFeCNbexlZEUh2HD1zdPkqOkBZKWIHIsoukaksWdjxVTsdLPSEsJ6eL
V0CGSg7SZQOjxxF+pt4Xv59WUmsXVa34rhF07BHBcMSOzHOy6SabH2MzT3UqBkxdKax8FZNy30ud
+k9Z++rIIyBg8wPvJlBOhStwtav23faTyLOc6lXnd8ihgTHz2mQ8QgiKKfxLKBDvKhhQrYBlvooW
BhjTpnWxvNOfKeOpSC7+scR3WvlXGsE8wKw/TmYYtfnP5kaBtybKTlGL/297pJUonlaQt0YyQGgL
Yyv54K72Y8C1z/wxXeNGypD3GK1dpWpADJgK6bJoZrgMaAs1sZymF55+vUfsx6d6ILXfH7p80uHq
iUuFtO1FzxZFsmewcP3TDasRDGUg7phuJBm7RZJja5knNq5umZ1LDJ81pO9FvONG4NsvyMq5Eqtm
BxdcQI2udg+c1cYcHPjdEQxODog2sxRuDNT/DDN3HTe1D1yEf4ekE+NvuO7D3Q0sJXZrKjLzdtOp
tqRZRjBE5dqrRxL5Ztq827cXC7a5LSLFIp4mxPuxTxjUbLP8C3Z7KO+rT4iQhAlD2cUdelPucxIR
rZlELXDSZYNGX7HUvNL/Rn7Qohq5EQy4ujvgWMZZH9iD//xb0BrmXUkG+8KIjVufTf8eGddiOHNk
uG9YzrK0GLT9s0kDzgHOn6jK27V3G6wYrkVkYWEzO0RWaddDEl3OHBL5XjOusGZ3J+NROsCCtYPU
8FMA5zGPNcMhEOjIkvW5b5VRfMLMxLimiA1uzsl8MXJ2fF1PYmKeMRWuES9d2LoGzJdUbALx0qNC
X4x38nvvciL6GvxTF2YmUwJz9VgDrmDlR1D9b0HGFgN24wg27JiWAIElmj88aiKpBCRQgefC5SxU
LVnccw09a6fBe3mlbvMip0Q+BAw3drxwps1mzm8qifWdA5DXS6BG6AR1wEIJSkZpQMR1r08IpHw0
pFpyd2X5xD3k+qRN9hP5qmUrJd1zvSuyTc2CDVebhIVkxa0k+SPPYNvnVdnGA6tgKgdX/u8vfyc8
foyQIYLx24JDqtbfef+elvQX+aZEqgxI0lO9ANzCKVBDPxiqy6nEfD8SifI+BqoYXXXdAOn/SqZ3
8dAxyk0s6+9vYq0K0wltFNg0dTuK7PG4oCWlWVtZEW84meqYPDKhIit4TnwGipGJrkmBqhcmAWB0
6/dBi5wDUWmUfbrrSKLJhCgqy0N0xV18mqv8LpbYdtuGeGcck7aoDgfKH8vVsYn2Z8/Nd+msLUlg
1QcCAXj3rMHH/hOKTqHohbprjXk2e8MB2ft0YpyE0K1vom4n4nwQ8cWGE3Q1+75Hq1WQ8t1kZ8GI
/vb+tnPrxLpslJ8pAWLGxbP69ART/e0dVZbjuOD0o/w2TRO23d28qsv06p78Bv4klsXXGJTTu44/
Qxb5Ja2hmT+Z8Cc7OSNtC0edcTNKHVvxKAW0wb1n+ysI99E5Bva262HvOWisQ76fcY57ytsDoOzT
4CilpQScCzjndGNRyi4MC+iYrXJpudWP1V1xkZw/e0xWbKiDGvBk8vxS03ggOG9jIoZAmTPhzblT
FoDG+wndu6o5KnlhrVkCt6PFFZrcjcQ3auVRFa1uGaAA51q1Hy0/jMVUqxFh+MoCUfZU8tLWus1t
d6JvJFxlKtXktvI5RMZKqXXF39FjW4Ujh4kSoxlXOZ2aWo6hWaMScmkdEgWPL7dd6uA/Ho8ecgv3
dRBnx4AHVcLhaalfiKDkJCyf/AmhucK/6y3R+3PoZFNynCuT8ArWLjCm30q/M5x7WZh6KY7hto8a
N7Z1Pkqkv5axV9u8LrQN/VI5XggC57+2mB9CbrARJBq8EPsHCl8SYtjXkeH8Ve84uyZVjdiZb1rp
qgdQ0R5YnclcjsXNz4YvLVfBwylVhCcVwJalKjz6vTncUFF5yfVYH1fAtbNmDLe7NMV4veSGbooB
9R2xiKe1NhjEmOaPdypJrQPZJrNKvNCMrIsFKo9K3hXK+Yjreyh2SGHfyIvb2n8VAe4cO7FTS17w
EJS+Slq7vh63AIttczJOJ4RsO7ZnipGBsz1/vuWDTsLnURAoL5fLcbgi6Uwlh6/ZTXcIlN+cG7i9
+1V762m24Ym/UiLRF/MhGYs7goL3/DFAlQ46ujH1J2yjvMT4pxAv4S9Jyfj1Qljo6cifdViwyc6o
DimJf16VwQt05KL2+mwNgSFK3vUypb8izxSTnQNnTPKZO1U4Q2LuFSt5dXKsrV+R9vs6Tukhp0Am
xYMm7BXNHNWZnGcyTrCqs8I4SLDc6BnPzQ/tKJY1lw+nLbxcMlAjI0SupDwJn9yYk3Qe4WVEcCtA
6kgqPa+nWld3hiRkLsJm5bia3+uoDWo7tB8AYfPY/WCKMD4pBG0+VPFP4djXakQDxqUQfMjC71qi
PqZGqkkHZaqKVFtIlU1cWuavSmFFaOifyhXXlFCZDq859Vs5l9Q7vs/VcTG5ngJ5updoXWYNU9eB
x3u+v6wYtS0cEcQj7pV9HVY0r0zRWIya22EVdI7eTeSfPiuv06+mLFleaCJPpiH/P3qV/vDvfB2F
obu3Xq/hMvmMZGA1ITMdOydTXkq/FhaEleP4XAdlWXuJw4Yr68GBGkOm26gbYhC5E4v0zdn/j8na
6Xc4rFqjNV8IdjWMT9q3MCYZc1cCb0wWEU2FgLC7/jRdDublbbMqoPFFUHqg9F6AmP/Zxg5VzVYK
sI4IMRsJDH3gEgsGLKKPIYjSyvfUIw46wROZcw7PrwPgMv4y3hS0Mls2LM8v+yG51Qepwg5jJkZ2
ECRehdkuwaGQNbf3Ftb3luIGWl9VjzWAv76rYIAdQhY/4JmKknVz5JSfLhzKchOGmSRllb+1syAo
HXoXIXKOqavjOHqeXBK577NM7XF/XBEW6tCVBtPUl6Su+7lvgn821nzIvdY2rrQvjOtJPBQZM+Z9
uIi0BGe16BGhXRZ1asxWM4Ahe44i23ahuXd5oWIhbb1IeIWOVznrbr1Jh1IdqRNbVYsPllaEwCOs
MCa8TjpZqb5EyZr/oeIc8GezpeqgY+rfEyeY+oIyv/YCA3XH2XxTktP2Hml5EayQ4pgev5gMEHcS
NNqAh73YloMN1vhzbJDcda4SdmeH3eCUr4erEjqPoWz6nElu4K7i+Akx7Lo7mNhIEXBcHMSKEvXo
rO51oS5qr0+3a29crP+ltsGB3T5OqEv4gRwRTgxTfgyqi9z7pHP0qZ6ZOXDpXcKBsZQ2IAgcDpVV
eFpuDN+NBB1MnN12csNh0kqsRukx7aGgwH+kx4pbEgQQkNSsDRIJzl+XuixEIUkhhe2njANkugl+
GKCU2yC6/RRk7C3cRCfnzj2fMZ5ZPtm+AMZuhOKbgSo0rEhT0AEtYCsM5lKeXS2D4bvv2YSQO52I
XCrtg66r6NVcKhJDvdFUmCdXbH9OP3IEyE4qreKLDYk9eCNze0HPBkZDdF3U3rxgJ5Q8+NVW9eG9
vQWcOK/lhV5AZ6DnRFUAJE+vSuKLJD8N1TxiWR0mEI2e/ZPzwvlMDa+1YQwwWOdyw3uzZe9IE7FJ
RYSKp7DMC6Ou6S49zTKgYaTeSBXRa8I3mfo8vjL4h0xuJaL0HpCHAg0gsvmayerfmiR9/mJx7hG6
Qw9YyP9dU1G0GSOhDXHvaYWSpg6kr6Occ2NM+h+xh/v2qL4JN4Fh9wv70nJ6vaP070fzi4I+nn2P
piuACw9RRAnU+sxEStDfBcI+b6nce0lCssJ5KUHMJchqbpPr1v6ChiD1dubSdaou8Vu1ao7XL1Tg
AzibtJowLW7d4uY6pDNfW/cm5ag03egrujwzFlOohTNBrx9ElcBLzYqFeH7K8JiqKVP1IZydP4yl
kQqIKGXU2725DW/0YG67LBAlMMWxl8/AGyNgTUXdBgXRyP7Me3qWyFeYFr3eGIdHgH4hz5JGFnXf
tmU6NOaGI41uP9GO5z6Sxr43HMrmMVc5pw9b7VEsceD/KIT+TWDuHOYvDlqGyaw47WhLCP3e5zIV
wtQHFkSzmdvX3dO9H1bTWIG5FuFMFPSqGE3gB95k9m/UrqCZgFrT+Hr3DLY/MlzHbsJZEgN4iEXL
+WnOiwlvt+KiJrPCQpKnb1TjqbDrWCHPrAHYsPF2CgUl1oZd0QLtB5WcwTsZjYCWY5Qa5t9mAM4p
+kkNqk7vbYvKrAo0iuHBtB4sMJXV2NA4FOZwZvnru7eztDa3/QUmeU6AgbUD2AUIGOHmJGBejLOP
Sm83C0I8unfo3BKiq7oy+C3bvnuTIcxYFu2Syw2z+Kjp+9Tc5WqK6890BI6P3iBPkjtZdpvcEWu/
RePEou6HaQvR3/1h5uaXU9wATNSvkGhawh1f/Juw87ul0imyeqAEL+hWP3p7U0QoXTBhqiRwEfav
+oxd5CZjhvdxRhT6xy2ziEvcX/Mrd0qDRN+BcWOYB7DKptoB7b6cRaqhL+/QsxnKn0HsJ9jLjzMc
MruVYR3PximlCZ01MgQHFK7nWIo57u6kdqd7uQgMuQ4WbZdGSDg1BITVsLcjgsC4mJxaI0hTgkr1
6RfPAoi5AfE6/3Kul+6tQgMauldaomChnINksA79TJKoHq2m4JCO3NmXwFH02FA6nb5Z+B/d9UmH
lgdY97FKgIHbpADxsyw8zUi5GEvmUh8icx5E+Q0spBFDZ+kbw9Kd/Dh3jCFX8DdBm4nxH4pwGH69
ECi16arnlyfpHohebnajQFQJX9vNYGImQ6GXp4kh2YOHDacYbmxuFZrPJIp4DYmozSJVIrYyI7xQ
il7CtKZu2f78BiSo6M4sgrnAdUhio4hpl9n1cLSPg0zgqUqofgC2o+zwzTaB5CxU/SuPRt8TWfOx
mUQ7Li6Qs/vtqcPRpvvAnW3ktkS93C9y1SoDcVkOExaBV4fTHBaU5gasE8rqu88PoEopBJJT5830
N2Y2BBN6lhSY03gAbSzcOZecR5V4o1OaY9CWWWz4nZUNemqTq3XaohEbC4HXo9zulaL6FzKHAtsJ
Rq0cZ7B6XAGEvrQu0Gfr/ZFNUiDnknMlSSb0nqTYN8LpCDhelr9cOntjFMTosUSibxH8ab6K+sO2
0gARh9oeFjWf4N/vOYEutrFWSdgKB9IQLv3A3zM4cEjqnJd41NSwdlgvlnjMYRsKB3OPwg9aqPA5
tAb+TVwlwhMNxl0twUW1Dbf+z8onHOO9frLllwKsxTUg9llcg3tydqUFrBev4LPIuJFgy/eBB5UD
MyTsXdMnbDevftRdJ2n/snxGwJNzibVofkij//O5qtADrMVJL2CQu2aA6Oc6xMYB/ut+fHAl0/A8
h2DpBMWqheyeb0W892Fx1uCHAJHNoRjKBGELBVDV+TxFU7wONLyKZaRRVv9+H1WTKS8fuxNZQ5R9
e01mFNsaEXmr1MTtz199ZnUKfCHDYlPZHTWjIt19+OdJNJ21fmJkFPuG2SRx8neQjSixAI7VMVVG
LF+cjliVoGdq9M3vemv+5a0M4ZxGZ4ykz4KGqzNhh+9QdHG/kZTQTl6NVQAjBQepUvfAAPoW5u0C
3vn8yR9JsdnHnVtlk5Fq1PxHrmgF/cTIWEmYSoIxH7M64J0jRzRvYMIdBvVIxVr22o7aj8OIXZ6p
7tr8R9hKR30a/QqeWfj/wfO78e+qcI0/cThDJ750Q1zamRNnRmRjJdBI9ytDOpO0YwYFbHLnXWgf
ElWAz13Elm09ZXeE9vUSIlEDO9/exOzrIyTN4Op7h5IwU9tXJN4UnguAiSUWquI38hpRcwkstT+/
iR9smnvg9YdUpuLJqLSrMZsEq/4loWKcGcG28xifrcePM54I+DoNgjONPN0B+tKzXL4JkuI0/Fnt
zsexulqHBMXJxank9SQJxyKjEO9vJt/d8+FL8cNoR6w51coLjSOH6cYU6/G/yQbwlLgT6UnZZOmx
7zzl8PES0bALKhiGk5zubWev7FUq8PSyusYbGKg7Kz0OVFVLEqtKG5xpMjf57qe2CUmpx5LzQhF0
+7/NBhJgZYXv7IrKHRbThveQMC3VA+Undax3pdtUcTFZe8TFofA6eNFOHhIF4VzeF9WARaMsZEhH
qdeneOggJ/Ca2hAymr4DBLau/2U4zlvX05D3ovl/auIP2iKdGhYO2KAfDjRr+7QhMyegc8T6gBY5
xRCwWAHg1Ee5cR/xcU7mIzTr9101ADZdMfo82g1NJlJQjKfQt5x6b3TGxf03w7M902kmjm4HRIqV
b7Y3c2FNXeA8mXTylflL1mvIKgzA+JSP1d8Oojh148vtlUJ4i/ipKbbqXGlGQo/Mw7cKljhhTI2s
vwYMTJFP9Q4wQ4Ojh6Vf2zKsuB2oIQdhWqbKRT/IcOvOw9wq6TzBX3KQy3jg5PJaSYyMge8p2l2L
tAchIKuRIsm/CHd9aqa3+xN7go2ZmrZ+n9HWqptZtoLTmRzmKxQ3IptRIqgaimqkomMPXSw4EUcW
v4/dRocOF1c3pvKSIOIGrneSieEz+ty9aFTBWBpfQJ225BNHc26pL1aXV/N3qiNXEd4vT178Hfgt
HHHoSRbBhdiI4ddTfHS43f5C6c6FCDYKKmLYsUymhgY8OnNcDEMYsmQgqC0TJ/ztPC8pQkzQwc5e
F/1MWSkeL7Rht5GIup2vNyNqDWXqglxBLsNAaVzmB1Dh5Yn9NPJhDP3HEnsmDJFq+tkLy0GF5bIN
y6EbfmR9vEekTFfLLdNS2p1BYPggWJt/TOAA5XFWiat5D/TO8P58GwStWfLp2BfP6ToKvQTDKWcW
OwLpCkBDs5wl30CaQKNdE8p2Xe/0cRlcMd86X7tuZPrTl2+uSUsKxcihRNyWMneSy5lLpJ/zDvi2
Rl+Z1O27W2U0m5z8r/OyooNlpbTrj0dRxOrRvSdnfObeubjF/AOkugxCGbbB57dKatnS3C0q9mdw
ziWQr9VfQ7r8/SjvrkVth5c/JNP1zV1XyNkdBodGUVgAz4vqYlINgK2eM3OCFhEcDIpGkC3GOxVY
eW02IKkqywHWbA5epAq1ypQAspujKpap5/WcT5C7fH/EaF5s6LeILxx/jrIknmgA/lIX8hlktErF
94q5BxGRKylrpFoviRs+h+H16CVFXnkkA3chK3ZUuRe1Xc5ZHHFy23iuMOaPlsrkWYCS12HClWa9
WE6qBhKHirl8vJ5ENAWcCKD9wed8T9sClF07rkpNAd9QioCsF+J89NCn2Fy7HI4GvcE/6N0jomOZ
jRP4PkOeHadV+b0WVICmKFrAqyBRdw1/TJD6SW8FR0nIkUhotLt9z/qEzixuYZGlZB92mTrid0sg
Bd/qQQFiXkie+FxNUNo4/CGD6VUVmHIellasB1tSwmS9TcAVIWrx+oFb3cYjW13zsdxu7ZOIyqYt
tnSGSj+rYsCD+EEZIpj/vJCV6WIGCubwXz02S/85jS2DIE5Q6X/U3EgG9yV3yJvy4skudKbwAKk5
A2bOPcYFyMGCnE1XG41i6MjcmAU3vWNPxFaEwKNNNxhs+vNqFrOJd+F1w0vr0TcLNQuuJ4jOW1U8
WLOGwea8NtUwvCO21kEJFs+5Z16If+/rLwsY45onigXb3Q6LPCiassBDGbKbMDb5QMjDf2Q1+9Uq
EcY+vmzL++dDAn0WDfkmct8HDgT81RUzNB5zEtNzannOu7u40fe+oZnSjC+Q5P4OZxqiKvUNSGmX
SvJEewI0nb3GIjcvCS9+Rf4kp8caXyWaYiiSkz1+efqNKdkEqVRxissBZeAlo2g2XHc641dVLFHa
TpLLsP6hVqvUUKoCT5Qbl270kKHiLvvZFrD4bfdGJHn3OzQbRYIA3yUjrDMlv+UXoDrSYv3gQXP9
DcFTLghLQMRyc+rLT7m+sHz/3wtVlTLHuKz5568ibX3QzGQqEqRgLoaCWWLKuBdx8dbwU7t5UL+A
YH4cgHILlOh0P6xipq74kpwQkBiDY51i377HcTbEhJk37jMmNm+M/N+83U9dyMwj/SiP6wNMyzC9
nWLT8Apu8Crg6QDAwpjxO308St6JqkFzt5r6QBEvzh0s/b9ERd/MUpXiNQkm/C2zGGB5h3zU0+k/
BM3szyx9ufXQ+s8hrxTmrsz/VRa60TWGXQ2FvaQxAnBT41YbiCJ1OdKpbIqEuDdp0h+Ktrx4CsIu
L5bgqYNyN7gajNLEQ5jeLbBYwm5Cw+9gaCKYtRBj240iCWj+26nLNU7esd57j+Cr9xtHVRRQxM4D
0BmqDb7g0wzzRf3QTSRIzI5d81d8f/IYEvENOZX012+dOSDfuOfAYwxtjiNupQ+e8iwRiruQ7v+E
rtmTGzVjZ2/Shi+korWWETKLi/CU69Qa91GBOqH8RRhjm7ht5axo6dQFPDc0KtXiiJmLflkT4odX
FfSqXPonufy3izDlgE+LQ6Q1j7sOTaLcmZA2w5GFtpea8uA9AIIQ7m1Icc+5M6yiymyUEpFZlFtB
qV8TfIz2DkV7iwDeHl6/QnC8CQmWLfgTDPyCx0wJWFAvcUQOBgOgCCv91mc1CV+cDcfktPxzlelK
Hyp9bPYEE0zCB7bI8kCzheFrQ/TDPemfJTyx1M+6envtZzM+6Yr+ZlCEn3tFVz10QRODEikM9D+G
OlMqQ7Nogb3eY12eWNZVwC3PaaTxUQmcUlbU2s7UkPJ207Oa+eG8EA72SSut2EMd9Gvt42IAH+Up
+rv7R0+oXyAg3DhD/g0wucKEB7l3dXHlrd7SilTguaqQPU2HnhZCLOAxX7i5z8Uw3ycaHzMah5R5
W9r0m+gNrJv6FmHu9GLSjI8/lOQfXXWgUYY/xV9ksjKFpCVAxhb/P7j8mohP1KJuLQ/dmPVqne5e
oZGOUW9L2yXcm59qjOWUuTh9S9oCAbYtBBqPs9gJoq5lGq12Uj3PmYZF0If5tVmDGsnAJn+9YvH9
kYiCNLEX8yTqqLcgVkYSiTukYJCJhMvzl7qWJSQRyL628QHpULFL22wyjk+NAhr3SMUe/ho9v4Gc
a+p8gLNhdk9QjYbbfUgl8I3wE+nI3UmggvRc+ZU2rR6kbH0wAAd9iL9qWcBkI3mJn+muaK6kZJow
DGxct0gMJNHLe+hHX+Db4VblHyP1HEirLke3W3rOLluJc5sBpbYWPgSn/YT5BXlkIZfLSEzma47P
vSdzpHv3Bxc5QhR6U79AmUx9FCnRIzqdgU1XBjU1Vv0KGuZfn32RHeGLvbE0GtZ7Aa73sqia9/L/
4IizaR2gokskIaeyS2FDZRRuDupMFkFtfmuzUjihx/1r0+WT0H1w1iitzHd+6Pazr+SRxhFDexJB
CU6mNQyzL5jkUPYwcKMMXwRLFTq+TESlxG/MJ5AcLxmFWt1pR51L9uc6vzA21Dt0lNzXWsC6cWqr
TLiAmTRJtVYR59d6vparaLGpLsGKcABwXWXLAYDQnCZWMRyvOCr2UZZXFTrB9Zb2q96pHIj3n5Kx
9U1UPqeK6t7qR03ry9uG3tx3Zt0Co71RQKiZTDRyYjQw8jeMIgJmJvwhb4bJpFtcKeevcyf2DE79
xAtNb3qT3W+LpaCCmI7d1mx57ggar2O/LVYmac9rLGp5oYvRk1LYthwNLXzXZG+k+BjzUboJUkRj
mP89gLRhPFV/zXL45T1/jggA5vj29/uR+RNKnSrGT90Ypy+kF5EpuCQnVHXlw6m7WEA/4LsX1uQU
AXpuOqouVf4uiyouq849PnF8aNdWs7Agyzdlv04fKxbGzRYD4EUpe/62ENqQePdt9NktPDHfr82U
+M/qKvDs7LB/H2hmT/++8H+vP7Pfefg+c/HputTAa6JG/nz4Hts/Enife9ZphCpOPyNGlzVcD8xJ
5k7rVfw8+ZtSfz1dbhOr/Ops3gAoXq24sLyFMIbSqkNjjQFHbPpxRJeBzbnHQFE+2wDJlAmKBt6Z
BYgByaK33N0G3rmpB28piv77DgfFrH97OabcM/D5iTKIgBnKajnlDNX07VSzvopmVBGMbf9RrsUS
mH8rchEjYty5+90JV338e68SWUJcq+BW6dredkuPMzn0HiQkGhQxNQIYDUQa3cq0ILG/nwkNY/tt
UBofdeNCJvgYV0GhoMM56jMZ2JyzZndZ/5LkmtW04aSgZZs2EZkb5yNsmoFJFIg+xC3I0zZ5NbSx
8j0A5ZlC75TTMmfDjiSzZFfXqYtJs+nZ1Yi8sIqgCDsah5jDIEzAXsT52+KMZF2D5EKRugeIkJVJ
UNvXHpCZ3K7jcl8PsTYItUIcAaCY9aShdFba6lbY0z3ypw5HcYe9eflPGXQ9rjwN8OZOM2jIH+H8
3v83CYvIj3eeTuSPkqeRcYv1AXU7RgRyURFNwOYG6+f/FnlxyT4ABrabzVBOqwloQRrZKA1L0MVR
z3pIEzqV6PmPXWx+JeiHnLY+7Q9HjBCJyd8hUaG246Y9OVp2+QQimAI4GFJ9w0pjgloMbO0fT0om
vl3QvGtzDJP4qCGfltvOCaVaNrgCWAJm3VlMhARaCsQMKjf+aT1SHx2bdlt4jZxYzSkFlOSRGc9m
EWg3/xaEjPnVH8eSmOmvPsypjUaXYctACIpMPrY7TBVnhjNLO9jF5cwMlDnj+uaKFNfC0jADmO1O
wrMMS26OmIt5ywEUt7BU0lLTidIGi2i1Tm8EckDltPZgVRRCzCMCXc3jbnIQlhAf6b4apNGRUmOj
lVqtDgD6QS7Gvmc8/sHlYS6U8SqkuADQ++PCBsxJMD4Z4zTRW9qiDTLxwgLXWkFzrhYVmVHa95i4
NEALJNwTDhirCavUIIw+gRSSEa8Tj5dr6i6g0yIbJaT7sWPCf9ERle9tS3blSuR+MejvNDKNlIO7
/b4b2xW/saBaawsdgLA0LhdIDu2xc9hmjDSMkzCRM2YFC1ijWvoMMfsVaS+gSM0WnzoN+hW7/CTt
jwkUf5HFct9/ihidKH6r7bIeN8uLxCes1qG+ARb+diRuOvC5h8317GQSlootrB5qUGR2XLV8S7c6
sqYSBMi/vSoAcda4Ie2tcMKdra5PtR018KYMz9BUiElRNcCp6wbsQQbQTmw2+gwznvwzcneh63up
ynUB1IWHHYYxIZIGHiVIzKrj8YGwXMjDvFqKdmX2t/D6k7jcctyNSLJtqpE8y9KEtYXsvSFzqrZL
N1wpDT97+3ZdFCd6FEh+Hne70glhCR3OL7T3SpJSHA0HK7Zo63oSkfP4Eug0jrBZScj8A4EIoX9Z
aq+EqbXDoR7vQ1o6yUWd6D8SqUgUo4B2JpyzMafoLNjvDQvTKfqEZzLjlmNPT5rmJgHut2LH9KmD
pVMzXASII0kESzH84fqjKYEemb2/PVVtUYw9caynZTjI2pXXhL7SCDvWsLHK09oOxSZCCZO5H44D
R2TSZo/4Zz5G7Ju/JpjvDfgY4f+o+CpLwuONgMtFwwYvPM7EidGwSzs2TWb6E+/W5rQ/h6WrdoTn
cq/qL3Luh99iB+5I7HVf4R6kTmPB2f0/AlocnhMLCfdNRNOmcR5nAieTE/obsDs1aTraDNrN2FEH
9kmAbfZWMi21U0/PXAg+AF4FgwItO1763rcbpa7uC8LRUMSl6GBTrt+zfZsqIX52EK3J9lRC55Ex
0nHh0gT2xAZkQ7pwCei/9g++gmr/GiRF/+NmQl+74xXgoF9xv0ej2mIEfegV1Sh/fRNCmuilzUe1
TQVsOQHTnDKevIsx/5ee4anEzI8lTfLN6LJHlv5q4d0mkwVAJh5shE6ZfWXdrhufz7c0svv0RgTz
SClAlBk3FxdnGidNasi+8cXWwllIiG22msorOsdRBTeKkZCslV4QvsJK9qn06kI/1fgHGEyZRxU8
urliHuG356qgjEXBZqqJDrnSKx26VrMNZYkfyv/eKTpEUPIutfHinJIqqXDz/gMuIyst3l0TiSVS
SAhAXqk7wa2E2eEPDQp9BU0yznNBtfWlg5NWumqCy15nmd4fe7pnmJKIxNEs1rlQAT01lDwDVBM6
lCYAymz0shTmD1ebbSyr+KGSOJFVtIEbbWpOiso/cftHvfzAa4c9M2enOVPzg/fAa/qTorViahLP
P4zLR+RHDGJc6rR3kGqz/kL6JfgBRuBwHaPM4312oYWup9sc9WicZ88AxYfWcXNxSEaiDPl1df+g
nX+CbQLOuqgjRBc3s81n9ScuiybvLy4T5t3aTouJICwCyKwSkiV94jmgA7Wcv2FxVr7ZIUmiuEqq
+2G5+WLomG+Coj27Kp/n2tCukM8LG6rZsXuuvKOb2A4UNFvFg18bnbHITx0XZFdfP1aTVOEW9lzq
RKj3c7EyAc/iQKfRdZimYSXySI9C7b0agtBlFuMnA/a88wZLIv+Ex9o6N/rLcNNrtYeWex6D6cq4
Ld5th3qY47NzUMPnxZtGZ8C1eXjDH5/hozXyC2Sdz6cAEF4Ahl4FVfG1tsDqWYkq1VQuLYGeDCGF
zR4qlybXT92y6lzuJzdaNZ7DNq0DPS1B2p5E1myOSypJap36GDeenVOTInEF6Kq4ZtaFLhPovoMM
Om029uYoG/JqL8QeYA2UGasFy9NN7x55SEuYGMvblR5GHaAfyJ6F19e2IqdHtzWqQB5/fFFyihqh
UW6yTpacOn5GCPHJlgAU5VOcuxcR3wPvrpt/AVD/4SQ/EWEc9odY8zD7369Z/KkAoV0RQx2DMdtN
+cBuf8akoGq3fRz4MkvK4ccH92B8rYVel0PZZr3n8TS216OU76cH2gUEulkT9PWwcLSfsU9UXC6f
z666FOUysCayXn77NvAGTPfoJc2GmrKLvndwQWnTLCE0PVjYt1A+5FkFkgboA4pgYJQ3qofgV+Sk
gmSgdLO1H6mL2Nw2Udu9D7yTegBq3rBCf0D9etBhDEhi4QxbiI2q3jSfzY/SEdbNEiLDdI4P/z/z
6UhHn+inV3XKihq4aIOQh89YZjQ2wTrq0IBu0lIciaDnWw5hNY6LqU6V3a4FjTDGKf/8EFvef+Zu
21h9TT8E33v+2CftUKA8Y4b+6UAY8q25lsXb3ahgHti63tv6ohu/7JwQPBs1abRgjlB4Ccewvb5e
sv9KtejGMiFpRtTBHG0bDGBJrnmgnnu0Fp4qlbluwrRTbBR7TEPzTwm2ieX7uQRdzyyWQ1p6Foh2
vz5JA0FU5qFp96Dtn/3Fubpc7o9dyca8Wc2PgU+2dJmRQCokXocF0PsFPXTrtJUOP/flLMDInLBj
4uniDWqsEJN+wpQpthouE2+4QNbAyGSA1stAsBqo6YG084nWiw2fUODhjDBI4wUgmAne4V0FcwBm
75IqQHXGwteFD0fFIF0GkojsNp1I0BUsMt/DkwHgYw1NwBHmIICAG4ZyGNKE+yozJQGvZ75zkm3s
lIqkXopYNGaDOyUUH394O+gnOPowqXzhn4ORdUIXqXhITec6Li3Oe/kh+RmaWVJ+x4cgaiBv5kGW
HGU6LNsZ8bzaiX/0fRGhE5I+ma9rItkNW3YH8uGatAwKjYuWho4dJxm/E/uf2dkHMJnRk68P6GXD
cnAdOOTTuO1bzpe5H+Web6+Z6wRCQMIGkFqyBItqYFu3QPwsFBhLGCqK34nNHbkHurQO/z5HhOe2
IdP7hwbozGfao0VAadYNbQu5RzE+/IyntyBOGav+RoT6gRc3GBQ2eUlFXCG/hPxwYe/rGE1BG7A3
D0ngK8x6fruTxL4CClwrC7vqhEqDebrKrhR49Dz3pMVTkG4vEBvS+oTAlecQTKnMIZkw2l8LoWM/
4v1Q70IYkCW082The711zga0rvcSqyneWEYxRIov3MbhxSV+3yqbx1rReHZlveWXyTz5QOVkzvv5
wygYc7k7XUGPltNUua/ki0zewrcI3jBtjLaOs8fOw9ansAfflMa2DPtotOJS0Itb0+FQJYtzftj4
At6tTNXl6+TwkbR+MjCcXCDxs46LD1usoIMO/GKbJjx4sVy7c/m43KE7aWS9BuvuuM3MJUoMzqa2
B00k9Z/lTB4tLD3igkztHEx9xHz0cbhJjrjYn8/RxXHDc0kdVI2Ht281l3yJYDhbX/nza4MyRjSl
2eCRDVC4fcow+lin0+ktWNRIU6nCa3cOjlZVTWYcGbuWWsvDTpuEUwQLs+AXWQBPherUBZXaj12A
KRgPzSMb7o+HhxIdecqPG7Qg1aYCyScihxn9JrOPWbWRIgAVeMwHHUXmGwsLLgqG4UVpMsaMXOPf
lQjqNGqq3lgPUWGixXeAfkAizjDg3jVgEghLW5kkTVugYpslkLWqLvbCFqL7Mc3UnjC6X1SVrqz9
aerrlmYRkQRs82lbxRG6fKBa8HdkOmK1xki/Qc8a//TXHZ7OY5dTy5moRLk4WdvcWXsjbAjM2+rr
DNfrh2WjJ4ukd1bXeYABrDzxzw4k2U5ZNU4Wx9A6uKlHG5SaqP23AyxuqHtatN60lQUaqx94n21N
5a0+IcYAd/U16Bozj41QKFN/4CvTTwpIMpuiUH0SGVxc7SxdODmFAipJcTZl/YU3HB4itZUPw2yP
ou/jwQ07uWGXl6a6aAyEIIMFMFg3SUTXWO5oTmAlKXTRdbfgvxaDPFPEvIPIzJFjTkiQEZhffw4x
WZ93piBZJ4NgVvQTfdk9woOsTI3wz5XSJNZWW1TUTSufeLJWRFjlOpi1EuqSmnc08tGu6EaRRJ3I
zcKwwhyj0e4m2YyZQSLCB3gg0owMqLcGzMZroRdVhKse9datvuwpA6XT4IT8xLJMH9D2juZJvmLe
OdKjT/SeLVrwrVQhm1WStu29hUbG+MGmhhgl9uUGAA5ps0Y7geC9bNRxZ/dXNw0nHmFHjCIpHPfm
LUvq5e7sMJLaVrqozBEhO3RIETKqBZ6tcdo7s13laO7wg4cstJARTsgjATTOomLRjzVnrRSxVyUx
qPBtk5tDugrISIZvrnkox0DekAQtjUI/5klcRUwuccHAiOQXAgSlOOUdUFVoTVAWD5UhgjjIq437
pO0/ky9KI3h4dPwvJ6AwLaciID5o2br+Hx3FZaIoVsCFMwTPuLZ/QtDPydWPvVoGcOmIITeCUzsI
AOygau8F22BGQg+sxApt5ms+4MR98BHWUgHeKiJccyWqU+QQHp5ETVHfRwj3yucPpkL+MSWR5U6g
qXnylAflkZuYvImcJr1KC6+g2IUEVZP3ar8b14+Hgg8eZ/xfjUEzgq+0tfw6NaXaHkgt+MNFOxM8
S9ZUtr5hc4df1b6EanQQsZVSKxp+BK7iTbhMKiBbpMmf0dBONZEitXIBSYN8vBSE9FhPUmSC61qU
Cffw20mMb9+f3dF9pv0sHhD+/spE1U01o/p2A4uMvgYCyl9bPe1uzl/uDl2I4yUNWQZyWRnh4meI
Kz6n9YU7F3BiqTM5Xi6gZpsdg4bYPDC3gWRS1uZiEVYJqyWJMVlDLAcBkSgFmsG7iW11G6UIy48r
3GkZl/irT/1jPClsF39LKxOufpF+2+IZaMlI4YS+DkyI52tGQgseBRIhYVsF0FUVcWGuOYntWot8
B9hPrQZaXc/QlwU/s4yLIYHQEdcuqnKEGRCTRx106UGhLyRUlnBHcan7sfqgCg8rvYQrnEMPmlPt
ZZyN3ugJhIyNsyIYWDQGdlN0yzmsVJO2vQgnJV8BfYQfRE/8B4A9pGJV5GJmEnRzO9p9RpEVqv5G
ruuazE9LSb8UzoQAsFeMKB8z7nwiwRe7b6zYKJj1CpOKeby8IuSzEE9DwQRT2RUpYgBrh1akG8BV
K4AXCi/9o24xtwgKKWAvUvbq6QWghQanHmwt9P1k+XEO6ysJYq2ee1rWnAtfRSzE/QA1OwO3Qkr7
C04os7fhaPbtArehmeeulQTdBSJ7eUq0Ywwq8jmIRwAr2NRdenUHv2Hw/DD5oK7JgqSq6f6WpzcP
9dEVvXYJ5GBJXNKLvBeuPnU+289QVyaxv3ZpUJfhDMNZ/aWv8Qs3RbwWjyPrTmImUcguU+GD8QBJ
FQs4ecD/lEx/B/aRM69nPPGCFBgX9/UdFKT2kYeHpiB07eo1o02b+1xHOYKZETqNq7ZlWPNSITx6
6xdoWtWWSsqHdh7rYAUOytzVtAmF1/HNdC4bjSqDVissMlReFufTiOIGjSLTQSEIdEHxO55M+6CI
5sthSEI3w72G30lEZU+Rm49gILP5OWLtoFJhc8cSEd2RrxVrmQfioQ36VIipmf0PeSF1IhqueJ1o
OMRpbHDpnZucJJvywBIV/Lm2pHOwaXRKj0oFAthN7XV9olYKfmuPfsxr/+8+7sm5J23F9z9d88ue
pN5Tl7JlAqUES0y/lxclgD0NqWuRt/j8TYUCUVBtp31z1Y4b4/t8rRIAQrBpW0yvz5eM1femirTU
V8MAYK+nKyuYcBfSzK0OYMGKd8E2KiO8+faHG21X7FXyxtDMgSeeG9ZxNzPn5u4kNekn1aPHG++p
cRK7GW15+HN8CWKO2ud8tlahso1uV2cG42GgpWiMO+tjbg2SUtyn7oORj5CgRcSPoyPoXplJJQTl
pwnVzaheqfoyd6hmT8zL6XDgPLkMBCutuwmkMEXUKc/9Ft7vyafj9V4a71Ms4gHc2FW6DpaCrrz1
yezlc50B4+OSZTTI3pJ07PC3F8Zy+zVDhak0/s2frw/jFKWX4iCqvppRkq4m5Lkg1p0j/y1hhuX3
ihOgM9kUeulGEutKVT8jf058iE0CxU+CCQvzE0qR6dH2qpDFZJqGcdPXTxxfqJwF9yQwy0tpEQS7
g7dWoYgdeXOgtd/ccpKwtYrvz7MiEdSRGfVxwPmT+fqDzBGgOqqvyb1PHVMvWAxfE+T92hBSbEls
WsYvmEnF95eX9aZHyUSvup2z2QpI7KzYaDDq2JB94fdiXNJiWtGS/8mafkoRHAVYzncku3jZ+QD7
QkNZ7JxMvWaSg0tVYr5EIDRnJ1+Xo77xQeZlgbVq5JTY9Vh5P+jQmQ0hIL6E/hxgKNDMnsBoIqkt
Qx09adK3mXc1K9o/kzzEKj3meosnRpFIQzUH2TIWdFy1ddI21YoPzga+zxqB7qCZMRzNi3Q6yb/O
TbzQCFsle3uCOJgGzsSY9exZoopTQNnSJQoRX9wzPuYLUeLyK6Xi6ytCZXizaXc8y5Bru+Txt11+
9ms23yWlSsIZ5u6D7sWzHzFdAFd9MsznMbMs9eXl1PHKGSb2whgW6jft1rhckYm9ezPqLhug53Ke
Q7zGllsCC43YzAr+tRtVv/2HxdVfWlE2H1rAKI+5KtOfMjSs7Rh67YFY1SiCVx75491R2VNCf1O1
AdWKkboH/IKYv0zBJeCgiCaaSGaQtw5uD92IgqSLiGiFHNwuwPOHl4OYBK73pMW8SZhJ/vZaK8Ov
NpNqlGMZN5cH5GzGhP08q3y4MWOKMto9Y6R2ntWMsCgmlkHYR9Wg18XBMAnDVty/CQM2htWu3Wgi
TBUt2gz/7BaekDAX9uZfjFjEp1c4XhC3vW5a+2eqcQSES9qaLNtDeq31f/c+X6xPkGiC9tIezYID
114kOugZzr8opCbFTmUWG37WwXinxEjy6YWbYgLmfUzDW/pkyfwoRUevEfR1BfOM10rdetL7Pxnf
CnEHwsIsTDg+qQtlbOp+vPBYZ8RjdgN2Kf+HxMp7/mpFjvi5qOfUE/QQXHZMjCoc4WYl4qj7sj8Q
JPPmQ6xquhoaX09RniUsVH1OzsYGGWaDCyTeXwgSbYbAIaSLQe8F1fNNZgXN3t7HHPCH5v3ySyQe
9eUUhsbC7pm0cOlwxd6KaqaFasl7P9d9dIPqoRp+V7mIEyRt+OPmnsi1pCgCF5BTZv/EpVaFHJEm
jRqNBBOj15Dmp5s8+PCMdyvkVcXRi4tAkYXUjh6+nP4TXNhORTJ9CwBq4mXzG3M2BF+65iMT933k
YR+VUzWBL95GH0hPcsDMUh0a6wCkG0NB/86RJFHvvPE90VtkAcRrDn268N6SBtIwz+99F8Ex4MWf
m5WGf0GR6wQ4RQJ3fIE6X2F63j/rjFlYqh2nhVHR4aV88u7XO99r6Ov7F6bKjbOFFvTWca9BWyUz
wFoTVtUxDRdJjUPd1dPi57vAZnWgCw2+IF51YwNB9Six/0hw7iytMyAofHGI6jklvyg73WmxPE/O
sdtQnvxdakPxcY93HnP+rlFg9zSwnCUMOIYvSdu+EssTCcPGzlcI95lvG6GKf6h1U74XjgUDqqwb
8Cv6yZsR+DkSVQn/FO2o9PWUdRAS7V9gyJxysaruEPjYASEXb4BJQJEX6CrlKTJ9aukMIddwZSTf
eOt3/3hocoyhJ2P7akNBQEFHMiUPsES3BFi5P9cVFhDv8CSk2WXTnPWy0mUhXURJ5YzlM0YXS+Rv
WISa8AjQ//F2Xe2PX++TTxlUSA33pgg5ggTDouvt2vEvsOmneotxqEBNDBzqDulDWcw9+idVQLBb
oUeL8KRCnkBbr1H0uHbL7ocT2OTzdjslHTwkXTKzixmU69Uq3qJOSrBvxZhE+MQWI72FcJOthP3+
NGaY4HZ1yGWMaF6uRUYz41tfnQcs+TqzByGRCgnMJS1asWrm7/rEDv5JLaG20S26QK5PewQ0C4Et
++qCMCgH0aUIfi0C+uSXYRCPb4pa0FnhZcfN3V8VHl3aENzCh+AqKOb/KkNN5Gr8mY/+vubxpY48
LrrWDnnzG6C4XiQsKyr7bhNG0UuXQgaH56Te31b1QElfcv231KpJ6d6gf/pmxAnvq+tyrM8wxJEk
hDanttxsigBFvq52j0NPMoZFxqoRhkc0bftSoN+Uc7N8YvBxVQw86UmRcA/pTw1Tylg7tcAFSX8V
x8sMNqNV7koHCdqC826EIpOKHsT2H8rXSNOe4+QMvmdQzGbFjiB6G88yuaCQNmQagfw+WKpWaZ5q
yJQ6Jl0oGYabtDbOYj3jQ4l7YezRCzzfUxMr7p5rFSorsS+kmxJpS6g/so4H9G3079VQZK8ufkel
fF4trx9aKsccfr6Dgk1I17w6jMfXpgHffRmGTy9dyv9bny6rJ09oI2FWwgNo6zIBqba92rATT1Ux
Zev6qczFJsqmIDbvBPhGjh8Q+CUzokyTiHFIjSUVmnEKFwbWPwBWj4JqS0cBKnefbycAeAPu9dca
sgrBF0fZWYoVdpAswJypLlN6ggQCwjRifL6jgRw4d9/Pu7msooCP4TO7tACZalS4a4t/pHldvXsk
uo6c7E0VADmEDSeEex3zOzdC2WXCHV4QOZfI51vrfiSQMpBRz7v8ILKUU2suArfx9FqGzHaVg8Ff
f2m6UyHQf3i9VmlZTqBp///d5AfO4wNhd66tffUAeTfYBDaGKZ3T9wmAFP2CVmoTqwQBg9dBZyoc
kT/U195sUDZPpDzh/pFmO+5Udf2rKkvwD7alAlPGfHCCih1rtv6nS7zCR3EalunJ8eTaKaKPK8i0
FkRfg91vZIuepw5u6OmYU1SoOwv9Q2fbPCN8aDRYx9QAMVnguXzBj1A1hRjKpRN7gZEhG/Hrxl9U
HJUn1U16i0etYUuA+Vyskm88Nr67euLM2dOF13bY9EMwRAfdqHiPxle5G2na0xzbRcAp1WBpOUkW
YPXC7z04Gim5l1VRgfIqr5BfjCtXc6yKQt3PIrtiZ1HMM2K7bE7zykGi70bb1U32TCFG2KtLNT/E
X90h37Gy9rsHVrTpK5bGTdyUcGGpbhSSpSVM+MwK1Qoy5+j/+6XB7L0aIQw19ZI0vY7G4FEyyALI
HY7wk8aNqNQfqi+IRZJ+MzK2BvQ+ayoeH1VqGUCJmEqRPl+iY5p0FGnwuc/NAx806HKtLauIpcuo
5ujYxRpTZTyFGyF1RWCPO1/wCfwG9+OVsj14EchwNHGKOB+4MYYENDIGzui7fjgjiuIPQA2tHoYf
QLQMHuET6s0XGWJf+KXagGwLvjTohe5MBf934pBj8Qm/d2LyYvHhwZ8Ore4um/VJQspHzzFIsRub
KmDkvVUUYtfU4WqrfZwJJaro2g4WydARbV3nzSMEAd6Od5JFA15Bm6EVpWBgx6KSfIAd0x3tHG04
F0Mm6dU78UFbK/U0tG2xq9zDb/Yq4af7km8C3LXW83IgAW3jw8vCcY3W3T0tTLzCStB2QyNVPx5y
/lw9rS1kLN59llq5RfFiELW2abXLGhvpTtwiirTkd8EQMOBsetfGQPsPyfR0nG3RTNrUxUuqbjue
o0AX102nlA5gNw1z2pYlDYZxmHMq7SiqfIzOcI4o3HA7nuFg7oK8gUnSFiA4dJLMYWVaFed33eeJ
fKVSZ9I4l01hposuUtcgSn0b8oejjMJFPp4Nnib+SAnt42Cy8cDwXeBljDfzIKeB/ZdIHDHoSHcD
3OPvWeuXSmBG24sohedzkPNNY1UyDZl4JNxN2T6PA6htaOscYK4oGFZBlFJWosG8umogQW8orQAF
GhFtXcKvo+RnljFiWutm+itZCdsAMOVcvhYjfZ8XcbjNUJNATRGa/gphIGD8fmLKRs6St+1zcLIi
44AO4adoSxo2fUW32Hx4yZZAPbomoMxoVKOjzZBpl4lSubadtoNgLspJp4G4Wps+nraNsq5+GVUb
wIsWEAwsOZwOod7qgXD1JVLP7fn9euANIAj5DxcPrI8q/hqrfKUMYWKwY5g/LO+AuYaVRBXf95g7
VKvqfN2cGiwfCiydVkdqotrsrzdgLLTMmSZ1z1O5GQzrVwKkxWG0DEmIhZfXUyz2eY4ek7lDjc8G
zQ5aFJsy7CrzIIxUhonLw8kDV7pQ68rqWcb4fqTF+9NWevNWwskM2NgVUNiCFG0404BtAeF6ciZJ
9VYy3/WXHV35ygHsmey7dZHEQ1urvzCrWOyEncfW0kccC3zKdyDxRwyekDP/XeheAgneH63kD2Um
uk4rAYFFLLQf++3weaaY8B/x8F/l8lMasciDzw7PqOpnj5E+tIDa3u4j4CcVmIXytp0X5OYq6bZJ
G/RZCeipq+Kw8E/uMl9iCeU7KZnRAq9l47qxLgipBx2fOkd+tq1ZcNIuAi786fbUK8LYWQqt0RSI
6WCs/JMNClpELhUE12DcUlcZ1xgUCX6NXlKMpM8HpLeVOykM4uO6SxRGnUiH8etngkhRJyupbVDd
2AlUf2uWBpCGIU0RVwnp+DxNq3yNPZmkMDPvafeXjkOWH2P7SHE3i2OvHrWqKmYo7sYlfn4cNPFU
h6m1dxolkw+ldWkzfnG9t1LR4CjIAooD28FgUEqoVRHXV/kYyAifaEG6XYLpigVAkTiAfSme4lDT
db7rxJoGOkflXK0KVooUT0opxvUrscGnZvrp0iow1dAULe1OTvSIVeVY2Lmh8qiUAHXBwuVHH3mG
QN3V7P6GtqDY734DNweN/taYbjHzXJx9CGz4mLYlDKrt/gYnKTEhPcTtZ/hv77dyjyIUXds3lP7Q
ZeOslnsIgD/xs+nhFImbVnyHOFeIPzw4YtbjPXB0X7EhUl7fOtHGxBYCCFbATRqBnWN4+6T8Elet
8Xx025A4+8AuaARkCO1FNPTI42YLRrQln3juxmcsHTnzkdauQZ55cLRRiEyFtoISq1wzE7BThap0
4AmbkBfGlPUJ548+UndKoVa6xi61kpwBsdZlYl0LjMzxYNd6nZeBVFIedtjNWJH0bV0CtPHrVpPB
3jNURroH2fNdVQjbgK63T7RMeHdzdVugpbJ3rOMZ0ptwsEPl/KZxoYB38Mi4OAVRxd+/u2Ra5QGm
8R3Ampz5hM4s+9Zx2ahQKO8nOsDO2fCb40NFpi+1zuOV9jd/VgsILNHl8tjGhV6Zos9PlNsuQsgw
AOHKRChZm8jSgwN09HIBxdkSrMwHZDD/8Mr/pRGHc5t/S3oSp1InSY/visL8UJm60dijc4dzjkUD
W5nyixrqlQ1bc0xEm+JfRVItgZ5oH5zTXdA1p4zVXZgW+2lMTosqt1gKBRaHEOakwHnRD9EfJlwi
WovKL3a7a9X6Em50O0DORRoHbQMyTH9lnwXJ+SHVMIqqaUvqpPl1C5hhKBPzZt+DQeJPVRB7ifN2
PsPVdOm1BQFU435cd2SxbZR0o9jbpw5ocQmvn4KMRm/ZF0yZEYQRAzukFiQH20UtiukI1OShkIa9
qLciPiqpS9JzSRfr6UBhkYGrl0wbYARq5pvXXWPMbmXMsewgdzLkluqru28sGKU+tcaCYXEOyHQ+
O8U5tSExtYPEz54CAmZhW88f2zOa20mxhA+LHFTM+Vo87TfbvcPMCBwHJaBIYQYXc6hLs6M4NqSD
N6qrHtwwZnxJ9UwFaAYFjP4gj9qV1JMTwOgJa8NBylHUIM6IIP7yKNQXxAkUh3Lk2L8FYqLx8Ctf
Cex45wM9v7z0bkluuT+16GhRKgBG41pdn9Fo8En/kkj5iKijJFZCsg1at2AFZ01qeOavRIt5Lv8B
hNXB3DRO7iBmF83lRE2bS5XMooVtSE1uOqSvaMvdRHyXOmr6xn6xPSPeW6NmVo/WyQYa1MiTo5Lr
fd9u7NX1LiaGO4/REWAib1IFVkKZl4X4HTOxa/WLs2/Qy8LljbZ3ZQ5+fK0g5mjyzXjNyCLMUmTd
wtd6pn00qWnnaYc7/+9JMOS/AA3y22FWhIBUnHICPArliczJPcEdU0emOHfnV4mMvRPRZ2D7Ea2a
ML77WEo7NnEhK1COtX1jig09lCW5uMNuNVGyyh+v0nMIY8arHr0jY16lSdMqpVFv/Abe1dcp4E3D
GVbkWOwTBrFjZvRgul0rnBDu374XJAaWVV93VNgnwWqVBDqhoilwmwAX6i9AtaJ8xj5VFOsGAVj6
ooHgRXjusgzV292OX0Ghk1zTsExrBfMZQigewH3IajUfyOqcoMLQdncbhvGf4C3FWw7a+Cuv0ldk
8AdoGBm1mo3MuNx6tKdtP1zEI49O4w7hdgAdG5ET4XjA6dgOpmngWCeMi9MWyp7wu/DUCBtToQI4
XJiyo0uQC5lFl09NI4PQRxUiMgOtzV0eSB1MFoTD43kcFtu0ZyZQx3lNZn97HljBIGRHRaWYFlnY
7vSUh6tNVImc/TY3hp+9UAmEXQnPc5v7TNtnyfB+ZO4LpxiJIDWIzMWCFpT+rgmnsgT108bXUdgf
rNnmsI2cHLCFIma+tc83lzZz6IOxcT+tBesbiEe4vwZu2x2nMlMeo117QeiiOT86b4mkwfv78uXO
CHziJKrgbDYwOZ741HeHAwbACAsBFLuNnesEXDLc8hy2H3DpWFU0V22+GWnNMVnhIzSLXJVkjOe7
Lc9qvaCUA4gkpuzFKGEJ/z23dc8S/38Q1s8BpIdGV9u7Bvxx+sEhebdrO/PZAxjTY11bww/PBKXb
i89v+xj0MZ0Q8PSwXbGwkaRlw2GQuao/yhehvbw9TAIMJ7ZTbvU7cE0P/wsaSEdCRvIA9VUNxnAO
51fKhS5SNsXN0l6LdSu59PjTKCzbB9If1aU21tRzocNXI0ll35s7h33XcEL3TFX5UfrP8NbMOyKs
CLucwNEsopEmN6PQ/UkE+icj2s9AFBlt/5wjh+ArnDwPbk/EfvtllwHN7TYNqWFUJbwtRwIv5McF
hAO1eoCIrtjVyzqxmY3Dm9CyeSDUihEEZBrBnVqPV+XEOUC5ucbJi3PACKIllvxhb4MO/tguoO0o
tON2kXvE/IDkoOyRmhdhXqkqsgI3/4vxkWzlmQWENd2EI3AFW8m17mxRmL598/FaR/Ii1lYlXYyu
Ed+M5cDUMIm2s0lvHmeu33kEHWn/nj+iPmA7dDoU5MvbAjXGJtQDVCWXWA7QxSgHihgzxjYfCfzN
88Ypn2QTEnWldE2vKw49OI4KTsZP1IJGDE6a0j4Cp6Hz8b0/a0jaQHgMMrLVZ0WtGowvqoAZRgBq
igoWUdUYDOqMbTT6IWiEZWB/Ucsg2xjXDOpTqYFvHUpzM9ZUu4tGI9BzXmw4bk2jqc/OpWzI9mgY
AgfBGn1nxWa5u7MHe0QRqpTAZ4pZY6BHDomnwTpuNx36VLlYrLhwzosW17FiPyoXEzRv1WwbZm5A
4Yr/w8TW4Q+Vz04Y/8J7ELiQNQ0Tk7YU01+0CFD4x0bRKw9aMFPsQHzNiIq/12Gbay9jlreE/K/w
One0fXt3bvxe0ng03yjgbaH2QgAWYJQcdNJBJAUazicU8Yqn2yG5KO/UiIw2X5QFinOQogRxO2qF
TPboj4WjCSWTm7262HIXps4nqPtZyY3jkXbElwsqXLTn6DImHBOUFDFRYFa5V7RaZ/Nt5pNBjhBk
w26dv0FZsDzT6Od3a/drGf6z7Sy37hnrQchhOGHYRuKPCfRuMkPc+75YutTjt9lOgOXraJAqiNHX
L9Wpu60i6moyRQh+ETJ0RiiBZ+dxPZOXLRsOpjQGr6pWeWOizywSt5e9DDo0UgzV9QzCHZ7sjelI
j6BdWHP+EudnEcvfsl7oJWQ6bAVq8ipZvugtYx8ynf6MRMp15iInx/PvzzBXQIgl5iz7AdamqSrg
Z2TifB7vwfyXsYPSqC/vm103TwP48N/7OLBGtQuFtY2t9m+infCDD9RzMU78dTb0F6h+1Pmwfb24
06Qqs8eGYiC9TBn7nugYLjd7Giml5l1P9uAxvnLkrdMcygPJXvS8JRcYyx6uvp+Upd32X0x6hjOu
GOcd1OMuh6bIUA8r7iODg9VX1sxw0EtJ0eERk++HIesi+flGnuhA2FXltvf9ADCWInpXlRH8Ude4
qx4RtFqTkS5tkCbMl0oIDk7PkS0k7knFXi7qrr0v2g3Jb+ZNnP85yaa7SK7SGSjguBwxzs7VWzBJ
DkHooov/OmVDdM/3pzlTdMY8uXemsflwCpb7gOBaJqOMc8P6LY42xWRjyUIvVl1KcTPIj5gdZt1r
uTXiPntoZxSrWIzSnnlWpLazWO89wDvwI+fR5D1trJ/CAtkoUy0kdKqRXnW2Amc6+ynCrfQZX9R8
30PTVCFBTYaMwhks8N4uxM91KgPWB38nUeHoSMW0FnDQKpTUhbscCAq9k+2hmYBhv7i59aY+deyt
gPwncYj3zCV8da0WojZlSlbO+YK3aCqwZcE+U5XkXbiErDuPbZ1npKXrZNi22DuNSXN0m+HP/C5v
E2vy3yG8xRPmmr4gil3zhgwVhJvU2St1jkCoiIJ7thDCZccY87hCqrD4x77U61lQGTERZO4CCQJ1
Wsm9A1dg/ncRTjRQKEAnTJGu/qZvAt26D+N49MUuAD/4oMjoZNcvspXBEgGvABYw+7sl7eJmXp7O
uboaCtTfsNGR6Hv2eWDXVyMXBa1k9vryBpzK2iW7T9ey3qOGrEqf9W2LV97w82KvmtiYP2fRipZO
RYFkiPezFqJ7MmzG4WoQXmFM+GX8dIhPB//qMe9+zSjYK/+YYSFQt6EVTHeGUOiYWgthP3Lovm/6
5KwE72TsLN5JuBuw/68h6V1m8M8codrKOl8VsfkEi+Zw86mCtarww1K92k7hJW0Rg2SbEnnOVEQV
OEVDAXcqk2Ic2uyGgGh6Jy96R1JZhXvAUX/omcWQ8t2Byt7zIMtOkcvSGQTSVaegl4yJdyhFWmDH
qUZU9vyvc6AVdmgblSD+p8Lhx8EzbTjt/EddAB+vZyRl6Ux3SqnbnMgCxewWbYU51JndfAZjvQ7W
cy5UVn3ByGZMiqFvvJK5If1tjVQP07D/BCFT89cfFfneRR7Lm4T8zxcNh+Fn4ILVlbuzF51lWxnx
1j3xm+a6c+j+cn1xFZGPDsjWBn+IjDVcTYPa6lxadXrFn8822AddFNfN1SKXk9LVYOqzyBWIQZIY
OPDN2scycVIANjobuA/r3YiM75F4PiKbvv6lZbbZsz8PJneOjIh/s1qbYuyrp196PDJ2guezx5YI
Hc0r8sDwuuGwbKd4vINx1TU+t0K4AkI0nJ6xc+FrOc0CCVgQJm4lubqa1RMFmcwNH9X901H8kkBa
9jKX28BY0OZMc85R1jOWeVsmSAwAU1kD5ULBPOzIeLR5Aod+ztBLVW2uBH9PqfvEA37iBTFPH4+E
KAif1JLudkkXHBYR8qn8gD1tVmcqF9KXl3uhCerYnrkxIxoKMLdFvOxr870C5g3W0CBLkLrSGCcE
RzlGiBB5swsYh0zL4LY2dlwTCVsiDrvTy7VgknJq9Lc9SDQTRmM4QBC3jn3Cnmk1RaoIjQBFev3X
Y3KuShQG9I6VnFA8x35NUn0p/TUvDF+HHdAsGx4I1+a7WC/1+3jz28nDf2IbdP2u7+yTA892Gohp
p2aN46huZJPNqv1/twWoQx5M/drW8SFZPXdWj/dBZnkPMoEKWtEoz1NOxGSYXUkerqupEOsDBKo2
lfXFCwA5MS0UPvZcnbNaFj5MT+hdyBGH0vMsIZFIYlVaPCix2u2+NZVN2SSYlk8yBPWyzLcHExjo
pQv3LQ0D+nTVpL84bItzKq2rIUc2vEPdRf8zhhDQOVnBlnAwID5cQKTYMcLNacqwPb6G4V+4XFBQ
lurCvLik67lvkgzkVoqXHNOWtPTJn9ytPuk6aizpyMuY+LI2oe1YjaOjrDxiXmY2pLO2w/jFFqOK
Tfhgorj6cVnNgNbAbEk+bZVBMdHmygu8UzAW6Qkf5AC1bi73hkhdWua1ra2bz6WS6wSOrQYKEVjq
SkO7LxTcDs9PsN2YLaTX7Q4R9zrM7B/utRvbrQA6OOPyrj0nD4Kn31BpzaD8Mu3hBaTsT8M7iLRd
SuT7jUMSb7nNFEtU+pzMy7OZM6256/k7QKXN8/PxgGFLOIFy4k42flwZi571yDO3qYfkgJDaIR1m
cC3/hlaju8R3Yd9i24gyrLtmwTIgAuw1d7QghV3MPxVrMOlshQau8Fg4jlEmbJYSmIkOjZA3NuIK
LVF1wpmsJWhebnZYLAY/x637TNyNf5AAG0twXhEuT6MOj+Bd7x3Mo2Yf88WsrsSHOQcd7p0i0x0w
sUFPSa+j9FVuqnZnXRtaSOrK3gWXzTdqog4VEjB4sp7cFgLwWLQBabLk+hfANBoyIl6yfxeXp63v
Gg7vXZSd0+2qEaiGyQElkV5A3wAKSnE6pZVCusVbVtd1JXAQBTLmkXWDNCdL3eBp0aHrFaK2T04B
ljFWBy4lEX22vdo9SOgv4U6+GM98LMZD8PMLwruxIg/OGGoCw2iDauvliEBxYfs5IGDf/fMHr6zC
JskwTBdHc/iioDn4lxZ+RVWRynrLpt/xuzqs64h9LFOy7l4h3TWT1fPvYY8yBJc064thN8HZ0gzQ
w82IuA2nBDTrvk6ssMZtOePh9P1Hyul12Xd/cGxTmbjCVcWBKbgYIXIZB3zwYOaxmm66oCEOhN8s
vESt34+u7eUlWMr3S1B1dOlJEJ1hsB/ONSsUWJNFmF3cTU5dCcgpKxYsknNboTnWQF+pZwUUNv2Z
Vdv5MqDWQF/c1i8ddV6jLsydhD3bVfrd9r7v5Vr9cPwVjqPUfisre7NmcEIvLwCutRNLVdk5JlHr
050T1iXI/g0qiOCtIv/8REKkvArbsB5d6G335ukydbckBl/qTn6GU4i2ejorp4S6HMF6I+V3MV8J
PyYSat2OUHoYSWC6db9Eq71VUuq8m9PA7WIoe+vNXp2uTSY5PZLSJocM2z3yoqwhb9wk4RiSaQU7
+pkKvu6rE7X5Jrvy3QYWVdRSOn5tyj7t5uD8H06dmGzl9nuELXRbrjZJ3LaM4Ma5TRtSmnaaurSt
APRTlsEohMRdiCfH3iVahCO9se2TvvFs36SbnHPmcoep+D0ZXwgu/6/8bdWfthkb+Cvna1oj9cQf
IiDvL1kZX2nVeK7/J5pwdK0GgZSMsENwKv5L/1H1O7U3wp9AVj0myO5fMe2aebP+OFo1weltCTBt
A288uZm4owNZ9ekLe4ZiSvytApYrGVOexqM1UIgSARcfzdTBF75Mxs4AlduIOEvQLbbqskyBAT95
u7NSXTfr1HRMNMXG2OFNRB83L6p5dhWECHzltuLimui4ZMWFpLX1+u19fkzYFinlgiJmWWnAFOQZ
JCSVOmR8KXZhOrWsIRc92hWLFJV14esi7LvFE25qhFAu0DbWGVbUQQpWgBG+K8pBhwIYPp8DM4le
cY0hN81KJU5e0sZu2RM2/e0LzoWbqPCh5t/dy19dciQ/HZj/NSX+qUml5jS5WYcsqDpGLA9gvkVG
0UDlTbTn2O75eOMy551zBofGCx+woawio+uKCdfy7FXBUPJo31LBENW+loTEMQ+A2GPnK47W2C6k
xerZWaSvRVzpHy2SQHrMgO10a7aPqOg0ejB5n+jdZTjgiRJ/RXQuWEycd6i0rJGXw+tsUQ5536U6
646OYIgBInI+hVBNXbeiSvefpNMId6ZTG/TKsklIztKFt019WlYNMG4/qL8n1iKmHme3Xz9fFOrb
jquPAyW/WhX8yQb3mB7PDHV5W7p52uTCijyAuC5JcvAdclV2+/MOICk0hlky/zdTe1bM3o+R3RTH
jemFtMn36A+qmssU57azXtSRACe9ZPrDLde/FZtHXKe+uqSCZYwy0NkzKuCg2YiPmY/bnEpAELxH
P/oivBPNKgUbZ/3D9q8Oz4VEeFTO90iLKXTfSvB6o63Qe8X0nVrUM4qBn/HSwlhM/gBXPxjtss9m
g48HrVuyXkFCSNbmZFxogpEVZHhGYT5HwHMqNBFO86jBZ9nZALnsy+OU1awuAqGAEBdKbuAmsNdO
UB+ikoLkKTCoKl2ZHCPhBwfGw/Sp4+S/CiBvgFUF4f2Xr1i7dmH3ccxq16kAxLicmAmVRo9dhsty
eK4YDx2gzcdpVZLvg/y/t/fVlobraEKjM5CLHnP0Det8ll+yLAS/qXQvRLmWLwX7QDHPsLBJMzfA
6qGUszyEVTCzVuaQv3gSQPohI03/LUtJ94gcCo9i1qRjE1TJbaANDGYTqdfosio3iyCFNvv6MlfN
ksyBb67p/M99WiYRyMkOm61DlcQCBfxi5207SPPErf7/LJyeupN6uJ26ASoC2EqxcsxfL3opfFcs
d+N/iufv6z97KUBNQ4Wsu5YBnjhYQHaLLqZhBzjwjh+FS2mmQpTEeIz7Jy3qb8WAMFKVzlqD1c55
gmBJX2yNQDcA0kS8Sft+OBqn8y3vSGZ+JoRmlC1jGJtBl+XhU+cP7Ero2cwcVBXdVhLQ8SaIemKc
8qYOOrSW14IvvMnDyYKKHNaIbckZIlTPMxXbSRrbJo9aAwb9ouVFW0Ebxcx++Fklr3qHROoLYRf5
4WkJOflSHWp9R0OdnJv1opzN9ZHmPjmQGZIuPYiHHj7c3HnePi/agflS6xc1aSUb+vThq/wM+g85
M/BncTlcHpXBGou2Lc+QuKV368NRprTR1Q1JG2BV8KpGtKJiwAwB9Nk+wOuwd5WDzE8DNCuVPIDr
3SHoJBsv97FN2A/uVyWpc54ReZ6REUbpQrrjsEcQbBRdpjenTj2FuzOXfdBdKzUSMOCgtTmFUYIe
y3vVRlfupJimscxjldK8BaFy+dMzqXpsw1Owu0yjCb0HOWnTVrbWW6QHiMvvUXuTcPQmL3ZWue4y
itGnV1OAtXtwwuoZPgLWod8qyaOncRmi4JQow3FTxOyUsX8SfbfM/EqvcHFNpOYW6VdIdZKZlihy
JPOdiIWgSexb5reaQfovYsbwUVZo9YU4/uqjfftpN9wqJoftQrAyid1stlGnProWupIzKyVTkcya
Utw2RENsiUNhQ8B2GGnztAkfODZZH0mhiQskOK1meMlOdjvH276hgFwjlFBqeuyASVog1DnuHvAt
y/GvJyMI63Mr2EcEgZcLDaS2uiiMSbZFd5+ychVtsCvcm7+XzRRA/AhpG+YJ/EPryC8USXVG4XrD
8G0r/mITX7n0EG/W7RPDjWo+K1gVqeUR7RoStRKzfzB8+MuZvlBGjNpFJBtNjq6UBAs/EHRmCSnH
7e0v9CDMiMfR557S7OCPb/aM5jFIY8FDb4rfvFoJufhuVFSrnBX0H/ztJvF2rthDCrgk1iQgtJU7
59vVlkcCDWgDq10WsAZjYMmisRjaH/5vdC2Kdua9GijORp7g7o+1/FDdysfx07gYufUX6Wh/HwlT
3WAYpam63MTszhUEk/13sWUeABw5QVSCdyp/NSGsDZHwH/u0jd0/rv/ItMcJSZtbxA3/vK8rNwba
WdMNesTEM5D/TVoZ4vajbQ8Qpg3X7Ukm44UBetG1zckzQF7SN+iauZB94T/TeKb+Fr+K0tddJt/H
2QEwowtlaY/DJtQvKHqV7WnEHn7025Ek/MknsV1Wqf6HRJF0MppVSbNYBRWT6LOc5Chd1EErv8Yo
GA8YI9swljtACVvT+H4ZpDmt7J25fnjhVGzAg9MldIwRTfcOjd72xFB1qQi8MXw1wu6bsLvhmScH
R3fHOZOz7o+fwDTeMzZ05mcAiduK8U7qQFsFfgIISFDTLtWNSvdR35jQSmCOzorAv0IZoj7mH6KT
NIVr/BYadrbVziAcvMC5WIEu8R/v6wUbB4P7d7oGo6cQemr/iO9a17AWtbwE1fP1UC+i+J6EdM9w
p9C1bMfhDK0i/YOHAbtlxRDTF++8Uz39OecxVOo5gvfJJ7fixQgUokkzkoFPF0oGG9KuuYX240qV
QCQW9y9C7KmN+yHfSnQZXpEup3ARctPtynMKKJ24ILqCFg1ZV8ybuisOC+KuQEFDPbswOwSOiqnz
dnjrLHquiFF9MySQK+kv9aO/SkHgmF/y0sD+76ivAWSq4P1Be2/mRHAQ91J/GF79t9rWKsEkY8Ut
PDeeqMf8sZGUnpVgkCX6XtaeF5Igom/3qnoJ/bm2h2MSzcQgGaMir97WtDPpjtXuD0Ozb2leXUgd
d/JWbpE9JIAHnIT0P9bb03D9J67F8Rsc1PuliaNbLkw7rDybO8pUtkAGAXCQAWjDZ68H1xKlVjq1
+G9fI5jKJBQTNr3V9d2Lxzq3+Y/R5trshTLyIueqQxky/yTkCkiu2e7skzjuvG2qfrDkNofwmlco
C8y/6h3WxK974UX2PGp6BfB5VdYG8i02ia0HbtlBsWCcTwT97L1jbooF+8Txc/uU9Dms/9spRMHV
3t4ko9lkudION6GmVleufxjaA8y/Wwo5le7kkqKmVRXxoKBijSF6Fiyp4mDFTceeHs+Kj+GmJipe
+IFY+sXzGlCa5y5pRhwd8cz0flfJ9K6X92rxcvh9qnaoPZoEgTbJxFSwSjQxtjXjLraPbb+NzCTT
xIwvtHA8gnRM6of3A1JR4i8G0TJ4wuYtU/sqXThSfSrsGbGyL35FGr93PP6GsLXtlK579hfJkq8V
WatsbBcvodgLkw2p236euV38Fv+kwcYrZzQZU6chPK/58xg6c15GMbWqUShcEcGKgVI2rlRmIRax
HW79ccPJBDhs2p7LB6sBUgjY6JWsDhraR7xyATPpdKcYTBmcHyxMlpRwSOme5VYqv4erTjY6q3Kp
2mGAzza9LzTB92OqIq5T5AzHgNzJM/PL3/lBFhYjUZWuzxDou1BfkKVWooxC1YV/ChuyqkBWa844
e9Z7Htlfmmgk+fOdpvQaS1JHVFWOc8UOwGcJ5Jaj4Xn/FwhKBPRZkeNqaCofRXZBE2MUg5YJZOay
wfpnEgVXho2mB3qXOcsrLmAeNckuUFiyRjLmwWR51vpVJM5c8MKJ5Ww9kHZkqispSlzJGZjGI3PT
uDrm5KCNdf2MnUhy7V64xrobS7Dwf67QYj5ZCrm3EeojNPgq2YRuJrHeUppjk7Q1dfGfQ1g9LJ8d
0nnPqIF2mw78/RwyRL6jN8lnqrWFX1qhF8Gh8DSNmbURhAHIAoJor37nbOxE+75unTG2vtV+TmVh
5eUH20rnznPnTJWQuhq7AscP93PR/rEDPDvlP4biVKX57rL1wWvc4nVUOmzWIW4FteVKKDBd0qQ/
JNLc28yWP58mx1BxOIEbNFKSqA9KAG7ptG89SMZEhN9K2toScV6vsQJwD8eBqEZC+HhaQfW8t67/
plyGzFoIk8eHO9RHDRhOa/rORzPxdbhehhMMU6ak8yACcUvim0IUbyoZJsN5ulJDnO6RFE1uDAiV
ogiJ4S3ChNDe9kzZrScltMCRIPheO+sanwzJanHE2Eu4bE1K3t59dqzGi61OkXudqiSq2Jii8mdo
0Oiss+PC3/LTV9jREmnH/P4xgYjLc2nomMi6o1wc3M90MylaXoa4Xio7tQI/rkWKHE1Y6IoRhQ2/
rdorrKj0mSncD98zSiRrgMg8dwJUbe9P5HJaAPZqW37C8McfjCgqfT/YlbQuTSCxKcnMdw2CSfm6
2xS19Lo7hMcAJ+CbrqiTBUhtHIXBn0jPaAlg7r/w6r49w9kFZ/75sXA0CDTjLCPkPBfav8WsIEOd
IEVc2P8dQoGY6LASZxvW3+07IjwPpOQHjzDxrLyUxLKAnXvcyY6aRPpTkgwZ1N2G+GGzIrWMB+vT
Dwvm3rNzujXIT3GYjsyJBVx8VxuuNGzUOw5OdvIQtDE/1Cflaf/3eAP43DgSTi59QL3HZp+5hbY4
U8s5/aWKXfl5jw/C0vDwK2L6FHz7U5F+/YEy58HCIMmFvLc1dDhCQxKMOVv/PisRRQeYzcBQgtTM
l4Rg1kwGuhSi7vaQrQ3ebyLpY8evZjKPkd7qMABxflyKg9H1/n6kulsfO1xWp2YssqYj2pAI9CVK
I65U3qgH3tMSVkuF5v9wcC7YYyXNvikm60MQDE5R1fPWO6LbTdQmoXB9KkeNkmv9mSB6aNExUIus
E6QHOcS2iqu/gEP7QqUSjy9j0V/HydKKSHH1/nwF5I755yB4emZ7otF8omIXkFmIGS3IXK9jv34U
cdP+7knLjNcCUMtL6i0KKXD7n6N1XBrVjRmMv56KOFRAFDxawwZeoLU7tudXyLFzjHLiXY+blMCJ
17aKeUl/9J/aKNcczsR3opOuOZSi5PmXVet5goYRIeV4JjV0L184r4sUczG+WkTkFW53HYG6cD2L
okYQZtnJKtkoKdUDFKLH/4BkztAm8juYfNUIkyZC30UzRNgPTSpkr5L/HeeykmjjoJ1C8ODRuCmH
yJGq9DDk8LYd3R3JAncjkOT7iHTCYt5i4poGxHEtB+MwtwaALKpUsxoT2wC7RI1JB5kTtl5J+fmA
HrxBsn1n2bUlvj85c4kNktD1YNA32GCBBoBWDlxZLmCLtD9mwI8unILUXrd/8zaMScRsS9ddE+74
6XtKlRMjU3cPt0ytHXs6xrHw1fkHsaYaut+rEmdSi7/wrE+ECqZZr2cNWm3UC7n2XtuVi3vsWun8
oc64SpUyigjoX0FLOXUhdRXsrfKJOxpVfdKUGULhaJYFUdO9Awbd0mmvPusLLs8qmG9TxorJ8mlK
ceoj5KAv5/4J5EU2qEuuXGzGD/mN/8g1dsXK82FZ8PVcK6w+k3wrH99cEq/fqoVhe4cD10xjY+1G
fIsFnIQcDZ/7Caqg1FbDkV4FxafBz78djEAHPcqLOYIrevsJ4pr7FioA/c2652CYOXL03xuvIif5
LVrUm7lWyNrsQqmka13lOTnkmzO9Eh2uXxvnsL3gyJ6qDarxgE47RPs0em3d1wfwhm6a7w+nhR0c
NB2NFw8jQMbvfLYys4r1RXreqK5wy91FEqGv8ZgpE0lCRY1Ofk5xUwaWQArRScXQB2P9xxeFvNH6
377BLv9YOSWZtgmxz7rC9IvYCOGa9plnOCSnFrMtsKBQHZKNw/A1KhTzETuM9F6JLU/isPDFLXUJ
KIlmXRkVhwQStnGkA0dXGzXAkFFL99ok+Cyrf6gT6khmtSOlX9rNzDqfBMp10g2403ngWppYdDqU
02a4k5R4NfxSR6hKG+wldWChrBB7byQryMsLAA4CXRKCkjHmfWBjcfCf0XFp8QoQyv9C87REaCrT
w0DxMpdTUQDdY9P7JOCQrMV/xQiEQzg55i/FjaeTFC0S5QjLhYCe0AwK9MTd/DWszIiochMVp1lX
J0v6WveBs+/4uoeGVSZJxY+pKQkozTsugYid+dLs4/YNFeVcq4DoYAsI0+X3/1kBUlW5I6SjUXqv
ie1pW6dJyFWm5SdZmp7HLt5XHboO7EIOd9d1kUDsqdrWv8wyvEU8+EzxvjBxhrWqR55Tgu81dvBy
y/Wn0D/Av0DjbIBzax/zvXu5K7oj4u0/JM97U6AtYhbCdESepMoI1ZRtCNt02cBTtsKioiG8UORc
GHAqf7SPYYEvjQZOVSdWZpuuA6HKnkqsdG+TGtA+yd6hg6VXxWRAoqLOObWylI6Ip8tIjrYu6G7n
FubrALpV/gm1Y5bVocL9Rt4RbUbQx/gMfUaE+jMN2TjQgtmqgZJZd7zFQh+pZjXGC4NrzY5ExvH3
vnQNAYSHMd+51wEcJT94wf6n0qtm8qwAmsS/A5mmdE3nXrXAcPQ137oRaykKIWDLuZeNroTS0j0l
JgRDEHS96mfNqQSv6gZUU8aZVx4v5iHOqmpsnHGYC/Wqox8MOgXMD2x5bhtXqdlmfTft8b+hkqfg
/dmQWCxjfVJojfzxQlmbKc0wtHgRtZH4/K+55c21v3SwH5AuIztnWwEfASJZSFptL62FtLwML8cU
hdtD4whwJ0iqAONcS7bZLPsQFtfnMZUkwNo52JihRheYI1NUyhJ4fp0yBz1eo54hDPzr+LbBe3lf
3bUNM7svPDswXY76NMuwH7srzwV6iUTX9ZirrQJpcuFlHCSNZP+yTToEo69ZHoGCOBYZTQD/mxb0
4N1xqONHFRKzEPkTqh1ol6miMEbhlUk/vjltb96BiX0NiQzMhLdagOPgZPa/09e92ID03pe305D8
slcdaodKU8W0Yotx9Ci56T7FPd0QIhTrYR+f1zSDLxR+jg8k70XLbGw6qosyt446FqKzmcEthMBR
DuSZsC01qlyoLMtGDBg6a3mo6dZ5PZYSwHFsN4wMd11ed99ETQiGiMCDH1KEUc6RxPAYJbtKZaVn
nb9qZAfSg0O9THOnSznLH6b5T/uIgFG6dEHYn2AQo/YDsTFcSxh0CLXCQfxatM3NeS/COqh3E6ek
UeLrCG86Bfscj2Z8B4huExaAaZEnf9W8q9e5qkXz+CJF5k4I7IYbGIezrJC+Sfds+RTMf1fmPGrb
tLCLS1ZPRStBR3IV6CqkmLxb8J6HjwvDGbd46WDHKFCMP6EWTszxxAUEsDdZu6YE8T1RqsexNP8O
ykiLGSNpZW/WVZU76SSvn1r3BpAiatqRlzPopLMugTNV6+2LAAUdxa4y9MyF+rN129rIS0PayBG2
Gs/xZM2p/BKpjmXT8jDMRJu8PpUTHBHKPM7UUxVLQVCWfWOORRwELjB9QMegu80BQQjXPGnnywjw
0jvqFf+wixrYXvh7zZnRxVUc2H9eRSxrniN3ymXVv8SSaqAe4xyiJxg9/aSAx/qZGbdeq4Wpb1HE
TxdMlF94/n/HnrI1PwvP+eP32fUcWtnP6eWuj5VXaFJ+W4b33XGP6NM8zD4GFfSxrZVHLZcezFn0
NOQfGDH4FSX+D5XfJlqd8ROk4dwx8WWjiNG5G2ikkXMe4KtRxZjwYxn6r93Hcg1yOCg/Ov35AzaD
IR7LuAYyfO6YWqDBhQ+aDYAjr5vtKutJlnFEoshX3Um2MwDsfMpNcZurmyTddrqaW1D9/7HkiQ6B
30TTmO77cQlpA1+Sak0LoUJo+H3qnAsSwwBZehxvU4qpxpWyfMQMVGURbA+aaLwpG0irXbg89D/l
LwOQ4UdAjNW79I7llSEvJY96xt6Jel7eK2BDPFZIQFwTzj14hICCMSb/qlPr7dtYtX64Wi9QWs9L
ug+bK6i8mfH0HipF//BfFg9icFqpTifk1BJtSiqVAZhBIhktD1upz528JmnW++CTC/iEz/ja0pNO
DDyaKgnutQ7dTm2W7Dzp7JR2ttSFtBGGjxYGjQG3IV9fCtNxTmUFdkYEuzvDsNJghJPuULuvK6p1
EpaifMNRUswySNteSqemyhYV0oFgr8uIvgsH+wplf3rU6DC/pOnE2t8rejEzwdgIn5mJM1ZAbRpV
cV0dVPyKI1jBlcjU0KGSpyDK6RGoBLW6a7GjX3Sx4hNKxjaiheAn2Q9ERKleqs/FMlrftSJDpcuW
d9UxVOsFto4R52xu7/2DavTvmgqL7G+5FE4pfYvI07moyez9l61n6gphaNA2O0KMdcrOfCOBfvi8
1Tfu7N79ErhkpKN5vNmHW/lKtYqwpDdXezVCWuwxveX8kakUWXzu+rZJuBubrr1dXE1VbhVufbX2
nexvcsUdzyqmukGB0hoe7+28F2i6kiBHcMSKvssPgbjTfDMUbLMUYWT/HvZo3Z2iqcnJLDWlHFzw
u0Z5FN0m7WFESu3/DwW1R5iWcEwHpu7hdMGPsRpRQhVTKB7AW9xFJFMEW8q56kKheHdfQ4EazrGM
twSxgqtIrhsQ919eORpWhvHq1+ehLq2YxtA5PQa9fV1RF8xLrFZ7q6U+zzBCvY8rWu8rgb43xrUS
cx9PU8wPoQcDANvpZklxJajR/W0+dCslJPF5vav1L6Dy1SFRGCXkff71cD1xDcyfMovJinSuyT6V
XgSJi2JOHSUT3v05ykKYN/tAVgtzeosSMd/ia0KLdbWujvDc6qXzDLbubKKcQuLFtOiN13ugZU9v
oH7qPypfduZGgZFlpS8jeukuN9aaow/rA75Ld7heh8uU0tsN43a1E+KYUmVARdrybry07Yikp/dn
soEzxn5NnGZ73qlerpOjGW7987mWiExjiSd7LPP8DkhHOP+euejbkYkniYm14d9H0no61+SA+fyX
kX0W4J+VZ0yBVCSdyh/sjUvIKRczAYjdz87UPE3WBwHrSR2MHl/k5ITlVIw3d7RSiqwU7TIUNKac
WYRYb4K9a+qoPdzh4IUR2+rTVJ4P8bG76qpUoRy5uwTmTSDTyJ9rMxAqL3IpT1iMf/dE1xKy/unm
ys+qxKmNN8GEw1u12S6MOoM+J1DLaI2tMeqVRSjtuFHRhP3LS6UU7pKRUZwos6tWBUjBgUJcBHQS
IOAyjR6/LjGPat2rXdGYQfbVtdyvy3SPeL/ai51DM4tKH2OS8q+5FZfSCshmwvvpGb/IbL63ywID
dKIG7e7NJx8hDKpwmUJvoeUKBUMNze+pzCe5CCjFwjcKAA1PtOtH967yNp9PZFIpROil1fLWtHP9
THJHgY3LUqEDatK5BkahDSct2kt7dralt+Ot//JxXnXGeNSqe4UC5/oyrWSkEw+FfiNeJ1A0E/zQ
FeovM5MTxpeJ7e0YjZ2jejtqXQeFwqGbP5sAz7lWmZtUPooOf8PgKr/7Da557pfoyxb25HiyEef6
Cz4dRfdMDhuD0jy++w8mLl960/6mmj3mfXCR/ksvpaBKfgFuyLpcw015nPMOeLXxDk7dxnqZLfWl
axcRjF4Rd5uW9wE3yk+cqdowZQ4BXdxQNs7/tG3deQZERnnjyjE7xMaSWXClWaY+Rwv5aI88HGFE
6W2c1FFSAULGtwyb39czextHXY1bWwwqfVaTR1MXLcvbAMhHE/7y5g06RVBxCcsPDIHZZt8zMrZ8
zgsoK+jzUtMWswbZAexFOqVBi6VtZ8rKQrI97fKNK/4UqBmvc/e9G8x/BKcVsexD1U+GneGtTXmH
lA2QLbyD966cK5lwCZwI76CV0Tb8+d5HAKc1WhvyLwJ5rr0isdxgl/IRztk0BRX2L2TD/+QVMy3R
pla6Y2o67cCb+p52LHfwm6JU+EKZwtS1GvfQXSin0QB/pp7fqvCUFgGO6eMvcYDt9VGBt6IkzuAI
58lfKjrmIVqEeYDZeV8HqptkuKvltwHp5esuiT7hv+jPIF4yOvISINwGyaMT7NojxuluPKnweKWu
BGhay/2ligklQ9nM+C+fM3+9FsKBZTd+tN8Wwz+csWSGHn6LiopUctC7VaOTIzJGMRTC07NQq/Lw
2UDdi7gUrFlLHpJLGwrMhQlYx3g7FHgXPbGhdl4mvmjUI6XVXxgJQWryXkd+fN2gFSCn7jg9uThS
UkWMQYrCnZXbPO1cNbVWGNz8ridNLOtpzOn8kEG9S56UeVShbwuDd9B5Bssl9rHskMqj0BmrcTfU
vGeG8ukEiNYhGQnDLdVoz1FldQPXlaFxXeeopyd/UucJO8bBd1eTRXov22vNstcHFM9jrAvZ9z5H
RdWJ2tCV5RWWA+bRTDHws0mLDA0X0wG6ZhmV4JUhgmA39o4v4ANlABsvA7/jLl4HPTMPtZ9QOtzx
Gf75+2a1Peusa/7k8W/AUi618A/FzT3Qse0I92+zc7IHLsIysuu2fx1peSh2mvbXC7UfOUmi7st7
HxtTAV7j9Xa0TGF6wbiv9f9S7cs5Wxe2PSuMsSJvKBv1b6oYA8Vrgh1MUIySXf/BvzhADeffON+v
Q3sFTHdE+gvMkWqmhBuOTGXOfTYVzO/9pCoxCFgb8zWsMMSJ7XzYcNozHBiJ32DhkkgSdqyhjG5E
V8YR5mVHc6o9w5uwGEt3qvgO4a12zkGJQXpXizuK6XQd7naZV6Au1ikN+xHFK8a4viCqmtPnaSw4
rZihNeVH+rdwRH0GL8TZ3en2IkHdS/CmNB+Ys2kzZMmY6Yx+Gc7i7OYzpdPGhnLBbmTPENAaDPcd
VaPQj3OzjzbRE1JTHjTK48UNCDaSv/nH6ei9uuA3FgVg8d+FmK5p7vcg1Cdo8VWu4sKNnagkk+2V
JQsxfGXAmFQ+6LIWxu/SzbGWE4zjrP9zYr6HsSfkMnyUAubWDR2Sc98V4xZbFDRo1eK8chCcDd3z
lOhC0c9SJAD/6InIuVPbqH3APW7St8iFYCH9LYX5HXvMkIo3UE52w88jvJbllLATYj/irgE6bj7t
nBUA1s3kBOof7XBELPYJiEpHYQvCoIIm3y8K4c2CH5PTyuMKBJMEf5FeXmdrJCAo/Gv6XTnh7Yt2
5H+vrVUsbE6GOf+3HG/sPD+rMDWW+5j94AAp4TYQ+5A2c1q6BT4McS2BUpv6FTLJPJoLL52oHUPV
PMc9lxTykuZVxQv21K+dXEMRj5bdrdTNYnHo09WQLNAg8QBK+y6R4aag2KArckaQCOD6C7Bw8/WL
ykbJ2g5fHNENODpKo7r2LIh7RsQ4fLpaYTWtk7g2JGCV43Vpxjz7hCcKoLydZmSePIkdPcrl5LQP
I/uqvmDZhvk2HvoeotCCHWhJTOcrX5hXCsjVfM7GborPN/gswY1a21Otx5yJIYqfza0K4fNjap8h
Ug1oNWiRqaLOohW+lAghxn73i3aEqWsDLHXdKbBv3DNu8cesrNAvJZXaDlNrC0WhW1jJaRwts4vU
sGUXQEAVSvvWaojqu2TvIqKkeW0/t575nMkF689OURdrxD7vz7XSBIZhr17DfPfpSH5cYzYhqiPD
prHBPf2/kJPdNOPQg8W17ttB/9rpYMl6DfVOyCjNGe2PzC+JK8ICnVC7sO1Gl1br0GWCf5CR7WYp
sDt31ZuPozR6rv4zEh0O7kdK+TW6GLLw4GXTHrCp5xVR+7q6tADyIuVqFx/O/lRhCF+C1Jw4cFjS
hWS53wRjZXE+IirMLCCum2lNwzxJ1JKEnpb0ozn8L0bKcRVinxnnPi8pUtfY5Vjdup+dMWj9xQWX
k8QHaOq4VXmENkAHv4IWr2HGoqWqhjbUIg47KXnANiESk2BbtNHVMrPets9iVOiwKQ41kveC7lSZ
HlEQd+/LTHvi8qbBnys//b2A78lBqGGfq/j4e5AH9xTuBgfYj1Vw7HOaUZuRUixMtcopg3Y70hME
SZMvxRhFMXNVizg3zyw8RnFE87tqfQke9UkD/BgtJf4Q94+wbPoYkf8j0ZLclc6UcW/k03MYdluc
G9rGylYi4GJGlP7dZ1BdUbwaTqZXnezIRYeVxLvxSUULBj9AKGDfctkVsPllmQtWvDzhqqpXRnWN
e/TYyMGISR4gQ5L9glDwMiROBicLAl2I4qTSBw470Bys9BwDPRPcp5/a/fPzDS8inBAQeDQjxFOi
g6sad7vI3pSWIzkh9ex7WmMXkEKRWbXKygRCGICI1FLiFEnHQEGm75v0am1+WAApoJUaFl184CEz
q7w2WIAtwAsMVkjL9ESqGAsW23RvD0IojS5+Of0tAys6qhv7wIXSXzClhfGEmYdgnroeFTRXrd8L
owWNoBv287U41Xkdt+nVWKNoXJF2nhVuYCiQdQnB4b7toqJ57ryzSD6ksUxwyDHxxk2xrSXsfJPx
gvNWjwkEHYwPSyFZL3nfknYX/EMCgH2qm/18bnrIn7l0fKJzIbqanDaw2SlzPLSBevMas0KIhqzi
nmI00E9Ve7zUNCIUhA1OJWl4SxIuqL/RcNOk/IkakTegzr1ftMGK4NgR0mkATEWa1CN/vEp0UjTM
F90x535aLKmoFTpEexGMEOeXJNKdXdQXia7PWCrHJnrr6O3cO/ex6kxOa7sufPJkpN5J66Wq3pYb
1ckEfyOXJ1yTxheAZiSVYdR1Ma3thYtL+/N6ZmmU8uiMo6ZDrUMo88CQTF6Dg2m2InLa39TK4WiO
Z6KlbZIv/0Z6jo9em4OrzJ1kOcsFgBVc0CukWHabdg5S0mgzZdzGogYVYqwsGKT2hDb/4Y8nNW/R
KiKjP0BftHeXbpdaoOig+2MomUBXIVrWd+5v4Fe48ubCPp0+IWx0mnaznIpVMW2U+tesxGddgsLI
PUctAlb1ZydpzvNRG8bjHJr/hangoL8MbkZCW9Agv+bJezWYDFF7j++6MhkMZpkXceQylN3WI+qj
wiU/S474nObJ7mFFfgSIUKCYON40eL4QZC/UfiidkOcUU3lSuHFLzpdUqO0+jVCkNN2ltIvbaDOQ
feN3TEj8dBi2GLR5ALkWLXa/t7cu7XB98NG9v8QgPIyJayYvDiSbiggDiUws2edQe5HXxU4Iwm3b
BQQog6vhlhLLlLDDxoikwKnM7r99Vj9QJRNhCg5PTnDE8g/pa/76x3lX1qGWOtnQj6WKUOH2Jbmn
afoKUrg5jMfT/RixO9VI50+XFK2qwl/gHt1jkVJzjkBuIPiEqvFVnqzuCtsxmIX21QCr/npYSxEF
IRUAxbKZqSpUT79pK/TgRDRxkiCWvMZDlsjASTl8DttSMlbO2rF0Dk3GSSv3b6iZoS2O62EnGpwB
Ix5SNpPYZ0SiXpE6TZujiqTar6Hf6fGZ857BJa62Qa7QhvuYTXJK3o0ESFWrwBeX6DF5KyUm420H
qFSvf1ZJV02Pm2SyDW4COvqFMEk5FjRBFBG9RGmS393hynTuTNAZ8lL9dvzdyA4N51pF1smgDBtz
YaiZTtpB3mWWXuUoWqV8oBFtgJ3SrbUtYl2Qm0Hok2niQBTQaRKgPH1FjaHjzxtNttvV6FuAnbkm
epoCY2X4Ank3Tf9/LoDFJPHteyh9gLShMQrwRdCqmiMtFeG8tTu7lNKMGW8SAKOXOEEKoie/8kMu
5EsKTHlkgu5KcfVWfnd9zH5pt9+Zodc50OeiJnmjsCx0/RY+04WxN+eEgqj95RDaf6c+VHJ46W2h
NYGSUT72/uTTRmsA9WXL4YxzQDqdJ9FPPof9uO5YuJwzbs6VDbJMuHd2xBVlmTsIWEYfu+2bSWaw
gjuS9GHzjA8vaKXys5k4Ss8WB0HCKq+Ukc6ubPZTZIv1zdr5Gj9AdvDlAAmsNcT5wboMKdR+FUHh
80JvpEOBXxhQdPgeG/niGAUbNOzTLWm8ZxKjlDp4TvXcGv5PK+AcdzjaKhODJmTjpcVA6cX31ne0
PIy2JYoXC9gdCCqoFtZCE1gQ0W1KdSGa4OMwrERC1voLKAVV2VHk5wZIUQgZtpAfd5BJ8tRKQIw/
3DUkJ9k8rjep+XxolTWMjSINCTe3ZZgqZ8Cf+qSYSuqiOvsS4teXVm7Jh00ubiSY7AOFXlQYvXlv
6fRW3mv5WvyglKqqx0eRpEQvOtMUkrvMgTDr8vkU/JLaG7xNFVC1XbD/qvozHUOd9m3JCcD7rxV8
6xmNW9zI9Y1KG2yEy0WAt2ubL4G4kXYf+e8Ava4iT3cvgT4B7YNt34uqfbZ1uzPcM0Tie/+xmsWZ
LYap8wWIdglLo35+Aidng0mIf7vpBndGIvkri6MEd6gI67vN+34f855kY4tOypHHS6Qs4l84EcXs
gQ7kgXIXWDwoY5usxXOd4VOivK/tRvgOc/9buwDYxuDhbVmwrAaQeIfl1DlDONBkR+En9x9uGX8R
DV0qc3mRThvB6FB9aQn/GmHVe7cNr4TyBEn3ik5xgNqDEVUYvbERNm+8vIcvQ9x6uc7Pg/YRzjVY
o+X+cEWKfzD53E9LYDCKDcB/lPJlcA7NI12lR3EM6iSQoiiqZCHPuUl/kWMZwapiK36oxDMJ+6E3
eHIgjXbEP0w4HmfbXAkUxWS0zXT7qxDQwiOqW1noOrF7QxW7LJ+AUouViy5GhAR8mnoLIC9WxvfG
ScE0BM0aRFkMDztph04Yvkw68ewdBmOIr3GUr2fnmzaUcyliSemc001HoSJagX4QwIqRJ84zG+Ry
fboXc8zXmK+76Ya9QH+ZLWpa2Bpj4bmzt3Zl7ZHwbOByppJ/Irz4TDdoEPcnCkFIfu3aCW70/rFP
sd7J6a3o9yeTcp6eYK2rCBfjURts/CxKwdmq40fiDSJ0oI4JZ4QDH7FM2mdxbNDvCMWBllilgMnu
A1YZ5yNWgrCj6/cSbXl1sY1RSz7zojgwx8PTstmYH9fD/DWOj3dp4d3SkTSHBpsKCYUgicCOQWk6
8UM6caGndQQu36pz4YL5sR0aPQ5G9PCbGaMcjmgiGpKRNqIr1byVP5iDJJc5MQGftzn7We5lfgJZ
0/ezgUWR8Q6RBKBXIPgBVrn0dtyW0/6pxiiOuCXsgZLM0bfWdkmR7ajL1XvUVDvdXCfEWqbdDNt+
Nlz0Hyx0mFTTLQhnHOqwQhBActkqFQ7VMjnR0FziCV+qcTkDwlhEqo4IxsTUj/kUM7e491Iz4+vJ
BgKSE/MhAR1GSTjoe9kXkKNY+Sx15mH/AKDynE5oSIMV49H6/KxsWT2m5dF8mW4125cxuajHt/D8
i+RgaRWk4xieFJyN/VqnZ2+XgQEH9IQCi0jkUM3ASrPPupI9fkuA4m5++02QRMHCldteWBTSctUK
PSAXAdbrFCrhIFf9uvYKJ77N0dEmqPsCVjpyhnB+Wv7p0l9aydMUkVfpV1dzFpq5DMipZPYXUZfR
HPZppBs4dmZ68XubILWLIrY5uFwpo2hPwbCuJXqHKxJfX6m64gNo55oVO0ZXGIIbXzlg1Ey6d8KF
OR1mB2u8GVULVY1RWeClkarHoRKI/K4oxcrDEUfB/LHuA2mH9LxAP/Q0kIbnUmKFgB6wQCqGU7jc
TXwlsPIJ5sGTH6kpfoEdcaga1cLteFBBOzUdu+Pd3sXJtSEhx4xPgWTsvEzuqQUdg4a61gmQqJB1
JrJBFVo3lkaqjH2nJB/XdAF8dGisT6fn0VE7QUwS1bs0EvyR4b0oHOlDYR5/V4XZseNaYKX+HxD4
+6wRkKZdo8p+WTV9EGrrzYXB4nN82iTm0koKXTG83S9MPOiMz2Eiosx6/YJNpH11ngk0haqqZjmR
m5feYFT5j8soqUSz/kZzYGSEVETgM05kGnuYJ61CEa3jSQ7bUuOv+vBWSsHdZ5pBstiufxxNCSFe
+cp/sXcahmdN+rCyohBbClxbPwLa7CGqPEa7NCA7pFIYYouj5STrHI8J2cWZkdY8YuhD0ja5+X9M
LR/TE9RVnANZB8FWVHWlvUQk3D1OmV7wX3Jx3MF+jSSXbUMLAjD49HzGe4v7rwLwa3mOum6bFM6U
c8l5jRRLs0R7IJ8s7/LbR4VSM9lyMf3eGT+Pdfke3oO/cM1dKURrNXs9JIrCkz11IUNMdcNk8USG
XtaiJLlD/ZseCQ2HZ1Uj60r8Py0Eb6/3Ty/iOFtDA2zUoSHmH+lcqmpQpfctEXOhxBr/h9/O5tKI
xFErIghMjsspZnTPARAgvOq1Vxf7jvHv3mYAWj2Cw/0lpgG3gz0mnznau4sjqWUdFUY04LB2nP5J
U7lIOcy40Y8EoOQ7IkM+AOApDayY/YM+lLjvpI3bApoT82Vj1tfU+bt3O1efrOOvTa2HvQxnq/JW
DnryTi5JoLMyOn5NKtzcm4oC4VAefk+L4AOm7G7y28jZVTW2XapgB0asOOcsq2k8kN2AXOFpdNIq
BuKQue1N2LAli70AKn8TnRy2vMh3pjeTlUwJBOLG6cha8bojcpBbaScdroHQ/Gc6rrJWsN01VsWp
y1UZTnLr9HK3XG3LW2UvPtzHynafx7lljgP/V9svO+9/dsV2WJvR2SZisdDJkhHXdIPa53JIZzs6
48h7ax3FbfJqGiXgIJiMPiAcJkvTmBYD6P79hfOZfOZTnzJ3YQIVVNPI0cfe9g9Uf6k5CxyFMI1A
IvkMjBaqq29BxqEvnHOBEhZBxULLrMT4zwyNnA0ZxnoJf6ZisAefRvaXs2hGiuVVwYcVcnbPa0dV
d2/AoLi0yEuxGJEDk2+kXtScVfnojEbahXF+IOj6vhTSqqFCTyOPXbFvkK2TiTKnYJwOh6nTktjU
o+zx3Y8J8n3cU/t/UqVCWxHjRzKyZ1+PpcI+HlmEULMjXjv21xddn7yADS0iypDObYRB8UBq4dle
oCtcOqUVp4HDcnT0uKr/TSu9XMLNTbS5onwKDD0jGfwuRCpdZZybARVgZQCKlQycuSVtSquNi9rH
iQqyCE5q2d8MDH5dFGX8BxCHbQ9IMovk8/v0iQLunZY7Fbalst+ZJo+DOUfgn/CNsrB98ZJKzsEK
lzR4nPapkOipnDMExsXBRkqH7TbFxI5Pvh1EcqPkRQjL4QvNWgORrmxvTNFQRMF1Vmuc9gH/gxS1
HN6rFOLGD1fvIslYrT8jn3TtEMfdHV1d4nZPPTVB4FyIIDoaeo4LP6oFhvWv8MKF3Jf372KG2T0F
Y9rukmXaPQhCsSbT7/03nCLPu4DLVTxGFGviLXbSo/5ve9rF/Ea8+opmc+NfP+FKzTl7znmttol9
N5mINnxF8ZmpoJubPcaf8DX7QP1QlnIa4Z/QgxhG0b0GoWyZdIpz+41UinhUKL191y0cSbofLZyU
dpFBWj3r9JHlhtSOhGA5yD6M0mzOAfvZwCT2f/x/XREf8iX1qaV22D8I5CoZ+J+LvKkY/iCj4K/i
kPxryDijITOjgWiiCzq8P8PWFxkKH0WZjcWI82aqg04qHc1WJTVnc618xGUz9QUMUVrfBhCx84Vz
SREXD9EmOk1+j5IP/+londmgBrLrygAdROvNwamXFMMxJ0UaQgQ7yEXW5DY+HRCKRam5EHvwW0v+
bo9I77lF222qYmTOVH88cUXJKy5cGWj+JYgmlNCpGTc0mPDYQImx8ia+HQIrU1zAKF/xhHWYgB39
s0ui6X1ucODYUojZd3664fHhXNg8kKj4GPoaWi5tu/quk1Q9u1CpiUvrE3Xn4MkTObR9nhoSxXw5
p3o35fwMMh72HO3UQtobgTJHPHnPNF4tQHzlO/SzhdIoQ5bpmcRYSUF+H8EfWdkmA7IhtKDoK23Z
k4fvGkW5QXHT38YzlbqzgEktD+WA70rqa3/0xCqFLseVI+4WJT+gIGVVLeDKolq/wk91GGrNURoR
LR9FIDyETXS49FyR5Q7/DzG3miYTeUGZOzA25H7cPkjGxsBVZU2grorsJxWqfc7yJb05TKbRBtA/
XwLh3IbUCWuj/B2mZYv9Xo8Jx70f2dVp6tp6oaepcLY4GDPwlHFgMac3mYLQi85ntHCfdOD3xFXr
7arAGBUlI+Trb53fZMUZF0bCVAZho+gw6EQ8y9u9j56gicwpdOtAEo4RK/jGa+rh8jJAlMO1NGYP
cIBxeUt1OSndkMM0qU5MfdrOH0aacDPTc944NBw0i/U91hviqLDZcHxwEnRBw+xV2VHNJYARFJXx
oybha0TXKNJLPKjZGTy5reh0MVtEmjOqYq6YcYaM5JoaBGWPObHHpv3aKeYBxz+0cv3S7oDoTYdB
l1RQW+d5vHsdqPfAAOaHVVE6pYDNz0rUFUvnItJLouiBwow61PaqMGrL3K1sATTk4cGb8Qt97cFY
58XN5oCIMDZWWfFZAjUHa82vcKI50MFzyjLbV5o3WkXM3TKsQmstRWnixzfCeRDk1fd5TbJSoNq0
bfMcaRXq9KwKDwqon8L02g0tokGgues13gGk8KVHUNYFEykgY5bt5tfx7NvNDSIPXXKbgB2dA/TX
N5gmt0eh1uuffbr9zKTPy8yf4pe41cZsKui29mP+UUkqTou35fXuUi/LFJmUCRdTUIagTMgiJst2
y+kfiHadVlp+zqmDT1H5bZNSqr25vO4UFQFRjkVBYXCJ7Dt6+Z8Yh2299VHfQ9wWxXT8GhEz9oFk
E8KZ195TUdJXsgOilv/lPo5qmZ6NuPJHryFqbby/SnxA/iJ8WxqRS6yob5tCrLCZoS7prcCr7z0u
o9dt+PijB4wYVBdwQ8/IyUprxL+i/rF6SD3Kxn0FlBGX7xSALMa0MPLLAC2FV6xwWMNUxBNszl1j
pjFP6gRDUIQHTG8X9sihuamqLuS6AJG2O14g3rrLWA1RHUde876Pced0oO+HeicuB0axMe26YJRJ
RcfrsG8/gG+H0lHCmwi5/7o3jM1ORuiWTxd1tHYKhGSehpAofTFLhWCqus+ZKE0RwsISStYJvI/i
HtBEnEBhm0Sc3AssA4mH8pnJEkZ6byyVeeYokcHEdptqoZf4HyUfihLp/qGe0+HSIGCB5PTc8elK
N/d6b7iZf30cZAV9geshkSp/Gso3riqPet8xmFL92+8W7RGZbjKyfAmCL0HmWN/8jsEKLR9cyOB9
D5Zq2rq0EXtZUs1hqmy6QNzWfRiAPuy+ruf6N1N6BvJx4XYNAUgFgKKwDviWaC9zisqsekj2LC8C
iQfdHw6cvBYB6vd8HK4VTsjp2MrUzPq/tfOi/EfcPKSrc2+IvzCBorgYXIybtHJW3ojr1zuXKLi8
inOxsQoy2VhoWBQzb3mzPaqah5GEptLZaz6M0D5qgusU3I5t4OABuq/I8yf9Wr09Fw+Hmid4/siy
qYWnAEtLT+zb77t9/1Yn1pPy9PrASTUnvtZYL4tiF98D1/X1FLUFCEjUdsM2snV600Q4RYBEDR9K
Rv9vOMBZ/NDDRgdl8Eb2rI74pfxSJPZVQayr3buSH5TH8B+LgbVcsf94VPLUCw7pJgeCrthXlQRb
R5gRedQzTu70tcSZURHeOI+mJCu1D6BHKpPCKGm+7xXS9FBQ7FaixZBHNKS7ApWN/ZNaWCVGSU8F
Il9JFpVKdCM/wRRvP3XglnocPInw9tj5LSzdM60Im1vNpz7BdsXZNvW4/vHToQ22PZRhYXncjA3d
djrQwQV5r7Fp9KIdSBwRiFAqeXfhHME7PDqvzoI7jZJzSfGcyUP4Urtpo0RRhBPTMtvTcjrRXg2l
nVtwS+U6qsi9FOWULag3ROsEaB0+9SpWL1+K/f6LUTSvx+iGMPjkiI9UpIbZqJ9avIM9TRdcf6FG
koMUnE/v4va442a1DGSV5Z6Ij40O3q9opZ3KYj7YTmSeMYJMWlwbHaQ41XfbaZdrNkh1tnOSuzwk
99dsKYhNwauiit7XYaOz0q+Ya6T5wfZFOz1AoGSA/N0QQGWCfNRqBWwpMb61qLQuyC6gH9yEFzsg
PuwGhQHFCeggz08ZM2vHW8U9cIv/q8H6cR0CSbkzs8u91eJuLo49adnpgRYv0Yyv7gXVLqDQ1MeJ
VPzFjjinHI8ce25LeFJ/AghUjLUeRpcGeSEgxvIkVW8OH9MEivkUtvgqfiGxQVsLQrIuVCHrHwoY
/+z90hIA2z3I2CR0mrkZ8gVOUi77bC3dFiiSmR0VPrfXCcQVF3IpagD+k20q1u6HdSvLS4Ws3BuF
jIgodswmpuhbhUmc8/4j12kIjnytZO/P89FwuJHZ0bOQ/t/ePBfENzQ6RXDZqFhtIZZaJzw8xUET
+Qyyr7YPVI0H/RQvKW92HiFd6gSOC9BIjq/oHXhfepiJJsAwLRyKUxmuh1oWMvF3INwdkWnZ08JN
cDaJW9EUm3bNm496QtRSYG/T5rchhmj527vSNCQHA++HvvV1paCTJiPjoGHFN2plp9gIYhtrU/cj
vcHDfnHEktfH8u+dtV/a7cOgo6qZw1Ob1Hr3yPvN785SwmvtHUDGZp+l3agBNxoUjTX+k0G6iTzF
ZarwA3XY4mRIkEjPtXhG9Dw4fIJ1ES+1kTktxUuFS6/u+JM5LroNdXNf7CFonTzMPfBxTiFe/ypY
S4JVbtuU3tL7/1iLkAJ+T8dPkLdiPylg/wYzKFG6NMPLvSPJD4Ya3cQp9ixPJtY2kuaTc350fmum
v3is1NBPughmHhtQzMCEj1crFsEhs3nAU9D5MkELC71gmPouJntWslkp1HknRUmSKvgc3QPJLVPl
jBc6MkQ32UvV3rmBwzqdKflfHN8WRviC3xt7Gx9UDIjuz4tlkA4FP8Se1X6t4VZib37SbV51HYj9
wHpYFfGF6onv6PsFl2u38Z21qnIxE60TEJntGaYEOMCvU4292tB/z2fzvuLz8OHPgSvLG6QQR6F8
zK36UxyqQw8rZIbQ+wM00blJ7mY9XuHhLKv7sqNisVLLCrz7VxdeMb1OLToqNVTWCC5UqPlGr9Ma
4u9WbcS7mS14/5VocE7tXKPC8htiluVcrOzseRQ6kuW0OPahGvwIRXJ5wEIT90+am10TnUqGD3Mg
pGajth+5iJyVGl0fRuto69SdYQ80prcL5RVWWDc7+cdxdVdIEQ9xX0x9Pby4nkw1RQQd+PFk4Ao8
zzO8JKwj7QuKZzMpFUT3RtSZ/A78tRjG46gwWwPBiIEB9Gi+ELrv6EHepqWfi5gBNUFMrZyXqh12
0C8j3UQDRzY5Wu/BYpD8ICVODGEGOp5AXCsr5wouEhz/2JMZQUeCzX373+6K8vJQGKcaKxwtPvGd
Nh3b+0niziXxg0rctSOKT2FatMP906xZaVITNyvuI/ccvLopevgevSuiuSGsIvz7AFj7zztMGNM5
vSOpkER3SKzAk0EJB7hP8S7JyKDpigFThE5wHr746hRZ140ZqtigwfVpWpCbKrgWmyimqUf8Tphx
N4keQEl9lm5h/bCWlyPbroMauWiGezxQCYySBx/O9MX7gD5aUuJp9HHZeNr9li/4A0cIYzn+BdS4
gbxByzaV6pCygnyn6dTHUdAHuppCgsb9ifQZWn4L1S0O6dga4qVnzclYpjgpBG3PBASkrPXLM4Cn
KzNixRwnxQyq/EmnbJvq8ddcCYd3hbZ56pwihsi3OIDmMp/wWwYx3ruNKub5ErVpEOwiG/6bFMul
dku8YgTWQC95GXQSkuADCOgT/t+5pWnGsc0kaSfZoNX8TXqve5h7ALQmV4dYiegWyXwK311DtXzp
sEh72J6NnqTwgDt2FfpWNYuzL5FxCONbj8Ds3ingXIOHytzHCHNCT6Tgq6lS5qUkBn+t0rCl2438
aLc23sYQ9X/q2gr0E3Q0ZRdhBtE2pA2sjSvfrOvN11DGmnuXY/TCiCUkSGaytgbSA9pmcaC5Sfbf
m3aPxDXrU6GQl0ZP+g/Q5kRyxCbmKk9pPQN8kf36KMvi3PrT0z/DIqbiyUQa+bjwOd984DrzEMSB
IJDLxXTe0XjgUGRdRwC4cWBhTo7KKUWbwptM5+kT9izy+tWbFN6NiMcWSP5cOD8QHCCB/3U56mQI
s4/4KERFy0PJtK6KoLzPA2kdEkfldtbQiUs8oBoXRNp4n0dfs6XrT2uHsCHey14UTeX6pyGEn3cl
OR0/1KnEiQO9unkprQ0u+NW4nRksrZhl+GL00HdKM2iad6P/8z5imj+k6AVzS7Ur7658wAKacxeg
KHn7TXLFIIA4Os/RX/0GEhn3Pke6i7ho3Qg1Wmb0gYINQnVzBdHIsl9OB+huYKFKwCKQsabsSinz
+2ToaCyJWZdSV12tlnwPNDvfyRKcGhU8Nt10sMXKN0Ldd72IVxKKTuxoeP/bfnP7sboX4haOZJQv
jk3Q6Jnnj1/oN+6Ymd8pTskzBrC73A8g5ll3WMTj1zBWRKYpiYA+joq3W8HYhSQ3bwiZ3IZ6UYfi
THglGUEPfFI4n9NuFu1DaUIh3l3ELbRrw8I4hzc6ZUzmB/l3NEnnlS997wE/6GOaPT5lwmyzZLwP
vcL9CtYhqWRlair14tLC2BEwUMhgQM0/K1bHGc8aj/N/x7vVJ4TPxCUi96VsI5W9To4Uf6fV8O96
NW9JdtluTNpn0dDXP0MLW3vnHk3CPzp+a7CZSLnVrEsXXM1Xp3pAvFOPK1AA2cha9rscpHEuX1FH
6F4ylQAg+Pp6XwLtIOUonY05U8DcWV7XAmY77uJcIBmImC/joMwgYVfyDrAOIaOJ77ixH+4DbH5E
fUDXoYJHamPUkMCDMxbolAm4YsMdngsE6fMSHQ1a3327AxsI/7SMEhgaApoachnJWKLCJbzJRXUl
NAuxQ1A92TUJ66IQIgEOC5nnCazftvqQgrumOAVuZ3r/u0sxYE6u4uWUUSad8+PF3mFbw6n5OxZE
hwdYbcwcU/LMX7eFQSZtkXYEfbGLg+0X/8pEbvYrh9pemzVUAOsgtM3J15Tr/wI2MEMJdhEcIiCw
cj2cSNeoWlOtXmdG4EhzGRJsE3v5nW3ycE6wEgO//AHSB0KpVk0W/lXPiuIqS9xxLW7NW+y1zCw1
GRG9brgOQwa5YlZ1pn5KkUVKJOtlB8xaefqcTFA9wGKa6TV85JBzHimJQ74k3LnN4hR/C1i8OOrw
9WclEhD7rVEKkIFAlKmK38pXzAhCvXiSYI+EkRSm0Z/55r96b0NiMl9U+2b4vCtlBE3oU0lOFn92
eaQF8oCt3KHi+rWowIByHlTTFQtaGgkUq2hj94sBsKnNg2eMR2EEFMdeA83zRjaUl9DLKiORL7os
aAgXJNx7WRkmPB3rTtHGINotn5jBZzPRz2nuk7RV6UMT+qNXjwcB8QDhLpFMOlOt49Ilq2ZTVXn2
Inik7BF0vGjp4iwUuuNmbnpvlqP8YHuwJhmDRSzpYxOfD1u1tbKqseB18hitS+KaZCR7mXRvN6Un
QkQzj1bosGb1gE4AUwWQwRpI8EuWZQHfWYKroEsUpSvcPorEqsxvkHSH6JxS8iVA+vsePXgLsDpM
/yYmU/XbhiF6876w2taAQ+ogzhLQugHO6SpfCezK4UntSuY27LF4QeI/rimXdSRqa8Sm+8wzEfDk
aGi5xJUvAzzBSJf0JoSI3Qf6n85rY2xEbxpsZ4uDZDUv+jeGPJcbLdaFpFVo6nmqoZQ6qbveO1Sy
GGt7yHzua0znxiBIXAEh4ENK8pgRcMaGuh0B/q37xVsoav/89Dbsq0eMsQjI++KKhPXPXy+E26nk
MbE1aQgfDr5yy9DJLAvH82NUaBromgBlDX4c0VHTIerC2opI7TUIxWptgPOv0orM5LYuQLL3gmFJ
8jNfE4dX9b0rskLnRzqB5Dvw0bh3MULpM2kXNCE4L+f4tMD6qGqiS8L8GENP2owQZMCHTHn0zbh3
CH4n8wshoIrLnNfFICinQzm5ap6ziyNrFZXWvYT9X2uIroeM95xKhwmx4PDst4Qs4sPjoyAW7H4A
enifzII/r2sbbEZRRj6jo0j/CbifzcrlCx5kqI40/W/qDhWb99vjt7KrJJyGO39DVOL8Geymx1bi
R+QKITNzTM0w/r1uLvrX6zOwU8Fu0KkwU1UufHYjVtQXmp621iXCfX6wbrrk4ml/dFX2GGKwi4/d
3EB5DF0N1kQAIDUzf6wpf0MMdxKnzHuIhmOJUdq49JRJRxC/dzC/rpqaEXhJMbxKNAxaBP4jx4nl
x7LnIQN1V8AA0SQryH5ymBDoc6gXW1XK647crjRHDd/kTET+n1wILlEJeuZ6QLYz4aYFoJEBWpDk
YXNvg2CXfwwz+SfZOaN/lPX5ksPQjNwMVmrXGNh1vkfv86mi77pG7w6LmvaBZpPQTmYzNqV8x20Q
nl3UYm8vP92W/vv1SDzfzTeJTYfLh5DgXJQEffvbg79oJaAj8nJk1s3CtADVPwUDOKcBva903H1b
/2ldLm0XVDZyQPNiRVODIJioEA2+nODm26+IdikqsJhrX+/iYFplVhMBEs77DWhAnyG3CKIKZpQr
Sp5Yy2jr4bP1XGTVrk4H3fQ45HNkH+SXrCBS+PE4enEP/RSuFO67MC1VntuLmp6RVwAT+IkYE5Ab
fq1vXvj1Tgxry6ZVIV+BIocw+FH+hQC0TUF3ho6BqnAF35clSCYoXUkcusWZ8fUxGORbTxg35Tpv
3drUtTwc0kLSMOjBOMXvTAp0w7I2TbqGQzXV0fpxsZ7l9yosEOZF/9yPlmjNTHHiJRxx907oC44P
48COAh3XdtwD+Pfhntk3kBSfepz8DujRbU5WIVcUdiE+NAUQgyadrdsBVFlI4JDXe5vRJI7EwIlK
E5Npac6xZv+W5Vq75CJLLvA7cYVkO8qFzzZsYpohJu2X+x5Hzq16ET2vP51ocHgJdwgALy7eFeqY
1cWHXAT/nIeMAGK/AKscSLXkQki+4iJJuBdH+0/2hHozy+2ZyaDwYoUk82/qKLYX6H4kTaEmc0ho
QpL9JvF3cMPaEYlEZ1HtszuLSJ6DT5Kqp+ZSS3f6qbDCnNqnyD3tD9qSHD1QSzsIIkDbsYjgE3Mu
EPIQUzbAjyziMLur7Dt7v5xLTW7/JWzeBfYeu4slzKG9+5uSxYvTXVF6osjIBNe8NoBc5i0CbekT
nFcotDgDT7+gcs3pHotFayEF07kk9kNFIuDdHsVIQXuB30mwnVlg0Jh/1AMgQ0A07aWpQ4xQS0UR
5WSFXgwDIGPT+tZ5DBC1Cx9xKf9Ov3Hu1v/LALT36Nr2wVUXpv9ShmVxD+qBK4DRPiWSiggiYp0h
r6onF+r+MtH7SjEFlo1/3jwYuszy1VNbqWmuieQR3FppGfR7MkqX2tKpCbx8Qw34/RBm/uPr3wFP
Q2wTVYfO1gtRAIwIWQ/69CZkQ8P9ze1mxuHOV6YHS9RuDWDTHduWjQTaJ7K9BmB5CeyjMLdUy5lG
4ZM5s7exN4PhBAawm6EkQ+nvddqyVxKQrEUCWs8/l47ygfJ8fyaqzUaPPovK/Gz1o03DFEobEkXc
8LBOV9iusc4014sehQQPQ1arp/5Osfb80ICx9HKdHQXHtDxrrEPhooZKkEBMxJuCqPuPcQyPEMkk
L2E+S7mZcUxRog9b6gcQZSNmnhTeydETfPV22cuw2K9tECQyc10n4AUHsDsivIRWrfZKIBvY+ugW
6sJqfkOKKzVd4KgJfdUBDmUj+usFigByteTVVzqH9GlLSe7nR0Kd4SscuWzAe4CH75v7y5zgSu7n
hxtTFtdJIr8XtqrpzE50SGeoranaUTtzihPjb7TzQeKFLvnqMPzjHryiynhEUNnf13+rKvZoeMff
R7W2c5sGvXUOahpWM8eie5DVb+pYc5xuWMZ2mq8Kdp5rNqEKcQ904lBbvL/STqVvCJVSePywY+Gm
q28ZlJTpTXgwl/eAe0kniFk5gCLgvsgIexrSLo+bVQApPFEL75xd9GlffW0TmXO1/RjASRHlzQy2
iHyRntEZLJZd7AwaWQ0DbqJVtoejXKzfy598sMwHyUiZgTJHWo9RouJMZlsfAFJ6ughJJqyCuuvv
0yf214RwBWVpDL5YUokKZ3Z22nSkfQxPJQ3fnWaMDWBbnf3nIQr29jCBGQ0uRbUMzWNaxurY3JmI
41wli587OV5hkAnzFShVIhLUaX/dW/GFfNcY8FDL8m94y4jnh2qiozPELzAlswUTsSMNImIwUeF4
R9b9ITKZL2zoWudSBR/V9ZyXheWv22kqpVZv3+F7JFqmjKGMiQ824ndLLarXV29CctO1g6EDBkru
keBdCg6ASO35upv9ll8bLsrx0blJUiSRR60BtdAm4iMG0E87EpSEFsNKv14EHT6Hk4FFqQA+Yih6
TbJLs0IDm/0Dsi6jwVDchnSHyxHtPfgbgMHWmfSbAkb4dS6O//xVbNsWzRWxFDOYDv/d5AXA6x9A
nsOTxonPy3mLskByEFXfBpToYpG5hOm4bDUmt8EEcgF+RlzBYlVkh3AWHzB96LhjeyAhouYz3dYM
rpGMNe3HJ5wDLu2vxCe/NTapxIUygUZ1Q9hUanNnzBRvpUtmk9i3YC6jRSlneEJfsY6W2XLgT/vg
pH6zQSpvA9GKoz4K09lxXIq90QrEqIf5LYOYDRLhkm5LD7YS0qbRUKct/G99Aolw6bKCmep921D3
E/Q8DFwPAmv3LCzxwcWUhzjV8NgJ0scsTZCtZE81VGdOEika1CBIAUoRPJt31ssvIU0EN3mWNsqe
bhpPdWd6/jbKVmiK/NpwYb5UKjli5Hdex9co2G8Bf29z7f+49fr2K9gsYW9WdSLdU+S+KVvxx1zZ
falTn4ktjnJXQ3fmcIBjNe3gVvW0mHLxs0SZDwG5/qRynpRadbrXLvlLqJ6U+wCnVtDuY7cTjW/M
8kcI4Nnbe1LJWB178yCF6gMtzw5pn+CGzeorR9KmrpyTEdLDPBqBYKzGS5VWBerA3eqfhmSQ8RWN
jsuFbF4OCyrL85UIO00M5L2D4+Hw8chN/ruz0gwBC7EVK4E6y2GEDXrkd6ua20QQyvt0x/4Jft4W
QOgMBAh1yhFYhjmhVQ78y8UDc0oQ8M/VLtNqXKm/3BLK7A/9FLt66lhi6J2THQtFnqD1qFWHmaLi
3FHAB9LKAWYoh6HLzjz4FGG3DsYCdIp69doxn7qhwifcLg3yts4HEa+1J20o7WZo73OdPyAuj14d
mP5jjjXLEPOLfmgsblslOdIJywPlwANCnQ6uW1fWiRNjJn0mQSULtRb2Ozv7/8U/6v0DrzMwPYA6
Rq5aq2sKif9r3CGzV56L48xvfWqy+Zp7ufqiEiIpK66Bbj+Ccu5RCSg2CiM/rbjzBRBgX9x4/yjH
vbrRMDo3m7BjIJ9FLu4jPVttwlU5Pli+maf9Ju/t4icVJ5x3lqqhbPoEt6bK/QuKccW4v/LZxp37
i5ak/UkODcbqoJQdVr4uGlu5MFPNwoDOB/84tZZ6HTWh43fbBrqrc85oJIMDq9/W8HTyCeregKks
BI8IX9YBmY+PXB/ENfT0IpGBrRm3bh3rz77IDBJ3MxCKiE9lbqVB4E7I2h7Y+rykiCyGpKXUZjgF
mChIY205wMnYuAEGaGtO0evLKPptVai9BVBRVQzr7Y6PhQH+H88khdMv1xffjMEPqyNeHgAuHv5h
wOhq9OcPTh6KljYNKDZKZYTiaQqX5oFIKobZUDyipf+95WDTRp3WNI2EMUocMwstBiZRQSVnwmba
xR/Id8/ZR7oztj1RfMcLVkW/qDeOsS6LefGe+HhH6Ln17lOlZeFsAN/ZhmBOE/Hnu0+WBXqXmBWg
uheDrq9+GElS7foSOWzoBofeAtWrAj6RZt09v6rEYVUp9ouuvQbUlqJUGIE4/BQQr0rF74HUhbyT
jvDPNwOQ8Qj0Wh3OEfZ5CTfZZ3iD5+9mfwV642pb7AxXQLvSCwyEJnBjM+d2E/ggCMybMA4qqcfb
caS2x6gfQbxLCbixYbNkjLg3qyGOnY3k0VhGBnuQF0DXHI2LaC/obBaeDIhgQl1QJmScA+/ruJ4e
aJltILtUhS3RR1PWnrtp0JAmdt7UgX05TfTc/TGplPpprj8WSgE4OZgcSLJSpR+olbrshtCYWHnI
suhF3GkKmfEWx0IzzVrVP7tZhnznD0MuI8rhqMiFrdS6P5mD9W8PSP80LPyuDvo8SMjTpe3bLycM
T5XaVAxcREaIdrQC8U2AHwMKfK8fsl6ZEwjiad35RvRvN5RejWO7PnpMX4aaii93G6wZYUhkyBih
pVTKKq+mWECxN6nQBOuT5nYwdYXpi+zuzsoavi92DUwojBDd5dvGwaUbcGJYiOJD9ldp56RHZ2qo
7fKDKGg2DGAn75N2/wewWUjxkGieNPj/G8NoTkc3pH0bNtNeuc8YiyffNB284pW8pYUWpzqUDiYk
gydrQysVg/+4afWhxVeZMi2bjw7vwzL0DlwG+pPX65QE9sVAIBlNXnbvoiQr+mWWYb79kUBnIv/j
QxfJxBONFrVJkKS1xOZnrqmk4e+pwy7oEeTuz/7YZqFiU4cQ44YLdTKAe5AvJB21UwbQEUwtvxY/
QkSagQsdRZCF7g9dDy/YttRdPR4bIfoSQRdVml02jK3IwXS120JvtaWIhRr570IPTyZRYLn08gvp
syNvdeFw5OLP6UGkXGRBcmzqmuQ4KozlQHEcwjpx5y1iKcKHA3uN/wlcoBSnkoMudIV/Yptf1DpJ
c3Wav9F7a10mANJKHnGGEHwF/S4zmojORYLPqx4qC4LFxkfAuB8EvVQvMD1vRwlqB/l0EVI0mtR1
Itnep2XXS1yGM6DacXFOuOQ+0H449CSfffyY1aRSlsxmGrngDnPEoTUwsX9cVoBzZUwwYx7W3c0Q
vo2uyoJxblGfPau0iSvfgMyjP2nmno3ZcqSqDq98hiJAKAGy8rILM1kBgUhgvvYFl02B7nkhLUc/
lki+6YKthvzC6UFk+pTeG7zOmFMDHuPvdRCTONeQoDz9cfH7UiKP8jDhQvk+RoQlAG+sxizW4aS9
1ODnydpPxxHVOc4+fQAPkoDoTyipvZ1fFNDGdcx3x9gjZzdzrG7/0K3K2HZE6qVEv5ZbUGktxgJE
82fvLXNJdCpiUH1O26w5uYjBs8jD9olTI6QSaEpW94fL0mEHpVu8VWVxmWnuUVYNeW3iD/79PD2q
8VOhwSM1CPbJ35q9cNO3jk61hjiIt4fwrGWdw6Gind3kQ6jcj5x/cSQQw9Mmh3gthQDlLnIA1D5t
4Ijhtg6tBWs3pFBufJ0wnKGcCuWcoZbsY3ifbNtOvF2SjrcdRTonLO08mKSqHLE9djzarSdbsVqA
8N9PgNshEW1tGzJ5M6cDWP/g745zacBLulSOtC27f0fVP82lInSNS5ko47rUirpbshO3Aps5vZlg
8xJ46XwuvAD0Jf5s2qAe6yNbyejbNBy+D0WLTi5BCEYwzcU1jQ6na3BwoNuHoNaVqKnq6Hh+wWxj
klFABNT15bbmVacSL+cY/cdij0wnytaNxLDniM6fZjfqE6bl9O8Rm6z2Wwn8vJgViDSqwV5/bUkC
I45mKz2+DsNOT7n9jZYHXyo4wRfme/EGDM5nT3FxFZm3Pz6PhceUGY6byNkhf8DaILsVB8szgALN
V9oXzVtBBkQfNCkgHvLB8FprdJGHKaoZuhekCMaYr89suweawbIknIB+LYtd/cKItLmchiGBxB+y
RrJY3m68Tpz59UVUjeWHedV6loi7Oodk5oRYks43qsdWJ8FheQA+8U8u1zh51+q5BEWsBLT5ir7u
87o9wn/SxsqxN+9lB70LMJPL2f0+aB1A8m5Os/657aO5j8kF8DgnTctvHSrbwUc0MeWZYgwU3419
3J4/5msYnDa8ydPo+oPCI/xvzSvP3yFGuc1X2Y3IZOENu9MVEKqai3PKSZ6ADX0N3oylReGaRnHa
xzZhGCW2ISIrAHUECYBJC9smQxCx5gLZggvEnuyidSWzOMItxRzyyKVS2tV+mVnyLdhdYBBsJV7n
HL6gLhiUpuv57NCVM30P6TV7sF4gbtHyQ9Klr7LxAsiRQXKUVDn2QGnEhki7yez/LmVegi8Oot+l
SGvoqhD1cM5p6tuXCqMnsEomJllMnWXA8aOHYbSAHeQAW9F9WADOG8HLdim6MvSAQ7yDgqvXe51Q
7Y7GXSDnqOBjGwupYaaB84hrNx/E/Nh7nIjyl11YEWUwxnn76j7AMKj8l8HhOOI8caCFmuGzZmFs
jAE7bAK9VMlIlqwzH687lHUmeHlIOc/5Zyizd6LCJFfaPQse/aL8slxC4WjUChdgg5Cmm8hfQPN8
0KDQkSPZHbuSxq6XtIjG8xZ/ezF6MNqSDM0LUm0991j2h046MmZMAj5mFAoNR/FPxvt7UQC9rQES
cc9VKLXjmxLw/Mtabfe+MfcwOCErcrxoV6Pv/XvpsHS/hdlINBXPsSSoWdbnPrgBBZ6+/IcX2cvU
jjCL1mJC6mHlMJXpAW5+M+0bIkMaMCn5O32ecbWm9l0A/fq1K9HAzKbEGb+z8CzFsXPNaZYX8U/v
oGzAd/fv/yyVEHzseBFJ2fg4VJCGA/l5SbQYgScH1AqIY32enyNYetq/70wchrgAeboXuezQXDat
yZWfmyjgFbCP/iHZ/JJMkE4SFCIW9MselBqZrmwqRwWckhn3iCVcjel8hzOEnkjC6KrD3xveoMwY
J6+Q3VCN3GJLq7YrgtcW8/OYIwXgA8rYxeZu+9kelqVasdoemt7njAwFPKHWLqQEFDrqCc2ioego
ObWCMQfrApfItR+ZYZ2xHLvw7HiZPmgbUSb8LGMnlvrudxzgV8K36eZJlIh/KZu0ZXWpmvMV8RZE
cjWsMmXA0C92WiIhayLDJXV8KohtgToNqZqPzYDpYgWhiZn4gwY73a6fgwK19tNvMH+wK7A151wn
+Wb13PCXygJ0k0p624/wT+NynICXxoGOWfTYUlrA/jYB4MdpDPWdz2KNRjHzePtEh7VeCu17bA7m
rK0dkncdvxx6f2fTFxvCc6jan02UT7doRqpAH40q+IQXnu4ZgtWJqAxVWn6VOrvR6LHLpVXIyUdL
BtfZjP5X1k6v52OtjGqBFbX7byOJR+ShcNuO5Nm3oBZFcso6qFSdjRXX0ysPPHGhHAaBG9N00nOo
O4GoqGLsGM+4EWw0EVEfAzbZJEBBdDg1w7nlV+z9hJgEVZA0C99a7Q78M2O01fqOUTzAiYR0va+H
gbjvdZaQxxXiMASAS3DyePGseb4/vY6nVDJZKnw8mPPeQ05lz4dIFOupDbu5oqAqYc6bhrlnD44a
MfbE/nEaAbP52z6ouxakcs2MQ3qdiboHsabWebuydwBdUmPYljLa9ROAPwZwERWDp8oo5Y9P6aWp
aqumT2Ifkot84WANxVgpq6/8J0EIq9Y4uMp+gRQIn94BeL0N3fCWjITTh30LrafIMzU4AK2XROS+
t4JvEwMaaz7QM9t/W60I8Gb5/hUf8UkpXpZLzMlIQhH3t+D+C+dZu/b6WqFKYcX8kJs/4fkgRrrG
/gvUMry2AehEuSwGwrh8vVF/Z8DbC1jmoUjiqaMDTQrFK/t8zcUqgmB2uFhDkr3xH6A4EQGGhtFt
2P9AdqkJ+0Rw1iXMdYdM52hbbC3rJ9AC9vyo/cRjPpRdO6wkqXhUGumEP2OOMxBNeh0+GeleKrtP
dkXmD4p7oVMi87KpAMRP2yIntS1aZg32zyS5iHMongMv3oaVj8IVBm1UiY7+pOPv8AFK8nye47S1
j6C1Dhu2W3VQIltTuo85my5lrgCu/hAUGmQVbmqDubAB3BeWbQSxJxu2bkCobNfo065J5MRRZD6t
Z8rFN7G6y+rn6dYdzbmJrUfMWoQ7vQJYKGB20VryXG+rWaC3qKLLLIroXbOHMshoB4c7sjofoH0Q
8zFN+M44o+SVsND+/2T3u8Hcv4ADwiJnuAJLhi/Btioqz0dTkdSeyTVFBkoZtP9a0ZR4F7Ir+R90
2LB/+/xZwtd91syCwEsaXYMqSqVKA7wAMv1ahuMgQp1fYnJ2100UgnGSWMUpfyA0yiQAdHjAKiw7
7ZYao92yzk9qVGH1g+kTMoRsrQcPA4gpw6aJ2wbFYFpx6GtsyRL4tkBBjvRQzTQYbEPhVnHL8CIQ
Gd3GL6A+1R4WiLp8YBwDKzMxTcQZw15D5lB5vCCbhg3fHmMMhk3OfD6LlPYQpyMpVs1hDgI9TT+E
4yZtTMLY6079sadztGrSRuThoPbF30Qz1GEplPkChHF+VlXoDI3W/kAj/T5rS9loNfRgesSY231P
UY0/nrvouMZ2BnfQlx4oha40NGYWSk1FqFl3mHNDInyoox0oQu+8qTB7/zY1JrqFZhcSLAeD9FtI
Nowu9nXVXUdIm+RJlco1t61Pc+FiGcQa1ij8Ifh2EVYfrynwoCy6SgT4SWqY9betsMPLs/LX4Bp3
uRHE7LQF22r0S7zotYIU+4oHOT/Ugc9/xAuWW3/l2AdveE8K9L3nqZxAGvfkINaEoCxj3tp4dIpv
1ynYTz5pNcrLDYDHhh8peatrExiUJNb6nvg1h15fedqzddFxlBPB9xRhxaFjn/CR9paU188ZVt22
zppTxU0w8OGDFhFLvETsRGTsjB0e0z6At8LArHVL4FGwx7APzJQ9NRdNR65KExZ+GvfMt2GG7WoV
M6zU1rQ+k7Hs89w4XxqFGcsLrLn6GzmHoH2lAwzjgMpf2GF/RdLAcKKcIT5Kge8YT41HNzLxRKa7
lLI3LA1Cy68k5RcK02c0EFBIHChBoK6thpPY8K1sEHjothPMX4oWCVfNQzS9Pc712MVOyYL4Yu8t
KAlh53kYXJgGMl17DwZLoTjuy+RjSPi2UROTHsMhzj4N5dE01dvu2cV+lbltd9WXt5ztwlu2yF4H
iZJFPV8tjTyJUakiO5Ys3pUTp6izaFvpoQuzaZv48ZCPR0Pq0ZtGnou4F48ibW0/s0tT6iDEs+yy
Wrn5hRgaOD+hrQTIgKndazF4Txw8YkjQFdd+qIOQD6IbQHxP9dM1M3oN+TeP5uORoBlFQeI+BMDW
mJ06bWNBgDgzJhLfax4ZJHznK7lMcblrRELuaYsnRR/CDOenW+YI/2o8MsYGbNRVyb2tH4dzy/J1
ftO8ReeujZ8A6jte3wijecyvjXq7XsHY6kLTBAVP57A6kvc5t64hODJpjNKr6xlEtLR7EWfp0LPo
0jg408PhFG76pMGPE7LQjfAxouSaYdpHXT+ZnDw+bzTbSgd6n2cfqgib6oUaN2BWfHx689MfAobF
p4qMgkyroB9kjr1iWIu2ZDwO532daP28qXFz06XYMCN7Bg56YwU8Am0Q6nj65cwMhlKj4u1Dxw5b
Z1SW9qNNgvWwt96Y/Co5iXQWZEaWI0YU6Y9vG6Ba5XPW83ZwFRSII/iIacYTZhVz0aqmJuG+zvqO
XlN/xW826aMoMeynY2Uc9wBoZoRGvdhxhG0emFoqZNzenD4XnK8QH/sBXoNtMEOO8oGya3aOnuRH
P1Yt5ABm1uoFyTXyhp4GwaL46EO4rqUuDUCPe4rnj7F43KqU8R5KRYwrkccJRbAYJIesvu+ggrdP
fP2JwEQX5EwBAc4g1qEhbpg2WpZ6QiMi5HgjOwOHagrpkRCQ3bZZYBa7IXqmkedWBmdofrdSuE3d
N/RAD+XGLYcZ/0x7cEnqvqTYx1XWEh/DTuEWuS7DoOmg/B/MpxPHwO77E2tiUIU6p+AjJw5jgqn4
RSNubrCX8pNaMEmrWoQhNpR38ThjTG8yWHyyVhloBtLSoe2RMwpXBlIeXszZuHVm2P44bPGMzsMV
FmGC/9kO1GR2iNVX4V3Dh32cmBGB8roGWj2Eh9YTBPNWfd4q+kMKM8V7wuRxF3M4gh6Ww3nIW5v0
FsSqYmWClBV+Wh+eB1YIzX1smiOm4kJUW+WJE0Y3/JD9tvYfhuZU0bpGrUppjpxo4u4D65J8C++k
fHFxFm/1JeO3MOb2Z+locZUb0nj/aDz79mU2bnXAux7IMfEdcueli2KhRgCmQvdNED9urio8XoHu
iTG+cv9fXQViXcvkJif0ylQI0wp3MJIjGQW2hJgisRTp0hBOeaRR2KoQZHxHhxRo9PUMRmLNCpZa
Nf3tPICmF4s+GUzkohJZ2wWoMgD0/BQdGg8VodZRmPbGTlL3MG8gNOOUJfQbPlDCQOSWcYkj2mPv
VyOuyiizoqy9fx0T1CzKOE5Kot4oYdbfCYnG4evJuqIfe8bQtBs7+xadPLU0Xvhi+Snr6Jv4ww2F
lvJ30Kn9QE2c4jv6StNffHu00neeygN5o7FTJHioritlKIoyZ6oMtQQuoEV/KK/yo4uAm8f9P8Nb
SRIFjgNp0tZNrnM5N1DphJrOpe0dxy6xZAu6CdAfIT7n6Txwe0SPf/04J1LycqwmxULqi0B19gQD
m3p+hxEWH6C9jxtGPQ+j6HQgsaRS2lt+ml8acmsoXmvbo4oKWqIaW+hjvX9UvAPFIwbeJL3dFOMf
A6/CMrySYCzE0EibhDMPT4VeMaEeeuEayu7/5OrR5EldRqW6ePZ7UbqaapdMX85wAUXeF+xk/+oP
lVtf4u5DxPLd0Ecfr8ypYumokeNbbSodsWfRwdcPBLADaCy9bj7z9UFzaDABbxHURaHR0aNUSCN3
b08KjB3THNps1xKyKhesIyrwARF3YhS9k/WbqS7auaEG0pK+QH74+84D4ubpvXvmYGAznU2bylxT
QHWEWq0NmkE7mu5EtbEZTav3DhvMrRIlgO2U+aUAQB2quY2JuMVjsn5BEXwpISaY1Ahli58fBGpi
7WhfqN/pMpzVWndY7svfoJE1717X/8qy9BohJz7LwL+31KbIMjFOWn/tSXaEQvspQnvAdFstFCCF
V1ejBSDC0xgDZ6HjEUIUMvzkmSCyMrQYF7GlNKjLSBzRvkGiMLgwj+8ct75tIhXUvSFD9trrSW4u
CuD3xdkPv84tLyNPU+KuVEbqtIbbu97jxaAbHmhStQaWZSd01X2Y8JGSQbYguJhLX+Xsun74kMpH
GlnVGY2rGORMDJrRD8y/O07mRTha/PaDvUFBgOAsdp6ZAGj8yZ4KJRJewpKjAGVsfd1187R2ywnt
lgGkoJkXXvhiut6MDL4uWmQHDs7ouyh5qx+a+tHC+C86yIrOOGYxPl/m2pUQ5tddbIsMae0UrxPx
IWJ4uBSY7Gn5npilfxwo0yKDUCrAj2noJVD+5LaDIrEwgopbJt2evWq75d3H1PLk6B5rc22xKsJt
9MjIBvzOrKd8F0/jMYj3jm3lXjCwb32FDQJw5OtnPCm0e8OtxzBOuh2pozDioO+8hRjS1H2eY4fR
T8tRcNnAxjv0PHeHllgdDupkrs9HFqJL3Wj5vo5Q0E+QsMYvg+vfFEkeKfYDHL0eGs7IGL3oAIyH
oj8pBIlWLDLeExJL5vYy8VgV/0sQ6YUMJdrrIYnIMzc0vfuv9vOefxIRjaO4JlauhccJPdazCDVt
fT26zQ0mitj9alzcfGnxU+0eS+JrTefqU/JdsWbTaJc1Wnxv8Fsz4Lx2DuUjPYOLYiArgLG2E9Pd
xSr/afXZYNL0L0yHV1UVCpFviTgWT4Ge3u3GAB9hpKlUr+JwtMgBVlOihrNmK4uUHRsTVQ5LsVyV
905SyNodO4FqsXFqvAjZW2d2ndfnWLaxGs62meLZVA5/6iOjGRX6Tdpc3ls5dAml4tIVh7CAw9Df
QCK7Gxawf2gNREPkhFjydi4lC4fctxdJpqKNR2FFs1L73XxKKOk9U3BT8mCsChY+VS5ZCmK82avm
cfz58se8SGgyK8wSZLtfAoyIcy86XnqAYVgla2vRUJNF//QxVXCdhOIygBaZjHp3PtCBz0P4jGEh
7VRmMvgmfTBckNHaxwAtin5gdiNsmPUJ2BAfP7Wd5Y4zYpWFVUlVqH5e0iumPZiqQBtj7TAI/Ogw
wcWVz0lhvTm0Nwg5NH0wnU5eCpieFYn7tls++LXBoDGf3geILn+M2HUjF7jzlA/KK3QSksD0ROGo
bFTUernD97gFM9oJoUqvqpwURbqr75cXikEA88e4dUNg3nCiIhymTrWHLMPDBXtsm2hQi9tfihH1
wLNicfXRZfCjt5F2p+08JUKEIL5gXe8FQn5FSWjPC1IRwnZGL5SaHcsidEhxyJlN8Keh6EADgAv1
075k0a39WhToYY02qeJHHHX6jly+yBIilqZjvnDj9hFePDTuZCCn3J/Krg2+LgJ+W/XSoccH6Dmd
uSjojDz5DbcYpKYy3LKZ5Qr08VU/RGfq2YbNepUUl7aCp86Ek2s7WtlmWC4cq5pItZqXKJfuMtTy
0otQ+c1kjH60nsJVDYEkTw7Pae7JAwwabRm8joBTBNY0ulG41mI91VTsMynto02Tnlf4mD9Xr1Wj
X0uhsiaap3fCoT7M/erzyWNk33QDnggesbhrdYQyu9DnG9eL72qH5fUpai67y2nGP6xDoDGKIi6C
eNs1HQuz/0Pk5Lyx2c0wQ+BKL9Vbk+JqsSjCyDy0ShKt6Sh9OMiu3tDDHwENaLu07x9ubfNcvbsI
B1M1cWzg3HZP3vE8LgIk4HkJImEYBoMS4+qcZmXplSBm2gmw1rF332aCX+8xB0RdPaZ1qI4B252j
zhoKpKnAmsWMz5A/ZHO9zlVaEnZBdH/PKv6B8EUz1xMgqkenDgSZyZos3FjLogVbLbyE/xrNkoh3
Wx1miiRT6sruFVVNJ0IW+qDXuZxRS3hixZoSVwzVTAK/wxpghNXt73uF8JzURCKDtDr1/jJUOgOq
idTirMw1wj6b68orv5NP22RklOLFCI8SDRYy9kr2DZ9lIioeMTY1m6uFLYIwBGSIXWyElqRxO4Yo
GWl4jOGvcphIBnJ/leCojWqEiyX2ewfKaj4hn72Nk6NDtE07MJ3C377R4C1tyCE8jH6mX1VU6A0j
b52gfaISRzj4Rop8i8rPoBlOLV0RidzEIElbMNPCPh4ZJfcHEE1YjufPb+SlVo4jvb/g4k5yHXRO
2tNHy/+/pqRPa/Nq3XQC5l2G7KjHB7KoXOkQYk9AV8aROp/ar3oe1/ZYxXWtUUj6UawU09R1tD65
iF8mp21f/ZqC6L1NFf/96MZqeKnllExhbigkSYappUi4cpHKY8H5ZMV//+EFCsf01w2eRMdhX6iM
Uo8lEyVniK+DPIEGgNozyfXjq/sqpEajpv0uupURFBOoRRCBqzJ+NaHkCaSEYfkd4DXqB8HUzYX7
rkcLpAtgXFDyh42Hd+WWJbJZ2IHH/9bNiWZ1tbodhxjbad4TruOkP9x7uqm9yPrM2y91FueJhwys
O2UI0Bxpsh3H09spjxQsW3zOFuKtZCgjmEkn0W8zVOBfgdqhlSF/0YB+PuLEtyuaAW2N+bADaUzO
5s1UHchXclOZ/uJn+q0Xz3IQ6vCshLh2nQKP1+NxKXSbO9evcX71a3+8fUETefdx209RPdFFeAaE
bJzcDqpAtuARPNd2cFH03M5RcZXgylgjvjJkk8omFVbG+6Pps9uG+cohhftiLDCGjWJoRestPnzC
03o8kJjjPdq6tQR+YHTi6/sTBhhRCBEPI1Swwj15US8qBKz4LPNjNmnGIRN7PkDrK/AV7+Gg9RMX
yh2oJthzYrzNkfnTQfXJJXyhzjQLYFpM+Izg3z+ZQNRjN88TjvY5Kn9kaEbJ2wXc+8EMtMQ6UXkr
HoG+eSxHicXC5uBUrtfU4B3TZyn+Er6iWuuAjNQz4CnnQzBcw6y66CynAkeTkGKbJJ8tZZB89qN7
KKDtPlb5ciJQPlEvdhsXjv+at6F/Z3Xzx+hCB39KD4hg0gYB9JWaM2HIJ1tQg0dz2XpQBC+ds4FE
qMZw2FDlKkqkvUJZAaoue2mn5kn31FFoBFsxfiM9OhcRa6nCuM6K7sp4rQdbaDmkTFCY1G6l7VcK
5NXRFfYEAxy1A8jqeU3XN/IwuZONNpB28WnewJmr+EotyCjEAZQEgU67zrpCSRcW5rx2jPsmbFF3
Y/OI5bbYwW+AnNimwgPd7HeA6KJl6wRpXtEnI2J+TPJs9J1qH4vQOkKsgqneZHBaRQExQMhXMZxZ
GmzUAB5M6/ZstKiA8zod5Wu6j7/eXHbeLsM16HRNFZyHxeo/IVm7b5ojuJKaSrJHAk2ofhxpoc/V
ApE9pKJy92U4EIYaB98rIdeQzTzDXhgNcM/qYOPPSHtOBhF0C7XtJ+1egtz76qx6DqREDQ9yyGuf
D5PDkzlj7mTeyMje5cj1unXEEo7Qh+YDLy4QKgCC4ZXvOEnFSZ5HUjvifQb6TCYctu4dg9/N2XPQ
wx9oRUJGVxF1LQ3pFU3McHP4iEp98bspKuzT7aY1lppufs3Pv/XOU/1mDZoI7KrxLfn6365l9Wip
JBB2ZFBu4vqw9x0sIp0R0aBFqxJaOfgHen9XuIfXfyNlZsMqRI47yyU30oDO/fIcFntcZAaxldEF
DxnJPE+/1HVo0RG1zSOX/0LabLaGkGp1ANrd+hrJky1DaTPkvbF3OUcxO7vWZkB2W1goxirOz2h2
QDWq0GmhYiV0k8aJe1P1rYpyLD/u1NDC+THMLz04NFJ9rViyi9Guu4rB+tCCJXD2RT6HEiXiFTkv
5GDhGMLXurfA4fbGQ0I86gytOwMhrSozAHdBRxPCfH+25zkkiZbkttpzts80wYqhpnTQkaL7xaUu
1g7PsF3L7a1BPZ2/p7xlHSZ065vAGHi2i4TJIp41OxMO/zlR+YWdTT9jrNy4wuj0Wx9ZQJcPExl9
900J0BzWXn7nPKPnrvoUGrAIPcqvsw/+9/Mc2/vB29Zp0iUlBX79vhwOLJ0oA+mnK0N03pdkG4X6
Krd4LuQGeQHFuwCipmbqUAdET8OPV6lL/LEtKKs6ZahyjG/3h98uXW+7xlQq9+EP37pcwrsSh0ed
ahOtdGqS7OO4DhICCmfS+GBCUSZVhFFuas8QB8utHUa0AYLC54+hw3Z6A484LXLEe994W3ov819V
K+/S35NKMG+N1Y8wmxs1Z/b3bOfvOpjyz04vF1GLjrR2JGDOEYrTMqtWLPSdgx/dlIygn42lvJ19
U5aL3847PvqF1p/WDMOv+V08WowWKjq6jMWhj5peTYdXMu2fyV9tR193tm1yYbiaODiVs2z4VC07
YaUXbPGCka781qs+OlgOscBl5zoNCM4D6jQ6+ao7EWyZA92ox6OavIp62vgvQp2HM2KzhXuSGG5p
72LXLx6nNn1mVzuaYpCCkZujHBNOnvZxQjKy69/HBqTh4w2D573JzHbdEwZlpxM9ipibibzhHnAe
0YaUeQjZ0ZQopWKcQ6ubg/MP8SpXXBe9M8ValYQ8Bhf5HmQCgLbPMawrknvunyBxCKrNJyQkIxZW
xrPKmvkfcjA4DK8Yk+nPVJw3G44MHuwxwzzKHE8wN3f6+1/4TbcFEaan9LSD/OOzcS7PAKrhqjZt
AToENKPagw/c4IsvE7B1FSuD2sd6VKgYsGytOl7ry+tNtcH0XGSfjaAoK8ISEjeqi5DtWeMM9Hov
jhsxTLete/yQUZJkBCjGn+mzN9tCQHnaZRZuZK8DVCZ/4dd2n09P2ZLlekfnkPe7PJ3FIpASoSTb
41p6HgB2zIqzsl2AWajrsogf1oEKcpwnXqD7jTgcbgV7v9SQ1w5Z+6T1aC8U3u3rwi5EZIOghxrf
qNFgQSCQVS1KFuQaiWcv5qHjgmpYNW43sdE8RHH3Q170RrAF5Y2gFQFDF4vlPeAveyPVwM1Xegzh
QqLC6Kc5tWkn7DxINgP3+S5h1lJq+6OkrOh8cWfPGRgTPjIJaQJZNscQsMVIPW1wi9rt5RMPrBmw
IQ5wAOHIp0iE7M6p86+QeaiZ3RxHOlzXn8rNjJKCfAkeYon7yH8Ua6CRyk/ekRgQ/Fg4x36fjQRy
wbLEWV59SNwhZwhApf3jfnJzFVjttkvoaIRuaAKnula48IGDYv53MfQ98MlhJ0/5SxC2rpud9UZA
JopyfpwBe0O0YD1bh0omXHPPNtrr3ty1EZyzvI6SymNJ2UOHdiD5zFb608HEniXlBzva5Mdm2YMj
6trBb2jcgaU0dM/JkVEMzpOZCBH/hBdHDw3ORdAJTe5PoXPLb1th9zezT4w+Hgr9FSGEZ9py8vcj
0HnHzDOb26MtAr4MxSDNljVkuDcjvidRUBf3VXdU58XftNJJYXl2cy8lYp4QtRJj7fKyy+EghrOh
jtqJ7IZfLklIuci6VE75iFbCK9AGYbRlb8lxA5Mz8Kwsaq8M7du/5pxIhrr9AtNuqUVkIwULPPs+
UwSHrZFEAOv673TNPYUNDtQeOg9Baev6g0UytHQfIHc7yHfoGDpoDidFiKJARSmLX7eI1n02MOBm
aLFWQ6LXJhbO2jbG/4cpirKmgtAcIsMsFuGlbcPczRx6UXsYYHa0Ig4CQyjtjiSsVJCtmfRtzPs1
91bMLnR3thssiZyuECYwund1cBgYBP5FKC3G9QfzR2+gnZmnePbgNhIDF8rpJyf6ermk+NheJE1S
mCx0xORxy2PMDLxCYX9mbExbSH06FMdzFFZZTIoA6yl+XcQdvExBkzbn40veLb64Tch0112Oq1dM
tPmrE+grgWwC5KgPhkN/h7c2H2WG4maPAC4vXv2HX03wgi7sYSsNd1uADaCukGEXAOm14hf6/4rE
lSeQcle/oFHziODBrdj4PQeKhp+hhuqF2Tr/3VCnu9CrkhNXTt3fPIpgV9KoY9oNbrEquJEJ3j02
t1aOvlGv2IWFmEGUdmCwN40vNIvcOFD98fAd6FVr4C7BDGZCbkrxmjYSA5S6gnVUcjqlZkCuVBX9
kXdcZeQIq2921qmpOfYAAxW6FowE9wHEibOkVm3HIn4M/BsbSKExhwdsMmdckeef6kgIOYcfPDBm
QpjXmrLhdtLKTJPUOYbXNjPxq3qvIpFlrr/w8Zt0+bX2hs2zrwSmeP/5z1OqHR2srMPb3s6jql4B
Q154gTy6rqQcicSFURCKhEUyUPN7QbrpO/bYNTPBL1a1xAylOJC1FgvDhdoEl7OIq3ZnzNsj63+R
hrKG65Or5Y+p7BUk9pCQzLgjGHnsCr4mPTZsBQiwnJ8D6O7Fh+t2O1spytjeAfPXORdwdYm0to81
SbzPK2D9thS9qgVFNW5pC1i67ZMhNnfiCX1XD3vA3oVPqxQKy3DVJKKtlTqtB1DzY/AIopJQ4dv8
KShrHOWTxZCnFnA7wFV9IuFeHCeu8HJBbWR1/wXhkzyjFXCzt3yF24ejFIqeCM11whf5A9xRIXEV
r+sqqAB0n63ZU0ywe2FZ6YLxUWhI4CL+QP9bEzOK6gBJ/aiz3QelElZFG+PzqGrl1ClyMDNfzQT3
rROSofDjmXaSiHBdj3bBhRClUPjvRBlIbC6dwSvfqEbWskf1HqLIdAixE1UvKfNS+eq1WppS8Zd+
vOOQ4C+JvLVPHRFDOk5u58ZZch6fXfqPpjVtmV/8Mrv6oRQCU2bT/SmlvHoyagWchv2zenrD+4Az
YLKzHqSl4t7C4Q6y5ZhtSEx9qIcabl4E+2OIl+KCOF2XgSr/VEBDElPbeONkwhPRzXphstnVnPs5
CS+DByFlYkFicxPhEorV2h0yKx6YBS0wTUO6nIgZaeBVBxDdkMaYgNhfyJgjT7yXYwZ3hRmWXUqa
9/IDJSuS0aS5AGhlw5C+P/TvIxeeytXUhp8qE6zvsQRSb8nFFvfAE/k0SWJNO5SMnzhnv2Jhv0Co
UTTgnOZ2VVBHk/vkPfS43f4ZrO0+ejOOCQBv5fZHcGr9jCLMNIkCCOMzHTa2nlzw2m4FqvHwG14m
g1YdElI7rfI6gyouFDPE/CXddxVlfZCepmXu7oHWcynpSdhcBc2l3VzGazx/RId2xUvqB4sX2xQg
A2rev1xBQG8hPNq7ee2vrtBE19u+8xNKOV7wTEYxufpA0HHFayL3d+YWnbo028MX+NeLT2DXexX4
cqDgAAw66g0f81v3vj7VNEXhYbB3z/vSTLwZRptD11LB07eILIwM4eywjfvK6HnLvZqc/8+KTmHG
aRzIYrdIxXmlIIFXhL12JNM5qfsNQkHpy8ocFYjjDeakeBa58M2kcF+5egQIJTa3CFdlNhHCz7ga
R56DB56Oiu/0uggBcOypPYiyAIrzGGnVNBZN0yNr2+P8oTwWQ7EID3UsICOGooxc0CedxgIAOMhj
v6GulDAUlf90TBoz0MbhoVDWR37dbieBWfsIv1a+zHufCDDyu1/+cADhoNer1AswvJyzzKoRUiuk
aOxa7XuDDtDj1mSe6FUlu6ptZr7FtdGH25YAEUorJkDDC8Q74BK/UqPiK6kseNDYwbpDHtDzQFli
gb/oyoEkB2A6v962mDPlQexnZN+g1JfgL4rKqe4J7x/dS0lEYfrajy2zJ7k57GjM4WFt29jKFxuy
XCxlMq80cd2dfhctC+qH9uIDTka7TzKUs6CvZTE5HYsj2VtP04ilOQSoQQ7vpL3De1a6KCz3wO+A
AjjvDRWGEZOQpxF3dh9fckYZCHOAuCaUGMkGAhWMuLCmqYvIgHoHj0a7JUpaxcz9TPw+It1BkUhm
YlzFfiUFo+aM+hvcqNWwT/wgpjBK5XNhKW5KoNvi5aGNDiyVoILAufrQl+vAkAYc6mAd7bqMDkaM
QGkPbAbDj+M9ultaraXGPohLBPlrETDBz6TWNe/sY4EtRSK066O3AxJdvrZWzqbwyAzo/ihHrycr
8ceNU+WMIJCV+Hhs1pC3p+lcpqvdHn8AiLIkZVk6Vu+qyOdRC6pc/EZqylMT4Ae08iljeUG7m6kY
Jr+H1DwSb/0xDdSL2sdr/FDqUeTGHSUH5VvwhyppQOUCb8wsJd13Uv421QQzNRhRQo4f2Mg0tgyb
XtfDtV6AHnB/x6+FSYhO/Egbfv/Gf8bc90V92XcplYORYCHZdBxc1L4tR4uqcuQqkvB6ohrL4cxe
UNAuOw0I8/kVlLGxjH3dq0nQg9RqtjW5494CUl5C0OXHTtogTXRMHAvnhyjU25GXodLhii3exm3M
Lgfl2/gecPDCB17PI6eF2CGSelvkC1mmGOwffl7B1ExF/mi0I1ktJ7ZfGHbnvXrOf2kcezEZAfcn
BVdyGAkmP8F0P5rV+HliOT1z+pXwvIoz7DnwTpQjQgrCsJ5919qnYwmIytEP5I7DLsfcVoYhScfs
vvuzIRvNJxK2B4sfQsbbunXpaO3S1WgE3ZXypQ48jH95Ju0HVfgEHMdTBsPNPhriMN7aJS4IudvS
FdIAh08NkcWC7rQ0zyzpPbaxsP5lGbmL0nLU18pNQtaSA8/ROlsT0NIeskVkRaADp5OFICSw7Idm
jpqdZ+hp336M3P1nBnf7JL18KknqVqQQvSltocwNtv4I3mh6R6v7ybJo3RT6nwPa6qj5X9OFAZWc
9lqgRZtKOxZienLD5wDPof4Cjd73/wkQtZqz0FIFWYzI0ECC6l9g0JNqtdZ/AdeVYb1S1SitQ5Bx
HWOIeJzy2hQcYLS6kvfLDlA6NpwY7ArUkE0b0ei/lEi7k/ux4TXXah1+DRzmgpXuHGDIFLwxUOUi
Jxh9hJqFWKqleJhcQwJj9REap26AyFKgU/J92tP7U9NkHKQHovkfJE0jLkvFfwIDOpr5E0ULtSOa
N6EQ2iLyYiwOZH9OCZDYpL0UupegkJ08w/45j5MjjIoznqeeBeLAJ04MyLuKc5ytsHMq8L2Wcsmc
Ws9OFyH8W62I55aBfG21XuFznWNeuU6z9OXzdVsanZ8yvYqjgOTIHEvHTSrTlORLC8aUoCD/iTvH
Yca2/5TihEVdH/npnggi7LeEMQMsV2DZCOB1B2IKaGSWPhsiywlKb2Mk5K2YekMdUJbgrveTgClv
dQl2mYuZrosh/PKWUI0ORMFIEHt3ZlvzqQOwpViAXQU083egkVGQIaal6UO5pwLg0yYRgmMOyee8
CXqEWZ75e4GREOXFmJ2uwyvsnGryZzIpdE89oVu2WBuaxRSauSI372vhy3oXUVuIsWSYy5pUbwVq
zmrFxdeflDQJtGTraFToY0Guq7fhBBfQbLBu+c5whXTTJ2v4w4SE+7TY8yHOnq13ltmKGtF2k/ea
AGTTjNHEXErbtZdqXhkFyJGacDAa6IuTVD9WaJ39+NFdDGrAQA4NnstbRVV3CL1toVThs9tev+n2
Irba0cq7+ADw7WeU8UvtM78GAOFgP2Eq4szB6ec7B3O/61woSCklsVJ4ca2QqmY2eAFgRv9UCpol
MYAvGNDHOIsugKwmnCGqib+bEgTjn1rHuq4psC2WoenQwjXG5HXK/Lf3yn0B9/EJRaSPFXBNUB9v
hpHtrh+cAJ9LL8IGFPLgRD2V0Fz0UPbPAQ4Jb1X7uDtaMZ/ljRW7YyrR2DKwxiZyRnyhoFHMXHWk
X2Sl4sU/JS8jXv/nLP8PcumkUYLcFqMQ8Q/iu4EqMUgw9FFTPd1Sc0pivTrZRZ5gCIcKIEmuzBtC
c/ZqrEhnvvFagK7biukVBaGL1BcHRRjtpTAaZJo6SDMOQVID8vwJ+zm+ThPbJce7AkLD/sxc0oNX
I9cqdzBn8qtVmwU9+hJmif7nJf9lY36ocpYX6Kly8LfF2zHeL1GWNOzJO0EdqkZHGbOdBVLwI07w
9GCLqnvKPR+ZgswZ2+VkNJH3BajuryhEJyFkuvxgAvuDduTgRF7faIF6oi3c+H+hU6VmUXrDVcZF
HCENxuEZaI/KNd2xQT2CkkhpiUl2fH6BZa99RDrrhMQv7hgm9LVORx4llrQcu7W7cFSSq2pr6hrP
GP+SI48FgyG+mfavQ4RIsdeAa7BjNbFYa+cbkrrFEc7v9IPKkQtXl4uvf9Bt1DqrmyL3Qa8Tbo8X
UdAWbwGZRc35n7bWFtRfGnQ6CRU1StOAlrKzd+EG6kynn7DvXGJL+3cly85kEXU0KeiiCeoMMGMU
OewaopqkYI5onM38DRyepcBGt7NQqOHVdnBpbgZdDg8gS87mUXzccEcLkqtxId+FcaY0ewz3c8vF
M6RASCUmjOa1HQ0rxRpY+RESKLRF7qZTdN9wexPljY/ZePoVgB3Ra3/P019HjLzhEtoSc2WCtydj
4hBoeoMmPdl37tJRmaYGpjEJfoDXieZLRQ698NZPKwh2Dp6f3rVUHvZ3XD0/Kt0X9CVNeJcV/oWu
vPYbd4IwDpQwAp3rPPkMq7w4Bduvq/IwrgbI1A/lkLcCU/P3nUNTRZWpM1Kx4H8n2bu1LAx/J8qA
uzDP5rp27YlLGvmNNNyAYeHPdFgnnhKHa4Q3zsE4Rzchwj+tiFHN5bphH9Xd9C8Ue5wEUoBR2dai
7FoHLliYpoAv4wrMLmmkfs5RVbW94h9SAakS896wurHqcvBkCVe6Hx32XjSu6CW3wKrLUWctmTZ7
JPTFgBGRnG3XF0mEbe7GFyRlfPxFun/frSrXh1BbQ8zxS6+rQChoAVE9zh7YZ7bCf80ZsGUnSwBS
/EUC7v0iKC9/cm9fjXswJ9n6CzfZmobGxu4vJKXBCtvQ0tD7h2RFBLydT6Uh1FopdPaZdS7HUN/r
MlFji53Btq2psDmNOW4ty4SPaiyvQJoLnh2eBYTOdU+obciWOdbp4LD81+KdxMFT/JlGfoCvIeHq
C3Tj5Js/ua22iO7dgYKZ6R/n+lRv/O8ZR9gCQ4BrZVdr+gYVOlqHadYBsKRnp0bxjPsWBLYY5Cqz
d/V7nSbfZbSxXzylm96bkfahtaQfaFAhgLA5M76AhClo0VL9wDc3GGVkXO/VEprtCjiVPQlX7ASl
aNZcsBO0tAOGkZW21Rax0zJzksfItzS6ssrGYDQKHUM5L/NhWBd2DRPk4QKH6pfjSjCWAF7ftY2B
9kz3ITmyhH3F3JVjcYmVtKVD9rkit4YYTefXLI41sFDHtpWd64uTlUJKF9ljsDqUvekJuUkqGLfA
OhnDm7GJIolIKETEHSQGg90YuO2iJyhTWe9IF1UtPaHFRKligT5VrIs04vOxsQcis8ML0rWQ0EUZ
SemBvkb6n+2SA2vcDQlwhX4J8FG82AKMl3w7dq5rrQdIllk5wDRSaqPWjbUfYHVkMudKLG/zKEuv
IKg5r9xFvoOXB0uB6RQqpjDHOBowGj4kxFR0NVBc2HjTXd8iuewerBvezpsOJ5zeaygbYLeHD0dq
sSDrI3+ls8CaThfAdFw8bV5SrhBbkRB030H4PopYE1uftsj0vUG1vqCgaJUUM2DIEyyXu8yTWXCW
GzvRg5maaDP+a7WLbdGl0AJG+Ezq7bxOm7S2fFAdv9tnoPnC3iHQOUjtk5KUtdpsFsWQ2GbSAsaG
5i0mpUP3cCb8ws0bkjNS6Um6fRfakVyU+8osdlibH29FnQXPyjwRJo39/5okfHxRh+CjS+yto9wA
2aMTdL9b43Fpn7nX/MzpqwzRP7SpbBNCCK7ioqhnZ6b8WIMa3PYPLVTWPvVvlsB1c997egQPNWcX
bTQrCgJJ3eoe3ky1YQV129ESEklHM5lnScaGKuy0z4SFN0L7k5vc2b+GMKqYt6v2gCC0IJ50MnxA
lc89gEZsw3cS1IBlHFpDm7GJfYIjKZoRo/l6sI8Jn0jVw9ymDy8pH6JJ2oIB46pttjZsuxXaDbmT
um+G+NEV8XqMjPXc5VL48kEAU1Hp8kNK4Qqo6HwSo5HDrdIptVsLlUxX9ReUPv7jjZEC79Heri6x
gAkZ+s1oNUyH5bWWZUELk2l9bHfIalKJpxQsu/RSNg8B0qD25VOClaEPNusrDa+uWmfM9NvwwRVy
rIsNNb0EVEWYcrfmnQoxkdhTXp7CAHQEr6+PXJsyCWJUrLM0AYmAzjJNJTGSHlcF57/vDjvaBP3L
8qqR+RbJgEviJLstyaMIkUxJMKrIMFGQ/osNpeRuakH0jeXifhUVy5P2In/ILSZHOnegmpagIIjB
mgyifO5mVtXkE+vVO9vCOreJLFKETEMdPKekrwN0D9DCVc1iZfckTgTJlFNMjOeZKhmYfYNPf4O8
/43D72dIH1un64Jy+9IeDI0gWDcgFU+hOQ//EJqkqLtlHumQiRQp2K1BrgCviGWH2a8JJJnqIjyA
OqocSUX99w0TragZgSrdOMzUXzqOrOuBfoYd+kGvane+Q6t1nAHzBAuFTrPFKBHoaQumedUA+wfU
6FC0cTZadRzHrrLK/LKFXv/p19Gch78udntuwRW6hPJXe58PLhdEA7HiSc5bJeRPykd3W+XmEgpj
g8g79w4g9+4JqdnAf4NIu+R5/sfUUQ8Bw1W13XAXVxcc6RqkHsUZEP50JKJU2nkMeV0hyugpv9af
C2/7BYa81gYtSkrT2WnhlYCLGg8TPeGoQ7uavCacqdaQOwx0e5lx4Wt2yKNMc2TEUgX4+8qgrsnz
riAqX2RG8melJuo5jsYhsU8QDBXqQgvO2AwJk/Y5WoCpIRg5ZKrwNenlQklmWg3sDgscfD4S8OxU
mNnh1fKKob2LntVtSPkCV/k9ka8Kai38ci/F+Yib3ue40XfBJBuXTOzbn/6jLbfpU29qkT2+HTc2
6J38+DErY4RgZ2SVke7F6cKTw3bF2wPAvkDydIJD8JPpOJHIk48dXDopEFy1VLTaN/83LmF8joOM
7Vqp+jKRzsUjgQCSACLdSR+zai6GmIG7KY4ETAQ3+5L4bUDMWMN9dDi6Tye1qHyO5n/evJCdiZtx
o/r4iTxaLSsGAQITMnK7dL2bnwCKjfA68QAZg535RHHfS8ZjAu5PGgELAzKpBnHi5tFHMGRt9/0o
Da/v/yHjSmaaHtq/7NQDDvYxfPrvkSAx/2zax9pVmlQOWdEDyCMUJi82tMm2wHqaOHX0kyMVKu0E
EOzr9Enza3CuNROmmDJJpRY5LyU63Ge+J10STL2T8e/Pl6+OxqD4KlW30n4F3PsvjlUmT6vR0oV1
K7sRg72tTatdUJsmyhXLwIqlZak3pkW6iH4MYp9se/VFD1CC5dOhPuaY77O1Z7ojVxOGYXHHYcm/
/Vst9RdnP7CSMq3unouEmnId9jAup6/ZKnSssc7OgagyJ5nXx1M6pHmyje2m66ht5+aJOxmmVN/3
dC0jCMmghp5lI5SWpLDDw0mTkFH6k8sjM0nnBWo+4SjGXVW2nGamY4Dqbqtigxf+HV29Pj0MC+9B
KA/3na8Iugl3lDY3srVyXNZDhXI48OCua7ixtw4aRngjGFZvwsLx6YIbAG9+UXbtx3PVbp5eqmpe
5jDyA+DN1GZwmiw+K6XnWvxr0GXi88+jR1D6WMxH/36qio1ttmbSueGvSZ4VMIaU556u6LuEZPpr
16ghHnSj24DlLcgHjfYjcm6AZQL5Y9U5LGhoBys+527V1BE3yXPCjyFGOpUugnYw8KK8tEuJtmDm
nS4pgO3pVQp/VKk/1aKgiiGbkFsR9OJVHdAP1OGN2D4x6PMH1jWMPWMXkXW48k5pw6K5baOvvEI+
rPXXIqFFX9sPUyFYkanhIyboe4FxckVU3iNDamubb7ZiB8TCzH3tZhNO/8xnieAKVALtwSFY/lq9
Uzk8u+DEnxCTEWIx1grhntm8Ui8Lfx1q2gbC5D84y1rnoqgtAGHk3gj+n8Nu2wkSnSau+wz/FDSB
cRxwAdshkjlyQJSEVCDOfsIKxCSkpSW9VCjdU3a7NemjCsU8BF3gt7JuAdCY+w8ZT2ZmBRBpDRWL
cxWMYU4xbIQyEAbAyG3D93jwGadbnBoXQJRBsf9zGRYJvFP8C9OMm//pikYGB59P3KdnBSavIWt/
a7hmM9k/NU0+nSSVnZ0hPIrG0oE6wx6jFWEcE02nA4Ij4Q/E4D3DL6XTw6uv7dZW3SHYOCDOlDdM
9AAkq62qXs4/86HU0WKtekbf/tOFlQUg5OfS1tXa64MSyWHELn7YJRYabWHGAKP61EFTWDOWyeS9
EzfGj+QT56ttOKCuoVXHw402G7+r/QR+Ro0lNID5sYCw7i1pXTewGOvMtkd3Bm761bW9MgFDwZ9R
2+CKMPeUdWeHkF9elZj7iQBCHnR+Z+Yj7GE1mpLD2AWKXMv85BG0blKyeCq1CR6jzDOvvJxgyv/f
H+lkkMy2RAUnowGt9zxnvhj9smoy8O7/9JbFI14PqAWXWU4v+ZIZnu9PWUU8z02sU8xq85lgZO4b
IsJnIVPIVA651yP1cKRetAl85AYRdSlP/SDKOhuGysnIUKnfe8zQQhMwBsuh+VIvDGNoIi7QbsQM
FEDDsxoUwhS1mghSDoUwfGQ9mHwT2H1cM7fhntMfQOnJi4JPIeFtLF8hCzm1jtz+fPQ2mBV99rEu
sodkwRwIXBaaVI8MnkcVucTG4zgB5hWGkUr7LgtIRnNuFGe8KcJzpSJyUAMdunv0BHvH9/uU0yPi
lICcPBtoguT+bs1+2yCIaXFt52cN6J36OcdA+Dt3l1LCF/Bx2tE6jMds+dPkwJtXIH6Jjf9vj46K
XS1jhWRvfPQTrp+ocrEInQBX3tGJgubQwBd7rqa/54pEIqRTHsjNedxF4tXubQQKqU38Gejcf5fd
CE2QMXE7emiQNl1eSyvzFfTluPrhSHFZwRd0StgnjU6jQfJEUfbOAwcmIkQt6gpaVExfyjWeWeiF
pkgNwe9cGBhhfVLHmUKzuAVDbYrTxe3s+OUpWQSv/2JwraawMQzQ90u7NsF2VqoVsLpsIgZHi4Va
KFg63rPJ4RZZ23LHLFfwtZao98ZzZfnn+3FdOdXzrz2JycwifDgAQF9dBrCOJZrWNTem84DaM9Up
ay9EdXIt3OWAMDEFx2qb0YICUw3U0/mn0IwG/Ig3EancqYbG5idwcmzAWYd7uUmaUCato+B6KNIE
W+L9a+8a52eZgyJaUZYEud9jB0Shfax/tYMT6uogCMfi3oYQmFQV1KmFigvo1RPBo8VgXfBYIbWk
WtfcCIuarL48LrZlG4JjXIpbF9c/dC4fufZh+KVI4J2uqT1CH2rPQFtEYjdneuPKj3HB3xMXryQJ
HcYixig3du4rx7vaGp2rScBcJvYVFntyZ3CzDBunwjeC2+iqXHY7iQHdVXnmRXv733UD+/qYp9/y
65qJvJC6CXFphSIfwAGeqjBQywM4xUQitVtTApiFr5nVQeq0LeHnGuaBFI8xoLP0mRhBfOCBtD2s
pqJ+CuB2D8NRAFBivx/+6JoBohLwutqdefPE2te50rg+5ipVV3DLkcQPQTpEz7Grr1t/wm0W859X
HOP7A5oBinFK7AizTi5gL9E5MQe/lGrhWJgoQPPryCeoXkjeG4MnwXDE36yCXNip+1rsfZeqTuK+
5VcNWis5b8/yDhUFsB0GN1Gx8q2HLlmNdGgEMVpN4KHsThKMsQ9dQijUL7ygrplmd422P5VQtMZt
MHJFMOTVktrzkeiCF6yz7MGFwDkFKsDT8co5hO6gLZDfC8/iQX6XS+7BJvurZS5SNiLtZisP6EWY
bgIS0upXKgNFDXTpGrL4fME6XMFNGsJgK8K2vR9IETMpxgD2sEdW1eMhTna/zoCQm2GchE+foOut
gh0kJ8AhD00fknGgE24ggdlrAnCkDR0sNpsaMItk6UIkoE443LyBs6uBSDW94ZqgEXgutKNhXvV5
L+Hd13ksSbGcFiH/X9Dm1BAV38oCwQyYnNfHGS802iMff3pYcdard87Wxh/A28sxtRmCcHArdohY
EZpcOyA3FCQERlaeIVUYtvYYNXA9ieSxdmaYN1ARXJW4bZw2ays1V3WWG7id4axmYt933evkUyrE
5pGwe0Z4yF3fMamM56C1UitaENC7Nbh1LP72o6lWrC6f/Bnjzg4spsoDMgAHauuy3UXKlbYSPYCH
M3ToPuuAKpSKL+qbb2sVzD1QRlGwqEOHOW0jxGxIX3/GyAN21jfB5czYABYBnUWzSvTxbsSbxTsa
cohVmpdHa9ecboTk/SVeom9NvZARWAf4KvSQZvsyo+IfIilT6tvomYoFvliH+XLumCYc64MS0orH
AvCN3OYKPJzh4NPxSw0JGgsqogR8QgpgjRHrXZ+9hCuL0ruaNKyCkx+vTcgVV3Ukjr87SHVKGuXT
btU8eskexA/tOHhjN2AAoOhh6GV2h5JgnixUEmO0UQNlrsYhYitJRttIsdXPAhpTdziN+HwS0uGd
xXPfgla9ccjfCzzlmYe5mxvkfkdicdI8xyCXwLLRzyMfDqhpj8bTFItCfgKyvI9S6Y5Ojxg76Mny
q9+oRq7tUggTXWlUadapf5F9CR30wmqqXsFSQHZ5fVpml3+efjwqwBnu4AJFzbZPjCohQ8fz8j+D
1jX3qhX3oRwW28bbwAi4w7BpZ/jtdHfTH0BuXcOyhlln3ekCSrCb4Hnv0IpWzNievp8pB2B6MXKg
O3+Y2I6sxj//52Wx3UJnJo7Z5WG4vNPYohcyQKZlVKOrdyuCOTCLeUmRA2jqFIZsnWvtieiv/6eG
Awz50CaY6KIJcRB+iEAmATnw7Hx/b7/dgBQLs/5I4eUkDqYSE8WKSFAPEEbt82u+hxNnb5JzUlfR
snPU9Q7vLCwtVrUaIpX/7vDCGe1u8oHup6bW/3/JMLCVA7xRR18SurBjA5ETeXODi/NxokRGNicf
ad0ESkl5GOorIjsVGi9y6j/9NnqK1Uvm7uOilk2d+6V1tVX1LgfUO/AdCY8y6DyfcJFBzHHYjri7
mNF+EaybYlq4CYC8zOnVwvRYF/aZcU4zcnLnKjrSvJ/UUSOLOj+dMwWj7GDm1WrXIpcK0BJ9pDqd
CdbiAr28l4tzaKyXYT1VbofH7cSwN+80kuqjnXFldjTWDhr7WVVPCl09zs9Nm6PvCwhR0hcg8z5R
8Im6XkDiwzo+TnW55guSODQaA1D4VmuYXt8Jp/TWOEM7AIc8+txuImFkuQ3J/V8O57/a4M3ouGsw
oPIcSZfRAljpRxwlEhcmnMQ78toFZxodj7woKB5JGVASyrSnoytZ9drDScUD9watfXRfoeZxFAdD
9T0l/fqtX6XoZIGeAnie4ZBfkHhfItIYgFbXNXyup6uQz4aqp0qogsXnbGFwp0mD3N9suZm0W7tM
dk0wDUxrIERVpXwQ+1mjDQx1nlxtQyEHu8YR4Q3D8b74tqoPgQFdhbXg0HdiIPfFfbfzeGGR0MLD
H+MMz/imKvEpOBrJVi4/d65a1Bfe1BPa90Om2kRIuNu0MtzoAFYhhfSM7nmkSgR2tjt0bhQBV3K2
kWTuH1AUi7KFmhcOEPJRqst/yd1bHBgDRFVY177yhtdi9I5BQCufI8A28AN0rzUj/NXfF9nETVkS
C9CMKTaK2Fcky5MoIpf42xMVPsNtjCw9AwOcadIODZvb1Wz4f8hHOCQB6u2l0VfrsV0SU3Wx5dAv
IxtzjQfBm29KHNKlGoXFVYLaJvCGiySS35XgB5DlUdgBiUaN1I+dggsMgPnxsurgxQC7jHMQu7LO
H3YoK39wSDqVBQ9hqpUz32RqGfgkftn6z/hAz0ElHo/7a0sqYoe7M6ofNFenRt2DMOMeDL3zfC6U
8WVAx+hSfe2cUibPqViUmzSP31Ww5BF9gShDBWRJA5Uim+IzZdC4If+3dU6P/WS3NtS7v3w2XMCb
OP1CHx0fuDPGe67BKqVwFeJ2ZcW+BlKreND8I8OgB2x6H26alTr+EaeXMjXICe4dSSTWGqLxuGO+
7ITxTqhvecOMT6YRHR5J3GHMSZjV8jH6zKDhngoZfeF1EzOzB2Siwuvp3t5Cbaz1gyas/NXhdvWU
6oUG2sTPr4MPnoklp7YodSMZUDRQs9J1QTHAQaym9Cr1SqYf1gHp8RisMfwNgyQUPR5qg3F3ThLc
yEMqykMe4qC61lNOLOzxOwDYh+qrdq2b0pQ8hlNzn3XTDQh+PyarRwqdMeCIRuOgyiNYKlc9tcC4
gMFrIfQyzcmnX91OGaSqoX/v5UNuzTpiTZNPDZ7Zm+4tUwEeNKttLY2cKoqVbU98EBAjAuC10MNk
/nUXFT6D2RpiRlqbTFtG6OpShM3p1dBN9yRLyQfDiiaxeLCN5OS6Q21xYMELlGujYtHgoi1dXSlc
H0csUsJ4s1HSyJQSQtzqpdPVTden1HKPKaeZSHuCEIgQ/ZXR1T6Re5Ujq46EwReByl1xRWJB0P8e
mVzpZ5VS8I6r1OWbSl8NnfiXhR3fKsHeFOsQBtS/MOKTHcIjskp7+u+/jadhF96dALWEguQ471E9
knXIuQ8ZVZVWLQRtcGjL1cFOSzfe1Z10HGoGxHsG/Eprp+eiUqZjxK8T+gFigsTjYdTZkdM/uS42
yQ02Sw7wzSasu0v3EmkLcCTLSjIlGeqeQDew6rH8xu1gKi6UU2xxcPxn4lQUAVEZDqbfZu9POoMI
1Uno38+3MEr3NjMmWpuyMoFFrffNB+5HDvfEgQmdENVLih0tG/ixp+6JqQOIe/wYWzJ6T3oZahoa
TRqeiYQOsEwZ8I2YigD2YdMQO6mqK+XTGclgOvUia+KGNZgoUY+cFQMUX4tNZXoZ3A8+FTD8O14V
1oSx4Om5zGheg24z//BV/XVmhTSnCvcVDO12cZdJZa9gxlTlS8g9MLUkKilwdPDw4IOnQWo2FxN/
ZczKAP6Ov4vyO+GB4s003le6rE7w3+ElE8WRwr2MoY551lFc1dZ637KYGiYAMroriXL9IHpU+hhk
+wo5JxXWM4oNQsc2fCAWk9+uHlnel3ySqf8sX3ZKgURZBUDO2WDL2VNBxMsG42+j9dQvQPKDtlAj
Et9WpbkZTqrFUR/ZNenuLB3fgxEJVDjGI2n2bFhgKRGrEUihDuNMmBt7ccIFrjSVA4s/RbfvHDiG
cQD1tzRYHej1Yv0itzLoEoMK2AIyoy0r+IwxlqQOsQIjY0XDj8rWnn8eM4Vg4QAjN0lfxxZtzLvy
0a6hIPSHqEBxvAodQ6i08zpYqrkuCUsqrsQyjeOrfYPFM76oCHfnUlFo6ImmXyEp7yeMqCYOwZ92
cNIFhaWwE799NovSh7iJv9JfDRetG5KAz9LLz6hGRiiZmsjU+OffPuMkgm/LHissry6aL613yMAG
6GOYOCl4iYDmweItmg+/tHXlzl0mQVnreDiE5AW1Nz92+SyEOh92nzrzNTc5PgeFTgIEot/F7+ue
upcFQwEfXQqoQF/zC8jR7cY5/JCIW2zC/kR1bhNNLEagfBC7d09YrphGpSMxNYXBUnHZ4IuPFU17
p5+EwlDbIVXoZoyHVQPF3gIwG+7EN/UcJLW/Ff83fp7UncXn4/0hLC47mWOG41UZTshj2C1UhK7d
ds017hOx3E/gtnaj8drnZfFzPeb3gv+I51JB5SBWHSR9Ig7QNvKyKLc6RF3C3nXl33bXAtbgl3fZ
FG9RIW06cdrwuwJUeiYcivgLKp5wYITAQtUY5WwhHfXF+6psm+9FZkjbANwkplucTqouR02F00HF
J7bLENndrDcOL3I12LWTMad4ZLmYw9nsyIb0iG3wsG1752wsKPVzUQlnDT6cksX7rDkPH4kYYyWH
2/HXLHWL7GvMs5PQJ6yoULsjrEu4SbjDJVdVQYui8S1pd0yh9enLoMf9009CV71KXR5dIGHNIzz6
JtmBBWGmG7qS1BJAJHmSzsVFJbUlwuwzotpVh7V4I3ob8x93/1mb5Z/PoLBuVZT1Ch5HByU+cYII
573lW690fsZym+qnlOkEX8OjDAcBo9C6mb1C5W8XFtx+SE0FKlll+OH5lt63gQNyOlXz03fxeo0L
gI1PorGWt7RN8+2JXmJXSo2XRJ4cts7UV1pL4mrwFXiwC1oOoX3qMHccSO5QOJgtv6hcKxOTiAMQ
PCjDnULZv6X+8k/qj9GHQnYxJRmI/HXRmvp9AVrhVwF4gpYD60pOnQKAz3KLSPy0/TzPGb1PJsY3
+24WcJlraLUvyQ1J+Ys/2jmxyKjpB8/cCVN/2KUcVbajLqrzAqcumnCIkfRA4vcEkhSWCzoVCpIk
Sezya9UHO2B0LzFE+Rchilr88VUWg+Qfm1jJ45F+HB6Te1PDiR3Ad2dPuJ+dcN6grIgtHuakNPVA
bmFdGwTN6RV1LmE5nXSO4BxSezby21OalHo16Qd00yWOJoy3rnWmiDdlDhZ5wJ/JoK+YtfjshhQr
JLaDhyKy3OHn3OBXRV6DvBO/srAmTewcn6FFPJj8a2FiR0+RjE+0simqfv+kFcjb4t45TpydHkA9
3tpV/dRD3OCJkzhmzU4c0gf11Aptl753UjD8MWEdRn/AiY1z34U/YaoJf9Jy0GSIwngSZcLlCROg
2qIwgIApft141SDkvSX2FzqjUZMBLaclO+T2H2X/iwXFq8b8K4+CZQ7DxJN1A1OyPu6SsIc/ZXHr
qqw0D5+/iZRmHVP1AKhhlOS5dQP77LRlSUoTLmeLy9UoOuQIlwvlfQArWZbjHtDxctc06P9Pfeho
NExaE7iYO1G2Lm7P8/W5BD44AM7NR20efrgXST4W/MTkvwWlE0p3Bo712yi66KOA1gtzGOa/K825
8tZdfArovo+UbiZiLAmxZbxhBLJhOs37aOjCiV3gDYRLJSPLngjPBR0Gto0cNqvovLgfrfygRtB8
QbT4b3Ln4/f/+RaySZKqNw56dWQidbKbY+84WfjttyAJ+Lw02MkWld1hk8cTVU8+cBuI5TyKIxn9
Z8JrNJ6NN4mgh5VQw5OVno41IxRHDQZN0tkmC11HoRM0I7DVyRUR4wtOISzPavBN7hWOUpeOqelQ
OclAD/L+bbaQcntwErf28CGzNK+c693ebonfByFUDql4D3lF9GJ0NMRRmvHOuhlu7gqfhBwTkjD8
CuMxEWT1vJgv2FCqSWnS8dpJK89ifiMEe7ls0iT/U5t1VhNdkNUgpTq7Emh7pN+JMviRHT3DyWZW
ZyEhscjsLHa0VQqsY1K1Is6ZHYHQz6p9+czebY9TingpMOa6sXS+d8Zy0FPURJtlz7XdIwfDfpS3
GIgmqAiVh5k7lSYejiAJRzhYtVuOU2lrBzf9s8nFynWRovWOfMKIvVHqUYt+HaDnkKu9X/GBP60t
w1g0ynysz/lWU2QcFCCjCL3UW8PnJDv57uFze7we4fAOGtG7wnQvgaEAvAiDAxh0cJhYU5M4BsqC
7qOHbYONAX+c6PwJ/pINILHux0msZaZQe/MTG/rZVMIKoibV/kue2xIK4wY+xcr/YpgRhpUYYzH8
tm8V4j3QDydfW+78/N7jq6EWM4Wt5M8Oky4UUJltlA3ehGtRWlpqYE6aT5e0/HFdGkYVcY2Lt28S
Q12Q/UaleHqGjjiH4pn/aMHsGohppvANuUtrGVj4TEs/G2O0REwIaTnCypOOGlbmHilDDHBA+QzI
qPUN767HnXm4V0Cgd9b6ICLfgUc702+XBmJFKxKdMYw+NYiCZyrIOberPSaxdGe7jFdasZohllXX
tOkXALuI/nehkFIiWokGjZ110WeG4L+thLC9MUcFGTuVqjzpf8bJeVFApfj52Il3c20L1pDpI/Hj
l1t8sArCjoproauIsRSY6J8oqH29IJygmOQoAOPENJPwEcTQiKOKNoLN2pqvfThaZQT70kemhgZY
wo2YKiIrwIEl9WVIlnXmOnA7wtRlXsa4XuYA2Do7ZnDhyeXRkphDHwfPhIcQUC9pvLjitBNeOuWG
FYFf0JV5+6Ced5e/pg3U27y0pwQUK5CNhKh5QQ7jcjTQoGC9CE1JXfVtSg34+mI1joNOc7JoKgNm
Or/s3Av/W6CP4Oq1D7dTNGKoyFpothGUCAPuDV0pTbY0WGXaerMmNprmXhX2c25HtCvyCwotW0DR
njodqq+ftupCSCfZf1NOc+IldF67xRKesItWcgW5LPjs0wXOMxFE1AzdUmOWW3ZHGzj9ug87svx7
4Gik55jitfKetUi80nBQW9ae4mKqUSoypHqVg4aBbOPCOzAak4HZzK2jN9Lu1Y2tJwDG5UTU2kxS
of/Iej9c6yjlsGiI9o+i+3prKFX5fL1sY+H72Ri7AkqUP0tePYQqVkyvNV6oS9JBKPebaGVs4PMF
sI8BrlLMNnBCpGuTPhZsxR9f68r0go0TeVRA9hHMYG3j1imBUyXlc6DbVo5rfn+UrHlTqXGCmEiM
YMZY1MvvRVqOSL4dCEfbx1ICBIljeqFZfws2Et+JpfgFaAEfS1NRCsYMIRWRf5iFuJyoZD6JuvSG
Dxshnpberumy1fSsi3SIoYUBrRCdBUtlsvPE6WIM3iLFzL10CWhihmCAzmMt+agjtsCkZM5WSe9w
ewVvv9hgp9O9dxt2D5Vhcf/WnphK9Y3ukDmd2ZKbe1I0T9zXvCydBoXbfFGV13qsd8ImpGoO22yZ
P96+3kALMgrKlknn31uZZCyuL9ca/fKy7r9YWLOxOqgYvYm17GpN7WdsQOk7sBFXIG2nFM68HE2t
ViVusQusRt3zpkhw6uoMm/06OrL/eOrFQKG6asjFwuxgWBZMQESBlzki/PKbbXhbwSzf2zULnqYQ
2QzBGOYS3n710NWn5TcV8OFmm+aKt9BQqeCpbhyBG35RcKFAwRmeStMrXfGGuq8k91Qr0sf2aryX
T5BqN8kvQFbg8vWSQtAn+OvEVBHz9eOa85rETgD5+NQtZL3Km0lbYg26cc7gJV1wuYPFaHnWVAa9
AgcKEdfbqv4/5JzTyALIeqbz9wWiP2t9f8wY/W5QqTjGYNNvsL3vHoa9fPhrrBrchnMCQdlGezXU
Kki5r5pBC3GOp93zsOln3S3c0ycVWM7sn2H8c8otqwteGYc1n+vgeYU3S/WGBRmXZEfzXHFC+YLv
Q7lv3VXKHR2ZedUOv7/fCfcfbufO9tjSN3HtzPBqrF0j2yJRGCHrse8dDvI28yZnOLRO30aZKOMC
GVfRP32PEBpcfD04dQ4hn7hpjMNeRwQh7zQAkncICqzPgSth2zDxZ38WDlIWWlFIIJC/z6Ytipeq
hs0COA3lJu2ascBJTWEs86DmezQ1ph8+/PF6jUAHN2s1i7p09KXAPg7pOwtpAoBFfbghZQJ8SQej
AM46IrnJuN1H0/WYzVMeOJrhhkpjkgzR7j+XQt/FO77lwufWlejeRf0iR6/gUFf1/AkeKT3XzMSU
mN/ZpJYatCfEvEzhW0EoaOxhA60GH6h2If3WT35Ta6TuK8+lGZAJEFgUZfrv3wqwZOT/1ZYqW049
mkfzubdbBxtoCbqL2p9VxiN+p2GmnPsgfu9JnB6mMp6/Yx4wTBbqMeurR3Evl8G2BgRxxP6UVyXs
mb6ZP4QkEDYfornjThjSRz8lMdmw6jTIuEJl59IZYQMJ2NREThu8IbXMI55B1/MyN1twFFQTRcLC
F9uTC8HnC9btMx4IKdFzZmyW0CNBMj0KuzYcEYbT6/Tl4LeVdy8e4CAYlZthhUobrfrihb+6NVUl
Kq7Kkbn80/TAFkG/vowtQypmq6ojs4cf1zJZAhJ9iwKg4yw3rRlxNJB0/BR9pdWXj8ZQtxaSLouk
TmgzKnkaB6LEXetRVqRhqsfBjVCS3r5PoSvSgpXIZ0t4RRJF+9alkD8fodp160myvzxLPTdaRGNm
vatHtMc8stm8SrzMSI8EBcatPiJKq9I6STGy2R+r0AdoGL8gau+fr5/c0zWd/JU9DyI6O9+5CoqQ
JL3fgq8vmWnFOqkLPaA7MsHsLWXmFdEya2m4G+BPUxBiOx+1rOwJQ1+WzadNUUw3ttK4X0/hPUdX
6prkRyHhBwPPXdsVJda7hMGkgMBrYOw5vwP0sphrtFbE4duqTpQxm2AsfqpQDFeMFQB449z1jkAT
ULM6+Hfp9RHnj/1E9bdR1lBCnzQnsSwMN1MLgrFWIunUtB4DoBV2T4WXsot1rAdaoEkp+X0sgMBM
0qhUvq+poQUXjFq8AzurNGm6izXCT5HlhNpQYvdDvY0cZ7JSTRFFi3OkcT+nYMExj+h4NZcdlADh
BnA9V6q+Yr8h57TxN9q2yR2B/AOR/0A5QuY13vXnMv3ZyJU0NtB4NjAPL1nT0vVQwmwlW3kEO60O
Taemxjp8sGFq+hKS129ep3NEeneayH+VHAM6h9XNwWipIAyD5jmxtzEbk1t8trySAKV4g0jnqTJl
cw9qpXMg/yfsnnYIbk0eUx2FwG5Auc6qTeiyyuzkAEwp004Zn3bp0awvun/YSwkPPL72IE+7Efwk
3yuKKQ8dDBWNhvirugHvOMD8owrokcixtR5DKoyiF8t7qHvIMExG2M088bFfQ9YUUH97Csi6QJPq
f9Zzw7H8sQP7Y2UqPg/Gc9fO3Z2WEKpIe2u8OOHIcuKJPINfr8dQ75tI+vydX8Upq2jaHVBw/UKI
+s9U1yHXJQxHLNEMVScpBedO4m9nWgwXxiGSU9e//Bj0BzhU8pi/WYWyDPXMoYG5+DwMAVG9ujSz
5gALoVHTx62oXDOB9vaV0WdBIh0TiZUcpJNw5/aq6oBeq5EdJXQm5OAbH5ynSYX5IVsX1PDIyCki
Fcj+i/KzBY/AcfLK736UPwhEx2e5hjwLk13a31FryltAfZTYci4cTC6LQJrDJCfpUmBCpRsfU0fg
HpJJF4AHLC1Eq0gQVzftviCjnKYuXvAfnOBTMhpDLNu65iyPYSruz2onxJQs2KIWomY9nab2z0dZ
wlQ1WOeWFiMYUWJX9a++IVxluojr0wANXjKNXfx7pqj5wT90BzqWvpWHlh6hhU8UMejSwWbcLQZd
X47ZexAzLZXGQlr/XDPE41qUNg8Ny1T25B3OZL66SC8PjuvBLq9+OsmxMf2iMVk0OC2rkRnc70OK
ajO7yuP0LSAe+x3t507AaNSxTVGYCUDiUSm1uK/y9WCc3gnMCHUFSv/q5qsu08nlejciMNl616XS
eYt/tXdleJKlJiyUCrn0cyOcer1IDRUGdY57QDxYhVPMP7wI4fhhmUL27QEW/3brhukD4NraMsdF
2iwWmw8PPRWeusGBvDlhS5ynTKw9+yzko4EIF79dc3LTp0H63F178RVgOoABAMBKgPD4OjiXhA5Q
CODHbbCqWlRqzZX9Gjwp2PlxUUPu+MyCbl69Guqa68ZKFAwlYbEMpp6ZuF6vLakS8wCxta2/4zdk
LbsDxS8uwhfBxSSBlik++RoZr7mg6ZBcqT5mftN/o9zdUsdXo5490ERnm09lHSh6EBIq45yGXLFw
dcHb2Mf/Pwr+iZ1qAgdkyg5O8qK+hXUHhWbF3sF4LZymkbHADuxXLEVFo0y1K71ePF3TAYvU98+f
D2TuSafzMg5P5IwLPeml77FwncvMnYVi7M63ynvDfJ6qAAnHcNpa6igljWFeXRv6UR6dBSWPcvUZ
sy7/Vcxq+7RJcfnlVQnIyM1Lbac7X/13d5B39QuJvdCLjjBiCk98d9QNgfQ0kGlzaycPVw+U8vuN
ncLR6VhnMgj16PArSW5UBW53GXpEirS6Vtxt0olZfjq3BTQ/g1Qay9ANAagXO/eTIxO5X3N8vRdU
6oXkZBoM1SAr145gwdxgq0/JopLI5cPKj4gRd2Lx/cV0BMBzmxJJ0XHa8Ds5vEIAryRly1QFnt0y
DO5kkjAw/J2by60zevDybCQv94qiW27Qv4PBlVCvgO0QWYwJ+RLmT9W+iyOZchKT4qhVjz4dTkh2
StWt76tvObBAqL9VL+x6lXZgocXJOZmaa/OXOrTTQXB0HkS2mO0BdJfjLxuiOc8+POMbCM1/3g9j
z0DsSdxgU06lnBLCvQwfWctcgrD2g+dtpdW3hEE5tmiNyCo0cADpEYaPenaocXqxVVc49f/d0ACT
34viqLzkF4B8RXIDvSlSuGa3Sw8HSYmnmcJejYRAhi09yv8CTE7METDrHYAEAZsA1Etkz5hXsz33
Tjs2BESFiU74D4p4yY4u6q5G+gqAZXbQJQPZ74EisUGt/rkqrAIXggaQKGgIeUxK6qhefeTvQKpR
V1ogko4qOeho26e341wF8yp+X8dd0jmO+WayCpymIMQ2xxcntHymQYNyUQLMJlX3rwdTQwuhob6v
l3tw17jDyqkxgXq5F7oJbcN+hogxMmyaulEmyBNjIAypqi1otVoQQO8fq7prIoMlFRrI+YhJXJCT
0SQTf65bjndhPoSYovXYirsyMDPlhKdcCvmGk3FbORUobCYnZd1+Xs/rfop+mYTk4I5OyJdTtazH
xqsv7ihGWyAP70+a4cSR2McKaj02EMkjclDz1iQcVQSo0z4PiFdzKNWqpi48slw4G7HevjnYzBpY
JTc/MO5rEH1ZmNB3Nc8Yhv4swYffTsIrxnhrU3bNLtYAN41z2ujXnefGCqJjoEZqD+g1iBBD6adY
pQJ62lYf7/xgNtgYAuytGXPYFGq/A3+wZBnv7sUzUrCZFontaGPPo5o19MOpTrRCsH5M7Qo7B7Sm
VgjuP8CQoHETHAunuOSGzdFpjVH9yBVjmJLB7E1nbXfcfoxxgvIDhRYmDSuz7rGaj4YItIv7LC9m
H3FZsOKlD18L0FPbNtHnG19tU8ntQ9guthzlh8cHYBV0FSq/xSy49Pqr9T9hQHdTOZUZxOg/wMz5
1fhg0eVENiGXvf2fh9zgybjlnocSjwaihg0/xp62lWWiswhh+tVIys6uFowyXy5TYPZLCxcusI7s
3J4au5t4WkdAYsuHdxYGQM/9xe5BWzB7eTamXdNkBW+cMPgc1sTqtLZ8ZdmZzfrMUJI6SEtNvx+w
qgCKZtq42ix53nbCqWztQtSU/xRyEmQ7dQpTyUerLBd/5nYPs3KQGAd03/X6+5ylGv5gh3lETGm1
ge/1uUs0mRPwv4x0R6bXBeuls66MXRe18UUpbxt2Ku1ltaMpCj62qmiRsZ55a51WsFzhcn5NfXQ5
ErXETy7B6504NY4VCIGdmtGsLX6+rXrk8oIuFg358CaxYAiyrFx9z51opnLVesGEN0kGxuCBb5kY
fIiqv7wqs3m0q29GGzwOVAlRZZ2aVOdzjmz2YkLdnOAmX+tGoeQ5/Od52jz7O0CTWwKNLirAdll4
i4zOljgh568H52FfRkvIeFKeYsW/Dwl5bVTf4P3TGLdCzP0m3P3MWwVuX3UW2Fy9TrvMZg9r/J7p
ZpdFTYi2iaFJYjY8s/bKm2alQKAoo5HNAMomvYZJgUe1Nznqr1yEzk4ebupW4XoGhrkekU9t66fC
sUeA8H81Zmb+l1brTiqoYXlZ3i3YnAKauIAUAgZnT56pL/qkxPvTlJK66qOZFHX0OQuCAQFQnUCk
XDTfG6yDfjO/r6etMY4suL9eAMAWjjB5i3LEFf8c4zy1o3aMFnijmuYKM0L6Azm9EoUBCq+OhMcM
ctAJB4VNwgBy17SyUo/V+c5CZ9XTokcq/rFS58Go7t/4RnPj9pv/zCKCqMID9NPAihE/KNMpCxaR
C4EbFgK/lh36s/UaLegkO+xQR+DPkso3IWTCcd0SgceInbx0QdlusuiEg77VFeibcgQvVDjGjlG4
2eZv3gv1bSfTaoioSoHhxzW8qJrF5o5Zgn+zNOKW9rJiBWWisoj21eEjzZ/ny+4ABDcu2jbS6owg
Sqo6y+bHr0++YPM14PkcHi3h0nESvdn6kQfP0rQFDVZDTFS9m4kf19dpJFWLIcDXplrcvsqoL7pt
mhTuiSPvZSMO+q3G1wex957YCCbaBhif91zBR3Em4pbEL805W2xOF2pzn9HevwDsSh8cyvkoCQFf
GiTARh+oeAy4AXWwYkKqZA4TtTgPcKNBuSriWhEGr15kcanIoeRzkEa0PJEDtmswXtaE/Xg3bIDt
RAhmDE6UkH9bhbCPRx4qwbBkY1vxxl79cDITe3GscK8b7meQghSgxsArdBbRI/K4CHhcz8Ti+ng1
rtqREhc8JsEDpvf2sE2zHkoJl9ZdiXtgQC/FXwjKqXGYaciTZuZSwZQ8EeVboE/dg398xUtYxuFb
sd+b/FWdg1Lto04tMUBxENcE+Dl339jkDxg6uWD3iHd37JyM0zybL/l1VUKkFyspj0PcIfqoVXRz
Tn600aEqSHRtP2ndNRclYvpo6McSotrwIjfjoGVMEboWVTZvBjd+Ov83OLC6RsZq3KshL1smBeas
LKe0zmGpstcZBd4oTXB2uVRG6AI/rQBDxZlBms97cdb7vbH6jXgrI66xQk7aADqMjMTHxFl7tL0U
2tR0UhUhuR+BNbWMTQzsOylnIlf3J3MXJAYGK8R9ZCqwbRjqsKZaDvrw261HY5uRSF3rdTFKrZm9
sUMhgeRQMNhePLzzScM0K2uZVgOjk590Zcu4H+rWTPEqI0SmGBUoUgg+54NGihcMZ/TUXsibEgY7
EHOjjA0cGXKYYbITgbEo6TXoqIeQWdA07jp8Gnj2/T+37HIkKzgyQhhCGz+5lNPnhbrSRbxm31KL
9JIJIAUfCTfS8nr8duu10JH+fErkCGidd9Yiqtw1BhchVg6lfR/rMENYRiPEqEB25CvcfPKUF/Ez
XSzEXKmKF2bE6wWYcKt5YtBzzcY0Nxk/Vxs665WTtQU67BVmwM4ZOVYq/gXB9lbn78YjNsU3dY80
6vsSdFgBuzs0b9/Tx6bodrG8Q80VepHbndGvZLC8IAHxhcTf21f+C67i6u4vSsqHfTIGFsKK05Ua
jqDof/PHbxcdfqHe1/lWTEu+j1IC8X2bdWC+7HRuiJEBc58eyQCJab18b+/zWXTaadIX+VMg4b3g
jqZmIxxVB06cEYCUwM12n0ui5F0NL3YjSndCkdLO7OHvlHHOiaEY4mJdMUMHnOlmnrahjsZ/vd+D
H0TxIeAeOXYdbETFlhLhgIVw7iA19ikO/ERRmBi4plroF4ae+wVREkEfM1NDTX+4Rxg/oJG9RZ3B
u3Nj/55JWov/nHBkyl6g/i2fsbRRtif1WzyyB66RlhwlUSxq1Fj2iw/ToUESL5QS6N6HzrbBzt8I
AJP0wrWoTIkHBgTKH1sz/HS1PtMYVDGFT9jriDaYaXBxwoO2BLDzqPYdrgzIgTOShE4lrrAWNeA3
FEaTHji2BwohJN5C7thxe/YigmHgEXptpZ9X6lnJQIqC5tOoikxZLZuwPbChUJVmGLLQF+DFdZXx
uTBCab4i2Q8bwfVy4RqPssaoUbPSExxsILOQDKPpFeB+Wi53KllAkvEbjFDa706x5dupkQqwOpKH
t284euD+9ksdVvYq+uS1rLYs4W/c3/9nU5WaEUIoOC3A5kT1uuhwEx9wpuJy2jH/ewvEfDw5io0Y
WCloppJIuMFjDmhI7ih/Zgwbx+b/qIbsRJbhaQx7E8TDmScotbJgokY59iDDa14d4zfftetm5HFZ
HbSNQs85N9OVEmhv2sS3aP9qcz8bdfYuuG4IaBzZa/yurECKf+IAlGtwSt+8uw0HTU+g36Z6eLjE
cI2qyRFl+qpf4MCM94OBAgzOU/or5rZXlSwzsu03+TAQawItKSdDErbzN6DMTDujq66KQOOdGr/T
HDxirRLy2UTd/5it7TmGmqiqedKFkDsKfBSucZFyEAdmR0yiNvTJSha7HzFz7EQ0wItocECp6ybc
IoEVmua8m0nqDqtj/gvsTfCcvpnkfpzAzc21VgFsX12f2jEAJnRrlyOxUBFO/yj+oPPCHXAypwp0
Tq0jK12Nb9OYJWYPGCAZqStWnrfAU9JzXae8Uq/68D9mGRuckLUnmaqCxa4a+TeKPB7+WVmxTQDi
lgFITefxQA6ofOhlpKzN11IKZ6rchG0N0tR8fVvay0w4th6y/4EA0SqRg8pwmQL+jcKDI6Qmtud8
ZdZIyfHyZijR0S86XFnUGvNHftyJGW9A781WUIu68almFN6TSIY770DFgju06C5p1Zm2oIJ8571X
WodBWs1+wQ4nyc8K4c0CaTkn4rXiZqEuOvkSRQCZ0JlUJHs8gmMZFrTrhEm+/JxJiDJl1StjkHm6
GRa7pe0JDHNNrex5mqnWpAEQz8/qUYgc/2bATRdAAZWlpr60XzAjlS6vFaFOge20O68Eie4HtAgA
AoLMurL1xIxUhLxEvYXWkYb7bRBiaFyzQp9MkckkomIKdwkJBA6e4+IY9GsVshameto6ahF+D3wJ
QxZdod9aEnmH2tgtY2/lVgnw1bOCTaJddVPCVWGjQNJ67ka79DMRbrr+pCEfBlu7PBEgEgRqcc7+
8xStURgWZHPWj9GQLBaHdPM4iE0//r8IUV9NQSTWsKRP/luuICoNXhUgiW6ofO9mV7X3um5QGseT
hMozKa3fmkKUsARP402Bbhn+fry3vSwcmubwj2vvfR5yc18ok+veSG/wxTcvuCCIljpefIPTwZel
o2VOCuyU/A+s4vCfCxd+OxGp3hl3u3/uiRmgvhJkhQkrPGAwar9BytiJDEVKU0QwiIAfCdrKaMra
OUKSmu7C93FEc2EUOkC4NWVudKFVah6yqb1eUhC608NoFxqCex6jyQctVWy8CWuSj1AregovgqLC
9WTy8z5CPr6YybKoJ9PMV+zADM9fFxD5ET7yumcnP43Tz3BxffAPUbs6ziScbKSvwpdw9X3HKvcY
PFKxT9qTQRkN1xnlHr5ddPNyjA+n1wx+Zi6DINmTOgj7mmWjiYPxzqy6NWiy6bzbyIMK7FQHrAIs
6ejIM3lhoNa8bG4Z5g/EzbGheXHGFJGKn+wZrYsxFk9JriBQ2Qw52zbtMfbdVs/cfL8AK2mlddcx
fdRhgLc/2EfgeDqjIAaFh8dCULcDSvMM+O/IOCeavob+TzkrSI97yMyw/25PKudkJ6STDmqMGTPt
fihvb1nG16zaqIXpKUxhfeZn69lRu4TaC2Cw+C+uAonRDJUKvXMioNPkaPeQ66Q5iH5EZA7vLbMv
X9Vwi0CuJ60d82M5rk+Yl0LOsYSf1NRa8IMBuTolTCkrndnJVT1GEkYu8872hPaEpG2Bnf8ZuXtX
3Sd52ouqD+3JbcTvb9KEJFT2CHk+A6Vy7k3RXr7qMwFdcutRtTaL9TXSGXWorEqZMiqJou2he8tV
p70SYXk05Ew0f2rykjU+WdjnbyMFKrfHAAJVb68Og5SHD0cXoC+sYCoYBqdWtoG3/9m9eQPkOnML
oMRXBK6qQJxhJ2EkcdcH336pvdOhRddRyFNguq1oNkOlepc7lHOqK66DrdC+a7nKSn0EKLbVSzVX
9xCWc/yVIJaR4pTYNCELbFZceKFqWSH+ebtVFKufS8vkcoiypAV8WBwEFV969idB6TLiRL+WYVWa
8TnaNovnT5ppAHA6uTvR1Pde5PjNv1yPqWRU5mLxNXe0/6DICvv5NQUodRGe6+WfXrFx2xfFPw87
gBKT3s9ieEsu9e/UuEE1e0z3u5iEMKf/zm5XMdfrnV7piApZ1RHooZW7nABTqCOfJIQI+QsEfFfn
HmTX7bRPkER5dp60KkrBjSKvCZa2vcx504oakLt3tRFDBhyRSl7v+FCuSrYpwOso3qtdh/YvAsoT
QxZMdZLHk+ObY9vEOBCw3x/M3YJiI7+IztqPFGTOQzp+HEch0x/C2FswYGfVdrY6MadJy4zr5TxA
QnS3vVhSdo121+OiDbUDycBqdX4tYEPJoun9cemmEqvtwEXPeLu1mKActJQamdRvgniI5LFiA1Nc
E0k6efdwshaXWyZPaXorZi0e0NGD/NzeS62aBnVxhODb804jBjij3aSbeZhE1ILKGJ+tUheDRKSC
olm6jAGQ4yQZ61UFvIIm3wLjugyqotjCMNA08b40F8I/OjZl7/D2J8d26YzT1Kh/9NvLOTOCnHj/
Tq0gcL5OxpIqoxdOcTBrs3KW5jhaWw3tMAAz5qcGCKN7QdQvTgBR73BXQwBVMlo0giNJq8zDuB1C
kh9uzTbkud3EsVHvvx9L9hCzLT83D6wNtoCbkheKZ3zFGvu2yPfLJntZgV3+mFuFjr2vPOqGfVUv
uUfYpWTfhz2k74RFbRPZyUP0YXw6vo1KugNsy7uAmtiwOopa4JBjBWlh7DPMxaJSei67jfiomfRf
L+P0zH8Z6K74jLFunMY27dKfXPKlnGJ16FxswNZUtAYv+Hjf44AcxqR/8DvJHZyM2qT4/TLLXn7q
+X8u9j5rs5hnsttwHQ+O3uyuo+0TvLcNal06a0545ZJR4tdqisaLtXzXDT27c0QZ/kyPnZnml7ld
03P6vwZ+e3SrYqREjl46cw3wY6JM89mDXSDQcFK2Jd9jghTgsDgyPWqesf887KTsM3Skdbn7gS5T
/uzKV4LZ7aiOL1t20Ww7lyK6jcaa5PZLyulAwoUvQi0HTpNBB/FqR5aZUXn5qkFYaUrohsbS2zIq
H9Nm0rtMYvZXYYQvzUr9pG4gHeJXo9cjj4bv3lXhoH3Tx0TZkGYiimstBaqin6XA8vX5QLIXEVP3
ZcD0yyTPgopdUdM+/Nry1lfyMnr7iq8F0NHsxCfuwMCIRgUySyRnl8PaJpheRcQX9DVJQj7KOpSm
OQeaSGge85HoBuOmaT7KAFBPaqcbl/2FNQpHv74DApbzd8lZF0R+6ZFxqfdHIRM1JIbOb4ruCaPc
reqv1BEW8d4fobykLTmzopsIDGFeWR9BevIWLN2Lnl6CRdOBQcka0/hPz+5oZdXhLBZ9+gRuDQxb
qQTtqkdp63de38M7dW+Vs9nByjD1sQSxI38Q5pkmbshty1j6YavJ4WGWUHxgDx3nEyWFz/4BpFTd
IKWN2UkJd3Xv8AdUngo4Bg82esdUjZu1adKRCW81oruXa28X/y15EJKkLtjjoHPvSN+Iun0gvz4M
XpPRtwmW9NzeFNW8eCHg2RfhaHK3uS8eJnY089sLbkHkPR/6ibhOjowpb+ECpWa8YzMG7TBRu6wK
++8+RdRk6x/WGHeEbZclDstsHqAKYOO7aFSQQKPYxDbYFHHeRL/YXKPl7TzAwu2lAJwCplQU6rGg
oTJEnqnqtPl4FYUfkTaThFXGjZOsiH6NokscIJNpnC45jXH//PgWoNXpisdIS8+KXxN9I7BtFKpG
HSM0qcTuSy1IFaWYHUk+ZJ3p/TigoK3muFW/ZjT7zk4D4g96KurWmY2xDb+cs0PmrcmObMR/JVVE
xKHUpQzAOYvvPQSwRmx2DVg4WHJa4Kg6+rWHZ+YQUOEJP3+ejh0eROFngolwBSurnilzTyxL1F0/
U9KbfJMoOdVdD1R1uVwdpc5VCg5w2Z/fxrYq2RXT9zl+W2XhwYM68OyPdr5ktlvxGCWtQyyKh2NN
al5/TipJzcL4Se1GfF+eWviytAkutmP7jDnLHJwJj2NUdo8cNbYH1sK6sjSrBXpadjebHoOz4zuN
JHSiYhrS4JkU3zdZ8jY5fRmn0LRTdDZmuvL06uCSLN6glcZr5A4mvEwSXpn/Mk7dZVrrAFfoXamB
IeDr4Znq2ldBCieajx1jrqjBziM6P6DOHZg4T1Odgl3eh4ogZops5ZFpGtoXeAq059ySvvqOtOWj
jf1kOR6KIVDEDHEsYRrokTHHvqMiEkdoI0D4vGYf6jyLIIAuYTs2PGYCsHlRBmG210Smarrb3SmV
mGn2q6UHkdKOh8a2uGQnWVOaajmbKb2X5S9YK8tCfuf/qAs1A4DZl8R/LX2C/POJUJok4qit2axh
j8z39xbtx3ezHvFPOqlBuv7GLGJ1UyGgb59GiAymj0HCi+omNmwekRJ0qPf+3CnnAExOQpt4Rrtq
6MErS8pqQUU8GFrIB/RL7z/hTJkEFgIahk+5/xH6zAmK9et2/DPfrnaWTSA7mTPby1nYcXCJe8U8
rkzc4JiBRk/toU94oW/CByQI1jaHkMt+vTFvcUAIBMXlD+0xN3WTeEnkk6sCB1Gv/Q31wiNr42YW
iNYgXmyJVQwmjfZ1nCqNphD5UhF69XPjs9EH9kUcJmml1TTcX4FWMgR25zJJSWPynqr4c/4WxpPi
03mg/clLJMUBK2/vTKmH9BfBbddgB/Rg5zwG1Jj3r31aW9wzgC4FkqPOZzHo6yeIWFLCk59pfwI4
l2kl3/VmsqJuB2r6Lyh1QDxa2uRTPHNVu8r1HAYd8s2PbVh4dMksUhQ403wi3408emOamLmr4vKg
3cmaHlXY99oOayGA6KHJsC24R/GoTsce9TfG6no+f57aADmlFZl9ZhGUuk+95lOwouTCi9GRghfJ
3zRxh+lsCuePwWp7AOpRfGnIZ3xecxmQhYiSHJRpnCdzIgdMkuw1c3dGfheIZPq7rhXV05pv79aK
BlPLb8yuQXCWug5IoRctagqlpbgziD/t/+T+OfUWg2y6lO/8hOkmFuAeaEes1Lhi6u5kMKCft0Px
3Gyw/2Xo4JQMIFSA2fKWCikKLQLEgP0gl3rTFI6YoGcpkTiXlD3uwfEXRJFvzW8m+ZuZiIpZ+6np
gQxxrlZD+ZmhEs/CJ/k7WhczEzb4AZQYg66A8xHyx4D7Gd+YCwLBHvHoFC14Fb4Lxk4lu30FnJWl
q/usDbsBCxyvevl6GpWblsYDrkFI65HsCsGJqB6WEvmd9hdbpYB7tyy0YUsWp7hoYVXHX2CWbEx4
+HjiSN4mnaMY8JVHombHI84ZEIB11+ptN8m0caLJgsCNylNJNZBZteel/M1rJ25A1Hr8t5veX+gY
whgTihHhgOYTHsoppYz3znWAZuD3JeL5RBe291uS+pl0zlif3hfOnFGHuVMqdjvTMaY7QxipdIH4
LpzqhHgIu3AF7I4mkcZtM3M4RKCxq78e6WauoknBDGSVGEh6ep8Od5RCUbS+R1kPqHevpDDAmUBS
JahlTd2MxppGEWEJHSiBLHUrU+N4ExVg00akGbA0SsiqMwo2SBTl6kTo90yRiDRb1vHvF70kjiKo
NWZvZcn3QTMhhCHVdIXUMqQn86Wxc6jx2qYvgw36ps2xQhS3ekKXJpilTm6c6Zm/NarMmrB9G+K/
/zHcd2iJzXLpdImIy0N7A+CwnixWWLQc2vGMCYAfpZVo4osSpVOiCyCxfT34pM4Iz0felCgquxFk
ocyDcnsn2jLUGYkYwEX23Crik+Sb1e4Et5cmXiLBjmxCf5dzpUpXpSSAGpsyfejRlZ+jPRazQf73
Jp/XV6cldPwK/++GgnKxbHJx/wgOm18dW8mzEms4wXUFaVL55CS8JMPNCiLnXPjAdbGeosx+nwGl
o6C/NrbqSOVIkuvNKT3j6NUbytROiKotSz0DSkD0NAagGbNaWMEuJEwMvMtfiVCP5152JsoxRtYa
CGltQAhgxx78x5oOEuIrC8e1RFuxYk/jGE6HhQDSYcPJcLAivvcM3fiblp1pOKkKl3knBDLvq/C3
JVH8aZBGvaursTz/GIiVqnnNs09diKklXl/pKhtm5mvD/4z8l/nEwU6wImNOrL+4C9srunrt9BOP
66sV3oezjGnQHsFV12zanCFQ5zXaoYS54qnr7QhQhV678RKTFVO6gkt79yVLFwG5viHO7dgNbRfa
9eShPWCHn4ZwHvKu+iNZgKG+ohLVk0eGG3//up5p13akhkI9K9Lj7heYRJGO5OsqTPxfwPeoz5ln
2XmpzpwTfu/+LBlP8B+GUH5I9H2C6U6UPfuhDKel6MnMph4F+YpRQzhJdZVXz4/93+mA+ZCsa2bO
OlyXZTqW+Y+nFgp3RiBVUSPTxYu0ONXfnrCpowD96aCFZnxiBKYb1yYgUO6FF3t2D45S0g8um4TD
u9mcTzAE7out68J0pburEJrcJ4yCOTLLoWK3KwwQG0cIYEdSVteh8/x0QO6+cWGX/Ao1JfQcSSFY
2KfQGdaoE9CHS/zxo/7LEecuBi2a1wEu+zqhvpLTsF9XKv5wmHQIxqTutXxn0PoYHZUhFA+GNlxL
Aqdrl8Vx9z/swXOpm55rTRTmlfUOpDxl7BKucffhLHrG+vsUitexA0oL9Y/xetRn0FdFw4Rzrx7K
s/NDPrMKWezlUvT+elD5NOEZ0J4Ul7CkkrdohkwwZAlvT3T3HA9cS+NLTnB9e8J83hxM+YXDxZE5
NPrPyg1PCl9HS0EUQ0Af/x67alPHZLPbmjdA8VXPEjEEQb+YNPbUoE6A4UC6NjImA9X/FLdty6Bd
TLImwXhCwivx/JXNAPpUUi76EK0rThfNro8evj3VagFAyOMYCLCElJrkSZuC/EvNX0NMESb5h253
SxJGGsuo9KRMSnfOU0xQaFCFMydlcjKxOPnuVGYL2exi9b23HM/6VwOsMr8XaV+YqpzetV47T1Dh
G03E7vMrADdFg+6SxqU691XqGk+BSfCwMr19M+aMcuBdawNqN7D8viuU+FDFWId2NA20gKTvWyuv
f0GIpN/vzRy4CVVNUs9ybtY7v2iJMjWRxFdUabcg3r67wwgDbKp1kBaM8brTPPxsN/VcLhmd5AQD
ejNGw2IChEw7gdXhVbfTYMAzHX/nHRx2Z+keS0+wasmtYT/yNK1ltkqFOk4cLE2APrCjey4RnZn4
OC7FVkO5JXayENukN4FmCfxYY3P+bltFm1++0LuNm8iFOqqy+t/gxcnPnZKq4oFYAkf57jYJ5PNE
ClL3Y7ZKM/SluPHMbDyxbdpyVM5IHE9ewjy5+7ndBVLvAFSTkWdUpO/C3DqDvIJJXNSdOjr4XCaO
0Zh0gfkBfaAs4g0oSp1SgRde/fOBOSqKqfbQntWUKhcs20oBGViCGOE4AkbHxfdWtmFjudQQGBOr
EuQz9G8ILCOSz6ThPcG6v42zKxJ2cPcGS7j8RpuQ16yndltY1B81OOQp7STBGUMGVRZTJryL0fK9
HVywP4ft13X2jnIgbKahO9red3f3GwUKzD7cyEzzMD0rx6X4cMjsSwWB4HwbEQ9+yP4cuSLzLYNK
xfwXaZ3RVsBUYVVTgY+MeP4NtRUlvHa8Gw6p9uP5xuvy+esOd0eKblU4joa/V6VnHbusuW51rF3e
ai66nqspOm0ErH0xf2La1QQa0BFn0YyZPMQKbN/9WiwH0CnChV9KOLHYU7oT6kn2UPjG5DmiXPw2
9YvaEgnDux/s2j+2JBLTHv2IyIoNJNvlEkZ1PsRv3GAigFCWSlepha8LQk7CmLY82qLEC6N1B5Bc
GGHKCCVl/DUDTryqijv5OVt1E8fIthRioUFHhDpSAHA2DTWyAZrHsEQK9jkgNTvUMvCxKy3Y4oaq
Y3edfy2mB9tdq2f2PkUrTLu7o2nCL7W2GTnZrMC2uui41g2GHMPzovjshT0gOHMao1lKSrGI7sXa
uqYZa5P1JU7Xz/WdLG/rVSpkkwR4RqPAdUEIEhBdqxaqcvAOqlTd2Ar44asy7H2evPfZVBlmPG+A
GeuhFdAADgxk7z/pjCdL7GXZWU6vp5/VaX1RofLXYzTI5XSEmQmWVfPi/lJGfO44evZeOsFgCUp2
Y0ouVVvJ5x5TEWPx53vL9AHP+4NPkLwA0eShry7NHw9eiD1eU0NWwWUpw5C0zUvBFjJubD5dRV3v
mZdOI/PjJZUMp4UgFE8trOESxVVgFD+FNqhvqVpUSU50SMWIV+hptB2pOwhh4q0SyU5gNaSMObjU
f2PCTwT9UHWlGuUQm+M5tQG64uJ1wzL+iDKHBAgWEZSQHTUqbYny68VDm+IfL1ROrd5uNdGCQrhc
O08GDur4g05w3AzSj+x7efgSrpC0AthM+d0LnLRlLEl4OZAsRZhpf/2ELoDDYUD7XKsIgus9zpD7
jF1yXdbX2xbhiYpJKGYeVAdvyCLkGwBjU35VURUfUp3PndYZp44eREwtTdTBoRPpore4VvoYEZFA
2MaHzVLrNfgrt/2dY8QKMmWIZNwFl6N+Lwh463gRy82ZnaDEdb+VFBB5/BtHsamI1ZbbHX0xr705
NQH5QsHJ2ND3OcCCEwqlEzv49UKKvRSUwy/YZD57PXBP+jwnCw3+Y4IX95M3PpqjKaJoIusAecjI
EXGzg7E+uvtO1jtCJtxJHdw1zTboIj4w0LExVJYCOL41mrJZ3A3BJODnFgoUb7apEDKIBxdVQafP
dZqrlylYWkP9iXN3XydGTOIZ5MU9jX1vn31En0rIBh55yVnk/hMtMvktfJJxechYMbwoSLsxqQQf
T2PSNMhue+GIQocfERC3oZxL6qxDzvOhNXPpyFMJR9v6DKfzb/yzry2psBJE1BWOupoNLbBhg0A5
u3jCfYLO/zSayYpBk69lrbG6sGD7Dzbq/Wf5tc5TTNtBdpERh7/g4+UVfNEyv3ry/arzuAJbQhFi
EmYWVVcPy+0ba32cLiCwfhih93e6CYMGo28NXlVXEobM1AmF7sf/dHnB7SCLxP40swSyyaFCMLyk
oqIm30v8SK/m7hkzLzrNqc4ojHkXDh6Zo9ibIdT8jWptmjbVdrTqskXjFrIssMPVDI75ToqFofqn
pcqDy0z630SkzLF7p9Yx7Fv+U0svtKL4AuyDaFcjHFeVMhtGtqXwfkJ+YUyJUZfrXpekgs9FHr/7
UA2Dgqnpc65RBFHq/6sAI3FlT57B488rMZ+itvca+ChPywbhYgWB4AY1/wojyLOWH3Cf5wChew/y
HETtgfkdRp0o2ktL7qBi+BIsjx4DKKbnhlk1GFvyc0ezEEF1i39Tx4g/WHpQ2BaVsQiBSm8SNgRa
sWQtuGrNBWmlVzX7P2phqojXy5PAwNhDmQOM1B065FihkOzFj9EYDlS9NJnBtiNWTltpWUSYpcBm
aXY13/uK+y9C1yZart+ow1MxQSeD5PkfjqQN915bc8grKzaytTSZSlfVQAe8/HmTOTtOorgN6Vgg
3/3vIqi6HKhPiBXqbsuQhQnO9216nL1C3mxZ9R7+A0Ip1Kq8YdXfdvC7WsnDYAZkpd6sdIKZ1uJ0
+DsVTtOwCqu+xGjIWjqPSVhS6Z7/pjFgCjdElGkR4zLkSad6oxo+/YbsVVqdCmxBOMS+iP76nLUY
8Fr3uEKM9d352+yOFi3J/8dG97691Rwtfg0yakqE5K0+7SihXU3yQBhzYdRfMHWMSr1sZBGUn4oL
uv/1fLkacOtLO0lqaEh2LzuLsZNvCm+9A3J8Mwb/HSwZN2HrrzywPmq4/PJ1V+mJUCkuoj8ThnD4
UNWjPxgVvgo1lGdr3fmgSmCA7C7ia05WxzUk3wCYSzyRHHoYZ2mFrKXyJvVP8gI1rkeRGnOUGoUy
pTTuxQTZ8uNopVCoid1PMhtvxBJHbIpUPgLZtXQdy4P1Z0PdzUolub1uwrGTsBFItqSFJQmKT8RF
I/cefTpHTlUCSb35KufCd4indWX2kcXgtbpSsWCVkBbaf5xZdAC6+nRyFto9CJEQVq4Yusgso3uB
w6XSTxEPF8agMLCk8F4CFqGeULMQB5KFt/3wz7s7lL4tTQTo+7mhurvQxN//2c4U1wDSUV3rm68t
HBqXDBnfQOGUxT9aPYWPjkZ3xZ+Yk7CWWgwRxXb+2jPwkNi0HtYeZlbxv69znt6DOEjim4KRBjag
XUHdUZ5DcEnHplM70u5AC+5K4PPwYAVSPXHW7JgmfP5+BCat2Jccp8P9XKrLdF/mBeQF3+YlVXSs
DIzO+u8yL1RLdKyjhheizbi+B9ok5N7bzD3pAhty6jFplGrlfhq+/n/o1h6waCf4EGS0HCXGHsw5
3s9e5Ir7P+X/u0rcNtkQUP+SzzP2aC23d6F/vLXNjnkMmROl7dGnR9V9lmk+pIRXI2jHN/btP82J
kF7/Gxy9GTzpK4TUBWbkvofth5J/R4PtBf/o7Cdb15CgCFe529fJSlYyv3whYqm7lT81vFgeZuQk
1+6TCVLKJd097fGDi7GRVOBpvr4fL4XkQDewkiS0KkkEtdKQ1OnJfeHBBwMq8XlpweaQoCnJEmD3
9KhxqwsYq9EJfrniAYtTsRCq4tkYh0h5vc8R840iQnCee61JOwce82jfKU3yUkPjBSEszDKUXD0v
cTJlzBTg4TZVq0I+CHoFos4IanGWAVnXB32MwTsu2erh5daQC662vYYiFRbCCmBbqyaipVRod4g7
L7GuZvifA5xN/VDmevUj89KZ55Mp3YYgEpJhNaSFxg1gIvV/+TNtBDwlMtsbD+uyGHEX6nO4pHDU
EA5G3PbX+CThr2h+QO9nPIjyDbzvx9bbGczhN2yyeQValcZTcfjK3tQmXG+R2bhJJvWEvs8X3AG5
WxHvEehsby3reEcynAJP0QmUyz8Mpk3FlX1xTx8IQF3NklsYwX7897N5ZJsMohWOVoVBS86UlJEd
twICj7fuAnEs1ltij1xZtw6/XoTL2RYi4hYKq5ZEEK4JPlsrOjLHvxAuQTTiqe6fuH5U9Mgvb/c5
AvtUE6DEoXAjEm3n6WbyKOtYZO3Fb0O0SiEhQdznCv/sETOFwQbqlzukM5cpR/draM9ErqUTK1IP
2EM2uR43Mg/jdu4shYne/BtPlKxLhD2SYuIzk28TRifwcZ4v1zOI6P9WprSFkOcElYvLDwnfdpS+
t5upmFMNfbp4Ya2QlPHgmIod4+rgq2yVj6AsuEeQ95xvttxynaahnnfor+bs36jtLCcVEJhpMwbC
oRk0mgAUQloZfEPKLV0GpUyT9vRtAJEBDRR16vrT3TXA0sN/L/wOguEigsUJ4FTOrnOkdKzzRw/r
OgEXhveNHO4wqNvQO92RCztB4wdzuMTaY46zPWVBIb9Tnx98dOIovst2EoExa5XZ0C43/vEKlSBp
eCiDD0r+uaxEQsdYuy9JaVBF29Q0At5gy3s9kdXFzdDCYEy4pN2Nup7Xtjj0FPsBVWuN4DGoVDjJ
HsNUdbrLJu729EIEeb87JlqdsGfFGcfUf1h/HFFiAlVagVLW8VLIb0ktPub3ZRZziBdMMO7yWWmS
Z/bK5RwlpCGS6WgECXJkGDObWHbxAaNrs7U650+JE5jvBb8Uasd34ZXC+LWw7Q+gLNMmzFdgnyKz
Y1KbgN/TKgeHgWbj4ISN2hgIK/xN+f6E735NYkl/dTUl8rsJHLNVY1rzGElgqfsClSrW/vFI5zGY
2Sc7u58+nXSCYtLCf+feekHH1h7iwK8mUYPVmanAhDXPGRBVpvCXDLdtbjbAQBmjnAqRkiXdpVtU
X7hsiJHiVCbGtxlPHFjcdrBd832Ijy9LuNxoc2kNJiIs5cUIBM9fgwoc4O22vANsqI3RBau+xsAQ
mVjd8H2AR04MH4GTKQELJvWF3+Y1i3h5P/6jawQeOKHvhReWScaerBqZOGU/1krHxtlmOQX6E5c+
Do4ayUXuYM/W2bXz9TpmZEpSZ8+5Ye6B+3icmhOirVr0xO9CTFGvh6Eo1iYtbBrey76mobA+4Jq9
tNG0zjtw52e2zOnzwdb1ABtTksUohzItfvP/nVJZY4Aw28RljHnmLf7Q2B6LSajoGlYArjb/6AYx
QbR0fXva4WitdR8VG/7wD930pJbQklsgGRXNTJW7tpeSstBM3QnCsYgsklNXcvRlnhgE+ZouNSGk
8Erninfz1vQjbJu+d9hDSZa5cYXYf3x7Ocw3XRp0INFmtVJxk4ADwpDlBg0L3TSJwSo+VQytf/9u
DFswxzvL1BedxasNXfkiOm+VCMRlch2uPL+w9Ni+Lgg42ihXPSUfUvaChTwP0LPZIFGPbnjSwLLC
el0hpmgfK8via1dd8dC7Qq6XA+wnLEsjF7QI0t6TfFeBVzv9jmqwImcnpSpIWXPRNRD35Kv2qklb
BQU0yD9Oe0QZnT+WlVqGarGFrwUc3sV0Z+8pZ5x72hyLLF9dXZ283GbgtOXJgecPJlhbkjAfZ09O
JNx+rXUEbbe1QJfbJMGOG+U1GvWAbrRqG9mUmmkDIZKaBGx5oipnPw6nU0HMtWFm1tNB0xQjLzrb
JfomUAswm7AmU8Igdcw7xZ74MhcGoYdtkaOGd/cJJgy05whqXlNJT9ScZwdpsD1gwqHtKhmJ2bsl
PVQijm6iCXPojXbPN5XLXT68j7ud+sSFztiU2LlSDPj5UAJi3GjVL3O1Rg94v6wszZ8Kh0IkwL/Y
4dHb8Hpj5sXNhPFnars6vuAVanNvCmphGqIAX984EADUq5keHuFsgl6I4iD3BDSZIhl/pMPJ9isj
8jp6PGSsWiur1RdYNWqD6KxvIH4/TJ2UwbeaVZOnC3fzKAZLDBhWfK2Ag61K6j3YbrgefAgqV+GU
iFCQL3fwVAV5TD3OOkABtp64zWZYlzZ8Ul1u5jT15iun2S3HBCAfQ2VNaigktcwd0QR+JfzE8/p6
Ks/Ght1sjAZmNKqJS+3mFb7sAzYvLpz2XMCe7UJO1bwmqs5SDmGUgF+eFooljiFGqxpZ8xmxI3SY
VYTIVRWzKXnujFRIROD0T06EKxt0NAEpcQ1fVI76URNSUQvS2fSH9ZgCCurROpTR+FKPB+59iCix
TeQ+YPS4zHXhDKpqAyJGgwB3kRz0oJJwup35khPO7H7wyqhvUWHRG0c757NlLmzepq+zj/yjZjTh
YKs1uv/MMTsM9pFrfzt540qbnqP0366XzAmNKqxF5D7b0Vyo/LpbEHI7PekO/b2ed+J+0a6E22iD
d1f8TQh2qwUxqUEuPmM4Rc1spLvadUA5FCo1vl853rlIBuaWKKqyRc0VyTq1xX+yKKxgu5S4QSco
ueMpjQngXncUMWx1thAerLPieybkqasdlYT06owMSFxBwio89NU4/+uLOB+Jc8bf5oNA2S4SeByt
+YkcR3JvyRfCcEJwle24HA7kGgzVDGpk7eZ8D812P5pcq7yaQJkAHJssa748Ru2GaNBZFNpG6yOX
Cke0lStTIKRP7ilFubp8zxbmBtDcjetiUCPPVbRyTaoFO2BpyfTwZlXl/8eKMhmLLGYMuCZqxXb2
hoNRuyyL4jff6j2y0cPt9I2tZIVpTHEcg6HDH/je5UQPGXEZ+2UFbexDr5p2jgUKwpqC+gHLtycg
U++uA7PQs7tudDZ9mFtsMOH64/psb5I5mf1et5u6VFv6SLOI+m/SwL4PFtQUbji7D6yI0Z4Xf92D
fpNVgmcwgvlHUaHIb0z8Xt8tlKvPUC9vr5z0IBWuuW1ssklONadxmpAm2Of/ePQf9n8FJzamd1eq
YQ2ygrPTioG6kECOe3dqHIFgUSrNrd8/E69J5R9qWJLtkvahm4b2RzQrWeYlpI0+HN5/t68uizR0
8RX97oZkru9xFlXKa6BJffszMvfY1S9A3xlDcaYnXBJsuwE0sw5hw1MLZ4JRxkbuBFZcIYl/nBVe
NYeLqpjgypBZAREkgHDJJBTTaQRF24XKThgwzvECY7+PaCLqPKDkHk0O5uagbmY4PpI/7ZXzsuHa
Y20Lbr/paIx16o0tn0ner1fle6MudZN6WvfAJJYgxkn7qhmkpnlIvk6pndn90oy/7qGePEFgZADX
suQLOAO1I6ZPvx8qkK3TTEIIE/SVBUX9X/nwx/YFJ2tO0t8yhTDUH75HQCvPn1YeH9MS4WY2gnBr
aJkbHIQ2BUMKrNA2ugF4V8oIgB9RcX1Gb/4wN1xHoOnXCJ2yjTUbxUwrESf2PWTp49+ZVFD21fmx
g0SoUPNlB6FpZLIYo+mbMW7vMz8vjP3H6C45IiDxIeU1SHEBgQ2IEJ02sfa3jIpJrgJsMKN/83AA
6tvV2LFc25guC0ImmCVIqOHFlfVqpC37CFhesX7HdcbEdgj3JiKpb3MSiznFE3hCnuPYR6ShtM4T
iUskcrb7Be4k19rKyrLrRbBhQecD0hbH5OjHSdEaH2GSE1avGkK+Uo/7AMeOy0lMHqKbnL0TxBdA
f6E+JafOoLMk/rEYUGQxvIIVCiwKG+zchGzWmwxf17mrOcvAoBqQ+JaJGNv+GOX8Ebeo1t42qnYs
QupD8927v9Adyrz++RYD0KlyaMWjt2r+frgV5cxe0L3SSXtLoHTMmrEzTyX7UsyTgEl1XbeBF8nC
1h6+vC2FArPIVZ3YTcRFLtsIt63mkF/AYKgbTelU9fX6GGSdG1WuUpKdB9dLr3hKFCg5uQNehnil
5zvcnmVvrVyQYfqEXADMLIgGmvIjFaTs3uPmjMHNcOfLi+QxHnfYE+/r3YDcWSppFjnfEEFQI/p8
QggOcx+vebU2ClPnkiiNnM7swTK4f9K/6DSmgv5a5uZeE8xzFZRH7E98XFKHQ4lSVGGmVnRIeQsM
NP8tJce4Ap0kMavAa8Yfx5Az0JsRg50f7/bU7+iIFIaEsOlabFH2iaMvri3wNLhSt8N76Tm3bZpt
+drgv1oN3n6WUR7h1hWjtWOa4NR6MHTwEsyNiytNDrB2dkAHyjeiJr1iGMmtWK+UBcqH24ZlYnOl
cZdnBRZD80iMkZF1YoRdvitxzGEZcRzx7vLYMy/aCi9ndWRuq84Q56L6GCYi6YQgaX+3+MP3GTCF
vkYaWcpv/PWEiYlGjz3IQCGKblEDZ3cwflIiP6Y800ujGhQClJMKyx+5HRB6CdngRm4S3BFqs25e
KhZ/YHRr4FuKQukPlmd95CnpS0qVvh/odV/oLudagabE5f2H7Mmfe3CE5dtVVQ17Pt6C/bLL+EYE
kp8Da8l0RcYZN/gYlcvoAtNk5FIhZjIfKqQffaYekhH0fGR9eeNPAsBVZiu1OzYqMpUKTygJ0pIN
f/l03RRjQtNZFE9Fbrser7qr69q6UtVN/tEqp66r1pQHnvO+K9zuzNCXZ93v/OS68YNpBs8/cTR0
xKBOisyBHxipsktCpdhLkKFe4ckdjXn/PEKtUEmoHhZCEDQoW70YdBCmQG4CkqxFH20Ca/DwRFVC
C6s3cn9LbDxpZuebhuU50XOf/lAsB5qcLFZR+3c29w0Xm0FDO9XqalvfPtK6aMGTcz9/tGMwNlnO
gXDDOHubGjPpbi1q7FHJ6oXT43YVzh21ZedvxhPOfo2FO16LSn+1cKXKJOsEZINOd+PNwq7GUvrE
m1X2x4m5ns8uRTXY/0GsHzjOSrQT0s8wrg/xG5MUQv4UKRVgPgOvnH7yd4Tujw0HugIruP00BxeQ
wPkfiNd7HzbkVcZbTali01MRDYQPMYxIRBuRHPFYt4xP9RvZqIbpFWnSV6cprCI3ZEz1Jc5705fT
EQx7KcntQs6nK8tzMaYLmnrGzjyKNT7yIuIeklNh+awLoFdpFeiXb5TQYLorVtqZPAmHQdvNJxxC
OVDFiwLX809mhxTq5qoautEns3yZ6Duw7oovnk6lA2WFULIfIZEU0NfJ1gfsbQisCIpjdvXg4DRn
LIMYYMX2aVDUWFMSc0AlDeHBuH4EN2NOiXV9Qwxl4K2d5RoMY9+cArkwMiPAyxUrgpjS/kiqviNb
WatkNX6S0RxaiQnY+d78pTuddZns6fTCY+pioXcdBkUSJf57kVHIz+x5b8rwCN6igKzGS1TNuVRc
/PD/SNS3HCoWlHn3XxGfYnkfM26nU9kOS6SDvYrHiejpRchzr0O+p/PjWgcb8Scr76jjy3Jmpo6b
Q0F68D4/7BqHLFEAT1MrK2u6Q1Ni18WgmIEpe436x+rVdBpQyrII6eFPKFN18kN+sKpjN843Jpsx
W/6PwVzdWBj8IBf/Qbpii+8Kj6gciZlr3CjFriZf9bt4Yh9vU9CRhn3bK3vaqcfv0fwISIHN6Ipb
0+2JexQfPeLNs33XdEKDKFP9G9/c3o1fnGAnUhAInWR9sWTirJrvDF659WyLHWoKJimAIjCZaq3m
ObnnRC7unJ2wnJiwI2rV3Av0JxCbP6wUz4qd1L4PrNlV9MnVKlVbOAAPb1t6SeE86t1eRJTlMwdO
9DEo0mkgdrv1QpH2zC1EDrhlAkUfQykh3yl6DEq9LdFhP6DB3y9YDR4im0vfG+JR/XRfptdid9tu
zVicMwNmtBxcmTAe5PDJ+1NC4VfPDbIm42WVXKeg+lT61CIuoq4BWv+ysMFJZUIfSvmWtgRo4KjB
3guzJSKA4334InFerv30O6SrtJJjXo4IhvJyZFM5VuKoxXz/DgamJkMK6cczVDXscBeZDI7Nzu5O
uyMsvoNugz1glGutY8A78+9TkqxdXXPSJYwpGqFUCJKzlqVs6HCiKEp250kDYnMle4MzzqgPcYME
Qw1MBRm6KMCL1mHa5BnE22sTSGJH7v4gjT2Jvayvt+YtmixMM/d/oXUitHcQOh3guaEMID38UFXn
kgeEo8uNGGSTDvWqMLeFmGrvY3CVUXyGZowwr3+KyqKL+Cns+4OiJq4oBhFR//b+gKbYbArnKCg7
2X1mGDl6u3fdMowB9t9XYIChRdxzcGromk03eyaAOzZjkIV6GG9fbfsBT6GjhfFfo4EwsDe/W6Fv
GIfO1pD5OVBsyZJLwRMVHmw95CyF5SJs5NtUngup8a9EFTPZfPHZEaKCnkONXhv8xuO/qBL5/4/t
vSUs3adLlWQucW7+tBdCxEHMf2axQGIFMcdJOjRO31lIqHPstWzzX6GHeYGqclhzbpup3cpwgc2N
0PsT6aVQqeqfdZT5F2VGER7nuG/I8FQ+v4pVCIBBbBMR+w0uR4IUXTFs6Vl95nwebOWu/emiMHD+
TMCDsOUbGlsGrLwJ5gfh2OXFN98QsglFwwezyeWGavWZwZxowfzmlS2UTDZKAXMsfiDgE4bx9n74
awC0WyP54Rr+P72MMmxMJYPLcJ4mW4MYfDcxsdUozcQNv41QM0RK0+GHZQ0bkox/JZ0IKoJhtQGh
qaA/hKDJRr3PJZNgxxMtoXPep+Gjjf7Qs7yPRLbBMaCV7UyvJL4iDU59dUHM0tJZFQLuP+JFMg7z
ttq0FgBU5ZUfyBWDNVqZLYMzYv9swHfXMwgJlN5sLCIeGATBsDKqs5NtSmhi0KwFijsJqPmZoYgk
6Ca5Jt94hQNCPMrXy6pJbOpG8sdEunpINN6a0jLy0K3LXDGY4VXHGKdVtw14Hhk/NRWu10M8FU8W
6QZQLlcBtixttZ5ATZwjaoSS1EmUFEvYcZaW1OaexvsTp0VBIGDcpOyzhHorC7TuuBcFuLStDXzM
iUhhKw56zuAYAcNe6+Z/KweLK4SVlFgsvbC15viNbraJ+/JUTuW64SegpRBYw+2Z1gGxSHTIvnrw
/VSKzXfKS8M7rgCLvivl1bgnwBRGxydKAuOV54YI7AhwAQngqeZTTvHQEADbI5Qh7UDVJZi+ThzK
r3fzeOcmWzhhM2VcHjXxD+zR/InaWnrr8KY49SAEV59Q1MaocGXYFZ3DU3D55SU+fDkq1rjBNIzb
f+1rlBfTvtUdCDTfqie11iQhGqLDlRA1+WnG67YooYyN/ndAfRQYm63Ep+MlVTwKK0/2gnjBq7zQ
cv91ijSMdstlOxE/pdcVlg5a0U4vC/u6ad240qzXQV6BSduBLZZpM96LMZPMYuE9q4FIeR7ezwkw
jaqWizaMz7yb9UZxPWHPWwZTdoMYzHUwTlTa2ExZgMPJL0tpc8ptCcMC9C/uk5KR6W0VhcVMSALJ
82HPu76NrL2lA/D3psVAPF6/HCIMgJZj4DFIB0HWfJthC5b3+l6OlQR/qMXi+s0GBWY9E/VK45L5
Mz6xLvsxoGFlM+jsLE9stj3B9tVcjrI+7Der5dfgVDwM5kKu3wLNGO6P/oNQ0z9pvOPPqXWQw4aV
Y10ooJTCRkDha2+/O5vVdIRLh99xG2gX9GkQS6RAeEoY3siterK53KYWAaq5XNUcaq4P/7KYLuNL
1whWAfYaTJBYBoY9+JIss4197dg1lYzepsVvNDddYDbCS7AYjn9vTD9oB5xXR+tsyPmUxOltEjho
CCgMvr8Ggnj7oGi9q97nNYVlrtxq28WsF4M7fctulupacX1u9o2VxnyUpc6Kj5oHY84RuIlzV2MC
toiUtEgbpda42sY17c1IORvlRTWUJUi/T9fLKtuWV4I3P0l7VXd2ojujcrPMiql3KxaaGCWvpdG4
+766bxZqGZk4DzDpU/3u7ZK5qGWaZEXDKY0Db0titJLY7BpS9KOv28iFD8xeu3Qnmh375zYJ30AG
A13GGZ9OrQOkmHn1ZewBNvq8NlcEpK/ivu+LCKOqbwOaf6z6UuL4c7KRnlynXUv+kzEalCsFowv4
fG68Rb3bbNlQiaig8yEFy91n2lh6MMgc1xTD+bSYOxhuJu/cDU/9KpOQd58YAFUo/fpuhvq86Q74
1HdX13gyJFkHX9BrLrSPxXuC9H5sUQEDEv2AuCBhnHGXdxwyBPM+F5XgbDWsiAxtVCukHbN1PO6H
JAE8qeOfNP9Tp3V5Wnxk8ItmBtHUawjdUs6YUiYoyynxnS5L7rWxYRQ46maDJgBXd97Sn6XCxRFK
NkBDkl9DO7yA1YBPiC1upwRbffZ3V+TJhxq8mGjFj5MvF40c9E+QPOKO4NOPI8KS3MMLb2rVHb0g
3pXJT0GuP0hj+XhigdkaLQjhX2PF5+w3W7O05oTh+PUfd+hNAqWfKawvuKF22028y7qjTbSIft8k
INldfJZD5OYoax+DRnA/xyeSkxtE5MuP9nmgMVxNaeMUTNCm6pREfj5CWZ1es7ol+sPYMUfw9+HR
ci89Y/tE81HTPJ0DW+l3jtfLfj/mNiHXlKBXFWgaz8d0vVOhh6MLRNft5hnlp4fGWh+BS9Qhjvhb
yxEJnx7iyCWsNVLxUfJULEITSj9afNjTRczMQ4DS0QbZYR+4t57HYN5Fr+O5O8Zi+a1wYo6GRuzS
AqigdPZK0niVjNab05plY/V6WMMWyHArl1Ov9KSYEyDMIqh0v4X+1H/1SZp6EXjU97dh34/4YkFJ
7suIsSujGLLUdJvK2KJYFWtl/HyKzcJXYkczy43gXsQsYl57MnL/15YUHaHj4GoAeCyCqV0ZU/5L
2/LKvHOKmnpXR2/Zg478jz+sv5NbQwyfQtfW0yOtrob6M8wAia/RnNXmhBKXTuHwDvjzxkNfIRVL
PPwyJ3tpgufmweULxyJarhcghqiz55wJZ0EeWrFnMw6dFVjPvLZtfyWQkgCazO1aRzEJbc2kNYFn
yIfkXCXOTLUcT91kpwPpL9WxIIkjWSVqsWgyZYxUTynzPeFy8KJOw0P3sE70OnfVZyTgFQqPfZjb
WYMQlvpAGEBi/6XjDc9Bp8wv/X4Lb+95t2SGD0INI6TeweRLd2Q0WoN5Ip54r1khItC2EK1/BoGh
3Ou9gHHlPTP9AaAmtS/Gpta6vzdyjIp++cPaKDvhdipBxLMHPjZzggDDXifCRPx70kmu3O82BGkP
ILLs8BcfC2tN5sftCUe+y5J9sjimo+phb2l6XQLKzcLybi9Yd14w5ocnAewk9Yttg+cDgSAfGc4a
0TCaZdkC5yjsdo5qSzUA9qCxHFg2HagUZCe3Gdrqj0uVYzvz83ahEyrn0c8w2a2BAdLkwc9NPBxO
bKQHKPLEwkBoaQWMp0aexbuJyqvxr5nJliEuRZ995lG70Y8NWy5cEachuOrKTkPn3VRcvovr+l9n
6oszGZDP1LNcVrFZH72PcATy5hJm+R8CClvWVkRIVSN7cOk19w1at491nbZqUDOhZC+uoZdJp9q4
6T8T/Gi8qkf68vJvzjJSQDT62G8l+MQaQZGOq6QgF4IuDP1nrUuQT+7wY0GZbdhGk8ycbE/PQ4Xt
j9+ieWAiQ1Lt5KjQ50h7o62xfEIbGwI59Jnl5vFaYnLDKh7dgtWhWpX/c1XWkI43YTWS8mwFPrbh
jCxljZz9ZOSdlak0X6aXGnqL/SwfOJlB4CGrTio6z4kwYTEN1BhhKhmweTvb4BgZ8Zqd7lXaWGcn
xsdOoOCNRL2WxzghCJ7rHlt8FvL5lIVs8OrdTfdjZKjeDV8+sBHGQNUsfdctJQsRZqIy5c5/TeDv
Nv6Sxxr0soFy8D2LqAPu8+KiDJ8rSUDWbBaXe1iNCkzhnGQIjPTdaCcdx5XQWXu/+OTjuMh5JBT2
tiw1e0KBvHf8X6JAYE+dzhyJNxpupqZnxe3H9ufWspE9JPZHNgGnLZyNCltGtoGUbPb4R9EgbIDS
Ufk+Sr/lXxEyCpsY2cDTUYS96Kn/qO1MNEW3Rz1EHLZrDqwmfFi5grKsPmykzhVvclugB/UH1kh/
rUYH3OoL5nZe+yc3DbyysCbyBmfYmZD/Spjuh9DBkxMBMQQ+VJG+0YrimisQgnDPKUqrIqO7/kRM
b+Z+9pNYc6tOjtD30QgbxT5zBiJayrTwD/LUsWOQJ6qVXe8H/Qy0amafrgGkDsqyCchKkTEltfbd
pHavQBAPM8CpObrIP4JjcXt5eTUhpMcav8eCxf0SbFeB6aWzvNT7f6BWKibA0H3aE9J1++EelJXt
hDxrrkPgQDNyZe/fQ2CfS65z17IlGiSnEahqUdEhWR7qXCFvXEORkrDfwD9H7LEZ99wgdX+R6tKG
lXHWJ2LgUfHt6ImNhxJbIfxdim3H3C3Ue1uXBHju2o4kk4VfIh82ab9bK+Ylw6Yeb4RdZRQmvS3E
2YvBFH9dV49PfF+KDlaeKRnSWrIEIPqkEGqg/v3nwPjNf9NkDBS2DfMvsC8VAbxDlAz1Gf7sHLbG
mt8gAr32W387BFQukDG5RyvANUNnmjdWC3Fvla6zckRUAFKdOm0tB8o6DP/ebw0QPscFdPXtya2h
7jxV5/TfigutEVWqmK/Llid/3+WFWDnHkDdpvBx4ZFQtK0//a8KIzEAiJY5kCyYiDFGwiGDHf8mo
67Lp6V7owZJZm2sYuFouB5GZkCoZ028KrDr+wO9IqRLiVV6ImLi3bIbCNyhoWuR+MXEejzykQtKy
XO2MIyoMAftLu9v42IvwF+8N2navouBtbEHH5b06SNLfkMimHpHnIsLHhLJikMVdGhyyKgGCSUKt
cIyNN9VPdzR//x44qVANH95tzTwCq3ML+iEkngzbnfP98dlG8jjRtSlV/dFGGZCeObforuKy3srL
cYPGyVjG2Kpeb0JM9vFlxpFcMNWSIaXIHwb/RKfsFEfptwKMoYSqGwc42pPCwsWEz+yh9Jt0F63t
6ckDkYuczmxTGqgbphs6yiiusbFzVnJLZbB+O61HRU5aBjno0x0ogQetWP3iLhML7w5wAnG+Wwsh
WZ621NOaPFchmUArWNXq8OtqDaaa0uEB3O48Y/9rn3+OPkJkxpBLtjApopNthIV+b3PDiwWqjPwv
EZo9/AlWZ+idAMmREiGHQ9MKCRCLcgSJHqMCMRoXop4SpoaeQ68xHqK59q52J1o7EC4W9rlUjhxL
zZfU44cyTxk0bA+Q6HK47av6LZ1dkkn15YkgWDm3XtndrA2xOJhWMwkXY4JpSaLSYIVPfoQcEPgP
CFmOvSrKiiABbTt/HmGosKjdeMH/zSpffs4LWAMc+6RgQ+wiyMwX/PpJY+JATb1LVB+r9Mj+zqOn
j6zGJZ2YiSgA4NjIMxo3NiYi29gtEBJG+N+ykqqQfTyM6A/Qb2yARbySBUkzwPBeZCF6K35s/zqg
dfi0pL/roCmrbS+JA/oBDI/daG7QEUF6x0Y5RQudbTQuPWAFJXNXO/P5B4oS83coLIbsxeKgVbX+
vfMG9FH4dI0kP25RbZo2CtzhRAwpcK4ePRpyCZU9joxYsMVs01CRxFy6+Yl1z+MKNfMEh5ImZTiB
I+vWYEnKwgF/yLgBe204Cingl8mTsIJxu6JxjT52xvRacwCANmoGJXRo9ediWL43yQ5G04rYfBr5
3I/Zg1uEkLCbVxDwtK9Zh6TO/SjrJ7Gnr+KACh/7D5G+QlaLGJK3HuqctFCrDayQRtwqphNIECk2
4Pgs1I6ikriOUK6sTzV1cWdPH5Ps++gtxB7fWVxSZdnZ4dk32qvEJ0fe7YsH5giiyKQnPI5mZwFr
+Hs9ttAOSSW+KGNelNS9IKndKYJE2sNLfnaQLCNRZyN9PAwt9+WoXhAO3/wUnBQY1vpyOQ97T0by
GmOYD5JIP9VN6DPsQfHCO0zUsOv23NW9CoGVlZ1UFXA/UdYdpWjIcs/31QRcBEAeNc+Nm17XeRPt
ICa8omrHPzHSpaHtyOjl9wWxWenaAgeiT5Qu7JXsY0C7syFM0yQpbm5/Ssoz8+AIHdbmftVW6aXe
8z60JACbCpCmTItCHGKGk1a0YSTyNodntuh7PsMwQkbpNBvKconV066dNgWg6peeeJtmEFTVWjgj
JitCmEXx9BDfTyHqfK5uhVgIAB1Yj+ldsiBJ/m8raLVF5l723AmwbRr7p4Mw/qxdLyhrnXwl2YsA
XxPdADC2voG2NrXU8SCaemv4Udt0Vj/Afz0NCPJf4Ka+y/ZjZP5jV7ZOGeSLwAq0S9DiJeplCjw+
SnIy2am0o5smC0tUXDdG/RBs1k7teYY/nc6kk3mtBcLfABsQU/bkuLtWIWfz+PFQ6rEhbbrDJLU+
34H58VMs/nCPc1KD+9QhbkIRTgtzCfcmAlv/6hqF7qsTGSaScmiFZeM2CI5euqxRpfgIzTa8+PLq
mJO/54yDG/tk2Cr8MK/zjGWGKgmL/kdFCtdyqEz4Zz6kOy1YaALU1KZFaoLMReY02rK+065A33xI
QHKwwgAYzTnWZajyG91Rg1TDzuD2W/ocos84Gxm5MfevJ2fG/i2YsuLjHwbDBkfYtZZiSU2G1F5l
8RMPyrOMetFPPyqFt1YO6dERW1XIOUNdooV8uXiXFm0WrZHSFoiwY0DDKghK5jBZlu5ENb9JSuSf
5X1AqMjjQDZD9jDeYY+5YlZLQvlY/+8zJGJYsTejhgFYURaiQZzlBjBlux4kUWF9a9Nus9411Bof
S1o0FuMHBirZVU6k2PUoDflQCER/RXqWzcRvfsOg5laSMSjJqL0naOJtYwlQD9EX1AWt8tg8rW6n
N7sh+LONyjt+dtxLvYnrj5PUfAtRgpOnwn/j68ZM5DVl97nXV5mdNs6PMN1NnztpWCDDImxAdbV0
ahCGTkN8U323XGYbym63mlqA6CqrQqlU8noc+JL6L+/JiXEFqN2UpTxnmCsf4R4Du7XVMHkFDVuJ
GJoGVFmkE39V+Rqa3Sd2eVXQZGDrgIivQHasQF9F3iVeVSmW3rcKzfwxzbsk8WZr++V6NJXIOhFF
hb4hRTA7NTdh6Qu4V7TpQS0LDGloGXuM1ih0IxBpMatJcVwyhzKn81nA4NMP24/yKblcggHn9WDV
rMV7Ef7G1V5t9cbqwhoXEjiCwX2nOZlca7H1kSZh3DddX992pZtdmDW9ydTek7Q3EDS3Scde1X3v
rqBw5+EXWMXVzUxZc/lH8cMqdgwKDdMP8CvVkXtlLOCZOMS0NPrdEI7WeKYxcXTue01mnN7CI7Hf
/HYPgcJBzR0VOhc3Wg9uJ+MCgescjiHafYKPsDaCLui68MOpTG+CxiW/Awv5XanX/XjyjEyzkuoy
Hw2ZnIzDBHYpQS+NmcHPu123ALByVcjDQ2J9H/KiK1I13IuztTExru1aih6yrcc4pdnb05rGzpVz
mTqp+4/5KBtV6vvQWT3syZ7TR+BbW7B/bC5/5AwPP6prQeNFVFPnsZM1oOBvYDlVIvWaMRMeid31
8mIrh8WrwVAuqR0PsTShUEy89GCxPXg9sHawmx9LF6tdson8Cpqe5gQ9tej/08tYn0pnHZSZZTxt
gW477bgSiQy8MqNWNywp1F2FU2BIqJtW+/RGKg7OL/ZFluB2KacjayqTOz1a7L4djGF0Xnm6pSdY
ohorWqQwWb5KfJU8WHrrYJGKSQVW9wBlaq9WQ5uWJbemvRUMMs7cLXYTzCjGSHTFPBTMJzKD4Ks4
ozSb5SFN3Q3fIwf5KYF/jpIrkQkYzSGW4VuMnwnjFmqG4+mnk7A/GwHpICktbzOxYzNVpI5x4jR1
y8oWEZAn6DeWGRBrHgIdiV1F+jczgRkYz3EtvEp2a8KJSSi8Zp4PZbCLHMOHXugoVnuP121OqQuR
/sA25baWhnikUf1glVkXqgjdu0+tmrUo+m/GJ48Z9Rtq8DM5q4c+CGJgwNHqiZOhb9zSAru9eF+/
bMsx+MOoyr4u+IzFo4KgRp2OGjcMRHi/CoTBrYGBWdLIPOiKsfwrCamgauaMWL2Htf2UZMVziu5a
iTQu6gjTTJZvO86Ha1C1IpAIqXK/4b626BWEFcIYBwMxZ+xx9Ag1+tfEkpezuAAGwN4jT0VU5DXe
D8EqpQSUL/H1p5FN/cIhOUowEIEEatqLR9KzWFK8F4r0hP+uEq85diilyD8FNS4OBoVv/uJ9q6BM
WXqQK0Ep645aNDz3zn2offyhMLLjZDUmvod/GYMyQ1gChb55ZHSQj+Do5Rjv1GNhbDRRGHOoR+hY
eT0bVYLZCmSAgDRas1UgF8FCeckSV+3TGHgxK+UOMH4CM/Jhnv9/DbwaG5es3G95T89bPrrEacgI
mO8ny8PktljP7ONYYVjGk/s2tQkA5hEV5L/XF10JNXbBJKM17Dwjor2L2aNE77/mbR3P/bxNB819
QbYAMr3w+bTV4OSkA1VxPstJWv6JrulVzILjbSFHp6+kXAgESWf5BZQ/CEBHI9kebJRFLTgUZfxs
DT5tkHKBeS3H1bBHq4Kxe+tCWipQPhMeq4K2F8k8FCQSofRCYTToKj1cGxNJ9UhHjZRvi+dXepun
pTJvFQR+gyob85hBVD73cFmKYFcggdVBqanxw9ud/twOBUDjTJR1QLCvbJM0ssH/YMZ/OQNdCBkm
9VLVOobftWvwevPdfbqyPBJDmAxo55MLPEQo8lKeJoj+KxmaFU6lPs92cuzuZI1ubgitugxEdiKh
5uiPet5GonZEoDBL/eE+Npx/MwPRlUMtMWCWhK/cudnZEeLbt0+KbMHGtHnbFpmpcF/QrndJ7d6W
XrpXfgY/X7yRzXCIQj6r8cd6NWrgX34Q3JiUhxttyD7UKqiPtA1Baaq9tfiNrCqYGGuJvqGoQy+j
/0QgX2iT4AvhHf8aWxmXY8CpnQNLVKvHRgKFtY6IhrifSdV6FgDyRVugb3e6Ww6NkrXzrCi8Jwok
ILhKKdI0ukv2sq5pjyhLbeO4JriHBJSBJ8cgEgPlOVh29lhFKKEvYK0P9cb42x2he2LfTpdMEUd0
ziz+5TIYrw6hoAD1lIObITb2RYcWaeE37RY0xDQAGq1ewFqK6peYl82MR9FRO3rUp57ufJeBQxYY
1DvxnOz9ZMCMjvBHl2Agl0yHK/M889A69oTC2HOyuR7+FYYg2lzVxlLaQRhnmEbSQfhE8i6Eh2Lt
gb5R+cPAqjsGOFuet0CV0vogctSgt6MU0eTqvZrMXCwTBb8NfapLV3yv+XlaDeW5c1XwXhDkj0y/
DVPCYocMihkEZx4dpE4JYmonSaPkgSy2aeVxHjrOTzGyOFzMdXUs7ytBWCe/RTJXQouE251k8Ypr
TnTnxFa5jIQqwAm4z7LmaNfilRsPBzoev7hKD9avMtiR+tMXAVE3Sj0R+ZnH/00S5xzI+dFOMK6Q
knrwVvg/5x733L4f5ggTZB4ucoQP3Lrcp5I2mWnmPSfOYxpWW2Iv0mKZ1m4BndnGjoMqv7sToWfk
Bm70/BDuctgKy4IAbMPhMQ0Nyxo5FPbUM7zvgr9XZXfAu0keyGw4QZenuknynbQV4Dse88xu1PJS
kq9BQiiYZFHAhqgdZTCf5kJxgpoVkwKOb1aInGLEeOIxkGJSAOjPjPVyS6Jm0ijG/Kvzx8k2pISq
WIoPvAGwhare6tGSssH105gY3Jn6c7jmrg+r+IkrJtVjPOMXqja12POkOtjz1xmfENPItJsyDxN0
CiR6aL9FcIUTbakQsaqYR0EX0D8htqOOeLXacxU9JN0/n+INKZ++p+nkNTI80EyhNOztcZKhVAPx
HXJhU+2iVRGytAPjpg43PIhkXx/1uLkNpRthTfo8bpfM3SVTmAd2wQLQF9o6FeXLN6xDaXvRqaUY
2n9Vr7bI87D5jV7gXjVajN9GcO+cAyTOijl4mjAvi5Co2uRqCUIs+RqzBAMz9fBvZgWvxZeQ2yXe
8GGwgEjuimbSNyxKmE5AvJzF69mnWwDvBx00GCzmBwzuZu7dPe0Mgdjx/nIsroIc9ETMImezJofG
WxnNF98qrW+bffQe5EZ/GwYM4J8hAgRH2uaxfOVgi5OtfAC2HmqVBGRi73l9WbKDv+XrnMnx/3Y7
h5SNNqDlH7MZzkYbl5dFU9xQKcxBkyxIZuX+PGCjjbc16d7M8sdLXTrwFF/+iij8Bb1kjZjm7LeZ
boFp0cb9+e99Na1kXUmFY54r8FqyQvE73sLHIzK8NsohESEsMIqoDflJbLZeSYhI1WkvNtyQPY6Y
Dj/m9c6vxrVhxyYumbwqwsTQx0cmIHAAt5oCJh60YFnaC1dmxTy7TcGS7WmaBZ9bnN2A2rAoqs4W
bUjTtryR9C/7ykmPTVOup5ujnVt8n9NY+b9om2iMfB4twT/qeBlofvh9v+yxd9hkGeyi0KKIqIGB
P3iOD0K12YAFo3e3MHTufkEGbvFk0AHX3ZvaWPVtKLhcDDP/VmAPCXcGZh2cvkxun4DwNmWVJzXA
pyGNi6McsH3dM4Y/ewW/3cr1LUqRJQTfihNyldil1Ix1sP7SEwNfHTcCSDqUJYvBrXaK2M/Kh4Lt
5KYhkxcG1xiJh5r5S5LC3//RHyW7sPPOyHSrp9uecwKhFg3h/07lOufpBd8nzJZ1TH23EjfzMoNZ
0qPLufF5aQzREPeBf3f2S1D5g3HDJqFcPTsvBYIsYRBSMn+KTsaWYFYRABihhrYoL5ZFS+5Wp2cV
6JDD8Y4ETaNhTCnfOGwkTxEa3PfyFlsvZ/kV3SNXMZhs7kr5fyWvVugO5LusM8NapxFmNUc1MBqn
jJe159VkUTEgMjAds7USY0rn4wN2sau4LT1yFuOzu5+E3+G05lJKDlv+PtKLfOz675o082Ojd77G
5QyY+LvKN0h4amSZXQabhfkbb1mMc9QOkglUvXMwyFqGIbS2Z4D9gVtavQ1757N3N6OX4NjAzDnd
PNbrUmt+Sk7gyZe72Tp4UN22X+PJfmTQhULzhKoCH+9lizoFnavYVEsEJtbQVqtfkwdU5PA4XYNZ
Q1twi49LtP2zvzc+W6rajud/8EiDfwDDJCQqKtE9Xt9yKzr+uZFyv2Fk/U3Xj4UBvurlMMU8OlLX
WnhsQd8hjPYjwMK/qBhk4FajZgnrryP2CUAJn0FmCNnsVo3ZKD6pFm8ajIQs9569ZwFsDUGFHmiJ
AzYQpo9ePZxn8U6OUxO0zeYXNyq2Knc82pi2t/mFjAtk7j9yO7osDWxO8CrvJoMANs6yNgXVbxaQ
6+6sDXgnTlBvuWK1l8CKrTtwEvDBfTarYPsDAEEB8OavH04Ox84YCqvJRxhmID35JtXkLA3wCgB1
yj2KsaUGE/0NajRCRVDiUbOyqzOyBlW4BseKTdFE/PB9QrLKhCsmds5jzF/oy+hkXovdfsA+iSQY
erP7ZmEIBVfdhTMKvrcylDOBAlDfTxcG2C/FWqdxNfciTxlt6c8g2JOVBJjgAFpBwTSjd5p5dUH+
TkMH/9s8KDlRSsOIidWNgYgmwsvxjgajjF48qeHfikU20s0hO1koXs6mXWxMcMzBkMSfYJUXszbg
UcnZ3w7oJBmbDqUWysw9WYq933v9g+77j41rQ72baYtrM42P+96p5Bv+/QW+zdjfIFfG1r6ahXsN
YDbIFAAyP9PI+SuGAM15SswfpGjtSePaIaq50K0wBwqN1JYkGFQTuK6kUYEcPLyTOE8XVFl1pCT9
Zksa0OquWJPGEGnFtQ6ESC8zkR8/KScslsGwwDfugHFpH2PRNXBqLolZZgp4rc1CN8SA08By4wzm
VXEYylB8mRhzFkhNAdC7s34n+A3ta7jS6/9uiYOZ73bxsk78+/BYdeVri9gRz3OOlNCgdLDvHMS/
6c2TvKPlDmVqXNNjdpytfiwXoFb2Mn9Ez8mJ8TEufwa5ZYd3eelxLSnTV4zQEThlR37ON7qi8P38
HB3C5XAKpNKHb8vf7OdprttUaXqJpIcGi2lk6x0dFWryWa+iClW+xtT2cwQNVB/BvCuoqMhR/2TK
VaD9oUdsOHXkVfS8YWXkO1Rd+P5Ixa/Ttb9MNTn5rInLxghNld1drj4jEyODdAjJ72n5gklOlGBe
T4C+hSE0mpS09ZAfegyyc/B1lYo49nshzfDwLgV7WLhgyFmyfVhV5ocSukhf3OaxDASctHOhUwmb
fkYwtJoeVVC48hbRhfnrB25TPNxAzRE2i25G5bNaF84FL0Ca/eZFslahXuhrnL+KH0ESK8FbACDK
zQBsvkW1g/xB2qQKwJ7gO3R+Oyxk+rqSeZLwhEXjzA3unsLe24YtxOnByrfpuepOihaRtgSWRRSB
glUZGCDP2m1R5Y9MfMIp4UvpTByGZHGREUFW/xuuJYLDWJfEWm2qVogIKMZ4v6ellMbQBKqZVUSK
cEY9rfv7lTPgSS6xMPOTdqVED5UUYmZ8tpajHgOCzzr8xE8+Mj9h9j8AhWGiX4UnzgX+2kk1XHe0
NXMCpIql0sDx+vYNvPYo4QReUhOznJaLVc05tXN6iT0kXHaRfM3YFb3r1YlPgyC3WM6YuwdDGh5q
4peCfNnBDRoBC5hOXfWcTvZO5wVIuuEiL7yRxtWMm8/VnSjf5MiVF5LSsjLakuBRhbZM6+0U8H6l
Yj76/A0nBA+ts9XoLjtVcaCHVWssuAJDRu7CtyQvF66FdZccoTedn2UXLB258zaW5+KumYVpa19C
4fJuOyJNlde+GIYpg8zjZhp7bEVpKV5jYRvR6VpCNgc6q+PQcPUROmDd2xs/DtvlDH5wJDWbfVMF
zljIt/CMwKOA4j5OfGLVrV2Uxg0aUEFoqAE+O9mwiLYUdkP335vogb6NWPtAu4KyxrnMfvREHONB
Minl12pgHmlBLDEIS6v+UPKclPUnqzaNStlipxoSjsQW6qFKmTQWJfdWiITZqVOVvxJKOK39Cj/K
68jKwupOo0bWCpIatXszLn9//fUR+7sOrlhFBhjKdXTObO6yVA2swyA5rl2zm9eDzcbCoujM5PZU
Rab26LyXPWNsh+XCwP+ro8GooA7hvki8dHn2/1RR0PCMNNNEfLDi0mMTSCl/Hu9Tp05T2EkFmz6V
3WbZFLtggDXTniHlsdHf26TzcnA3sDFCBqnOiNYAkYAmOlSXPIZs6wYrlms6/pyFFDba9BsgxOx4
+bE0s7Qt7awUvU9L5mc2iv2ot86OoMoH7j3K/OJHMGEahfJf+GJ81dckAQzkIdRPcq/feAhkTjhR
eMlCrwNGfD053imyvnpUxHmMJQJFUS73bbgYTUgsYuTB5Vr/fI4dpxQT51uruQ7B3iuJ4qKSZgTz
vvtunCOIVuPnFR5AVJ2n/PqKVXNyUkPuNh98g/Yn+3nvr71o31St3kDo3caukw7mt0lY1YVTTo+l
SaLv0szy3XfcSwqyqOP/eblFf//5vNca7JBSQl9nOWcpvI+0ayUso+nMg1t/qlXO4P97MganeTGH
gsM6XPlej/MnbMjszOk80q6ROSBWUAKjXe4icoaXp4aVA2K3Jq01PzFyS1hKXEUAEQg0UADSVQKi
/FFP169NJG1pS32ns40w3xczJy9qzat0HOVbt1oTEXOswSTznbjsWp1ex36IN5oGXLJgjuJxz9Wb
TZMql5CO2Qc5f0wyzl/fBBib0tiMzAIxtcQfcBV/K3bbDdFvIl7l0YwZ8YkZ174NZvrA2lhixO9F
RKIwPViYdIxPLt8Tmjg4Q0ZB+sX8UzPFF/hYzBkJ6YcmTSvbUyj1ww44Bd7WDBQG5EtoeomSHvYE
Z84hRQcmOvTkhLXA3dzANe1g/1pybVb3omji6Ul5RweiwFU8Wlg1+ncB9xtc/81KIJX+v8vEOSlm
ITgVauLoaWvCZrYsBB+wygzrhj/zxabPdWOwtSnmDjqMJpP7kqktdz4qdtw/dkvdnrlH81GGvCFX
rXFHS/k21ibGs4rPLJZSjX6hq3ond/StgAjgsSm+kUJ1Pf0SnTv6cP73/dATi0QUHG17ax8LyBzT
rgHM32gydMvdRqeiWuJ0qsGdyWjNNLb8tVqQM01w0CZ+OWYl7ng8Xg0KI9AwgiC6nWIo4CW3Dwdu
SZbEsx4GboHDJjpLsOCJDfjYaJByOKBG+PipLtTQ419SWDri7NCZUoqSx92l4RyJSFTgQZ7pfDOa
Yf2Yl9M2OS7S25IlLMBiB3LLE9grdcyrPPU+9xK1XW22wqLQei+Poaw8rQXbf5+n1Xd+jVnlHHLP
6c9RBGXZtyWcY5SP8AlXweojp+pfdEKFHjaNrTK/ogXn3cmlqpymJYcwxZIjRgPcvt5tZT7r8aRn
zdvsQYYY6tMTFQ+67kT3gl1PmyQzr3Z0iWVrpCY5XsjIfKjSlkViz5YMykKkdpYtYo2shq5beMfQ
djfrroY6Fzim8b8UbEXycwcg4MRbt/1IrnLUgsBs4XqZU5VxSQYi8TU6uinjkkR1LXjc514SPSdH
BaZswXsrcOqeOgZdnUVz5l0UonE0QQjUImWSX5OzJHosWCB2xmFP904IdJfwLIgBj7hKm1rldAB3
YXpiTxiljeVzQoWLPN7PWyX9bzNoZE0EWv7Ap2BY/lhULUXSteK1RpugZlWZZZmYqOfx63u0T9Yv
iGA6JSWiYf4E2WPWM+YFblmv0hXTwSKpFRxqfo5H50BEqsxUzXpW3o7bX4Hvv0OZ60KfcS1VkTdy
vQlXQttg4UwOuG1Gv5MNxmduyUKBoyQIJziJHW+eAKRkFuzpw45VyE8dmEmrGC7q2EeDo9F1k6lm
9ylfK1MKsBngrAcg/gHVrwl8vcmmGeibfmrztLsC4LXJv24yGY54AWCiXz5Ct/uwC39Jlo5tCzmW
U+s/TD5GzAph1DIE8T5j9mBzOkl4xR/ziV0CoMYUKwp+ZQa1JZs7OMUktHDip7oXNF73Qmds6HZV
zLi03HfdGX5sqBt0/iyRTFZLU5GcVoP3UUD7FRWmbZwsmH7d/kXRpIDEqb1fRJyGQt2rRPkvoyNo
IxY6OHcW8o7uXMtpFLcBs+Sqn14FX3f3bBsQYUZKgPoAofZvkf4fyhJEUIzZ5u9RSsP1OMnMHkPV
4e9yTfnNk5KayaRDaz6XZft9ANEqFAS6pcSogyBfzG1/+hMt95/FvJSTFPVpLzKgDQRACzpDBL5K
8B2Q554ZHMRdZVRYf8dcJklI5VkJZPwJ0tkKM3YMtqNQw6Y4vUZOJk3AFkZtR/Y78ioh3rN0fR40
h5ee2cDJ9xc29WS4ub0JgvSOHXH+QHENTlzAkZA6Ma5kkzAquu6r5BfRh4fShPff5wlUPAhLklfS
aPrukDsGXnrTUIfhcU7dQIn5Wpg/9g2CjXMiSIWrzrjCWYh4iFR4Go4VCN5d2LT5lornx/k2Zfxd
ujVtMzCVqyBgXJBg/UvqpBLYbNvWRjHoZMAZnlSnxs0RgNCGIoisnQrdy1RSqFT9KHK4dfKMomJk
w6NonXnXmCQRyVoQWSeiPbjkzop7tvGtaZ82cWVkXIHlwaPSKe2WJ7jNDpiov0+81wHDXvduMioM
edI8ZGpTR9Inqb8F3dbTjNDSYZsfPjwc3T3JJY6IzQYN/7szlFu2HwKbn7WOPEXgAlTDmyiILsTq
n19L1iTkN9WfIZOcSuYsDDi07XPDqWkM7VTlNym7hjRY8ir2QE1TGkRd5ciqnc0ypanAuuHED6Gm
9weEUEcG62bqz1Ueq+cHw668Ap24/r0RlHM1jVrg/JwlMCaVFQhksM6dSbtq2aYblDzAuADxwDvm
d1sddwLOcRq2mz5EFyjAF+xB8+AU4ESu82lRUSwImJbxgu9uWUNoxUrP185ikNlDWrLPdylce2dp
kNNgqqSadmxXavm83KhozDcZtaWpU1DWfwxfLYO4hwzEUPd7lEsc7OQPHvSt2hwvZAU6qt++EQT7
DcNyh0vLaxvEWEHe6Z/KE3GkAfz7p0FiC+/AjZpYO0oRbx/oBZ4P+vF0HhyZ6TUWEvw5tjjb6bQy
S0oqUmK5M5bbJwHqZBncNKRnbYpzmSKTgk88AK7DcY2n9BT/ZEHQpK7RIH7Qw2pVnlRn72CJr83k
mFavQoKY+RNbqZu2fMrc9CWPtLXiM9ZYrN9ks5H3/N+nsTvc8gEU4BUUyuAOrDJgUawV5fBLNn/3
KCLgES2ksbhfCPZyNNuLM6DcTKQDe9RDh7R32n2B1fYokIaxJJdSvC9ktNpVtvtQHMgix9AEuE/I
xWCLAXnhBMKCrm32vQcuSzwaV8sBKp6IvanzZ0FPiNk7a2pWWrsLNGSfVP3nM2FRsy/YAy+x8rjn
TKixF/dYo34vjmJwAURMrSMigqyU9iuN6bus8wWpHICOkQCt7P1Nf87yTjOylG82QeQDcKAyyv9z
GIW93nIBp5EK9WA38Z5UDUjT4YIIICmlxyzn31+lpPTqQH3xRSGMnLwCFc0ejL17GgoLdHUtAd8B
lM29cmLqII8ziDzwPEH6BZLhzLTJUKSp5ANbwYr+DNB78s/CNjHhrNyxpTEWruxrxwVBGJCZ0qtd
jWD/+LSRIh2UO7PsKu5BmzVWPSGC4MyOZfD4KebOlxgR108uQV0mioO3kgKwnK2GhmbwvZW/2FRo
+BDDLbgbhZN+U8gCtuO0dP9Fb3urrBp+Og1m/42scN2VTgB0PSEy8eUVYEBo98PHqAFRxvkm7cOx
Ig8Qmwv1sGM8wibEc8VuasJ+mW1VfYjtRkPklIMIMwFAxDBMV9YSlR1+pJOVacBO4TNB1ujxrN1U
cKR1YtjEE1jCrF6izVoVt7dbVs7GY7+ZGnlkjTzF9Jt796EAoxvEjx9SW+zpsf7UjAcqcDDbtylh
ZaoXQub/SkRhlgjEGQ2o7MOwl57SkJRA/HkpBayboI2TE9la3o8CVtpRsKSlMq+VQEQsW/k5JycV
nphcJU3SOb7YPyxD6ZreX5cmid8q5I+r48L31MRzjJgX0IkZtDjXXIv3kC5C9/YgBTxR/9kMlFNQ
cSqds83jw2GL++e7PTjBPmR11koGzAmbIpDXiBvNp4ELxrUwe/e++NRl2yV/gDWKb9s2lkh7O02U
vl/cjTXVGsfK1HWVk0zBREGR0fThvpl+3Nt+pCJdaijS4/lHwCZF6rccd9lMH4c6+O0r6yOAaan4
uioT9hOHbCfJZgMITSdwTniv03npJjFDTgwrv/pzV/t0uiz1IH86IeNeBSqrI8NdkXww8QXoVacd
CNqL4vZQYhDD/zozlrehlu0RcEU4eaLWUvXOeVA+gFA1UxUYi9VKjfq2Y2VEUqvrlsgK+Z8rCIss
tp2SzNjH5hbwWzPflEGl79oBbmAYzxHagPkVvf2OdF+ZmhlOEZkswcP6svN7347YtyCmReu4B2/f
GcCJl8t3v9J0Vl9fWdjSjkV4qmChrPlar/cnGaaDPJbvJqT3zxagHWcNcCwUfHDAOPVJVHlEFAYJ
qUyg+iIiIHS5jlApyivyn/t5JR1M6Tly9XUhmcmQRfsf53RREW7GZnZumcO1wCbL/ALgMXPEC+YA
ZXWHr4L4xwqyoqPCS09noNhNEv5qHRgyp7dDgKxC6ylTi5hRio2TN537eBj8zN7RszU/TX7DFqYP
1HiwKCtXVcazFeEUgoAZT+q7tM9WnrMeY/JRsQ/AlkdlprFYLFqXN/gSYaX7gQmJ15LboFZMpuJW
45fUmVVage+EVP3mfw5/J7cT1XdQKesbhyo/NWEqXx++AgExywhMi93339vZA6K3Z4ZOCzPZK/9A
1wzKl2VTJWYUrYJDRxqWj45zu4I8ebmaPcTR6oqYKROGaMVKj/ZAyp/hvbJbw6Rzh3zAy7CpgPWj
4gHj5Yn+ODo9q9JCAgTO4LEo5RyHWPVThJlV5UT1+VflMzUDXH7uszcCMZDLUiIeA9YWvAbj7nhu
bQjIgX8B9RV/oiZG0nBNh1TML4wWzZlP3eUIBe2uEDNykkICO3E4e5007Ttv2ff8N16iX51jEUC9
r9cE2WJmvAMqrcr7cZHu8Rsn/4mv0KHw4bK269F5UBROZYS4QIWDb0RImvF/XF8ubABTWTZSE3yM
EpUE82nNj+pbeYHtLZnOIjTrXBjDPpSMkJUuzu08ZOPmWvKL6UDWrPzwIqRakV/v8dI4hg8UUoTu
GK9qaMI3d6HEVubWcylXE1cVff7M+aIOcOUkYjqUJHXuCMgr9rhxaliGWlJfHG6OReWDq7ls0ENh
ZzIvmRMxTVPTKxcat5j42pxKZzI+giclHlCk4Glkcni7CE5pjOblqze/yVCxE+jFY0KAYPS7n8fj
/KFDhFGq0Vhb/sPwiYzibkO3zyfi/5PxO85HKNwmy3frOHN8sSBbjh7XSY5uJ57iyhsDaOJaVZSR
+pdveEg5TKU6QKIBvqGrwENgr8E4ZkXnxq5cWNNbo20GhTD4sAFN7JRBvnpcb+F9xDSEP7vlTi0k
KqFYAv50os6Aesosy+yNX9Opj+pOKOk6llFJB8/pwaOqC2gkCre2pJK5MBJtpe6MJ+mQ5lMyfDWM
AVEZubXmjl/1thMmREYRPgmnB6JT2pcPgbNx7lalmXO1QRN6UePbBwIJR9iIBBdW26AW64BJZtfS
ma0NerkfP6VWCWrfarkKQvsaDxAHWg2Zef6gywdT5QsCmw+3IIF7tuAwdGJV+RYxGyufeaJtDb3B
/SBkjAfksFLr6S4JxG9mlvMkusZmZM8MLtc06WNIdX9/8sUEDaEPwzDIJLsfxQCpKuSKlq5z89al
UvG6dQXPlUfEOMU1oyr+JLxSCDDl3Rd1n2F3dIYepIxzpytKt4EdcuopT8k0Xe3TPDmDlZvFep6F
X/HAHjQtaciLEUtiXZ5cE2a9a8Pq2xiYMPSrEDpkR6+u0WHry0ZYUw3arWfDVGNa8cOVFwzEsVS/
KFLaxaIT12CzDnlpJiEwT48YGd5ZUNGMS6XFowOOBnC5RIZuZjOxkRV/CIFLJ35IQpqTTcUh6Eyk
yGYQR1r3Q84+ZwqBfO7ZR+xJUwq5BFRS0A1iCyOgqkwyo0LJsIL3fbSubPoLS6N0ZvAVMxQBe6hf
VSYYZ5pxO+k3WhR9Ftcx1M8gqhMvqTHMVzTxslrP2Y1xaL82K7PBYFGKoNHUddHlr6KZhS7t505j
TmMiXKbhecTCbsAyDSXfdKMILk817t37QrM6xVrW+WjohiMwFpNKubrPJb3fDnYzALL9ZDhTnblA
4dy2z9GJJ+k6iVevSSg/XZrZFU1gnguEdte/UgCRV7VYIHtw3dqVdFjKj23KjjZKY/8xBboGw6zM
bQgKAAxtmYluxCDqsbyJFyI8xKWOpv9gmYMnoNDQcAuGLukbrYwnPYYoV0frprN4QgGjuwaH5WYe
jBYc09iCDVTvawp4aBHDZRXMb6AqJxx3fEgfsoCnRCyFqwLa8euVt3UoRB9FUHQZpyz7sRh5cYkJ
9+KdPslamDndU6QbEdU9XXMrJtuZVKB/XPMOHLTFOQT2Wvka92y9CViWzPWLZ3HzCXpKEv+ni/jR
ww38MQMdOMXyWvu8D/s1XCH1KX5sCuteQj2QoK3ARqQ4wVX21fei8A226E8CHvwcDTlv/VoopFZj
17exaaJ6CdyvrbWl/FsIGB/CgfCeEqg6oVjdKMqpqnVxzsmMrP+5Lp1JOvknuVw7j8FoIRU3AN+q
tmNuD3sCvOQLcL1+AuorzdHNurMj5XdtbMt0yqwauZ08buvpp1xBlhSJMkcpOawI/qmWDBfulLFb
KAm5Jh80yakblQDoF9aMFlo5a8VVnH+LZ02FqzDP6t81gzyVQnO8eibXfH0CIZtHP1SPioJ3Ube6
zpR1gW0l7HUjMaJ/2+EEPScwi6qcBV4Ck/FSVuaDQCWWvl4wz5e7KGDTqVS7v0N0Gp8N7tTXBd4k
hnn4+E3kbljJZXsCUhLPUKdP7YU9pDJmd/lB/r9IHWdUkLTzcXCDtSRZ78RxRIK/+ms75t+iN4XI
zgoeHAwJB5wg6ccZRO0GfV2aS0OQpwwfgmLfOIdSdd0I3q5IWutZ9AOWfmSrakn/jPNr1Vf8mWf3
rORLXfFPDbkSFEoIFqoR89TJt0aVzXWlABA0XdZuh1ekf+3ag5RGzVltWT1+evUHuU+J5/Mj3lID
VlgZIqH+1I/k9tbIoWVPe+mtihCmt1fw7/7h7j6AR9TnB5GBUAsB6ttI51l1o+HS4ZxdsZnCW9bz
G/5dfm5bjBIkVE7jMtzqnrMT4gGJq3pvhN5zJB47glLz8u+xRJT/nUCVqi7fnH4BGZjkEoq5E+KT
J6U1FR4nJ2tngpME1fGgwne1gI0+lus35oy1LNbgG4vKRcUFaeHxgnumxIYofWzjVVP2X2V0g+G3
cREeCb2jt2RUBAZ87f1olpwQwHjMRBPhZVxFYDkRWGxlNGJEWFk+qj71BPSIxyCuxbKhHJsfWPJ7
g6tmuNu1pG5v03SvUYxmLhhGR+wcn18uv5/DHrczyNCrR0w8Iez+CQcyHRTruc5gEtnVuIzEsdP1
R06wmETtqxhREiDH4K81KNSgPBgoosG3Pld1GyJ/QAMtvm9Zaqb9vm8UOtVa2PiYQoBtjFi9D7/E
g08CHE6/lQ2fYPj9wgRiH8xtr9QyqQ7E7ti+ufvxJpeXy7rIxPeYOMW8TrhV3OFmO5aCvsQCNdTY
TdCfNZEChYQqa2BjljISkpsWmBpFnXXbqKtaNvVhMvqE59wva5qS3HrEZm0gWkZhHOfaLX3VB5IA
j2PIiwRup0RiYWtN/zw4kmEtQ9w7Uyybax35pEe/t0ayn3Tg+FLkyoMPCuUnB4nrwAwes5ftPVNb
NT5wceSUbdjEgdH5G+7oXSxZ3DpokXA1JKe/Lz1sOln7Yk7vdOc90Z82awp+zsoaJxWocTBt9TCs
qIr6PLymvK4YBD7IfwpuJgGozWdAMIx60e6ckpIv+d1EPSlyVtoHXgdbfhJrDHixY45o6H04bLBw
xrP5DKJenBH7r0fLaYOgh/8HEYihDdGyR/6yN8D45yFqzRPowuBAtEybwxEhLDjDzG9qjcdzcuMq
Ktq1+IVy6lB+ojcsthPuT5Y4pMeKElcBBvn3mx3i+HDIXqAggaoMUubKqX/TBP7hAh/DRnxTjtFd
9t9CaTKaK+e9lcXo2GcfsBq6ZV9KDgQPPnaxLhYRVET31CjVsRsyiYX34Tlx48CfY55h8kIyP8E7
gP+z+rweDLPClmNNFhyFN9YGSE07AbwHNFm7XXXZkR6s+m8PKWbQu6PfGJqKWmQu1tx8fia37i8d
z687aUck8UMd9wuiCWTdRJlWUnXqrobcX8FUs/26cChr1KkuAjUeKXFL3mWZXrdb5OOq+fhL9GRg
3zfUVHrKYsHFM2lDWpoUwJkFVRe1U2ptvWSaljd4rkU61XKULxtvsEId8T12mEyTG+c9EobCUT+N
HwE7qcz2Fmzi2t/KJRPNp/NI8WYl3NwqUky9cb+69+q+y3VT7/RtdAZ5c0i4YNydkK6BZleJwTcz
71gmOoPx4RsBT5+Z/gwL33+fSZ8nX7KUDC9wJ4QpPQjZFpGSmNPiZ6DgkZjEXGJcHz3iyPhhU9qX
Fk46V4z/TbDQVzedgOBDnnCjW5QB2wPveCyVhuD+9xIcM3aQsA+tcxpetURb+7lXRgAVJNWxyis3
d74Xf9WrajIlGjyCeZnoD1+mVXWd/4Z4VH+I7aeCKCIoV41RkrxdhAfzp1BoWSYmsxQKVG5hT0Qq
PMK+yXXQ5AzgBdNp4/4t6WKsnol34ZcGeDHE+PVqDDS2UuG4uMa3N1bfuKxLoMxps9nFxLh1Y4Z5
bKrMDstRTlaESj3xxJg4QRz4enye8zXKqfhK84QHTQ7Jv02krztlvyQwGTrdX1lVHJR4CzeEOO4C
wTqHk5gCweZyiylpstYIT9XGLCPgQrI4JrNpPKL4Ks8R1VOjuj+9fmMWnU+KoL51h+ztNA9Gjz1B
CX0dBq+fz4ENBH6LGMJPA8QxHSlAmwn1NlcXiGte+vIzx6yrQCPs3th7Z9yKQ9Mt3rJl8y0RhPCU
YaLUts0CqGL/ruvc5IpFRLPJc8frphXFMC4yWMrJKsmu3r3MrA10gDq9aaUqe/fR3C7qBYELOBXa
0KLbh0EAHt7w2y8LqEVYFR2Y0aNCOof35b/s9eZk7FYLx+fKuQoLJTV0e5FIiBK93c862ovPAra1
XAv7mxfZwwyrLttv4qoiBEsakAvLJHfdMPBaOo/3SAQzAJu+cbcmckQuLSWmllUoJhczLGj4KIWC
ttYmrgZXv2ZPMrVAfa1uEAVwhm3+NYdJcbXSscn7Iz3F6B1Xk39oLaCtKDJdcWn03yh7ybHeMXkk
sGbJJh9E9KMmmuys8NEUpish0QIhF6QD1YPd5+D8M6o/uKlkTRb/oeVsm9UM0x6TW0jrMYxdMKDv
ZVDBmRVZumErxpQnw9OOC01iAWw1S0ULbxwILutpxqDV4g2tH7TuPsB9TPNlWDlfsouUIllKmSkR
0UdhUwaVVq+kcPdwz0nEqZ2LM6eemmizXYuA9vcxuKT5TYQ2sYZ1DgnxQvxSxyAMFcPisTVRIOPy
IRZWyvKJtAzbzMPZuO4QvmN0jDMUkqoiECt+b6sM4l9jrJQgIyE0GfNsQyH7wbwbs2MrgK+la8Pq
gcGHdMBgUJ+vSgYp1QJRfhnUkuNPtp9aIfs4zs7QQ/LDABAI932U1pxKhQHI9xp+GccjoxWqhBw9
DkL+cDwWfZTyshV9VIYJOCKWb/EHz0Ug1zVXIyq0I1R7jJv1tVSKZ+onvclToKxvwCg38v3Giwy7
s3qSsxoBARTjYlyNCDIZV5skLAxNTXAiw2XxHUxbo0i/umUJLoOQAVjEnOZciHR7xnNhWpYaRHJg
tMi9tS24xYxHCLPuw41ezFuJZIgvLyagknYdUx5YgGMzdZiqTAVwGd2XpNpxfZ0GBJ7axCk+YahI
RlWl9ac1cOWFRTD1L2omDsbZxTzhnNiTYlEXa0e2QqcHU+3+zMAxHeorzK/uNzGEgzWD42+BA2sk
4b7LU2dl4y6Jzzloshdc2TJjzHRdZ2ksQSOQwNyxU2pzUCjbjEAkXGZqwN+nfvyNBE1L54hx4lhQ
6bjxJ4CWFK4LO4IW+F0AH1r6452tobWjeF++1kRYO17xjNxFIGxNcE4pd5DUHfoKajPbPNhG72Ir
WcKQl5DM6aO5eAakTqui8C5zHdJvZTSLO10W3uStvcXqfWEqmGMwT3T9NNjP1LHExV64Csg8krir
69dyy8aih+xmUxcTEhYjCheDZT55u/T+Na3saLFh/2sSwOC6nXLW0HNZmEZq3iBwSr3LkOl0niDG
Wj0tX4eDko5So5h3wB3/6kh+12TfJB4aQwX583bk3H2TdOyH4Aj6X0//2FUdMXqf7m2/eJHw7Oz8
KZiZxgZ+u9Ie3w70jf43ohqaCgRRtWef+Pz7aGk2UHLFtrETSOAgraLtgkcCNfTYuAUVcNnGYLDR
S5fBWpIgXMBYbFLuYdkpffCn1U3hbNRihsogfc25fdtWeVkuT5VRagwkBJr+f0NuSYeiB4t0jq78
+3ThywdCIpooA7y3cnVzkyzbb8h8u1z6kuWsjVgHJogGuRUuK+UMLCatIpAne+DBLawIW/sjbgoP
gnrcgsgapqAf6sXaRdFOECPzkaf+lmAvSnktxRZRWHbPH2ruN6O8V1qEo0A0q3lzVvW+A9l1CP/Y
hN1pR80Cc/YZljSGTcBjGUhqc2jhrrZhpxPYNQs72dgIHRNKsN5g1esc7uPUIce3nGu2Eg95Z9VF
nDBjrepHj8xS+IFbKnOcWlXXKMvOm8BK9Ag51Fd4120OxjCE1qHxvo+T4kUrYFFIbwLGlQLS/6Fn
0PlY83eZRnEB6jFDNB9Op7R9T2uTsJFwdUtDAQWtHcYZVkuH3gI4xlTSVD5ssg+X6akutp4DglQx
vMIGFkwYLKXxvjRqYIRklziBisxQ21IeLHbWsbrDLzdQFQNPsl1mg4MAh9Tmnl6RZI4xy809TCdk
RVReqZGwwVTi38q1oGgsMq4wxnCEsCS0h/P7+sultbNKKl/vH94BEDsHea/qHBIdA+Thok23F51w
emTWtIdcX9HZu7W8lB+mpWXVF4nFTtM7++mHURcBmfyPIlUDVwqlVq40uUSAI4VWAlsMzfsv8C3s
+iSXpl1dSokjO0Vk4s9Lq1F6KjKOfnsIy40+WNC39DwbQSufmbG3Jm+HLryp+hJ4LqMyhfo/PCt1
UzWkcfbSCtr+UohED0dxRHCiAzzfjZLZktjOQWI1afMHhot4JGIXtZRZAneGP7L23BLCkQcTqVS2
u4EpKvCq/T9UY08155bZ5+4mfDP+0rwz5Xab3wBytRgNfoAQZn1P4C6XXw30l3Y1tFiVl0EiTdbS
XOufU/rulutGsVxNNN+pB2yJq1JyKSZ22DfHTgxZ0eEzgRCsy4PfbYNppQDZfy+4PA8zS/1m01MX
aRXw6XHRhGBOgJMryzmhdB1eZQPLCwzzabXvr1P6wU+UvbscaCqpYv9YZWjl/yhBcl3s+Nj/TjPd
0lM9hNFNYGbn2FklevpGGL3YtX/QFczsB5DsG/GheVFImMw5SjtgXOten4OJ4Wh/6tdRYDkIjFQ9
L9aEGIFvCtvRnz2DeSeFtVE194aNMM7DhoRkT6VGL4fF61kLP9O4iEWJ7QTTQfYfwfAWnxfvF23c
y2KUWNUBt11smDVUvEpB3OscjQm86i1I46szmbW+tNH2ozOFrGKPlF2LuBAAod5uDwKn1jYeFMIM
kZsUGW5gwnpJKxrGYNSZfKIKY7dakpce6ijpS+hLNrFM7lPFR35f9Fmlu7lv/VCq5PHs1yg1R4DT
eIDJJXO+nCGvrWyh80TSBSrnWnxwVGQ8ySCit3b7SFUEw768sw36+3kHMjMUYT8uFt51SY2biPSk
r8k2SLaYgunp3U1vfD2xT9peQdQ0dHh9XPzt9+DNNH11WbtJ6AaSjKiVLZeCHzNiHntvSlFRDi+6
7lfLZtBhXHDOWOKvYMD4iiAadf+P6IfCUl89yKJtgd8fiUj/FrnTk8sCXMvJpT5l/29490L1wyp6
UEYB3CQsNtrwGOrZCdb1vf8dNNpxH/p6EeHPaVObgwS//kDikrELYUxMp8ekTQLg6+baIBS4HL/4
pHqdBj0yNxUbUbx/o9EBf/ZOLyQVo0tRyTziw1lD6J+N9wL/eJnitMvDKNRuPVGOBqTNx6Wa/kQq
tPr6a4duGXE7blknsLWai7Sft1X4br+VEUrTuRIrnfHC2PQTJkf6/N+BVOxLg3nQ7VcwUuB84ekG
9/TYRq/upjmeLW99TtR//gF6fH4CEBaGDNts9xwl4M3+banAqz0ywZG9EuRTSa5H2JydtbCHUq6z
m61oNLR60aQbmp1UKmuG/+MbzrQfTnwyIcvu7dH4Oa6OiJOQGYgigsQGMHlB4bLZ3MvO4vUEJOc3
pS8PXE3a2KKRTZdJga+EtdF0o/fi3/2JvoT56N5NWYJKTwgocIz0b5Kc865qnF/5Gmn0yLfPJGa9
xIaxtdzlWmG71xyLO+c+9lgT5BsMtA/lO/AyRGwYA9/83Ypf14U7ZcHcK8hg1QsJs4LK895GRGFz
FHeJt4VxDzWv4JtyLCTykisoDuzj+tV8wnkChSsae38FV/pdVlIuhhmuq328reji4i0+hwz3BWc1
CldFF5YxinJ7Ux2wp+EYjFJQKO5WNtA86p08yavI82JRX/heUM3IQIuM3OHYCq12mfZZ6oLkt/AR
JPnElT60Fd1lj7MRQADbdoIyzmnDjO2tL6PpDJuxyO/CsBAjO30Ee+TotjzevGRpXHFYn09/IOLd
8yM2YeRAUdgMo1CYP4KLX8B56ChxnxQYtcWUF2EJkA9hDlFU1lOOSdGtaR//Gj3YQxyS9u1rw0aX
r/FWydC5btfR3dfFFYHmsfywbRo9esWwXGBBXRP2W2JdUTKxk5EeDs/iwsRy7+J+QvB4U7CgVnGZ
+iKwwAM+v8iSpae0/O/iCdFD9QjC0/BTo91MnkkE5Dgm1uBc1mgpmDzoVwWSu8Ni4GU/FW4NpfN8
WzImID5WaTiP5+NPfnComb68ULsNhX1uCJX55JE+Guz3R3UtuLyjUgFlqU8I9eTxzCLAIVHcJXVF
/1NpBV3+ac7hKtXUJPkfld/eO1oPEYeZVPk7Gs4UK0yQX3qkc8mIKZweCSIzRt83aROcZhp59nvI
f557jjb4GxQhDDSegTHGSFOuNFThTXcwDtt8y0vb2aIhqHMDWbEQcTAiExbXU49yyIBdUeVvojRT
islcDKfR4Mqrsfs7pw5y3n0GR4MYhiBViEw2ZPi+y0Ja4xZ3TbMGiwyEVZ9R2GbmxcUSjrdgObY8
/3H4DOrsMNVe5fThoeNYb/2NNFX9yjzn5OW5Np6lSHXFo7mz9G5URAx4xp0gaj359IYe7OyoKqY9
tU3xkoUXMitwffhj7i1AucRGSdaRlWct3QtKBJwOvex//dLbr5ncdCngo1RN+I60GM/XXLBAODmy
kfjIzV6IRdvi7ED0l5jw8EVTpk9YchvFCVboVTE4DgR3aixtg4bfsAaDml4H2LOAsP0wxEaejyJc
LaUoZpU4VAO8f+w8bIQd26H05PPVPawsaLGsBQnoGE+CchEKoATRtA0cCu6kBopWNtcXcK4F8VST
QasOrZe9YJNBz4oEWufC0m1tHdXfK5fB8pQYatyGLrFw+F4KcFC+FbbifH8XRoEEis/XIl/6tR7b
a1qfdr08u9TwT/kIsZN9zIEnyIUHQr7wfkLH4vzu3PLaIQaCEu4b9o6MXAoi6vcFL08rqyVzXNAn
eVNVdEU88SF1pYwtaBSCgbMSqvGxGsd8Jc3nZuLGhbPbeJaDR3uZ2jqhcrChEzuD+SFh9yEFGBat
Tpci+/ZBSQw+VXMZEXf2pt37ANgjxJt+OI/xN2laAK91ez5VvcFVLOwU4Vi6GI0xbslakpqZvsGL
i4m0H4Eww9z0Qc4g+vEG2ZesEOV1lIH1D4kopiajNJgYp3JeN8LMYZobLA+NlDNCGs49B8X7wf3N
lU85ZLQ9faUzNeY3Z0dP+IYgmYsV/+lItWR15wjYxLBhSlk8TVBvLZcu+prtgdGcSpFEbmEHdD+g
TLIgWx6XTdTIY4IZKI/f5a8sjGco0YkPZRfAS6Ac2l40YnwzSNcb7VjU37nA+tNNO1bf6+uYl2QZ
DToJLyejX5nCxr3Hsj6VgTKfTvAn8EExgoCoAmW3Fakh49z3+Nw20OJOfur5UCQG6J9LWJlmQyzG
rD6LOgD1hdHLOMjAdVopVP4SWsDhBagIIgd9sbYXPTj32Q98ROGEEr0ZdPxqfGF4SxY9/qQG0zoi
S+zmJ0w23RtYPbinP3RNyGDuP5gGcCj5Ymo6H51TH9IPSIw54aimoTAElKfWi4d8gv7uUBMyP4Jh
GATXkAWQ09XKX6m6eQ6fJqNywWMiZ4R6IkxpVUnrcyGiZfQdwCXEN5Ell5xMELtmmgt+bI+SSLiK
WsaM/2qUV6C6gwP5lrRA6VXL1x24Oggm+b0mwMb47sIeWvZXO0wUFodmqFcEJOvuaHONBOykjftk
2NV0JmZVrfWGPXFKRdt3WpJD+WhQIVl5WHmPhHIAAv+OjTQlVGUxAYMpm/w3KT60fD6LwFK/U7Ly
9WUkksQNUiWnzsNS3KiXztDPhG7Td0U3jkzCuqI7n0V+2V0FuqeVYaml2uOeCPL45NXVGizt35cy
ojH/YMMV7lxrKUMOqR/3JizZkWH6Wu/2EVFxu5vHtRl4M7SXszI9LM2MrxEE5B8lbfVMsKUQGqHd
p6SIOgg8gZtu4WkDX0qvWwstajZOd1+KSPKKC34C0UfVclPPuAEYfGZumMXeE9FDK1YLe5WPBA4N
8sKEWzn6Z8Ko1to9D4lx36aZ4LYv8r1US3ndxkjtQBh0W3fsOZWoQGqv5AEwmYy7+Y0QKnwjGwpl
kr+9d4zPtHa9VSZ5AcvOZtQgh6w0+21fqAlfguy7jS3R1BoIogVHPYFo97LoBJ2UuFgszfT7nCah
82Xhhz0tlgMK73ci2IGOu2ItgNUTokQOwWdmznthDRFV0DXxNohzTr1DwwDQhvzLrUgbLLve+a3m
n/SBHk1cYR8t2kZ5KdQZa6ac0Cp2OwwHZSZe2nImmtHISNv/Wrweiahp7qejVHdwJaW/h30E3nwr
dlYGfD78gSxf3fJ7pNVOsFqIyJQvrBLRbRp/d/xFyUEwrJbNbcn/x+BhvjKAfir4MVGFhbOF5O95
z6PMrShwK9cORuzPg8xRytXM0AEEc7rpPd+J08CDzuMeJ8m988OzYuCQj690UoyA7EIsY34DHUSm
K/sHom+ySMokCMGVhXTw7yDDze5/UByKXzaIKwXPNh+0UEx1q04giZi5re16U0RkRLTdQbYbtx4L
NE4UbtLJUJg788srgQxjKjAFeN1sZLjNbxGYwsswHQrDv+MY0nXbtnlC16hCBVMUoFdeWq+UgStc
kWAMTwHQVyrwuBZC/nJqRu6fmQMWj1jhsKKiHdAOTnI3jW4+JdxbtHOuQV5JMpHEXzscNoI5RJKX
N/7ffjhPyShifFfJgAhDqwsnh4NExCEZLhzwI49+hJwk87RHLbHRPhy674KGOlKELnP/8rz3Zpkl
ATOlftZr62+3C7qRTN0APM57/1i90gIpmNAMc2LYXRQ/61yUmePPfVTQId7QZiJhbrWd/sFkJoCJ
y24KDd2JWQx1cRWx/KriD54vOn36OPiqaUSEduH+c+mwtXNAF9EJ7SvIrm17yfEgsIbVe23ev0/D
Axnv0qDrcqQh8yp62MAP5q72l6slnum3WR3T1iHBRRjiK/SggUtqYUWqzK8q3AZ3PEFGINy3FzIc
8KjlSIM2txXAVFxHvi8Yhgsm+bFTsj66aDFyJIOmUk1DYs6xPij3vvPUIRSkahAJB1bM1saoY9Bj
VATD3YT/akPmbIIJCOwA3aOCFzomgxiBrYWLfjSzkPhvv2qCCpBibEFW3i1K1EEIg+FTq4IgPm1b
coTSLewGe2wQWzP0LmuU/HSpGmr3i1E/iOmhWNhmGyCx1lMlDRCbrVoH9lOZgbcJrrdwVCBKq0b6
puJkkh65/ugELdGuDT3ND6YTe7BlrvDS8sVEZ04LhJ57fPxceMW2oE39+uVlqWozH0BGUzHFE1Hh
sdefy1lmyimRmHfEmz2nl1YwrTT3hOzrI7hPhc8eFR9AxKUvhGeT09yHF2RyHqCfXQZZlRdWNno+
ZWdgx9QekrS66oSEOaTIEGHcMS2Ee0BEldC6zorNQcaORxVaRTkl0Z8XkDimdauGBeL9tkRuvJuT
NB47x6cDx3Ro8uA/TQx1PmAODiWBrnDQxbkQYnUa4hH3X9cPOJK1QM6IONt46mRAgBIp/iYMsiV+
keUR6RI7PT2E/ScVQRhMzpuMjWl299XhULNcJOSEZADCDhE2HUlLCPl/S5jp7GYR6naW4qR2FEHo
gcjjZuEZR4xEfGDUyb9L9uMvHwLy1R74dpEfPYrdcX+3WYFSISoyaqA7OjqaJrNe+wjBRwrhWJim
YYKskqgEQGDeNGr0+oIOCAzPj0T43Tlt/ZsR50yhN4Zgp8Zk+rmCKU6pT6+Mz3P4sa4CpQUxCO3Q
i6uNoGHqs+bpjKzZ0GXkc3YQZ3DSD2i0iH3B+4qwPdXexlEfvD3J+z5BMVFsi3EScq505+E0/xgB
BYyUwLNveGqdt3NQoFtp0UviFsXI/sakCejcq6HOywl3ri3TLJF0HgotQHaYlHm0i6F+ZfgcO8M9
B4SMflpnpMUEHv8xyDopF5uCp6jYsU3TzQAiNH7h2YIO8DpFH+huedztX524KmuGWH/sGBCCEeSC
9txxh8WyoWAT/xMBJibPcU+KxF6v7f7qwOCRXRGIRIMUu3Uj869j6HE905V9erzWYAjBpLVzgkuj
pC+n9VMoiSP1ifpuZ0CE+CEqcNRinVNEN8HqEVUR37STo4cnJ/v2t0DTJj0yTedENUBueHP9w0Lu
lZmody+06tTkTcphnRtDYShLK2sMZXlzkcJqqx3ds5xUH2MK2eDP12I7BgKgiMT29X1M2ck5uHbe
CTIiy5qWpLyu7YovUqKd/BMzws9S/PrsgnOigjSl7ZKtiUuF8C1lMI3dy2JcPYTJVMDUdAG3YVXI
ICBp6qF5B0olo6CVY/+uqbd5wG0El2agLzIaFCVoH0H4CvIdS7UA1KseEGYn2o6BOVUqDb3g/1Rq
IjEbkdv/jJpeZZFxZddlNBEpWA3q3mrORBdtvNFUry42zevcfnTM2+Yts5pUPpkRKFWK0yfI+i4e
VbxtCj+Qyghonwyo027yzKKV4E4k9/XxMsnadBWKvvvPkcgxD55Nm09qP4WQjK//hpHnieDoOlqQ
01x/udgpa1NUm2v6SSRTZTk1m1HJdq0ArvH+mBKnS9nPNIBdWOG+mVin8ne+GRKjQSHPRdycdXYC
pdaRXe8AJsNSXM+vj6MjsE2Kkr4QTvGgMs4qlQtuWtH+ygBJBgHB0GgfJ2UT7nX4B11v3UOP86gD
nnrOayou7VgMJAX39GlFknANZwmyw6CMGdf2buAAcay3tjA1dbiimAKgzEiXZURZYpFt9/KsuajA
Wp+l2saGCvR0FbTR6z/qUC/nDJHSuTqVjDO9MhpIOo3dkWOi12ehtUfs+AjOZEkCQmmA7JP1xNrW
IDXNlIkR9JUDhJ2XCmawmC65TzjDlGHS8Sp1Y0+WNYvBfyp2WJJk8isA1iSybqX/+UQTkiGpy8jX
tIvh3jkQRjbSnlTDw05UaS9DEIJSghWaC7IoRRIj20tfR2CEZcXl/fURr7LPNb0efuodbbS0JhYx
ogrDmLCwU6KqSS9lqRawmC2n1J+I3/Jh+Sgqk1FYvBq5D0EidXwUd1IEQ27YZvCzcSO4acTAYRUA
MV4Sx+kCMMpW+aczbFBUN/o0TKVDKGvJBBmxTqt11FCpce51ucJXnqfEr9TJy4/Ya5r7jzcRLinE
wdIwL7QxYkgUNdOedTWj68Ul7QNG+07PTYHUHmMX+cs+W+RbPjiM2z42VVqYSFpeDPQJKfnJE7V6
1/iKIO/yReT9QXjkpNrGaIkkR1tjvADa62vgWjfX19EyPT5J0scL16HZ30sh3wNZD+gNJDO9OiOa
uB9lM4GtdTV2xWfc1G54j8L0DHFePQFyMCXiXsZjtv5A43dNptUUpmMotVZg9e8aAcmIIpWVfQfD
CxWzSA7srlaY5fPCXtB1BpEePASGgRWDNoXLa0jtm6Wt89XOW2TvIhCLjor6rv/HC3dXX/6JG9hf
vRRYiLhvi9ND513ZdK1p1DqCYdcnKVmaQywM3cDCyfjLNQ+jIfI2DiuctUfNPhCdS/ZqfYSRjEet
lRvVwtqgMJqJbCnCPLshmlur9KkiEySUPygiMMYQRZRp4dsVJi1aMix3g9j9b3lk0xHnbE+KEuxR
PobYHeSoXoyLuGbzs39c+NDW9FCWWorFUoExEghS8Zn1Gx1R6/FOds/QHgqi8Q+qyLwGpyVe5R16
NcyxQG8mdbE2jwefnR30mU2afyKryEOpzg4JHIOUzGkneuqye9qbNL9ahezzjGGW8mDXbNsR1Iho
gKpglPPD8q4WiOjmUS2fAl19lIhGkF5K95/XOlx+sQbF3AVY8Ls0pwAjWzXveG8R4jslb0ruqVCF
IcreU8xLJOtgb/mAIldmA6Jff+GAwxNbQYi+CBI8AL8XM9/l9xqzx2j0oqzwJBKl7c0Ddsrn6Kuv
Z/7dLFqpU1Sm1hIoOTw0IPGO0ITOZ433dDkWRcdDurrGl8/vnFLdENEmrn1oBVKfv3nO/+2Zrbz2
M3Y7+5U/yL0myGRmC0bBDovxqjZHDo6NPg+WShrOoHHqBUyY333SKqThGa1kzhA882uSP5G3pyVT
qx8//NA7gE+8ZqBcwRlXAqCXcHiWu9+P20kCT/wqYOEQL36/wkWz9mFviS87zJNaCGrcAA5ZWS+i
jAziJuh0x2vuXNmJTBrAvgTsVuTAY47kQj5OAlgVby/7chMSW4hTqnkPzoeRNf3FjTVw14xW4VGX
QvSJSWfuIFAk46EioimQ2lp1nLlzCrbhMPTL5Ry1UWjsxz1LxwEdRi6PPfRY3g0/HKM6uves+BUn
48iAqBCqCqO7WXt42z3F3qOz6yK+eViiSwrDJFSKqXZ7ZI9iaG8o6NGjuG6BcHSkO/oCtR919OzR
HiSgNQGv64wB1pYCBLxn+8y0wNB3HWzWSQJ1sHPnOQNrfSA9vcKRqzSvVpWcNksmZu2USh7VFSN7
4A7PZJ61h5OMZo1Qlp1SRGmdPpfLroJSw+2E5r4VOsLLEl3VkIgltwJ6KViwGBIfvG064Pe+wO3U
WzEnO0/gbmrnMTJQ9bnLwkaTvNx/PNtoI7R5wNFLUy1HKAvj/h4lexHcmHV23vRWYMT9KS2aghN7
fj001Ji2EkqCrMvIU+fx9ZoaYvCXvMDqf4bkF+M1gYXnMoFOQ5dX7Vy+UZpCEC6OXQjb1s8mLKQT
o877EPlmS/LezFmisxya0auNeGEp5oELts+1A8FRdBSNGNBDk3p1zFZ5U25QUW95JkNAP/H4M0qK
fsbmffBEnIKJsuw+c4Vf/WxEkeChV/R33lNWBJe42hFv0oNOeYKs2DQVVEbpBRMVJkRaRDrwXYRn
e4Rdeq3Rl/EbMLYoBS75IZmaG1Zo8zUx5Axf4+8YjMva16D2RL0aYVXKNzvfoBGLG3onLcwgVoKw
X8ZQLbjaCzEpOrHOdR0o5Cc4Rod5qe/AMwujdsY3ZQExboJP3NAEjqjQQQy+YXd36HD8XwFxcdu+
29TN/tcK3TBrC84s3i4ctSeQOZ+U31O3K6G4mWBj3wzPYhUvUvLmGqDZsljtyhPLLYDqbTuxNwZP
SdmvI6jdGJYxBGtH0jVkADpB00z+j+nL9vo8luK3rNakIoRbD9+1AZeKt8opNTS0h7z0CWQkop/Q
i8s4M2KsHqe3faMVIZxaT6w2aM/Wykoo5ANljZN2M974z2rh2xl/heQw89NicrPuPTduHbNHAbrD
w0b3oVR74TKeLdTYorluDNU+fdpqDHo2yCLuCA9bNBrl5XtCwk0zrRXzLpEJGFopjAaB+QNb52Ms
caHW7pI1JtVcXFpCDA0WNXigG5Oz9l1c4FvZyKIk19C6I7g4l3iCh1f3l8SwV9hxIt4tIJD9WZCx
U11wyPaxaDFsHgVi9AChwU5RxismJwz51u6y4wxfi04NJeycAK5AYebz1Ec1GwSRgdqchu/z4EN+
InsxOFJqqPxBgkSzS5+fB9FduQESBOc3A+LoNczoAXRssfy4ZRBN7R0j4cPBLHzM+2gQ5gvuwesW
ggq+0MhCtyqtOKsVAaIKvJ2TP5zg1t8KgJLuI3nWHOawdMhe+ln7Sev5/WeQmY0zWCIiRbsWw2Lh
Nhtt5Jf22w8tIbULqn9zxce1+jZXigBTiM9b1m8VN+ntT4O7ppo1zuo9FPq4spmzCnbx8DVpcO3h
d8w1TCl0Zs8wuZmsgBz7aYXNJ1EfDnaRw+fmA7TYtgqyAExA6QGcQrnJ4uionMrfspp2ui+bvwzc
BFP0KQsFJbjNAwveLWAjpSyG/k+kkvFOLgYUG1NLfQY5cITDptDX8zL5RII2Tnewbiq3oRyuzdyE
enmRH8bkeYY8mLojiIZjPkMmrwGW2q9ctTE5O8nvYIU4jgYzbhsHrYSmx73/bC8eozD3wqs3GVSi
YGv/LPRa6/9AHh6pZ5v2fUdPaOaZCfSpEvMWnMyKRJSyz8x3EAcTPoqxQuiucG/RT2Ux5hydzHDX
kv5bQ0nb8nX7qM8Dmhoer7j9HKlZNNepchrJX8lna7t50j4a5+lewE3qqAxOZrwwGZFRmbNALFXO
4JjnWjJoQR+kBMSc1gNoRNS9sYxaAmZcC69k4BpTtbeZOOXvPn3HFuLxQPm/z3/8TvGhe8yvFoIJ
DzmIbjE4BqyyqzrgHp7Sqwe/flq1y66CDPcPQqzMwWZiKEufuLtzi9JEv7oyFAtyHdg5EkjeACSm
KQt5oLOzXcEAmiFylASnOZNqWYQRB2+nS8fqhNS9qPhUcmyHY1dXwNr7ectr/Ub55HwR22Cm93NE
TwIgEmGXZhPH3iNGWWVjS6mYiqwLeHLPLXXSXQDpU8ihus3a+UUGAWkw1TAcZFB58vySxBzI8MxE
skDbKARmKJbEYxyxCWbTT5+OeAnZwq1eKhU7bEcCNwVJGOiuS6vVfN7aT7vkvx3v7kCU8bpexbW0
tanhDk34qocZzgxSsrlkEBdpaoavZYnjHjRuMHfLGhugSItJQ0JMCIDtub+fRfYEPZd3cXgFVv+c
GYtvIHpc2qe9MeIWtFkWq4gjcpvxXfXS0iKywvhi4UAOVFO65+fj94fsDX46NxepEWatRckgJ2dc
m89u3MV/G6mUPMIbh0TAXggF9nUz0BS0Y1IPT4N4IQ/F3jFdVH+p899z/4nIxL2J/6fRWUwpg0b5
SlNwSsR+WfB4ey77/z3tZh+KX5wC1OW+MEuQdHKqj22iXXWzAeWDmFvEAym1GAwOuLscx1TrsFUE
bZIpILigYTlSs+yLhp0NevIM05VU3+FADnaavusv63HVm9p2dw0uajBNO2rACOg+miGFedYtp4BD
qTCMgUNQ8/31qVNvP74GpIM0++jOLjwaWeqcIN2x+9bvJ28FBG2mwQfhshpAWim0XttcGpHxCdBT
9NDBjnW3SFWiIw8mL29BWpNYOiTS8ms6j0VRJHIt2QQp74naS9Y/nRu2tlaR9uNuoEz2zx38Yyfv
ZJ917NEQKjyHXr+mYumXXt3svyGAnvTQ1vICRyxrCkgbEzyrIo18olAYmEmxtXx6lZBEh5I5jFFW
XIonjjJ1G/Y+5g+cb/El4kNRKmYLGmcbzETIIHjsZTmf6nv973JBtgo4IbRmLQxqoxPGbGx07Ugx
X3o1UImTOxmo3+XlfJzug8WiaA5fG0EBO2IQyF5A2cTZr/7Vc97/kIDIvomBVvXuNyMczXQ2NC82
Snj5VcQBBdpUao3hwHqFFCTfT6B6ejz1um72ZYAePJRBM+YbHp2K1nQIQoG5fkHU5zY/lYOWeM9I
4zXT+J0QS/jSw6td1x/JGmHr/05s5YUHEhmOSR2opmPSteWw8CldGRf56BV4U+MGmnwhde7a3Aml
q0JEwSL3VAhEPvsLa3UdOqZta2TflsdQLWzV08tTT92BIISPuV0jDUMng82xpXaY1wrgox2Di8eS
K1EOCVd+Cr5UtFGnJ+63MPw28ieriVapdFDu6kZYVgmmPQlRLlKhku+wIq4QSaObngjmXR8pNsbV
1bzQAHuNeXZoYRf76o5pDvPEfxU+HdrBhPKt8cE8QBHzfLMax71atV/J099/jOzJvRhYKXdHpwNh
p0HyG7Q6UP7SFLMSqrbP/v3UEOJahBp/qsuwWLcEd2CMws8PtcJTDYVg9k2dIt1yyDfxe8bT5rm+
+4ynwLmBvonwIoH6H17Kw7Dwlbe9fFznevQNFTHq8ZVM2Y6LlCNdM6f5ntrHNqWRG5lIlCkodE5A
6phu6yOduQBTSCDiXKJMSgd9vxBs+H1pBjbcmtUOelYg7IcLa3j//h+i3hhkQoILM5mm5Mr6HHh0
ITMNfFn9a7+l7qWoTwzpG7w45U6VRUISXBf+FYFfLBIEyd+Pk9Dor7QCbo0K7lja1/VZJGK9xu+4
ai5CivUI08nCSaUc/51l9sLw+yiceAVZo9OeMXQMzLL75q0L2i08sOHt1f7+xNWy7gZjM732SfSV
iJq4+s3ior1zeyCy5cb7dr7z+rPAKxj2zc/qGJr4mZSOAHGC01sthNan27FgzWvwdpUGR4ftgKMX
OSuAAnGXlszx14WmhFjrN3hOh31VbTRQF41WTTUQzlduokI41OqVqFWtlOGbEJyxOZERn8t+se9s
CvrpZqE2pOjFZ7Kc+NYIpS7olqp94fQRgAXbO9D4dIqxjTiDskvHvRLezI3h46vUX3xt3utgvBIy
bne183Zrb1LUXSEq8EABeyjh4V3iZx1SIkhK9kQWQkJPKuhKzD2ItPVf6au+gmLLwUwjEUUUIjIB
ASb3YOFehsYike4YGqNNXgKJihYH+pVkxZx+yghHx4Ipgo4NyGo/2ZVJ07a6bKP6zl6D4pHLZ2fW
ReQAMtE0By2iuoSdr5UqZqGsQxlsaH9aiyJ4yhHUyjMlx09jZNrvaSE7SxGA+zXXN3qhsF7WZGFA
OKPvTEWR2VrmJIbEh5mxiq70RVCKvudHw/cLXs+F8iTjUeQHpuBLaUE5T/YOevBgi2110E2bNF5S
RD2ufH57335zQ2YiZvmetAfKs+xiqtP3qu++EcBskazu7WeANpSx0226MxPnvdPIrHIJyrR2l//Z
EYLoEuAPh0DaeltNHewtk5mZVWKloRS+3uzwKUTx6FMPC07I0NGSK6cB9Q3qd7NTNE14Z7mI89qb
BWeHhttm+3h7GubBvBE1Wc7qtUhJ/dNC3zBJJtEGQAO2v52siIVFIORvkl6c9+Qr2a18zN0ATgho
nQgv6ylTETooQNL8FIMYRiuD1n9+Hxbdob1/yFCx752F9cfeYzvtE+ltfRGBvSC8wDSScG1Nue2Y
U9QncRGFJNfI4faFm/fjx9FzGhBgt6/QkBJ3ZJsqFuANfSt3CQNVxecXfqlecneR7mQ0jhPMVGJO
oqmrFaUwE1Bbe8wUhkVQzPEqJhE+D8psJ170bE1rtxc1Ynhnmv2lt+ntzD6Ot6IYagwjdGUyJUHu
Bn/4OWpOQMTXsZTAZIJBCyQiOeMo2Y20LDBOI8ac5GTiOe7TKIT9/l5wYScG8/AreyBuxSpPqdwy
e4Fvxzao/SmzRaaf8YYGFmKiV8IhXOQijt1VUvKoCukNVPWMOPOGOlpRPtwO5Usl2brs3t+rxmfv
DlEbK/GYjjDZcwMOUim+KK69IJmYp1o130BA8BhxI69VYa6IaFTulw7lSb3QkC3HTB/zCHELeN31
7s9HjbmsPUzhoAytniqfbR9Ad3Ef+N8jP+KLkhZFYhSV80YIvvk/HwR5qBPqpuJ8i4zUru222SAS
z7l7oOHDx7CtDySyVbrS6uiiKIJX21GyqEawYRTYM8Pn7Uo8UFXBDJffOPLxWNFKaXhENxOMVsiR
tiibJjjs5WU1Cp2uf0cvjwEZMxhIGiUpQ02LPdSE6fVuC3pHHGzKnSJlQEpy0sFcOpTwChJbmo3H
PGvXFunKyGnm4OOAdLLDtxLBVu4vKlYVIse5CxYFbaAvX77ShoL/eBdui44/DH2n9XfSu3CLEWbG
D+jbJzBCwvcUqoPf+H9o2o7F5IWnl6F4sCYkbokzjksoAMuTcZ2CvtcVMxaN66MhLekV9wQr/+rv
DzxsU56dkbPqCSURg6H9Ze4d4lEqfgwy8yzcQqjobc5C9VISaSf9+cl8WbGs2VuUp4Ebg/XxY9sS
UOn6gMe+et60WFajTUr/QwnWPYYMSd7uvOb2+kmcMGBaRz4D5gzeKovmlR6dZAEZ/77w7C8SmuiN
GApZM7w06VhajiNT4oDF2il0ArmQQ4+ScMj702e+i4KVjJM/sJiPyASkkzwjm3VnWOm3NkF4hIo0
2gS/rXwzV1Znx0hsRIlQf34EQd9mD/ytDUeCWRKOjxCBeyMpt3Vr52TcqL9KMON/0HKuz19quWp1
RJLOM5NmCR7CqWAYyA6t76zjGZRrSSj7rpXVogbr187PIzv3hZQMhE1eXFEOULGxHxIS4oIROSFx
CkFDX4DmcsPHtKuDlEPfqGIwQnw4oiOE+564TrBRE8NIrfLO8IAPY595JC/5MevZlFygQc3ntvIW
WnRv9jRQscm0zfQTPwrQRuzUEMOF+zfBxdTDODpzCR2G0VErPJdrs3GGSP7/ufnSx3A7KH74usoY
Hg45pjUdO8LL8ALEQEk37FkZHWRcs1zMrVZSg7/2Yq8xPMmKVH8CoJ9Ik/KdgFwI1xYJcvdAIHpW
PfhE9Tu8psqyJeFJDpmYJ0DDsklB6AY4YvTYzI6RIM6Id7MImu8vOcaN8zmsoWm+NKnB+3WvTtod
PWGdrVFN7/uMjdcus7MycYRFldDNboK+/GpAvniIaVrcGe+8dOlRMCZ+gTei4/8mZptfuZMecY28
kQsDA6PvHbUYeQliOyjGoUcwvTv9L4SZ2+jq9pjKgJjuUKl6w0k+z71F4mNP/wfEPcC7uJz1s1O6
wucVpHwfD2511gx1ODDSvQCB6QxihgiWRRDOJubl7KPxMcckqSq5DuyAAOSbU+dV1iHZKOUTWC+d
VaTiz3sib/kCM5+4gqi3Pw3M9kh614Vu5JQOfFcQtP0t7TsqQOo+FBhxF/WWWfZ+RQCpbeBWAUP2
XRcrTsDaDhlhIC+/4UjH1fHKl1s0p2lrmcQn/AKKjQmebp2x7EWuO0eQSsBApGMPX1CQc8SvuFFi
HYBamLJdp6ffHjCM1f6IUy6o5IyJD209RHwmWHyVYT5Fk+3FuXAVmHqWUnU7MI3y1JNf7SJ8iAI1
aOk0F6gswEqHWTCUap4gHac+n7XZxltJSdm88FjHSQ0IZ8CzHMmyPaIJQ9iQIdzUS+R2jS7V+prc
Q3NhC2yJws60q9TiMbxFJlVymOhigink3yhO7de8LlcKvNpu6n37AiQ7TVnu24EB04c05nLCkHzU
Neco2d5NqOOcgqcP83UdBSv95RPDrz1Pr+4tPWiYewRSGxpaZAh6aWZPU7e7LP/CZd/D5KROGJGW
lOgaTclgFmeNMf5csqoDDJjBcjRBEzrYHCDYWMSw/KkDKmzll52TUQdYqd6pAJwc5o6uYyWUOWD5
JfySqXVAzbaMMGT9Pnkw40PVUkxUNNP0hBjdstl89f9rFx2J4e48FHyKmaBTUuc+ZH/kuYa/Q98W
KeMQmRHOfUVD5HPvlJigABZNFBeJWKYdp+QRLig727GnwtLl11OXCqKCCUMLpBk/P0uoziGoflCX
NGs9YOrQiA4Hzo8y0B/DCzIm9r3XM6XuIi5O9bLrDFG0oXOP882EcElA9zYjTIF/CqzhKEObHHgu
+MM3B+2ANaCRcn+CJHOeEY1GSr1YnTjOMO4la2qaQjMj4C4cq7nSZtR0vsu15LuZxubITDBAcXhz
hT6Lkw/K+brhe7DmS6DWVmUOHx2aA7WVoKVVd5XFFolhHmfF1RXPi1QBJx+D1HFHrGWKqS+GydPq
VeOCYxKzXSc9JBhn4G4s3kPO+N3u5tXOvX8QprmpD9cxI36LsasqWViBgs9h2KmH8izuu04HZ0OF
d5L5yXHRHSMx0KxDqS0j/2a296qRU0/R+ozhjzC/OMjSFRIYMVfXJfDVnGEYIyT/+SmxX641GVMv
tOUC4MiSk1E3egeOWuU7gk7/zyVZBqZcu+nuu87KlyrZ1qgsGzVpYu93ZSoLGYYY0EbgVf79GbR1
NhLJqmMvAqQgh0q+SrWKWijOj1Yw8knogfQp7s0SkqOgH9QCyGZrUdDT7dcXjECvRJVXKzQkxsoa
srl1rQKFPQXfHsTb/G8HUrSxL2OFw8dNTvc8B4cKu8ZjQ23MeDf4VNVZBrp48+zO50nKlFYoVOWU
b6xGIyrrYZ3BhekV8+mdCGzd7dLugEjbYs28j/AKlMt8neLU/P5vdqwJzKnyoacMxcmgAHCQAhPO
ax6uEMccVc/TMrn3OKBdGsfv7y+qW03gJrYMqwrq/Q5e1THgOT5VzhzKX9ZMj8HRbOvgvu+Sc5hx
nq4VA5MfRvv0O/guFyfosDyBRCGrndmkzcUVEnj87W0XcmR2RNJ5aN7DNs/ZEAxyQd35bJnLe2iA
eYXvMQQQqUV2+SvCG5o0A74aWZ6jil3hEoww06n049PQZqUiLyTM9O7VoVQr+Lm2Hx7GozNt3Dd4
SDhORIcZaDB3Bjea/LPABrbrhVb8a+3x9/SuzdrJ2bFxJTKEgDHS/GcgxPXdkNX35ACq3k0QRHBE
6NLe+BkeRlI4KvWeqvL/nFZoZZkxeGD7yYe0ukEpWvjFk0OO0+X+pWpMzsux0UA4FtLve95wIuIn
YxElqMpZt0MfsxbZ/kPQUkSOlReFoKLFWhjLG207S/Sa8m1qNExnAKt2kOed7VJ/2urPQg1Owcc8
4lhUVfojztALkNUHTy6YlpbQqFFgezQf2uFb/1DzgaQrcEd6SyMMrLtkydj82FXViwoa/bVHceRt
hS7YC535sAKx8Akc3wzqQD3x4U0tLfLX5AVHNlN2Z08EHt8d6+hEja7uLaywtZAa1QD16FC+Zdfg
8KeO4pcKztXDMJ8xe8o3rsZ08BN5qCU1ZSIZLIfWNfhFw4PQUb8DgcpZEqWjf4NUmeam3DHIs5AL
zYQSbx2jYySukzoApe3T1D0K5hbJD0zGzF0/VMiMUaeUrLibyihRLbBqOT7y1eKW1EkJrx+pRt2q
+V0tTVLN528SYOjLLNye/fOtWrNBxDHm5W3CIIwMFJugPpfJMEXliqXOMbY1S5fQJWv7WnLIRoRJ
8nE4ep4hFN6FmKPAUhi0yHB/oFVE5bafChnYYRLtLzAbhlO7RRsr0PBQARcIRvs81AhNyhyVbx4N
SbLyWrw5K6X2AFFRydpaa+9S0q4miB7KD4fhCliZeOqXQjdyMWgIJGFBfwsdApaV0rzw+SOONvG1
vHWNHPLPhtkIcvTVb6KDLwigsuglhK5LSeLqJJV8o5Y0Nl/0EEhohRFWsTb3zyPzmPvTCt+nzyFV
dlW1jqL82QjWHPyd4NDWK4KsL2wujNySDYgSZ4QPAOXGJjqLpB9bRIAtEhAbKlrwLtvkSfdlMaCW
76ZkfUW83glVkM9RfT7qSrH3UpKnq/EpWctrtnb8hD1g5+QkvNEiINMYMBjonQrBOxGVnx1eHLTH
+9EdNGRvt6V8q0d4iIHZ9Cv70GSKyZT1sBMZAN4FjBAYC5jKxEKfddzmFLmiRmC6elHfXrEzIW5n
Q2WgtEsS0NJ4g+iWZhiFQYP53nhvwmDnAHtLWaMzUsnQm3WMCWQcLvAKvcVWC4fdfIojFYjldk6N
PG70O4Tzct0IU2gJqu8DW1qe4BP5BfGEcHh5pcRXDa7/8RvHM8XMZknfxXm+CKBWgPgpJ7/o46LQ
YhXA5Yrib4SOO2opKAGRxDcjRO3+zikRh54pVG0Jo5tXAD1vQHtgGub/6e+X47Atg61yNopTDAQt
JVSnLgh4DrhmgWjllwMu+zYcG6pzsOsb/OtKVyg+oNVMghlfGhiObiI0R5KezJSb52gwJXc5ckOy
Eozw3hdkjiEogfV9ij6NjERXN5cfLqxK7lEbHIRBuEI9ECbFJA3dIj2zokic6rR5tVO8SnhQWXKp
WyFBjNK6HGVaq4/ktk7h0OqSmI7T03QviTHKRyIe7GATDNmExvk23F/HsvlSD8FIO/04v3zfivfJ
9hhNRPTtf3AgftbwFH/96OpUvMqhY0VviI356NpVDV5kOdGf64jh+kPVlUO8F1QfflJuFUFI/N5n
ZdS/KEY8BbV+HCvz2qUxyxPAB1Gj60PjY54hD3D7nzuKiXzX+44VoGk8NsaliFIOLlIinazS7ifL
16GOlgmFDNkG+vmGWt661J9JHvl8KeQfTR0CDclICp5ssXE0aszQF2B28nUghLuMzUN5k9zrb7Ng
T6Hb2zrrqrOvaccuNs6gce/wFJ+Trf37cz2CJw+Ic6ZjyNsblwcHsdYK24sG9bsbmFdRXXvIqrPk
0tTfdmLEyxo6XZPUdUizCyenBJOw+V1pzev8BVrznMYGHEXQM+ILPnTmFBqvjpmjqEmeZ72bTxqq
HTLbwAB5ImAcDObxRNLBjgSVo+h49tM41lccT5e7OPuSEUoe0RnnLnGhqPi6OTrCoo4QrUBm85P3
T0BsypWAOtliPQzQp39OJ+/ZjMgGAR0KVU88O8nwOxB8JEVJunsRmnRDsPYo3sdHcz6OLSYysCpi
TGl0ufVuRTkPBBoqbD1txteBHeDLDcOTT1wqrVRPhPqkGLSkavFOqLoZ5W904wZXPxWSudu4NbCp
vuAGtNm+6V/eaHjYxgxFBEreRCdz0TGADSyukkFGo3k0/WG61XemDtG5+SJd9PKMEN5V+oHda4HI
zMEIAkADLMYNVmHW6uqeglCGx0vni2H/CCUgInChX4BhiIZ1AmdcDR5Yan9BL+m0/9pxIH5Soopg
/CcevEbnkdNec4kABK0lN6H0+TIyWz804xZ8G5JB6VCjaBVLosX+0b2dCCry+ET8O3BfDc+cZ3sv
tH6AxzbqmZRNe7BZT/eRh1h0ju2PKO1lKFG33Be2njaw8QM3zg2qDhbrySBFxHfnj5cdY7qPdlJZ
/RsEehbgzXFs6GNQs0Q4G0tDpveL/W7BHq8SRTaGEl50PfzMW1q96csLhRnKLHJ/lRsEfJAMqOzb
HjJAjmg6Iqg+JUTZZ66Pic7XIrgve1CHeJeXUVsJH1kBwckPSoZrBvM+JgLZ51d9GvxgW5bXZUTZ
WlnX6K7pPUhmdGrzO2my9rWTI5dwT/O7n0YpzjCpHqCrw5W33m3RsHPXNHqRQy4DEzZMpK6CXnKm
U95xZVhdKhWZGA0x3kcXgmuswJwrzfMG2cDzzx54P25lGsXqraRXx/HvUqc9zymhpv1PHW5tEOu4
UEIFJPknfejk41pC8J2Rr7IAXsVCKqu89CNPPLac4HyyRkvCTOvJfqdRRZ7NeHQTNiJTfUtpqQLm
dO3mgKp4P/Xd3j3uPvjcDmDr4Hgf5ZA313XoSoVwrmBcfOur0UgKCnCJyv0vfcyL/7NXl3PRmPf/
ZLvjOAOvQutfjroouMTicpK+qX6lm/Vnz0XrLH3rrZDV4SuJ4peJCNHJxLy2LaxGmEJmnT2DWtJb
G4NhwQfu4u2MDN9BcePGs25HKDT279NeZ50Bz3MA/QCt3wClmCxc10j2ZexaW+zlilR5gCzzMRh2
23qhcOjFKVV1nSL8hXvFu51BjUm+ACuP+wNlXalKkucYw14a/sk/A7nSjjvwOrqQecXG38NLcUrW
ku1ILx0zo1GL6Y3VVRSRAn1UzIZx2S4Jvc/j2i+H0T7WcmScmLit/PLpubvvYHav8M4e0uhlGMNx
Mj+dut9aK6HHLI4apHlLhfwN/qehgZK3PC/ZDMTlfGyH6gMPxQedX7ewyBNA/Jxkk8DiskyyByME
cy6Z1iRlpAIwKIBig0QHnphA+v8n9qwXHTruYUJUT21sv9cVbgj/M+2Ot8S1yeeOmd49qW6OBN23
X264FwC6WsXS5m/8mdTjGVoQmQ3eEJTLOUK7bapfllzbu4ihpmgNBop7yZpnK5QCAa4ozunga8ly
J/G/xVItuv34uGFydNmQIqVJgXrdl8oHhAOJZlo/zmoifqcgKoiuSNbTwmuU40FLnqwKRZAtXu4v
5zhieosq9esBI3KQO52zwl1A/mSm2woPRG04iz4mhuper1sZlp8iwuPlGjUy1pF+CEuQD8be6sTY
raAX9EoWMz+m7XfIsqZ7/46uyQSfhs89Mbtteg1zH+Rn3ocvMb/jh53yYakoKhugIP3U08Dr1ypU
6HKJaSbPK7hy3DFACmonrDrLgE2m4dL552c+tDlcn9VcEIvfWpDqTs6OqVJfpiVU44Dv+YZmR46J
HpUp+yjhtP3pepUplAPobAuwq6z9kwri0a8fWxEce6eTvcFmXrkvvpY4dMsuIrCDtgUK6kmLC89r
XRD5GhcYVCeO+DqX01G3I8YreWnSsTTYO/++xP+y+3V3KEHJKcW5Q8Ee9NXCA1ROIgh2nmNkdId1
KC6W/foaau9EWgSiqVBmVaZ7X40MdumiRmeN3dmZLnaqOqam8obYlDSE7be3GcVloc+E3qtUTlJs
WRFh1gLXL3Kupfvc3G46mFDf/Xdz/ZWjwNvwKy+ZwYkKk26im6MKJqCiGMJrzBWuMLwW4d30GBmL
ahsG5hACF7KJn5BiPW2YyL9J5cTxIX4t4ZuR044lF0GZcADjX21HOYwuQVkQWHrvihMlvErvAcUf
LMuIbWq0r/+kdL/UnGylwk/5cD8CWQNVS3hHV5KxbTofW8Gw5p68uAF4o3zGGLM5Il9qndjP65ZN
xVnAlqp2kntuRPw5aeXbKoNCxvKF79SA1VL4gEjIG1cFaZAQ2B/iWTshfKJjPSb4r8dhxgys1r8R
EUs3CB8YpEHOCsEgd0O/ITXH6ESwDX3HaxFsI3Ly0reYtMoPJ8W/dFHNswr1nYZQT12Xp/nybVE4
57OHR+oDESDzvK69eLzYMOYeEaNA4np9PMAyWDB2Fr8U5yNtTRyFJBe3LCk6+jQwK9VNq80jzu8N
VXh9rqx7jDbAyNtjbCK9O7lpq5WLjidYbnIPkjKXaIa1jdzL8j9ampW70Qm9ykPoZbm+d4qOO83j
d1XwLspngqnufcQ9SPd0TPMplYNzjIZqSmDgZS1W5SCd7+CQ3xxVlHU/IqqC+0qHddwULMMhN+2i
yAOBlA4YusvAfAYNo1IfWviDRuKoriNEylqhJyya74XBTUjWieM2qDSJlBYTnseG39AjQ6XOpA2p
w1hcXYmGwbXdjhvqyo+qbcBMbI/rSAozxsRP+NCSh5Go7W2RKKmLa5yE6w01z70BLK6GoS3XFfZR
gQMTyfLmsf/ShyOLmPbX1n++iqo76WErb8p/oi4U+gqV9/aopKJmGEoPrGcu2FjF8MsGnqBLpXzf
si+8+lzCATAAuQ0eClslrMQvNA0UfLomc4NlCnu7upA+8Gt5fU8WzA+ufQmYMj9Z5bWd1DIZIYNw
dn1xO6FNzpn1IXF9tS9JfLhgMQAoWxcRAbVu86sMQEB9SrReO05A+HB0aq6kgm/VEmmnWmAosozv
JT1sFzE2uiCs8x5mHqI3uBs3E6cXrFvhGh7bEjPSRjDBTHwHGyF1ZsuohPAdLixhQ9tIYecxgVZu
Jc2+bWgFGQ9L/JCzI/h+rsSqzGvVTcFIRE0o8CjY/46lga6KcI4qwq1aEpu0FSiuzi+Rj2/9FMaI
PFtq9X5DE1Wu6+as/PLaBWFsYyfEtEB0pKTS/CkDR0dZ/OcLmqvsGFZBzePjYKDLvGpf3WyY033s
hu44y+bZ1xZM4ZwJ2tQa8Fwq+dJQgWKVGK+foQkHua9RTkqerbkFM71qKDLqe1JQNDRKiUdFYAPE
9LFaKUWF/O/P91h+QfejlaziDIvh8R0ws1gohHh/iN1YheGnjpubTRk0F4p6VYcGaG9cNEWdg7aH
RTSt4veYU/oDph2FSClL04yXDK8rEBctjQu3hIiOjmzw4K4X9YKL2FbETMEZ8ik/0Y30is9ZPVUn
m5+IXiSLQNlJYIrIpvgFeVG9omrA6ffrqcdU4UUR9PjQJTG7aOLIOm3C18KP3qIAKVQQFHPSNAQa
C1aLRzyZ0+uxGmNIQ/Png3rweKwwacupVGD0xBXk77te+2+cQT6nwReZnnp4OREkRSf/cn/4ijcK
0Y69rFZFOf5SRq56Np1zfRsvmjaE0j0klqNIQmh/CJ9mXpViwTMj7g3J+viI3hVM9eV+VVivzLis
Fp+nGbkJ2/t852drWaDhWdPVMXa9e6sYgOobgQqa4165TUd0LFJJFrxUIZMFxhqUh8HSo5ikF45v
/quoDCW+aPx1NMxM8REHBKTHtGakyPkx9LpN6/ztCnZxHaE0bE0b0+ZHb7JK7T77S0YJD8P7iqT/
6z5bdSNAuDpKR2w21mzwHlDVZRx8VL1uPFOpRQNn5NNm6kH0BgXYZxUuZmSF7gX2KMe24m53NmEG
VMtg+yWg2+JpZ273Q5agcZzZK2bW9Cko2GlaRSm2xjErIBb/j3mTtAdh3l5EP9140NQTE2wwbKTK
1eq4WPRgBdGkBujBSf+VbcfxuiQd+/XDdPcwc06IarGHLGIr+01VpAtYOYbfP2XhgdBFL7Cnx6BS
FdNwTyAv0EL4IHmRVvSpornVBGElOteWzyOJ3xpYkxc+PJE69BveG4wBrhA/j7ouCMZjmiURVMZQ
kXi7rmliFPttLvmBAN35WR9n2oDBYAAvSjcZGtPCK0Z3lAfTBLp9o/oVxJeBvTsOWMZFvo+WpBmQ
ZCSS3+NXX4XQu3h1DAxwVnztdM7H+E5hBVI7bn4qn2k7KF5tTtDfAAboVgrCxXo63RJwLPd/ci/o
RT9A2nyzMzgo+YCkkvSY2xy7hoIl7DWszyXuLkB+460EhYmewbKZ8gjPfX+XMK8P8ZF2oKyz9Sq4
drxQu4lrikZNqNj7PJQ6jbpoem4USq89NIsJ3X+wQu86o74xQIPHynmrJlUeU4Y3hQFpHad0VUHE
xF1zn9wXN2NwLYXW5r79ztZOe6KFmGWbLK+KnmNHg9MciNN9pX9I1TTyRrBc3ogHK9tsaGxBreTR
NA6ORLPdjhv8Pc3byQ2jw51lmZmEaJU1hFQjocPdC9dexFdqPdu1HwQWifm028JsRFhd0xE55OiC
Wm7L4w2Y0ETlqWn3Nrx5uw33YjzgLjX9FeVw2cQzJ6X9FYg93axVwvY7KY0Ft/WfA96K8c/7U353
8gguBq0F+BabqtUP+lyI10c8Nlu8AdgNk2JcGgTXXsPMU2EdRhEQ9b26W6ewBUAv4VD8gY2NJPCY
WTZ8QStUUHaRGtZX5LA2Wrlo1mTs0AI+cKi8rPfRAwrD4nb86J90+3heLNC0iTdqtXoCIVZBDf7b
1BGcxJbqzg4xR3WP1AiCmJqn+VOKqCyQEmHo+7REEadiaiIUfOGda1WuRigG371f0JXp25e+LFFA
hZKEQz9FY3J0I+8m2WX5KwCXjoPeIKmHKnvktg0dOt1GmAOmuhotp3v1iSwdBASzgVHnIr0kbVzJ
TwOfooCD8gWcVT9uqwf6yuaLBBUPfpsCBihAVBOEFS7fMc03Ur3ZqtmpuQV/VNFhXucVAvpeuFT+
uoWMaYLcukm//8I0uoC65NzJT7VKLmiLazkfWTse7wLkWeq++j/lsMVHN7NozhiAtNP7i4FJLB9L
EEJzIM4PCBJz9bbOWzdkzo2vOkA2n+qN4NOocAHzsCfNlz4KIiGA1rATapjdB05w/+cSOmMFkYQ0
C64OOyfl5W4tmmWGwFWjAm9lH953bLDE9YqcmI+gyok4UAeCpACpQcARdS2Qb73yCG+ChfxjUab5
2dZJOKkeQrYKT7jHvEK/mYjQRt9dTC6FZX8wMd4OMbe1P3K4qodfo/rXUYOzF43EjFMtCVKS/Wik
LIfmJI6RtXj6WKhLZI57OIqJnO8mYf6Voyh8/RIj0qIhTmJkUc1Zk6vxuhMA3fvlileQNcb7CVGs
wvT2DfxHlT18Q3PZEELMv8HtH3DOCvEyk7DFzQuBWZ9IALniUD4l3UaWEpUsjj0hX2aTQy3XTHCj
6LOtKbIOfMrLBmYl+sPU4wBYP1S0U06Yg2zurQYO9URkfVj85a1jf/rWpGBvsj/eF6/oXFA3YXsD
pEGG8zrL8GQEgVaDEwwIUBT74gHvTAvpVkzmebikdZjOj2l8sHZblPbh2wmbNu1FJC7uD7io1LZZ
Xxg4rHsBPKmkHnCTL0LPnTb0XJXLjCca5lXTgLcZt1czbVf6fNT4ApakQIx4GGSp4r+fdCUUoyBM
k8OE498S5UC/TxwuqtCQi361xN2ioWSu0AW4x905xdsS9cyKCW4VbSYShFOM4urksARTBLLsPVDE
HrtotjxBN1GM356InVY8aFYXc5JEcX/O9JCZSX8vdAwu/JYHSEEyih+4UjmjE7mDnZZFnezTPyJB
9QKpwAX0KmZ9v8yAAqnZcTdFs005mgm/KYrlu4mGJpxymJ768jtYc3yBCVEIhMqmSbunQ2A3OEqC
2bUhyxob5v5MdLBI9uJ5HAE0RnP7fnDqygm12skXGm/kCEd0mJh2QQVvBHgve+CzB5zJFP/+7v/u
nEb9fR9vAA8qe5lRBxej76olEhC9r/RoStZpS6h/KhdHnu6EKKnd203F+QOmN1PXeHh9MhPO0G6Y
tjfpqIN9eJZbVWSigAIg+intR1MKLBdtdB3PT/I6nal3oxjbpb0Ul6VhXjpF4nLFoYpOAwiFjzp4
zmqGl2KxKQwGXLAkezPRK36BnL+FhD0hSVwFwBuETLnytmVNL3aPnzqkNHTdy4Y4UDu8YphQmY9+
MjUmEEt+3vfXHK4gx0Ov+8AvyhAg2YIj0o+8szh/hJikeqZ+5PAzWan3eRBgMJo8qUonKOz+NyRI
dryfFyGQmTcorF67wSLlaqBs9r70u9xJldr0Lod2WUzdYl63++syrw7PCeePWoe7ewicTYRDMcol
nWjfxm9xMQmFmqOCiKilonFTMdBY/OGAh5G+N0VU/E8zsytApf61XZ7aWh5tbHn3rRH/wpoMb70B
jB4jBP1M0pLZ4ZfmUNdqAohkyDfBlWzD8361CCJlMDCoPg/tHlwdqVIOt7EZopWiO15WRwOItz8L
KhH6Sq/KwdkdAXYTop4fOdy7uQImikUlzYrCbQq467mg1qy/x6zNTZxfeQBiQ2SZwoiAMA7JLY3M
+z8Wgjiq2HKJt9z/rtI7hVi20oVZn8IrYTffywz/uAlLZtTr5vXEtSnqGKb3/BGe0vbgemSrAY1W
4ZbAUWXjGAQ/HnfoqNqtrmpBkoFY1lUwTcv7vqhRsrH0nWgf/14mikZozEuVev/hFvxhfnYiW5I3
wKCae8ujTOeiNm7jbTc/rEY8ABtXx9mjER4iDEn5dJ6d1M+9HTdjjx7r9i+JSNpnqat3pgFmga2Y
p9LXvW8AYuz3w9FJHmiLB6mRQbn1xVcDdWdQbeCEJCdQSQLKXzGwUTsvZHd7Ox3rZhHhxV10psfc
HPtTMGMx8wTlEaymZoyC1/76kOfIhA5cxV8gf+pajCRegWYfyruwZoddreDjxVKXuRzGfzblY4WZ
ShYUxjtRUbRLzTDyL/jJ3t5ni05H4AVJAV1tCdkfQMOpPnwPSErQVVVYcSQRRFFPbSqveExpva5s
RQ3qR25isY0ROnKAE/4Lduw64KdNw6GjgcKD178sbDPR6h1GBHDUXZ4jFdLLtnUZ1TvRwQVnQRyc
dPB7tHpR3bAnBMFikJleXsMfYp/dyEQnAXpAkuOZiKsUgosLJH7iLj6e/p95MiXpHJDEfZGsov61
3DsI7mZvZz35WW3qbZswzlLynaAKYSAf8yJ+ug0n4JVFjmiv5u/c+IB+UlvOcdD9T00qx6UOMXgs
LoVKeasj3gw+4+Cd5aUp/1qtv75nURG8L377h2Sw28D/Upb15mSyXpYIez2P2x5zwDuyXoVbfNwW
CnPIP8TkTktj4oBY7dyLJbwsqMm5VuyeeII5WA711Kdge88j2fk0wuMa/6zGLS9mMoiL6BVm6hGe
T/SU3qoJTmp36qEz47p4YXd1v5Kk2CR82mZaFcdcSSNVtVtnYLR53v3OLYTwaVpBDjn/9e+wFdo1
OwZ8QmD0UVC+CC3mUcIUbEYTJEk6vYkMigYO7HnDmyjz6d6t1jp863T6V2lGKZB9mLqhMVdbE7J2
eWzAIErkQsEVPwgq8TJRlgiQXbL09kjEOxWIeNOU69XT4xgYlvZx6+BKK6Abf+MUbZvAYDm03uob
FMbXVijxCsn31E1qTvdrdzMcMHdFuIV1eNYpFyGUggY7/1XhqWwjEvAt1yYOOft8smakfwAJRNT0
+fz/7wl4d1yio9X6TqMhHpR/GhgUiEuMu7k5RVxmr4jIIDcYEjXccNvjV81FWqKwyz3BeD94I5BY
b4IrD8sN4mQrNbgjMqaX43oXQXAtgg2sXipt3TY6Z65r6MSNLBNcZ0NMVMQqp292HllV7grJEPFg
K5UJu39wZ215mzFWuNWDmrqcSPpX5dVMJh3pIn90XKPfkyE7dp8HQIxTQxRtJMghcgjoeW9OrGZj
rPai2iIs3ZwAFTFW96be61ivpstCf3Byxx288KJ/6Xt+3E+RjJQ37QMk0ATBoC1sms0jflZtkH9a
V94oXPiS0tXnvOG0Z8Rpe8CllTAcpDhHX9D/6iZI6DRPnQwAD89hRbji+hZlNks0V392KoPEY+9t
rwiVbtSABYxOKkhl0nuE69WQRGV0k5TxvKgp8Kvs0ZQjKN7C/Gi3B3rXduTIe/GXdEqYuOMfI2bm
UxxsMrRUdOp30l81zP6vENVIbhN2tJLb9DoR0ajpPZs6dmcPKyjY/1IhoAKRMglvnpks59PjceO/
4BfOscuuBT03FQ0cC0TK0ake4IqYnK54lwcDgs18ExCsBwogi3EggBetKRCZhNnQJ0h/EjTcr9nX
Kqx4dvYMGwevKvcc66gsadMhyOJIhvDyDGT+5vMDAIfREIElAvMMsyRt5RcHZMCvP3PGR4z42/eT
Wmy1mHu+qQ0gPZIJRgoua/zXy0m60WSpuXVs5DljYmkGHkYqaloPqWBtICMQOZMHOzGtl3KndWlT
iwvMATyDK/bVuJ1C0llaYPzZDkUD5BbcmoZWJa+vPheW/qOFDHuDNF9AmbUiuLF+t9K/tESjmcu4
JtZ7Tf2Lu2LIJkhkPfUO8EAdqEADUKMDjEUDliXVH5feDFDE2CGoloUp/n1GXgZoZj7/dZwdYqoY
GPMhGeLwq8aC21uOWsDIZDSYtsTKq1U6m3O7BiYUXyDqqOB2vdHQKia4OuCjBy+lHaeGEQkIAXF/
s6+GPGeugkGiG/xmM/tGygkyCBG/mq10dgaEQw0eLOq1JOjZinl6r08EZp8aagAGl7E+oU0ycgqI
qyp6qD51qG+omThZ8vOuoIU1proxpsBCMMcSHwsVEPFo4IgXGfug6dMiaNulsjzOUVIgXBEs3F68
lUIoxInvS9f7bZsdu+rV7GxM1UdgmUCav0sZudfwpf2akFrd/68/8GxPg+Ngs78Te3FAEQ9Id45Y
F1Q3ekLHadCX3VJdm0o6cUjtJ1Xn1qRMKECUJ/t37OaUUpKjQ/EDCqY+3LfX41fu09PttbBlguJU
Hwat9xw9+ozZz7hjyevvMPXm3Mfzgie0XHMUYEvE16uWQMgFIjVjNfvw0nF4+S+SuusfMxrBi3AJ
Qwi/ETKj8rENEDzwb+rAevramfd1hSorWh2htbmgHdxs7NFVAITq3UXX5Ptqg5lhQTsT5S2QBAwV
EVXFoLqukfxTe72meFcGHPDOmzWAoxjB0rUkWj+7B5Bp3zFv1cq7GdcbMa9/gAr33xH8MNFoziDf
shcbxlf3SucMj2DrWp72zB4l/OpG/fVojNf80c/BWAWPSjhx4wHrJPBUfQgGNuLCwgVrFI5qCFwa
miYHm+bRXivIxMPrffmPjuhfRZQE8vKSxJ/tbBBbwMGdNTdWpnjaVkZo2y6Xlaf1edlAn+xpT0AG
BZlBNCLt3XER+AAT7BGFdX3Ewp+80GJQUqvUmdSaXlSCCojchglimpY7pEhyjRDdtwQD2+jdIB3H
VV9nHn/m8sFfuo1G7ZpcgOjKXUXXroEDR/WHkpXhhZUE8p+cSdF2I9sZYjJh0MiV3OA6mjz3g1i2
/oA7KTlJODCyhs/MsF3h4G0qJpRJTrot9ZfW2xtArhZyz8HNmmsMnjF2YSQbZ8DYdxsudT8AhI2N
4j83e6HRmeiQ6VqJhiVbnbh2CqZIxxB6yVouMsmrVbus+pAzLVVOBrEm7nhS6T1/HVh8EcOQifbc
WgfkDkeONRkBs/IMqlG6iT6I8Stj91HiUtpOhmf2Mufm2LvP1iS0kUn5J6rh9xv5FyBd7imaFB+Q
ap6Iyq1qyv9uu3bCuGshvvqRWwX/Zas2I8HA6q0atQc59IS+t8Ayr+EXmYQ9C0mTUi8D2DKR7zuF
KTvItp4z0nB7XM4ZAovAKlgyE3xBZYrJGA90uBAgWfArx3oC6cjEdluPlg5fR7JVQGiHi/EX7wjf
RXHORUURiCiBGaqkBAZw9pAfUMo/IAPlBBSsClGW1J2PAphB1ZNMWVBtZ+RnPAovJg4xkZqof35g
zRJJvLk+11HfQe3gW2/3JchipnqT54gPPLLQGCogbH5Vgw+2A/ndQqeFL3GTVC0W23BOtighi3QH
fZeLmoIJoCU+T6tPcsL3p9oYDHa2mN4vQGydW/PP6qlbtC6A7bGvY4uembTWtVLHnFs000whfWqG
HorzfVfMVOs08sHlnHDRSevda9xpZ/cn4BdpUvRg/+ORiPYIjrvdyBucr70lwNOcWHDiwbG+MFo0
/bnto8vdtAvWSHYrQh+RNLyElXPhYu/YR3IvFByuny7iJu+UGbM2vHi5OORjxRezfVbkWsm4mtF5
JuxqrHUfUhPSlu4ud1uW1STH7HqBbJEoofIKQ45tf/pJvPiN4QILjckGkwZr3BHbQEbxDzQkMZaI
AAdCdkbmvLx2x+CMKbdTE+nOj7ZQJjiQy/RAO11FF9Y5shTWgGoUmeqafIHChTFNd/vO4C6xmv0L
SNWfX4Zipdz5qELe29Riq3WKkZojJhtVUXu89M0sNHHsnygu+wr4nul8dy1fvQzK1v2smglTF2+J
v4qjxeA4fg3BmfbPUJQaQBtq9H/uFBepQ7+ZIcmE8fiJsDOoOTUgLXB6MXJO28uCq1mV/hlFTH5X
GexRwmmA3mtlwC24lRa+4/HYFDvgsNC+wVh/oLdtBEg9RyH3k3jkgeHkodBzw2+23EYkHZu9H4/Y
VMgZbA0TTscH7ZhfnuNKFzmOWokAHI6Dlsr6f5sdf6tVky8iHsAHb53HrWQSirBfNZZLZneMEgjw
wxaRyvRzF/eRBQwuC+CNAE57Irw8KhtKPGCUf44hDDmq3Ky/QAf2awsHd4Ww/iX+xO//+hRlOJHM
i8yif1w2JrKqBTUBBjRbgnyUJ4Ox7rTra20V8Qb+v6ywk/Uqcv9FprlJrsrPeDpg7kFQmbH3+Vb5
n26csq5uWuaHoDPNRYeb2binVHiXBn5TbIGLQ/9xTfm11uiwwlk6j64TtVMSrj5ipr8Z7U3JvL1b
8Kh1nivim4okLsJoekJAH8W6Nv9psRihdCJdK1eTfUAkdoFcPURujZQP8Fj9nCMjpjYjZlIG7PdH
2+wwFn3QiXV2OatqDM/h/0IgX79IXRFZH77BOssKytO9Nb2fiDafHxc+05NWagAnJeKcs5ppYnSL
GLaPgZYWdSKLAapY/5ejeJsTz20WoLFhShaXzomPJpHY1QeFwCBAGi4hf209RepqUjdCLhhYNQNj
jk2/UAycjwvpGK6UoUEuhLRHrxsHTaheRWJ+axE54hkqDaE0OnPg5mXVc5dKvkCHuVaNxDOn1Nzo
fFeQa0Jve0mvYpZguFmvOBD/3ltMX1Hs19FFrdT5AzLqqqo7Jr7PN9QerfRqBXQ80FWpELQsdy+3
/LoXfcxTPQ1Ll9xsccqIkqf8o2e5jDQ9vrJhUSvs/XXtAmzduJo6XTEwsMBXvbkNqWS+iA0zbhW7
f1FdJstgfwZiaawMKEwG0CLlAZrPy892Q2LtpxchoG3ApOMrPX4SDxmHhHvskfv+juLRx7rMzFfJ
D3s0q21ZCW5eyGLKmYswokUKheMi0fbmg6vCDJ8uoVi0k4NZF9BCmAoKNo8hK9NgljkdK5eByMSQ
gP/yD97Y9INGkh2UAss4nSI500+Qy/CFQH8zsCdUb/wReViD0VzRpckEEV7uLmeT0YSskWQZ8x2d
H9E5rPsZaWMkHVgM/fVYZg2wgW1IVPRpExDjXLBsVLfzy5R+2tuOvpbT3qQHekYwtwBECgMUoFda
qWShZhST/xSC/sv1LBub3h0wmUEU78lHRNIpeJ+yejknuoL6mKlV/nJ2lVILHxTJf91vbsKx5I9d
FRlVsl/36LiTaXJnzh1MeEpVlZvXz4qKjIJ2Huo5YOD8lnkz6NLK8kZTHsaGnsv9Wyje1gcDCquF
UgCUhx3LJNIJOjInJ8KkptQmPuXyaIF5EO19EpHU1ZPKi3nUMtChi6pHSNhX3SrunmGasp6LEYH/
B+h73CPFjsI3c95NNVq19rx3mzj/cdgATQ33ukzsR3NhMnAqrUUiBW/g2ycWTuSMflbH62rAiLV8
I8u+raIFOxgTU2Iuzf3bS8JzDI1agQzaMl4xDMqnCyDfMiMee/L42CmYX5OM3bKErRW2bp7XMGQd
UiiiLqZpc/U618nZ0Nm4vfdMmQ5Cu2Z1VeHcs05DgdLHUMFP38OaxiE71J1LKxL9gJLwUlmLzl/E
l4Xm07fgA1V1YHt6J65eb2SWp4mKUwBuW+VkmjyaQnB0ruErxvt0ec1aRfWUfqS7uJlassVDl8/E
mv9ggZykqLh7XgujmjOzYB/oTXXU0rMND0d+inVvGfJAuE+kAsI/kEf+9k30x7l/vz/6JWMBHnIe
cDvu+WcWvkaDuQprA4bvk+yQXxHihSJTiXXT4vE3z5PittYjbOiLBfU4M00Mk6hEgBfzu4nfY+oH
PHkt8XTrWvMBkOMF3aLfeHdEmgW2bTD3pP13Az31JeQ5UpemBe4T7OGN3p6SBwcVnK95RnPEi94e
xR+u/TNvTVL8jgjFIRp/idhgi5W4VJvDcng2vhV80ntMoBylwIsnDxAut17Z639NoksosPyy4BZW
jIcjYE+JINosRm4tNa5lfZJWnaGNbijmeBXKUf6QBOdt5Xuy2bNC5mH3v0bS7eE2SiLLz8zCzyJ+
WpoFDCfrzwq9yEcnviJAxohkEXktNf08wGiZLOTrpi2YDwP5AObdk4MkE6uPzJLoYm8Cih2cAORU
QsITWU147fvxsVBMuJH03zFeqLrG1NVhYEK0amz0BnklHfqz8ZKDDnd/OZhCr3tibQ/0rMLHiQC4
yIPSDkx+x9meNOC4go6XLcX4b1wplzTcovxgYOp1tKsujTD1KMkdmUGLAtzMeyPPvaVdJnxsoHHa
WiUJglT2u4aAH/5ecqkgkmheS6Rn3/GEb6y6wn5SRW3GLDKWo/MFi8CYQpY3z6Gyu82Z59+qMSd6
JACGyQfGkLJjiPPnvInZFiJD4tnR7BMInWs7txT35OW8cNee3Faa9rz2ePzifg3gZufNufk2dGQ3
ilpgoaw5HLuKx/T/dGJPhUPhK8UdbLIelPasJyJegdopIKTrewRMZN1pL7YVDKHe351yccLbgt3M
LDGOnG1w/JsB5V4xFrwGZcH337oCQwzL4ePRQ2DXSYqnXyY4SdJV/kYxKhvoTOLZz2ixmmkdn4bd
hnkB43oKlJRz5bJOW62idI4jQ43b1pATnKCdZtkV27zkWYw3ITIOEtSegZllrx8uqMsltQF6FDFH
agtOgME38s5ssQRJm54vxerQvB8ua9boqAXJr4MpoX8muSTTVRXPU5OxwKbXxx7+VsMWbKi9r/vl
ke9aeK+9T+ZI9R/NlUdgE6jVpp5jZjjeGrdKvQJTWVc9lBOT6YUp2JYhLJaDRzW7du4+MUPzNQgH
tKRycNH610R/cB9zdv+tbqAWWqq/qzXjG4XsE03oh30Na/0KXuMnfPKEFIH1eDLWSDTQEar4ezlM
GmdZtL3pavzwctoMuAkJU+MMG8YNBedsWrj6Ei8GJgmQiq/KDJ27RPAbyDAn/kLbM2AwVSeRZyUj
sqjQJEJSu/alvxA1s0tPLDIaHXOR4jHsJRIO6k92pvAo6TV/wSm3FL3m9rRI7GUY6yH4FzU+5bm1
vgayU6Tfq11CXSh1J1VRhKtSQQaVIr6gNYc1Vy9xr330hABfk1t1YZH7TEyZiBBta4HZf3hxgfSV
zzjW+fO4GpkXYfsoyW+nsw/du38zS9fnOpmSwzG1D3IMrm4ddRUGPpJ8I6EoGY3QJuWWqxmDcOM3
Tqgk+yc4Xg4s6F5g+TZTp43mmKdn4nqu1kOdwF176+GDaZx7y5s7H5/t2DB69rjyy19N0rpmd894
NAbXbha2u/6R9gbAlBQAepfqSXtMaRG72kfJYK/K4ml2rhbApQI7KzU16CgxasvxEUqD+toeZ5S4
0Ozopf2aFUw/pCabPOrCHPRfEOpweY8Fprx3o1s4PVx9I1kxPXgE1jUx+9AuX7jHY7odUkymaj8o
Z29v5xrOz0dN0e2/t7Qw+ai8QU8C6n8MkGJsSFzxMIu7OdLaIwXkLoYKkCI5Bq8K44iPelC52Yc+
i/PKmwRWIM+ui7CI2YPNjwzrdOO7kjTxrV/Oloh8FH/OVvsAkbUtb4LXVSVJFhvmBGbV5+t5ZoL0
jBCIRddOclsXlYWnNHXFmeXxpLFcQjAcjgVfQqq7YZWAcEU4ehUKlt1f4z7DL2dl87dZFthgH4oL
bNQoj4PhQuiPdJvgniDLV6pyX6IRdPOiDQ7C17w9WPBQMXmXKnoG7Ucmd7js8peQnPAPJzIuMBdH
953HUTHC3rG1T8/epLVaRe0Bjrysw1n2lcSB0qvo6nyUYoxR+KCet6LuApQxY1ASSAND65kBPIKI
uTnj/uE3bx5CbffQ6c/XsCGFMvouOHeZQgbJeXUPkg+4Shw+GkdooIjpqSbpA5zcMtQ3Ezf8Z6nv
FdMeddOq+FGZN4K4KPD/3CaW7JSBrf2IugamZlC8+SBUU8WIph49kzXdVweBCsIJaiUNpI5jHJiD
WMHunUlIkPAnkVv0BQIYySnCJaHyXjufgwinIuFbqXCnOyFnqLAo+3M2qJ1siw1CBw9pQ1Ogn/62
FXWTT4QGryLZ7ngtxUB5GyMIailzMNUg5qTesP0wlCCulEnRjGOdsKILNnlbtFnuXUpry4Fwkg7w
Rn51PfsFqa93aKTPJrSIdfUQYUHL6rqsoDfGakbnWwS5ONUPA294EE+DEufislNEzuSFGSXh2OtN
XaZIYS/JnxuxsbWqlHpqqCR5sYVirREJyQDbiTwJHGbETc6ZF/x7ax2O9TP7ql8o23insQnMPf+Q
l816Lj/H8lUTmutpuX+9dBCyMaOzXtoVXSGPt9Iu+uFpD6xyke2UzlIix0aLfyiWZ2xQ/y/5Ed1X
+PQ5WHYfFzTcdIZaPgRNClut7pXI7nJ+TjZSCf4OViHmyitPBn0719U33hN5UsHKgL1lq42HDZds
8bNRZu1LIby4FjAApTXtSd9kaHJRE6VosS6j8r00UpDIfldBqDnR3yfspkNV2r8FBEUjg3BaBxSY
hR5ZBhSDb7IKGg2d8eMKysyyqr3+Xkg4OFbPhLz1u0B5qABMOHXehYRaWGue/tAki5Ygl7NrIcq6
suDWjfQigejBXp2mJkAtry8AeY7U8Nmsp9brxfs48STFwjoGyeH4gwiKqzHZnSobXrmn2/X4CDYD
lPevttdQt6Wco4+yMxC7V+I7h9oBBnFjthsXRazPLdr6ONsp1jilnl0+hMts24S2hSeqXtB+B4on
ZJ5yQQXJA50G0Cgdx49eA74Gv5HVjA6etQxB1AnT6VMHwi8Md8W8P7zyJ67JORNnVdsIQRfiEC7m
0zrhl2GM/fJFsdkg1478e3ZLt0p813FqcFRPJi3s8hfrQI1MyQ/TlHQmtoPsBByryeZG15H1sZeb
MtL9DshJbJxF7tCX+c0eQ1EFdWB1WhvKvh5MlyKORZY9qbZpVv2egO2BEALkMPYvFsnvjngOwypp
ANCp7jqs+ol2PSR+BRWsoi35BcE1OR4HfYP6tyjppuhIvHz+1+Say3S0ntHCBX3wkvvaejYSSB5q
LXOl4UW6Tdad2RVQMcNm6SmszPaqD/JCybVIwAn7m1QdoBVMzcnpZavcl8Bg03meA0hfeOgmr6Pr
C+Simt7yGpahbPshi4MiGobLO81EX1t7m0STpJB817IYTTFmEIR626jvzdubqYpL3ueATFgz7X7q
sSgsi4Ybidpp/RV8Ycf+6xkXhevjYMPa2W9OdZp7iQsyZ6/NX84ZnZLbtZpbq6MawnzrWLSx0O3c
J7qnYhy1ACJQuXGSkFEoIcTsjSENVEberSl6Xv+j6qDN3cw6L6+vgygMyMt1PiEZBrhSWCXDrIS9
gC7heBqdtDmVFwULQ+T1MMGTW1Sk/CINO0XbGXKHrHzq9EGD3pOQqyTE4BkPwQvFjg32bzQUsVXh
nsonPSze4oOWwyu9ImpH5NctbYizEw49ZCVLq3sfwL+0v8ZufVTudRDac2rTa4tzliDIV9rPu/Db
CXtsNCubEGG0t0xChezGvpxqGFPtXT7ltFjCOy4R3854T1AIxTCNAPXBmSAYsSTDf69CT5I2bzXh
MCT3Cv+ssKALITeClDaeNk9F3kZqCFzHSSl70wQhj/xZHIQsMuOKDzrj72PNzqIMlM0TLNZ6lZp6
Yl7TkdE5IQ/3q6xxIRGtknnGrC6eN3FsmhQGj7gPmXcZCx4TgNT3NbYX7cex07CuL2s3EL9SnpmG
HwVRAd66NjXRDkBDcgJNGi6Hh32lp2Qw2hpBp8qaqNr1xgRs/HmuaINsxcHej5IpdJv6OddLKLsn
lCvXDY1RwLCWNyFUfta53W7P9vhRVOhhhFvhbryfVn6RNCzXuCw21ZkE6FZ4za97hFdwJa41grU4
C0fRMXTGSKDolht8+sbGxsnqoLhC5Kjw8uG8aWxOi85vYj6zPpQXC+ahuheSU1AXOPp3BWTz0KYT
lmlwWhdQG6BfXzS6XNGkhN86J99/AlW8oIykdKDIj+5bnSpl5UpY/zC9kfGZTsSXTd6klz9PHpFx
B1g6I8q3vozKGRJQ2CyTc9m4w+Vr0CdCadfJeG1k97p238r8QKmoZgYIDd71Msr/SsNIoOpEg5PF
P1DrX9V4J93/bVeZtkzwcySu7rLK1QT/cTOEjG/xC6sk82kXRPURrPdg/jEuNn58Gz+zxb0MWOEm
7nRzYqpy021ro2ZiQ4SHM2D7TCRhnLPBy/3T/WaBHHg2BoPkOAO8oHvChUDkcscwNobyr5YvJuYk
3uHlRbWFSwg1hsgaNb2xFmM7jGPrWvc85uNY/F2RMprzKq6nuzTKFOP+3y9hgz1JphSbcAumAHjn
4y30gVvAXawJOx98yVuzRm2tkgyjNAlaxhhoZk19JnQJKnAMJpriVtD1nIkEmjRpd6SGUobEWiiG
5JBZU00BPy3XxdT7FtHMaI5NcVRIvrWNolkzHmjZhkPpSBBYWaLI5+Odu+7aVLFijTqK53iAqONU
Pzy1PDhU/vKTUGN3TYcGOX8vvfA7GmhaZm/Y8NlNYE2HOnp5JK6ApFLdCsAKrGssKQAbSZMFIFAE
oRwM9diPmU0wYhRMSgilSQkmqdhc4vXZsrVhATCPAuVuLfhh+7Lruo/ohRUWHR+eb1VR2Sww+vH4
d3vIonimlqVUdaEFk/vNEbWjWQLGzjyajL7fC5QVNZMTwuLnoPBtvIvhu0hs+oWbJtMCycgmOT2v
ofhB5AUNdqvsAg/OL2ee5DIyeHpEy+P6z889XDaRqKTjK7VjZwsr9D+vSpji27MoKnSxKfnT7feC
t6Y0GNiS/crpX9f8LX0tzSv33gcxuf74Tje2YrTVf54HjrkXDKNE30nc/vrmrwsfg9P8L6CdjPER
8YRA4rphnr8LMoriMEFm33ulCbEyulIOdvQVBzzQwyNoi7a3bUFqhbgjNSsBbis9x9kF30Yp036B
8HtpX2lo06vu66LYzlKgm1BUgkRXcn/G4EOYpQyqngOer41l9foo2xXqxLoW5ct3FlSK1OTrYnzA
D0RevmS9jNtLHE5jqufnQruH08CnmB29Tz4slNujQZ9DjxssX4vjPsXou6z2mexyKuXqHuzE/uzC
z2oikNIZneHwebEmTwgiacthsFCJ6fydmBqpNylz171l7miIzEP4XmxB2w5nx1U11qH5FnZuvg8h
PL1tLKtlwNga6dRpKzsEsieXbY+5xETkALKd2ky6uZe4OJ1K8r13RWU0O1RVpdoRdddsrjMmbYyF
nv9jeaooeyO4/rjVzFJdFiEXSvBcTSUE6wuFbo9YG5nqMcapBEFCnyn5JAZ/i9m7a/ViJVt+cKoo
ZEQsznLFxNGJOPJncpEaVg0tkH+PbS7AGl0kObcfPgdUkRmo7kLywLGB7d6iRL5o3YLrF3B30wUL
n7OX84X2X37MfAxER0waTe21MkSaQVv0V0FYKV3wExtuHj8BBRVbQSfDa/W7IcSD5H+nbJOSgsww
VwwIJ7nQ8jNUp8KWSdaW7J2Tpl+oiazumg9gl6MKDmJTtNSHzqyBEIjs/zhQhUH6/Blq3l4gRGWn
rN8doND1y87CsxNupj44P+LgHcIUIFVDgYUzS3iWeODZAGBAmm+Flyl2pz+OCo7tKF5JjZv07a9m
NXF+7jR88196VhTOatNc4LPPFLMoU7K1dCJLSqzvAOeVT8E0rWSvgSQxt7WKMO9M+sU9f84rbe65
k3oIhmhpif0lXQ9VyJB+IR0pG7aggNoQWPvoMq6DkVSybdbvC8mJcpZ48A8wkRZNi/XodsbKl9aS
MkvD3Dvg4jd3vK0YSUGOGNLNxkhonYC1KcYE7eLxXHZ9lGRwYrQObn76YGn+4tkDYP9WryrGqrGv
6tAN1f61jdklVRjlv3hI2CtInbw4VOSZjWVs0sDgokJiPI0Nt76/tl7do/qfzBFc8L9xEW41kwoW
tUxGVGn4406+/F4Fok7PEXtPGbnp2/VpqA6i9ZDnjNEoalVu9zO7yI8DI81kOco0rxt1e+9n900v
+N9Op50oAa+GLnxZXhdJN8xsxTYTiUwGyPTfw/l7Lx/Q7xgifVFOcmfa443n7LAC0kkqX6WRr7xh
p5Rrsc1a7Q/IFp8N0nDUTUBotTEVBjYZl8RbZTqHW35HnVPo5ACRyPOBMc1trUcrZ13zB4nCdTbP
XP9Xcf9S8E9AlMKXLWBa6S073ScCNDmsmo7X0JUD0UM1M8Vb15q8CQdrtXMPxb/H7XGCeW5ckUiQ
JiwBREGLXOMK920iEX/nVV+oBKTQaiFJkjNJztx39yj/+akGgd8XEh8C5VBhuKLOkP+KMjqa4n9+
Rh2QtoXRm1A4h3jcguT5bQJJ+l2UUsT8KZxTrlnka95sWoeo8jaMh9mT7rFt6X8le9p+CPsfbyBN
+mNMANPx3hL0Zg/nlWjjgwZBK982wzq+Eob63eEWaHvOpbyVQkX6Pq/gxIU2ImWPCUlwJsbFBwqE
FMGY1xt/4AU+wtlEEpde685ZY5e0zRcjsygQ2bpStDXeFwwHRfecv8Zhbb0WtG8gZT0B9V9r7UU5
svmu0Dmh5woqutQ3pfJBz5+HKf0Aj6ruhIU++BJR76i4FBK6sFmLSM+HZZrjCJKRqiwrB0lLxOnZ
TkLqfNgewdSmcs79YnEO7mN8X8fk8kiCydQo/K3UvbG7OVkNqL761t4U0xMqHo4P0iOJxCj4pmlW
3ORKO1JftWzDlll7gqtDvcImD2+ZYc6c5yEC+MkgWz2bFlYPU30k/b+JN9CxPpUDLuc8xzu0Y1K+
tx3E0Hqkf8QemMyEHSzCw7bKm8SXDOYJtg109g9gocZ1m8A2hvu+lFtByo7miY0wJkDWZYR2i4PQ
+Uv50u1OvOaKMaixJqaFsGIi9PUFuRjmRnUOyqgdChJB8YIAvp9M9oTpfYFyBi3GfHD9b596/vr0
Q8+dgmA7kWmCvMxwUowH0TWtlOHQBxdzbBAAwRif62iVgkTgOMcbRlPkLPScmAsDUsjmIHKXrbje
Fgqxe11TXpkFOdycVV1vgij9uVsbfxJOloTFTTuzNfRN5K6f0NDyCWnSMkWXplWX4YHDE7EOC2ON
U0rXaMqZ/fG1qvRnANQt2my2RVmYVo6N0juEvukjFS4qFhRBY+Xb+nGaQDYSSzBQvN+PTnyiBIU3
1pTV9KFwakcF4KP/WXeXEjvuY4dqf2VHWH774H29e4fLYHj+6mECxLUwQG8Uo6lkRDpSMGt01HNn
FsndKDqA2Y5XXLCJMFvd71v2WGELVPJrCdmWRr2Vs6nX4xFxmGPfJO08xXPW3ipQ3Jt6r56l0vWl
QHOEmuaQWbZNc7xVWqW63sp9i5FwzuAck2pxMkLaHXqbDBnNU91NdknFrCrr0NlL8mr15uEt59pr
QXaucvbnE8u7uenqpxbHyW3TYaYJwFY6teNqUxhCF3Qyl17TKlL8l/Ex8Q4+9Bno2C6zlWnpWAQg
kbqG5Eh8ukYB6KQItIKF9YuHpCnvfKnFF0TZxieqpiEKbHj2VH3VeyQScCrTfkAVUyJSBVxEL7jx
t6+MANBGfDswI8pRj6AUy6JhtKJ2HoJZmnczxwJWZuBx6i6rqdJXXu8WB9DZjt09tsImWH/3nJZ4
TEaWLt/LDX5BRaiYOG1cmRBSoZFo+eUdcG6JTm25foH9dMFrRyO7JOTXmwvDi6txG1xYljqC7WF+
p/42+umovPATuIZbdcZeJAkxqfdNIBuR+bvPBBv8/BGb07YiBTkrZC2wFubMh87L28QBUyt4rIT5
s7ADQk3E3/LS2dzer7E+FCvIcgZjK47FmAqVqSEjW+P/VdmISL1rTaw6mDseJ3b7bNhX9So5cbo6
DG+Q49ywSb5pfgvrFJHqU1UWFZzlEn4HNl1s3+V/yJRQzpB15gKyR1XfvpKyK3t6ej5kPDpdHQ+5
r6LcW2RvYOGL5KVV6vuWZW1pzOgZhB+burWoIRcI7M0Rpwiajoh3XigfO2qySShGkJ12mMbWDqWY
Ej7LacXu+WndU/MksahYcBHoEvVotebtak/EHKj6+xuuMfhE4iBCWZRPNc/+35qaX7u4VVa4kVlt
7lBycswWowIwzHk2zCt4CSXl5AzAFRz0oZCYEZh7ADOdhr4DCOV4hofhSrVXaHKWmVfbXjQ6gHHB
NW8ZQBl6klt+oIR5tn7D/0YJYMpQio+zbp9V5Dz8BMnQ8gGmnCen7oh+rkMPH5Whaeyrhm0cOgKY
hk0Gfl2frJ1XBQyJ1HeypiJ1ER4MBQStoDxSqk6UYjB/SDL+vkak2vMRDlBzGYCgheUNfmjs+xsU
SNzxgEdW2u5L+nIqSkwYaRC8dVSZF7aBPKCYD+KVzzX0mUvgevoJ/yNLc7WpBl9b1Id/LOnbA+i4
s/mpquUsWj+v1wEhK2XNkveD0fRnVMvezG6nLmOdXLVlxkSRxIaYMIIcfJYAFJTcgnmxp1X+46Yo
+mwkXEfcRpGU5G6h0uTB7UBLzf9jw2fzOHf14+6nYxPsNT6+yEsJq9VyrW938eGoyAN+XYiIsV/O
aB26kd15ZYbN5kbJgvt58euC1MYwW7Hp++xuIOHxv8o0GYZp+w1Zn0JrH++EEPSiuB7VDOwyzLOw
59+udF0pfKj/vSjU3kAUddX0r1tL4SpFpIdbl7DFDFyod3/6+sdsYc+c9cBbEqEhyDXPXE45xnh7
Nz3gFc/74CLLsuGKbgT/0K3XNABh8Y+EJjx0q87jzMHbFRdWFIP9/aSzI3hiAWJf6fl4Hawdlsg5
FFtTlCg5TMV65tDmOrf16HSRRyHTRKL+NstdJyINjBgUbQZ6AJTLhGrueY87fqrgQALgRjhGwzx4
kWFs0zfTftMrX5xuBabDvSO5PPy7XtjPOIbWKgrb36r/jXKldz3Rnv8HjwiKC+FhvAy/3J7U4AVR
5sPfN9BIVUb0kIa/0pqZIwuXbv3/+xpJLFaTjjaO3rWFogWIeKf2dh0fns8SCqQkLKPrdG21WkYZ
3l+KiiddEaUhUPAuFZHZTEgDeZh0Eqs82rJFrvdvmGLffi6/dr5a+av0OrukKSZuDqe8C5D0Cbxz
wsUlgNrwjwJ01VsyOzxf201kEr1VTxNg9hb1wOhAouFazMnytBMAWikf5tPRvpnfdYd75wlrPppM
CqTbmBul/GAwsHzqhz1r7L83+FEYXyN2p+MIqpEy7pFHDzKVuCcEUeD/KX7OMVSe28EJ/gD8kXfz
Nz/hoqKhpeFvtqDRwINR5JwEbeXJsC5KXM8zU56/5TiBHn8YQ7T86bKCu/2T660qjnSNHzh8YaMt
3RPET1gmmlP5CKU9juxnr+eh1Tgj2OUdzNHIykxpd8IrrjGq7D4lyWNAvlvPIe143wCZlvE0BM0d
agTCujBsVYV8/hqSUpK0zDxQqSvsRpJOszxBuI4yEDTp2npnSslFE5dtfP+BfgKefN2D7DznbqFj
vLKIpOMQTmsXg0M2JamDYrjmocaTNvCG0u/Y6UJoYfIlVvszO+MrndFOiYMKXAGZvGyqdX/2kfg3
5P5VViyylfbXVk6kXLNfSWmw05dDfyXnjE+o4w6/pgNG3EG3Q0uIPSXsZt1h+QYjzXCvmjckhJ4D
FToRmNiaUx7qcZ/oEcrCfATI1iZ+zr0mTxZEQu39NlY/z7R/t9z2gJWVXKidpj0BUwE0WRsptC2L
MKQE4T7PVOQD0/X6om94aRBhAQM9qkmAzL1kGkKHBWy1N8rTeEVudlCczu07jw4Wnv/whbwLgLz/
QCu1DIxWtoQ2IatyD+0MqDaA8bQFEr6ULCEFZETiqSR6MbJqU/xBSIiU58BQhfY8fUdKqIE9dGBp
Rg4kMTG0JR3Aq6tweofOe9vA9ZMlzIgahJ4edVschkrP7oBtZ9QDazmbuVJbVKcauBneC19whi9I
jNl10eNE98LuZ0qXTJugBtZF7Ga3J5OerHBcqTwZ83e79t7FZIp55C7U/xPS7Y64QouQiyUOwVoT
ylETvfZA6ZnEa9xFHdocGq5rxGBjgsC7w/1rHH6OdF1oriSX1Gl2GHqFAGombjYK0er548MZa8xW
UT/kJVLrTw0Qy73syp5oOzR4qeScBxVo1kHwL4y0vq5/8hj+y5ypo1bv1IWBryylY12BNHEQ5G5N
M2oXB2RhBAstsZTk422qzTNiNdxXJ3+qrfJ8nNs79ktb7R+0fhUxhTLgRWtyd3Ht8xTMfuYfY0L7
0hAnzCFpLrFqYrW0YmtmOR7CeD/WYc7SPGDU26HbWz/TyUbOOoJnTMbBp757432lHY30GiyTaiWl
BhzGmRg3z2ptoJ8pbKYI0kwS/Ftnmq3aGI8WYqdkVdX0iyj8S86lOmR+N5e5Ypg2Y/jnEqrb8KJJ
+2tytmiEWeGLOymiw/gcNXw/NQFrLn18YkahdDyyQYePB2s+byMB5GivJei7dxBgjLuk7hTXCwoM
CV1MPA3eLEk1sLhPoIP+s30C7m1ircSZ3vIpKTQLv8vAcX7sEC7tL4NdeYOLEtP/vulpKeG44Dst
ARSfe/BZTyKR1SB7Uj3qXJ+tSFM/EYooErJEp3xf0xw0P2rMqoW17LK5yKtqJ+cJ5Rsj27L7kBSg
Pi9qDjQiSxhD/9XAXzcvL5ZTyfa0/t3G8SgPrT7X3WwARibovDeEim2TkOLUsxhOcm+wmOb+mzp7
YjTxkuKxfEvN++621d/hHeYLVSgtsnJftztIsRhBvhVG2jGnYsJNAg0F2OOAaEb0Kf6vHx5GiGy4
5zEAWaRjlt2o2r6Oaa7SquQTXf5cc6znnrA7mFDwGdlMy80QUkPo0NGIPaIVIHx/GBSgRRbbfGn0
GrtLT/QHJxfBgo6j7UpY5ttzAuVbLqrLzQSXNqoMcOjaSiqoERAjszr6RAEPOlKlCrhmWE6D4nwj
K5phsnVdsE2ue3mpMPhsA72mA4YKX+5W2rcsvKe2olzu89TXRVh5xxP5nPJ22rahQeUrppLxeA78
MlM8DPftcTS2QT2wfkS185lk64DrBBz9d2Em9TQ5BfbrI55QQLVHvqefgkF9XAkO8OrkW8SQW0aP
nW0oHrQEaGtagwSJwQo3B0KZyTkwuERYefiyn05zwg8lXMOFx+r6e2Ss1o1JsJ97Odp2V3/n2DfN
hYf5GFz3/1rZ5MF/0+SMp/x15kgiNNalG8iGSjDoY2pPJNlcgE2BKaPhryLkbnwp0LKyPaklZbqu
BIn0XCurF13miQCg7kzoQ8jTE+sGXJZ7k9LrKYN10B/KdIbNdOv5lWURWib28NHGWPlYkCkqfWr7
SKnYPGOa6+4cdVRq3tKFMXgrw3MzxzTca5yOAY2x7cGe5nFh2hkOO7JJCLbYtjmUseQhPENKHOn5
FFJZymAblVuBP1R8ztxOgLYrDbTq33lMgFHUwynj5vqqIHDpBjGHudcf0STYCK7QpnMEnWcbsSVl
hqkW+jlOHphUtiaibZcvZc6VxC024QsEVIhYP2P8S1b9wtWlvmh4DFpnNoruDy2wC1U3ijT9bigs
IPU3NdNOwgIZgWVzUGKsuhE4oQLBcJH2sauJtXiIAWl7AlRhAinBEIH8c8BNiUjsUUeZMB4pk2U5
hu57VLLk2cutG8sOQA2NZic4S4LbrVg0w68IIi5t/VB3Y1hv9E2l6gcbGoo8lXZlCFp6q/RJQzm1
HnF7jow5393Vwy2dVbNf18O+eBIH/zk+Ck+X7ryVDp3vOK3IQkHLDyCbDPHR3uimQGRkYoDAinii
GSg4YPsFpJ0ZgU121r79C/7IccJc/IZNNHyqnt1z4TTHpvlUtvsajEM29YAdyxeoE7QR8GqGVwdg
UebNSQzLoXpmBhbVvXahnCfeCYlXsFBWAVaOh4vu4x0++j6DY7hOhA9hGtfEzHTbyWOsEpcVRpYK
bTbLOrMT1bKoLgAbfs2IomrLa/LhQ22YJrY8x1tMVoTPjoE+jeCq5xAO64X959fQOmvJyoRMcyYq
JrkpELbIH2mF7mzGYDc83YhI0npwIcUdkl9dM076fA7hrQtki25qJJdg732t2shQxH9GtHIPUrFB
jYbTztEcrMum7BxC2Q7aA6zQqPonkz+l4uhWSI1si1aEd3YtWCSvarXd1KpXjV9RXs0Qkq5SuBsS
Zi7eJ487RjU/PHy7kedu2pcmudyVpWkuoXikriU44Zy2RccxOziUNRTkCUr4bxF5yXcLJDPi5qbx
MVR/7HAUTsgYIAKSuPy1gUtNCVD66Po3Gke7uJDAc4FwJ2/3U7RCs2O5UiFUWY9/64BuztJhLNTx
ZnaELRgSEjOzJy/wy/NeQ2/6HwMpelVG0cw+Zc8TJ+CgliyiAZFZWttl6D4sgnDpjyHUStzgUl4h
vCUforhG9kV59iaBK0retommHyKwsy5OzXjLf+xthznQIWr2gNxhFwD5GDZAwQFJwk+QRU0hHRla
dj/g8uwcag4yxPv5+/wWaj7fDsTQwjNRjTfEEgV1W2X1nkTnWJZz50AkwuPlbtb8bf0YeBSPKv2o
hQvEjdhyi7SQJulbpdRhwB/vKwzUZj6RMLUUtIYX8WzzPC/gMgoQ1DvREpV4wWkD3wFRU/2GsX7t
kroxrwN5XNQ1BHO5TN/ndBio6362PjvaoC6SREHjvAOqnn1oVNi2IsQSadyohkMW4ZkXbmlRyQbv
Fjv5KZ1e3PRztDYjTWN28Wv4Lvy/HCWpG21a45EgHQMpbM9McRkfcW/wfCtuzYqOP27O4nE+yFAC
9EPtYxOblPOneWz7pO29JSETQSEt6d+v2GX9rVRk+gcgSbGQ4JiKhmrtkXUhjxKNUt/BKOaMmNRi
aK95WmJszGXl+abtGPiMOnj/k3zwykN/XDFlZF9BHGTMPvhY+R0ncj0VN0SvopAghiry7WfWfmZh
o277I2el6PQW2kbSiqW/tr2VbTZYT4/mMMLiTIwGeEubUdzrGYp9k0rG0bHIVkMrkFYPeZrLmDCb
xOknC0WNZ0gXAGCMd41JUktH4/ZiyqCjNOEMRx2f+lHIzgEi+WKnQgH+nCMJQF3UHUQeYjwACkgX
CODzKGitOc3x2JZ9H1MkRF39BiUskCt4lm1W+q6Me7RwN25uWQ6SbHc3Q3hkOWtJK3ENaXTZkgsi
SGsYKHFdZjohMNZ0mNXILKYpOkPqArZVIxiUkF7/oMSCXdctnckEMzg4hcdO/nefvQsufq/Y0cew
amjf5O2Kb0yMGpFOCnczDVxD+DIr/jYjcEFhf9O866te2X246elPWxcQtMyAsM5M3VrQk76gzZB4
vumLZLci9JG4YePldnn0Rel7aVzjp4f+kWutpi2Qj2sPge3NF0/BAHzuWL3bz/orqh2wcW952zZx
4Ds3cTcQh60ouMwyLmHlWV9QXlVpJl8/+WoUESzsKq8rjcQYdoVTqp3nj9CagYRhivrghxmomyr/
YbSHAksMcPfMzgSylGId/ft7HXDIUc4Tcsg904snBUlScRxngkWguofXRTjm94qyj6mRp9we6MZO
6xygCKcfTm4ecKAk8nOAhcOLaXp7q9G8lxKO96obLONZ5dpQy+jjuyCxYTna4GT05EtujiqjyNf7
oRNtyZD0SRowXVZJZ0Q0zFFsaijQx6Ttog93pDyPUfexzw5YVlpqpf2P+ciejT7xYJUXOjIZt7El
7ld8Y753HfIGu8gv+1c/sHJo2oUC9ARZ5HCQxPTUVrVTQ8MUZiK+eOut4vjUXxvjUGDP9Q69Oacj
tI7S0uxE++TUUMeXtWJaURTgANkaWHkap3itX1G0EtgZ4A7ObKJduIVifsfn4TEbEk9lvl8oBw3A
Sn+d6va8LMO1DV3RBAPjQPwOiqazkhg9CHj0ywhhtEP3scDSnFd0KEMRMbRZN86BS9ouIfkbTjTJ
TknHTTgVx29rmB6PFGgzqQi16+Z097j2NDVsSDNkYgW3lq89dnRyGrPh+lep07EuT8cOh4VtzFyA
Df3W4e4dOwQbLiV8TWJO2WPdeoXorJNwJZXud8NxtcJlXM4yj7TMypG0rxotPq1xyYft+0tN1FRz
NI9ktUpjUV4EdEsjFRObmtkrrBUujNlcbZQkXqhsFKY9UEDePr/myYnj/eusOW7lQ10HHh8+rT1B
uBN/vt5f3jBnlSEba1a+yrRj/XShC2QuR44+ZtFgtSSmcS2jlzi4Qavb+MsTIr5L10/IT2q1PFSA
vfHoILai4u+DR8cXW7WxnGld3YW4MrG+ebJeM5jX/ZW+gsGL1DCenH43GurSWJ6NQYy/X4S+SUaG
Gxns1JYxkzyaunqrSuqkJH7L4mccWhUQYkZE3u/glYTNK1sP3R19GbO1wa1Pw2vdzjEeVQQMFgwK
KWmqNIoJnzAbf+HLdCTnZ7OHq7gn51cyg4yAuBryr9LJPttjp22cfHATxF+/2S/hNp72aHoDIcJl
Hp9kw9OpzYrIinUT6HvU6G84d/aEyM7YE1yG3y3tuaHeRdP9A9YHoT7deML/0tmF+H45Z8MQcYv1
y55Ho/qypLx7Qt+8KhW2ZB5lvLNC2G0R5jqpWJUMdRoXLKOtFggjrsrw9Hd0uohGCbc7k50lB/TF
zO68fO8SMUjvyjyIAjfjBicn9jNgcckbk7pF2BZItiuFB7GDteq6do0TAn5Pvy7oPS7K6+hgDUN7
MbUaLDF3VCuAPpcAyqjGCoq9Ij12pT040+lHcNxJAIr7XN+EEM95r6M1f989xb8yv56Fw8V+gVOm
Vz0JeYzAcG4zj8vMRCmWeaZJqLA+JzdA0dIfxgmi5AwKRtU09CvnwYZFxwKlneNAaxvZH4SEif4r
SjTXVoTskze7Uxw+MHxfzpDne3Nj6DCTddd+Abw9D39YEKdBdx1TnlqVriR2rI58dQB5cwFBeGRb
dcNLROzvWqIr8WawSgREEeCU7yDLnrJwZwmwXieQ7CUZ7FX35ruaycD+DjmpL8WGmSP9/n6NDnBF
MnXl6wf7j/dvHncp5NKOIIxr3OaFsN1tRa4y3sx3m1q4Tw9xPSyZZVH4iFbl1MQe/hWwQltw6YVT
kVQkadnT2TryjEmPvFCKTpTPa0zrP4Ldzy6mvTB0y/jmUvuj5udeev/ZxRQYJLdhe+b1ZxJZsgFB
O6GTdOxtkRY75SIMqwYji1ZEld1ygNLO8hZMumwlxEfbOcL2hfqniIBFQBpo2toDnnQDhpTAyR9G
lxTqIxYefo6jgxfg4o+14Z1Ns7U5cX+UI0U0tfPXFuX6vdNJq6f5AgBdldIPbzpgKvubIL5kDQMN
SY/WTE30r2lxXzUhbfVh/qxzQBiRI3SQP9vClPoQHgiKV4aqbAvEpeq6ycVmT8t/zXUcimtcR8Rg
hZC91mKVE4nA3dbb2ZAqqDLhNYPnkrcaJRcyFkFGG2NRD7XaddnfIXy/DyPsztQ8z2OIXuLtswK5
MBHwDtc2igY/GUl49DygdsvR+sGdMnwc31fijI4FlxLv5pWMP7Ls6Qvaf/COwbyeAFDOZRSJ0mzD
HHBcLyuqE9r3RYIL/8XPrjAHgJmDRJ1ujVvLeUsMd5SS3GeesQ8qnTkOW2w2VOJicXCzjfNdBXLc
inE+Dk30e9zWJZbz5TMvMyYWaHbVPygHEsl6xKQAjj2hBKPFWf5LY4Q0Wgh3uHvk2oIdXnu4NAXw
dgLsfDufzAdaCLhOeKzRpdegzHCxthaOxQ2U6PIeCbVehmR6fl7kgaiScBpv3utAmtg47K5ySp+R
jhh7k8D835pKkkocHKJxwtyxdzw1Htijo3vv43LGqgsKAY/RRjCmrmlXUFKpig/RpTVlhtnL5Yfv
SAgNdJOIKLmI8K8d6tsj87S1Hrm4cvSg3Y1R9lOosupHZeicC/xwRSFUAEu6CoyRMqdug5dbONbx
QYnO0Dd/UBbaxygtFlQ1CzwgCwvXSiTD56cKgxtyOLYyMJSuUUDAx4SuZHStXfcTTkdQyfPUou4g
SV1P3zy9xZPJ8BKi+WfXGGBcqPaxloLEy/FrQbW4nd2PHTGpJ0W8ZlOHOoQYimnBI26gq8CW3t+W
XezIy9ChGKQ8FxjnXGJ0YEc/FMhOrEZT/ILRkAgqOJ0Dw08U9D57kYz9fM+XBUvhoPHvYN/HAWps
Y8XUpAUM1sjmcpJd6ON5dOQsC2JAwEy66TJXzX8cTi7CnTXeWGH0r3Eq4Or+vmWNWtVS6hGisvVx
GgoP5deWhJtbcVWuND3rpq2h2EzuR/lfhOod0faHPWqQzbwhYqRVbT+eR58QjeIxxfBGZMmqJzvr
Q05flB9shqva2CN5Oa7ehTOGzd7dTzWbIgUazk0IwKeEFk2jRvqyDlovR7Z3vaqzJQsIqsXzHlqc
sUtVCzRSCd9fL1n2gSr0jVAvDVrMOI7MFUt+fjEItW1pd+Jr4YVzmU40aNSYAvm1zvim08SN7ttx
YHae1M1EMPodx0iw75u8N/4gSsG9Ztn92E02y1b7qoqaA/LAtEk3QQKNCh6BRqxtRESSHUTGt2k1
O5VDoq4RqzbZhj8a3YoDq6UqydeD8lEHpOp94+HusI4B3fEoixlN0WQbTWA/JZcSMzfmNIjl2Blu
hamN9b28a2s79BUJBA/XVbLmmpsSw0edMsd0dlEaLxj/hCsNNLAXNkUv7dIpQ8IlZdGizw13ZC95
+6qLNEoMZAHGAroNOANt4F207wjBtu7kaPU8YLLhcDcjX+ntWkt6AcA2rFRo1e4jETZNIAwnDqT+
dZYgow18mTQerpFpOZOBaLYXW93Ni5KNezHkU4PQ45NLrsrkdnQc6IqgTB0kynn3sxLAfbpD5Wrp
R9EWhzv+dP+nrK/UdLC7fmh1/5a+UDVx5+ekr6Z66+JfmNh9yvQV7Uya4WuX6AN4WIn8ooIQsRtL
SKdZwsUujEezdkNJ79oIKAIDd0BdSXJtKBuz6H/JV7TY72b0tSwCqoaYfqa9XQgpmq6xy+qYOK3m
PeGCDkR3g2xk/Bko9UUE4vKXqXwI37t7E0o1s/uw9wfLOrBN/rSq2/yRx/WhhkHkpbiq8TkERMuV
A39vN+kS0BojnMuUx0M1KRtOOeHAvQzTcuF18CxNx6oplZWuScqiu6UI7bVcrqokrq5hMYEWdUXF
emUBpj5E+Mr4jPB8xDf7GwqzibrEWqgs6o+B4UnZOeWADFldeWHBBgTvmpnDlX+kE2NBK35fjaZh
/08MAqcCBtEyyo8XOuWJSAdd9HKTayUvHOAPQRzpL/1RCbHSVCxbph/3aOL+PUeFB3xOFGmXmqrC
HQdXrrCDehiD4mZpxX64PL/54rWMCmhJhxKUAq6xIOP/CbxuievfF5fqiuhDVz5lcIwBQsKJOO18
aU8KQTtxxTGixcL97MY5owjUw3Gx4h8JOHthbJ3xWa97Ue+fuVvHh/pN+wUBzNtK0e8t8m4P4EyJ
twCTh0YZnDBkO3hxSEYYu9i3qJupr/BmKZlZKBRQrzDLaeTRX1mFnOC2R+W/hkG4dxvZwyemOszi
sWpI/xCshLwX1tcbWLPEGl4To6mzp+uSFe2XeX6hVVQewEIbrhCgLULmXSDli6xnuwv+lhTbPdnt
KhdGlqVFSVgHP88f/xym1+sDF/4qNBoQtN3Gnt3hR8Ivw1rYiMO4XVe0Sf3fpHDRpfOZMxCwzObk
4dpQ+vr1Kys8Oxv5Fb6I13CyQp1oK4QV5sW/1oYAm7pOyjJPYGl2u2u2Yrh8EVzfmASvTZHrgbvj
s0y6n8rQFJKMDDO4UwFYbEc4BQrz3KV4w4WnTcUSBZa9F1duwFhHp80n1SbeBTvUriBTlqxH6x8C
ao4en19PtCLf3uxOvdKX/xRW6obLJLauV6S5tdbLmGTIsfEFNs/4vGnhFKaEU/e+otyOH0OpEiLs
KsL9VFU92auNPIiPD2wQpsoY+YwCobmX41gccPjSP8ll4a5Nr1U/LdQReh6NvcwK8siqvRSceHGU
Md5XJggVB1IAUQmg2V/KtPfTSuushXpFWKZeFujBJpItd4uvqu3+gMo7P2vhCWf1vvAnnmTkTMj0
MPH57soRbFtEHeipUE3on/dKEIKaeE6yqjbZiUa0k7jylvuKujbVmmtVyszDq4kYUQ5XbtCsNQcG
g6px8bKt/dC6r8B2JSKKFhMi9EEEvCDlLZKVK9Lm6mrJZBqvNaO2rNGMm0Co/5fkd7b1fXnmpK8z
UxKGRUlgx1P0VaNsCD6jeeT4MZf0UwK64zmEXNubkCN9dJ5c6iMHCFApKt8kiOSucSaWcN4FE1hU
Dn5LBHndV9J9M1XzlfIvVd7pPgn0/RWiVDobeBVUqT7DzQqRq9cIYbGymWg5egTjoRvGYdwsuqwX
kJ4PpouP3gqcp1w3PSeawuayCjiy+wVj5ucTaTHby2A9jOw4CG3LQd9trXSxZ9YlU5AoLlVakMbF
y0vtB8t00kHxQl0OQEV+FDK/7X0M/zEx02ARJg00Xh0aT82S54rGmZnEbd9di509ITg3cF136pre
Ng79fyG3m9Yqkqib4qej15W0ZFGB+mmUWYDOHvFtwS9Y/NEjFh5Sjc+npjYi4eDRaQUV9V/Mn7JT
CFjIcdQTZou532h/dZRLrdHyG9UuKZQKdOKlCO7/Vwmxn+jPeCfqUSYNWr/CL2YR2Un+KkhJe5sZ
zu7qNd+saWQV51phvtc8j6Z4WRJ2rpAaoKENhXFHBUKeJPGgi4n4mep+2b/EY8n5HatnwNvnecce
rY0bfwCTqvR/WU91QoYPGoheNuH17Aw8yVokaZDJaX806+4b6a6i8mJ6rYMgOK34kOtNQAoKN6mm
WqL/QVVM+ybHqHKZCkEMxRedKMCUBLjWXaB45YEPYc6aJsr/UFT5jNDh6JNlwgIw20SGzCLLNDTV
Nnpr+xB7B7B2AavTHhLBfjJcR2bPKaCZdLE0u/GvJg1ci9p4hCUOj5EiuBqN+a/bVTEMPnGtibCN
Hia9yupac5nr7e9ZCia67yFkx5S+C0tJrscx0sTUWsIRhgwoNfqzjA+kdYDawpQOTgmN54xX+doq
wGwF/5S84mwEr5dOgZNlgYUvS/iL1eV+BMC7obUGaHssaBpQL8WBimW+Cv7i5EYWbE4xH5bgCAaP
PxoTdcCMVcj9XYMtLGv2T6bO4ZLM8Re5gPGQ2QE5NoQX8nsbg83Et/XUTxlrCa3/WNvS+MR0yAlx
vZ4ZcT7COO3W0Qxgaf1N6wBFWsFma2xXv4iCMW38Ts12MrfxjUdx2UutH78j6K0VPww1EBEMXBy3
HyCqb3kwonnuB9FLR34TGANr9SJ7sn/a57EpoXCxVR/EEqT0J0QTmiF4DO8RGwNWC7yqB0nvfzBB
Q8o7jQbhTPXJoeEz91vRN3hfEFu+7N2DacwQDEeptOprxOdBig4c5HQX+87APGs/0+uZhMfkCPlx
QwKHfeygSGc4dMvhNMHGCTdlvtpnL8DHYSRcUtsLD7EOCo5XN+izAAZBppCDQbOP/E0A4myWmQ87
TKjpE5RbuQv/mHth/klvlIgFiYQlkEtk1aJwMbOqCUEM1H8VVtUdvO+ac78lWG4eBoDmb0Kbf4RU
5/HmQ7Fbvbv2WJOTCgwEOQiO4BMnArpj6wWi3VMipIsUSWa4QdBOt5ghZd1Sr/dsG6tTyMcwmyIa
F8bKgioU7eJ2NZYqZ4jgifeVUbwA6QPOczhxnOg2dd496MGVx1GXeX0v0Ir5HovucQhYEq4+UIi2
H539hYAshALBnM8mcBGt+AokgLmOJCtdbzDAmBMFPRhiioO9CcP4DDMJV+7u9eIGBry4AF5xbEsb
m6XMgoVW9MgZaTImw9n8RtAt2uEJI//2kgQuE18rLW84ri38IBxXKtccd2eBh6cfYpemCyobI5bG
+bYhjYLno3iTIAO13l1TtWqVTq2BN15OUn0jt0ZCj5posevLsuf5D3WiyeYvuxebHDCUJRxg176i
d39nTjNN1pX85M1QSE4gzqLAOqRvqlVimYzuT1WeaRlw6H/8YHyatATI7Kzr7XAyt7Bz1Fe+RUR2
1Yada70rutkPLu+Vr2sJxxWqsLGfCMuFRiOHoEF/u5Qnt47FqwmxBXTwATSP2LlrAovD8FOng7jJ
O+p7iCfITQOrP9+axe7Ce/LiczTa+WWgKvPCmBg6MeH5+1/iBog3U4T1VR4uvUtxMoSksceyYKfp
k+6r58ox/KqYLwG1jES5gjzuc0kuJigzVT6OaR3OIFQeMmlXT14nDnyhaAm6XXrR4yQhBsc8CXLP
X11EXkuMiYab9ubNCxbIbTUDQVl/TyYmGjv+56licYWY/qvuV8NPTjwoJDb7pUvSR2GlTuyNATOU
hlewpP3YpJX/xTuLjWT56iN1AitTBdOaZGekO94DUIemfDravB13jWEfIs1VI4BZ0GB4B+qlDHXq
lL0QQ6gAZAGR43WkV4X90ZG3krtKbfBrisTeGeRXCchdKziPpbVeAAeyO5GMVL8j6ZcIS9wbWTei
omV7FpV/E7xtmrQUzftr/4TvBDr1ZlYHHbJtQO98nCkJW3Ekuu3YPgz4blFzKybX80e+hgrLQmpX
XJKQNrEtmcD4Ao6h0so1/DkAqNDb46K8qKG2LtGparq3OUxeSTyq6RJEjvNuMBxgldUcX5WDWVcw
8fS9pHt/M5BmopXM0Pp2/lLW08BZoo+x/LWvVu2Jb1c2/GHFt4S0zloI+lm6l+f/lcwziOJJdPQk
7OYx7WRdAPGzpxlOJ1YmsO43+eD6Ca+inX4sMMFArBIQldceCpJb2wNyXLcBLjUy1pH2/6wPwbry
3V2ndsghDo4vwDBe51jfDutt2ife7NA9LlxdNZFc192zjVzm2gaYTpmeBG9CbsI2EGgcfAchkL1a
KLDtxnyWwr+V97o0XFXhTUx8kItrwVcDlzxY+qZgAHh59dI9zH0pKkhrDelKAd+wLVqS8sCARaUU
+lyMYRY5M2D/IkaOugHp09vMUZ71YjbjJ+L3tE+6lN44kOzntIzgWfaK0gsPwExCdQOwBZ2x5757
/GRs0lGMhXhVrhrLkjNvNMCtkzfVo9EEiKPfepRXB477dky2fdEeSAjf10sZs8guQn8zvCFBFX1z
RqSFqt2FHjhHrqhUxaEWsRPeycRZsLjWq9NgLVHs6FHfcTKNFzpgXBwGo2r/h5EUwVU4ZWqzhEcA
NowXv0OZi/wImMs1r3K/CbDSZniv1zqK5usMDEzQdp+8LWrcwZBj+0krzs8C2EAFrMBqe9JeUJl1
w74oQliGMiSYjt/BDZKcBcAQjqTFMUKyFG/RS9NAZslK816e/64uB5KMKUOKFPJUqnV5cAwAuvki
YG1n8h2SAM4buW/T9nXdXZw0zFCUgS4FJsbf/4YCodDXy9/xt3DbWvKcfr5GtmeWzKEpVtFYheoG
vuOH5h1MKiYU7CzdRvAVj+sXP8te6CMH1d3QnXv/XVyaoac8a45Zxjm+49fIL54ZzeKIk9xXOXl6
RJEQhtoyrhNxa9cD91wgfx7zh4HdTk+mn0oIQkIv13Y6gbTAQDnebWHCra85GP7zzCxPF9uZj00k
Nb1xgldsU3Vw8zRaDdyU/wGyXK0TPsNt8WuqA8uQG4PM5SpP/iZ2UujMA2O8vwTLQHfdNVGmHN5K
dqPAj/MhdUPMj4jRcEQYvwSDPjUcY1Ghg7Ci0INAkUK6DOl2YFse+jlOygmzvLRSV4gMFD4pobPk
eP5ekeSZCu0/XlyCubHdqbMv5KvJwz0k1BcMoRKryK25AZ/WSoZMMX+cOeFXyjQDwHnqYQuH9GET
ysi6DEMsXlBdmUFCk4U9r845OFVn9UPXnRWVdqKwT1zmwxthxw/HdAsWLxVMjYV5DFPwi1HfySJ8
n9+iFUzXvjGOXLhsl4H5lQbIehFsh2KmYUnzN8RFtLInVgdEDEIy/kQw7IZXOETDEMwPkn7M6eCs
A1ONEjSb0i2ZYhni6AX9OYlUiwMxNt9/DFRJmosGnpnsLV2otJu1ZOY40xR8w8xGdgGtnIgZddBV
Gz2yYy+lfotIjPo5K5tIYfAIy02mWPjVAaZ7iV6GdcbcJnQH7n/Vgw7s2Ge/v45fnvVOLLY912/W
TL31Q9NbACaLzUa2v/aQg+7PGlTzjhcbtRVAPkmDHwWD1uOQDabQP3xMYSkEmGmAYdl+u/wB3/p5
lNkSI6XHWkyha3SIYEPUQfMj6wxjjPJ8xsB7PXNU7jgm4chlfK+dTt4+azMYZ/RhXtJ0wZp7Kzdi
pl3zaBRB74sB0qEkJcaJZYZic7i6dOM/Q5ziuaS5GqFNvmdQZNsGhlgJWlq/cm9jLm8zSvNw4AUd
HiOfGnw7KDwR28oxW6d334JT0Ce8ebsK75fYoyu0jrkykMaNvu3Pg2RPeG5oBv1O6mlpPCe+SIO+
zym59xZTEgCMHvfr0dJ4B100aWbPMLs73k+HDzyIv/r9UMEYBkNjBvus1MdGsFZ/fVNQw2Rg8uWt
Wj3Zf6cnVIChzUBylag7pwP6dxey7dAvXGf9EJvUNmUyU5Ucrfnbkxll8F5c6wWo6NEVz5AxfFkj
KoACC4J966Z5StVmULvzavwAP7Nxh80Bqz8bhIkoMrjI+WROj2vZ1islqCX8Hi3OU3fghHAvkgC8
/WmNp1L5e68Lwc7CSNBAUxufAzJgYj0chIMM4+ZPWHL5Kul4CIocCGmUhnwshNz8J3VGLrPhnsKc
IlN7LW3vH8cBgW0Bea8h2uhVf+nqFTuRgAbW7WsU2QpKP0R6vgZJVRYrjxQgz4sEOKcdS0th+E8t
Rpm6Ai7U/shWGOOlYOFNEcxr2kXIb53X/Gx48f5sVUbXA0ENmaey/Dg6tt+Pfcj+x7/kLaHuJ0Tw
OYpiMAwpPze5ESeX/VkAPRECelq76zTLd/JHGx1VhiU5BZPVGYemkAOyFGvNd/Zbwmq0yqngXLQo
CchyBcqutQ0HoAvhs6AzbIC5VUDrSeQCmZ+Pz/qbEyvWD2fEJmp7L3rdbY252G8SkWf1w05wHYRG
4xS2piNoQALM/dA1arOfoBNIUgAQQcqLjWB+d//2usQ5ptEQArZUdlDHw4J4vaIbbggAG1c33Z+j
UMZOuEmqR2E2f/bgaX+U4tR7dxXBYFEA/+KX5gLZjqdhz74t7vbbRP7y6hokQa9w9wcESn/GvKNv
RazE2LuGWpzy5jcXG2h8UQ1RP0OpbOjCkiR6q6PB+ngp/8JWEtI5qcwXgMrSf3gs2lqWP09qJQXi
Tf5bM5Y+nesSkJUAikcrzfcWaY7cHWMqKFgXCrnfSNb0tQ9hQZXteDo1K77Q4ZW2JFUfvPADGjhQ
6p1SFAUhBIgvFbyC6CTH+bpODvwFbshk3JWlHEgaTUymFd3tiEY1Q1VsQNQ6xF8TEG0zE9GBVwme
nMM/ibxWc/BK+fBVsL+bhln69WK5PBowaTavHwDZ2Fn/O3snI+KysWQxdujqh1+6HWpGweEqyiXQ
1ABEz3W46+GIo/sERw0JwQx54bKBLzjhIPWS0RzuGnYevidzRtrP933xNCje9Modb3U99UmUnxU7
NTd9jQ5wHGIiaIESokn4sHscWI90uI8zzF3509f7h/w78miNjDrjvcVBf40NV1XFIp7fcRYU3aVA
+l1tXlewX0dAXO+GpcGEXkTl+5X6cLdCc6LnR+/YR89wkMMvNoY3DtFmA7WehlJyOjWDPGQw0eWY
a6W8ic3p/dW9ymao67SxbPOXhQOnQLXXUmPLdud455SqXDP8RaoaidaVZQe65MmrnUJiGRXJnuB0
f0XlVWslniK7tQ5mb/Yob6BmypfeTx0q+ALWRrPBFqM64HhRSUnS3aGWSQxVwxIFMowHhmGXm63L
JkULieS2tzAQc9PP3DpDSXm0khXsbc81ZJsks4bd0VAe2+/LYiSTJbU4dtJG9VEI40PLH1Y3w6ZX
G95jm6swvPlzwaMDOr7fcKNuMi7BJBUy1GHpe5B3s7nhDpJ6qgw13KYjEJzFPEZN+RVmdTvG5jJY
iU00mlScUkFz4ex9JqWMp8hfUnAHEsoeUHV05NKc6xlBeYryMb95pNPLIpEvS2K+1iGT85FKCSZz
NSFjVlePM7x96JJ6FptgNaFuIhsjtxEc2J/AFYjx8a5t6Al6xEc6OXSelAzb1EqSnlxPgB8hdLlW
t+idLxhgyk9iqK0kVkclE39TRdHX9bqiUyXJfRvOYvyZjZH8D3WfN9RonCzqQS9sOsknVpRVhTlX
xTVuEImrKKb3bavlGj22nvmhBRjzCkKE0SyS+H0PE0nnhsfXPR7p/TjJz7pasxcfXNgmKPAdBR0y
GNxOhgQT64JyTsN2FM1Dpd63xGZ7grgtup+9QQhqVH2JgiKeGGTpoueuZVUTtLjlNnnrSGrKKV+w
YqR6Ycc6YWa4Rfrhc+APOEGFU6RFlUhJK2uEypH0x16SzimXxOUjDGEZYLUKGZUqTKLa3Lz4Yln7
vIhuTZQ3nxR2VrLuLXYu1CIQk6iVghc2+yNEQpTQ2XmTNpXwqHJGslxHAqz1TQ7oJMa34MYndYmH
tj+IAfr62S5VZpU3DRE+nxeZWHsv8Js5XHkEOz5Eom6K56qPIRLfZPwnUEnJZ6mVpho/1nwSOnSp
OZmocMafc2nGwxkLTfrw8fRlPOq7SFHUo28BhfFmifvKL+K7g8aNCJ4lWCCYp9s6e497/QY6iDnE
RavoN+U3ZtXtPSbFrR/9tdjaZJE56g2Hkb00nFgkxXT7T+KmCpEcK/4uFCxUQm5P1xjBz7E2HMgz
7vjUhjvroHDnfgwclO45uHeskXBBwKO+rxUe2u6B02d6UbMYC5dtpIp5kVezd500faH4M7hfeMML
ONAJyZ3CDUG0s/RmGW6G3G+oMgrRZufVsheb4GmyqmwyFEU7xD5ljHPgDIrgNYj5FC0KIBh0bnDe
blqs9WnMceVYNw+a3GhH6JR6UxU2vBL9PzDQ9nx322MgELM0MY4b8o5xPvdz0cwE91CpTcI53ipJ
rlFectgGDU/FE9heVquACPBhmSSWel/Q0kQP/m310DKyhzA8tg3O+zIUN6AjgKVW6P+UGyxbMIik
ABgppvvBdCVv2p3HyA+XDNLPI8K9Fk8w+Te6VbiSWF0oYyrsu6zn31L7naJfW2dFb9ToBVvkPl6k
eqDCkmpEo8MY5hT5sAXAyuiEuYx/FtDFvkHNEaMa2yxZbD2c/HAOCAoC3ERd7HHH79jUw6v+OeKC
hWKbh8rpuTtKP2ecPfPGgUB0Fe4aGuButM19swWh9NdT9B4pgBVgKMyg+z1QhO0HWh5z1XUNL5rd
VNaEtx7v45vPWhwVk+XHP4vCY+bDFtiu9hPNIkWg0OHQqDcwOfS5YkijFoLYoDAZJ2tezy5vlfJl
tje+fTaQ/c+r7CRRFzE2bLXb3lTj5z/WYiJa4GZuFfV5UWV7vS7IVjCHF3d0eHCuYbDLY0fILYYg
G7kzLja+x+6U+FKwI5tKlAE+0YVfhSJ7Cd8zaGAu9uK+tBb+gERkPIsjdguVPkZRQDasyf45oG5B
c8lX8osGPVAdQnW9Qxf4x/FLGYv6SpYUUToOX++JnsTYdtXf3Thh0626PaWPfCt2TK+hmfuGKDte
o7dXz6tdemAUgTgrcEnQGD0d3eAdui2T5VK/pYsFX2rOR+NCzikdZrRCtM/Uxsud7ZH8i1C2wMEU
EBMnrOjySGwdgODml79LmaxiFbVIjOBEWO87lTB9J0ao63PsFO+8JhaCZy2XpxaUaWZWObYbDtrn
e+GBreMc4bEKaQ8+mEjyHwxqakuBaiUw9kZhz0geTJzcbIH/3lNVPSwhRm6I3T+S4r+0iNr+Ug45
SW9+ubTeZUK59OB+HbDrsdcPVVLzc5EdwcaSPX/Y9wRvpIHKe5BBa4xycD9w0K4zqFuUREzLX5N3
EuxRfDeYungvZZ/OsORiJIHLtMgwER1rJ0UKmLX7Ek1zao825lgZf2LDLiDy0rWMvsNos+nct42I
hlgV71XOr+eBiGfOPeVNVnNg/pPiaK8QIQdqThCbsou8jZvBJ1S0q/66NLeXFsefywHJkzBoFLg8
ubBzRRYxY392Hs6N52LdKcPJjFklS/iScB2ABWz2nl9YuiJ4vND67qAhMZ6iDDmvPlLw4O23bNqf
eG9BBOvGO8SOHGKFCZsGhSLAvIHxOgMe9SssY5i2u2L7Oi3R6E0iZ47WDAwbd0iKN3JdAYWMvbns
4hYB5PRX4nqHUleuYCTx4BuLm3srTInGaWfKPtLQrm6+M5kDACkwQdoNcklJ6YBO0XAG1ymFmpbe
jkJd3cg3opzUrLuiVwhmg21ebaUVKd0pHzwUzgmhIGTlF1sBAJifEnJYU7L537yrp4+USALtj5Gp
417x+PwCSzqMDhQKjS0SGjIB6hfNYZ69SQ1b87zbP8BNfSNkga9vLdWxCHPzXfeogFosCHM9dHGF
tmyRfhLzP48Q8QWzeW+25SaliK7rX8Gffh7NOdaHRmSUfwGhgo31KUCnDBiKT/+GnBDNt34NH0KK
31IP4mBfoW1weZ3v1xZHaedymE8h3Wjtk73zAMwaa72WJHKPNexSjqbuLAffN2j4MBj0DyLOYDDn
JCIjgAPguY/Udz71CAuMaHZ3UMUlZ3djUp9tzJ+kQyydEaEp+gy8u8orucZRiHc8BPjUD4qEwKYs
K6kx0fAezmXZ4/x2/Rtv2SiAbHKIKxPkkX3D6JVuin3vLnjb9Im9tEbjzwF4nYuwHWu5kEQRNzfS
gNQ9tfs3C0AC28VrZRfIP1xcnSGXWzJjSL43ae57RT6LOOjo6z4Ltsm72vB3/JNLRhiWAAHHpt0t
dGBHkpeiWvFyZCMr1hSpP9lK6eqVyZZ8z5BssZuywvi5rRCszTjeGY5ffIaLh3fICpJaUj6AhE/i
c6KGdRfeKLX04lzsueW97HU9ha0DJ4KkdoiZ5nwVRE9PZ6LhNZ1xKYO5Yx+vZLH5K6srIGdgEVDF
3eF0RuCcsVDOXbgaoBGp/vshxNY6ONofg1kk198GHRL3NU890XUmllHuhazMQqxckJjZ7EqCobVm
skkyTpz2YqvgdPCtFKowXUg4Nm7T5suxSNIKTf8vPe40O8WNv2abrneSRH8WHIBDZVzRAb0Z3UmR
RbydlXaSpMyQx2TWbTwBzbHzbwXO8et3rFFZelUvykdCvdThHVHJ2Opom1gEAOH/7aEUmga+RBJf
jFt4fFlvmo7zPCW2jJBpA4t9emHcLwO8Gsa38TLGsrnUopkrs7uDxIXqVp5FJWL0boSbRfBJwTS7
BWOmnAfzszLmXq2A1XNp0IKa4XhPQgcCZDwVUw+Bry9PxoQhdE8JoeZFBO8MBPRbx7jzI49zyOJ3
3DzcM1ZA9hFTlUDqZqOtmYax+LNDoyiJGuqafhPJQVfhlYC/gns606RPc7vmttgavldaEc9aS473
O337/n+Bppom4DhpljF0FNIiNyDzUN8Pi72U/jkE/yto/evlnJvoLMPPV0bvmHPwsP591KwQW9+V
kYDkiGCqDRzM0AiYMnp0Gw3XbDLA4ncVCmW2nJ9H/Xo805mfEQzGgiyRv4QS+q/aN1fIwBuEVsO/
icWOAQRWspN9KOSCGWKpyBdGlSPKLHBnUCHOSTElA8Fs88KovXKyPXgvWo/DMt1TAzop7puMD5Vw
4lKHU3HOjEnctBI9UNFQI3PwteO2HekrV/IH38I555iJp1Q1QmYaTiFg8J8QY062FpKDk+yJvmD2
ZWYCa7DJxLxxchO1ujPP54dr+cLhEM9wLyTpvcoThMTTMEm0wrDiFddspWkjPIUnz+1asF08SEos
WrOb5W6ViH+SN+/al9vF+TfU2RYoDJqJTYgdzW567j2PxNSTsStLYj49aVroeaGZV8FN9b52HXgo
aaCjw6WtvvnikLDkQoa92vRnwQ0jGlUr6moBnRotS9Ar9zoYdvc5banKADuNtwFgWW+5p0ohm1ln
o1Ai6ywkslFEjlUJJu/j8jrk94/XHMAophzc1r0qVmj3PZ0+ODd/X6Spxu5aKVi4eHu6Z8SHoSqG
2WanINfP1hswi5dvNR2oqrHIR7s1HWBGzp07LRhfTGzbkjtqHetwNQbmBmj67tsp7atYSRTRoFcW
jedu0qkW7y4WIDSDmHCOqrQTOdoZyIf+hj9BZqew2Io9BKYUoyvQI5cjaTJEKYnov2BhBRv5rJpz
DK2FftbiuiVryPtfC0hzDVACgsgd+jUCieaxibz4RsKoksCpSG6FaqLeS5ryJR5OUUtro85FjGyL
aENOtYKazIsdS74+acdT7hEQbdlb2dAWDN7HFoJAESf3qa7Ix2XfVGtbqKArHfXqeVC/cUpZ03wq
4wgp5SHsbVkPqDg1TuqBFOgBMUCx9CM9MkICXBgNbsgTJRpD2PrAeVXyBXwOGQuyUUBzwA6iUapm
V8TTVmwlefTfCb90mA7WDBofCMst9/AAsUC1DT+lChrZN9k5GuS9IKVzqpiZjsfdJgkogSJ80Osv
YkEP1r09ZIzXCuqo//tywhUrUE8ncu/2D/aliQkdojfpETVpE4+SOaKkGFmoNfl3wKXtUO97WDbs
JkNCzTs4KA+oNUQH2XTQn+h0/na+7H3l7rs+u9yBRyLnIRuDSXUBEL756h4lZuPzSbNp+Gt6iaKN
WeV0KmXPGBSg3w4ATG/jkAjy0TL6/9Ep+CHLl2aZazmpVdvVIUxiMuBapeQupp3aZZaAymXZ/mfp
+DKn+nfkmz/NrfigdDNklUuORJ97JDt5+3GvObwIOcoB+k3AhHjmt1SHldzt/BF2i0cvJBb5VgeN
wSKagxnSc+OjthxiWg4JadS2rjCGW1cdwyNb3HuFwKyfBBj3GeHUCijZD0VBDxvuFo/NkT7sRTyq
czqeJjDwdfLkJrk59osTjU3g4AVc7E/0vWG8I0ZfPgdyhqpZ23ojEvh0MrPRvYG4Y0glRNUoX0fh
e/4HevwzDArQKDwl4K62Gkz7t7roj4mVZKUK48VxFIyEaxFhmcOJRFFr/cY6z3WBImg4K2QPaNlC
RxcDLfkI/LB8822RkDCkpq0CfLh3PcKshynDI9hCTldk2QYx5yVhZ+S8enXnr0U6N8uvZkRmfW0S
9CZtQ2abs3lzDXdpPDyB2s0ZegFgugyGe2KAZNqQ2bWD3mOexVJNWOQJkZXzmz/glPBuX0oNYX1m
sDNlwObqpwM4JKK/QTVtGSqSnxnh9Mrdg4IwE2z1KyEp153dKngKKSCN73SYwSVZW+YeATQ6GFOu
Md321NxvqjeVzuB1Dv5nT/3ynLtpe/WktPrZHixfLclWL1mR+kKMW3fs6/BCNlmdpbyvIL+NNeK/
Vxw/MvqpXX11ltDDQmZ5/zyH4tP08zzr9ZzPHewkYgdOiWHkwQpVLHAq2BMBsEajyRzATBwFOTOS
2ztBFFb8gPHjsRX5pJ5mDaZhBkr9/8FFPT/xisgGePVjhLYw06cYBL8zZxY9xRt5rQ/FCZDWu7CJ
qoj6Um9z9UXl4yRsNnMKNcDxP7klO9dMT0YxUhXz/XS6bPqHCuIgHPs5xd6F2uCe1i/lrZ841tkG
2UA/8oN1zPdFqybCO4TA2HSRuR80FeABNbtFSUDWWU7qbm8Nyp3dV45G2vt3V+WDYQPvYHoRACy0
glOZ7TzQmRKs4uj/f0p0n3ceik8MsB2SSQywK6GUk17GGUduCBo6H0/MP+IBHyw7RFdddxc7V65M
xIM4mEO6aepB/zEXNXARhLCEfV3E+EpQc2S7DcouJvAyI6b/mQhC8n7GRboACDLqCL0LGT5lnf9S
iq+Oev/pQN0mJ56IZNE0NPMd0dXYtQ9iPVrrw4HNLZ2SPBvRk38L38v3YlI7fnx+6nJVq4+gO4RC
5ihjDgEbsBgaiDxKRIXnlujOFiSNFQVruLA5U/w84vUurb0A/cSrq8H7mN2qlJjnOc4piL/swpdY
2PfIzvVCLrkwoefl7mBETQ7qu46xi0mohFnYhzkxTaGRu4sPLAKVd75ul51rSRmcY2NKowmBv7vH
1TXb4zZa5MoIc5ouJsFZGZoLPFipyapWtrJmolof1NRJkiq6qGjXBL5s/5x+qk37bZ2iSjVjy4f9
6Wy+IOpl7Z30Frg2+m5dz7IesxWMxFv0FEBMPVqaY8RX2EeG6w/tKvK/uvWNXj+UDeBbjGL0Gv9m
036Iq0nXdv3FynzCYaBsRrGdpmFJ931bM2tsKnXx1kwgKRe91by5hpCk3+HQZrFBtGUSxiDMHESx
yUDJ/N0uuNnp6f6eWbE7Hhdp4qtEtg0XInCpf+Y7k5PC9YzTM7MKRj/peRkfW6sxc58txRUY0SrZ
r82GvXzRg/V0VuxsGJe5319w/Emb0TxzYt/XQRnh76QDkQb3Limk+Y8F6s3+KP5KnKNvqatF8FVj
/hpseM/mGHItJvKxOJyAt4gpLPwHkIrvcrK4HQFs3UNRtJV9A2f1Z1bVveBS+MCTxSjmNaZ2QRYq
m7NiYZk01mreAVo9NrfbFJyO/djYInfqLyfKdaCmNGn/1nthLj/4Gsg7c+YcdPflZ+Mtdn2rjCaW
UbXqOfOyiMEWhntoS5MJ5+VAIQf1nyBa049+kF2mAXgxmym0dgh8ZCgPA2aajDxoE5gKGSukoLJC
pQR6E4TQ1ETRg08OOkZUptzSOC7yXhIH3WgJrVuSZxXKGMsNMRi4QS/iMTePHk9O29u6zUmX4Adf
uK0308aLmD0cZPW4+7OXuIL0qgWre3oQCd5LvU0KrjM//qFMs3Qctffd78iHTXCSarAtgKsKmGBj
7O6VrUXaj2qWgTlWEpxPm/AMYU6uV6toWl5rCLpr02Zr7HgyGQK0yViO4aO8p/mYpKtuXSj1xDdC
NabD/cVxtJrIYpdvF0KcnQ+PxlJ9KpQD+Lwilv/X3J8Y82HZBeiMMQSuYhvlxfdi/5OWz21YLKPa
+xkoGANQSso7MeEGejmnfhW4TRlRgQyYr64FDkvwkm3fVz5Mitm8G7c0QVwJ0Su3ar0maSjucLUq
8Znx00obbuwxP2g+LU4lZIPBg+169uelwhJS/szSjgKM0L7Acpdsq+KbNSyllssHAEVpoRoga56H
jk75hAPWBTXUFupci9DqIMw2ZQx5K9SqdFoatPtKubRbx+TZuS2Ntav5gJU3CLdhtR+4XYdGXssK
d7uRCoGocYryVxyWb+2ANAFTjtN6y9eucbM7gVoG0qPuMV3pdSDc5BXpSXmRxZUYQw16/sfy7sXz
7a/rVAv865MJjo3wm7zPJtJ/PVKTGEqQ5DZLh/v2ERlf1XserzdU6prYhtZ02aFwkbs91NXp3YQw
SkbPvvRNnW9TsR++YZIubB14btpeg8zehA9wVb3fMAoJVtNIszTPUOHmoaIzaPKoXGPWG6xgTBJZ
YqUmfnOg7s84bkFyxfUhFjPLbxnxK8DaZHwns02Onc9yD/2qHo2FteeIyiKflX/X1YiRLThyh6IB
3bINoldiQCM6HFnAKq2CMV61B+yy8ycf8O3AnBrHdRGQ9IrJh1ONVxfyJ6bnjJDS1lSGQe4dLV2S
nSzmv6KYnjAJKEFsgLnAHtHtn3MC4AeNFeqTk+M2hQ0UfAz8VdccCTD3N0ClEajGUwSQsV7O3IXr
8J9Q9BiQcDt96xsdgqLdS9OCdY6y9BLNYEmiqfL6GR+TOnB/20AOQo5BQADd/oyEypfOLJNI/xrn
KfDgVG5Yt2IgFElQ+Edyw4H8WstjbL01Q/R1/8+WYLkcOXQpjtOm9u+KTJiltx7vpe4L5BrHhv4D
ajGEfefxo6rcK1SRzUfxLd6D6ezWAPs6JpxZcsKmCI7SrSvXiwuhGdlSnUeTCByyMeaDOxUUsM3J
/ejL1kV0+Io1Mhp+JVK3oSM/NBPldihMkKYPoivw5a6z2ZL5fzg1qYLP2BRjht6ePunzN9MXQraZ
b6qTTmwMbZV1hp47XfyGgl8wUJVYrhxgE0d+QtRsSB09zARlLZuOVpqm8T5q6tr28zEcgZ4BM/q0
mq/ts3N0ZGD7dhf0URBl85u/51QiM/fD7iUGoAJYsrYBQsFkCmkAExh/X46HI7c4rRIaXaNYCmsf
VHwpTLxmig1dtFHzFeOyEDSJYu5AIF3zA6KuOUkQKCrGGOXA+n9k9AXzPncWe2ATvoBizJZbG2c4
LqWOEO6LZXH+ZazAL4/iXlyzC9bR1weDY7siN69fajG9gXu9TJYShdfLhFtYM0epmwsOmEDGSEbm
2ritf6IJL7kzqSJCaw/kkgsUHiZtnHRfVeZYcd8kRP2+Z2ZkDp5MCLDO77N7kNnY4NXNXfq8yz2f
lIQBJdx2qgiedY9wD2v0bSx5l1N8a+MRpeBU1MlpeUc5bHJoTrswRMgVXsgoMWRCnDDy4sCyeuEI
GqqYDtp8GwpWSXCqvubOBhykeq7yQxf6l7qzprb9Qw5YID5mjEa2D3zPqZpjFwuGFgspJv/uhKb2
qFQl8aPX8F/fVaBTuiXIpPSV2Mhb0EmRDE/qG9dEg6I34ydlu2KNqYJEfLDF4EAuLWPj5HZm/UCD
bl0idN7MK3pp0rD9Bfg8+U/3NiacRODJH2NyY4IneO4pmxV0KV7EIUg06Kry3JGHtMiY+kvm9fSb
NP4xzlDMsMXRobW7WZv7ExEN9SLT1/jdiIRmhzxPHuoP5NOY5JKhTwn/AfMC2N1y12pI6tbPJsyu
9HToQY/mBBjxqCOb4cW07a2Oh+DuPQo99mG8/MkwaTW86xacu/cGFRf6VFSA4Rw2w0yE8sQ8pHAq
9f+9S0ih+ByeGA7jsHVSGcn807NdD/jlaf6zq74yJI3BlMxrnhmkW5/LyBdlUyE4hARI01tHzyC9
B/ka807SKs+CkClto5jg+7uGh3ZQ83DEUki0swjqJqzwche5wT7WZCCF6Dd7JYOfjytH11xihhd2
+IBIEW8yS0bG5Z8dalYJJ5CulNflMclH/MRUKo8R323mKoDCrLsYBnHEQSNpvpS4UnMcVOIzW2aX
WJypx8NG90P6ZvCR8ghqkh28P7gTVmaPhgRGgRVKv/5PRGY723xqIPHYJFF1WOxbhOQWvKnQ5TdC
Zg5R5rzVpFs9L3RT6+31FsbhiljKgrs9VWJSGqa8fYcS6pdGJVXDtCORuZrzmacw2mznm5dIRZPa
VwCrMvpnmv/ATzwcZYqAEy36y1TqiM07h0DjeegRKNgBfrp2qpENMPTYLufm7wezGbBIL5D7cbrs
xhwJlq9G7rbGXoLPCy2c7GxphKOC7CzwkQeW4zr5z7DqECOhafAXXtwS7erpXbEGMHfnev3lx7Z9
LkSH0SDiGo8C50QREKWlL/8TXP8QlgrJuvjjYy9q5x64SGgMt85syFqwraa4d5Q5YHBAXOl00PCn
R5wtj4uGqc04DBi5CIuddZDkJGxMuAqqVG4cey3bois4LfBRAY+JMlngwYDp0s7jsziO7BNI0DZ3
tlsRRyLz/mUwSOTwX0tBbYL3uj4pC8mAJz1DqZGZTi3B6mrCVZJ9GAzkQ/B34FrHxCJW9xz5SHvI
GLBTFyUxh3LcShSqY4nZ2nIPaW4544oHrpFZE5y3Svs7FsK8fvgqIzobQHybs3OADoucHOSBY6/c
lAxvgqQ3J1qu5Ag6piLbWAeaxkGQ5SXGmiFG5+WpOsyxkUIy9fQP4fQTysIjlkZSJmSxBR+SxegQ
msSty5Rie91V0DM7D4hxEWZIckISKEsxn8tLvGDvi4EnoNmSuqopTYYPu2zj6q1uZXjvMvHfQfS2
em5kTR74NkTaoYOGKIIHxvHmzHJ3cjxx8Tip+i9+HhQIBW2t1wgiNEB7NyIXDFqwVdNpjqNT6Or1
34lAZonFZsGYkuJE+tGDYlrazF0lnHsbFeeI525Zp4192Zn/BmaZgA4uSfYOaw8Mj0I9xluNS6mw
saHPpZp86BGHu6gIZ0s4lTfqORFVuJ917gnnOaIAn+61zUjKX4Nf/0juZnpGCjz+E0fHrUUf8UV2
Vpz2zcU6bQxqsjFto3eBc+e3AGgTMa3tF5lqh993vE+qCjvNU5X1Hvv9yv58hBTqm/Ff6cSfEVVE
Yr1miQABd4j9cegzMTQW0UvFtSn4Rs36IpqjJAOiwq4lnsZglKzYggbB/56M6xMkDtB8XhJ9bB8Q
sKYvezQMN18XENmZudxF4V9q927vP1x9EdSgmPytp4w9nhsgoVP+Jp/LGYl0VNiINaZLzy8IsZmZ
jZJQs8c4VKqc1Wpm4P4jxrvwirLCx3Jj7+7u7S8vkhKrWc824b6RSyh/GQWhhocJPM8EBlSHtMx/
j41u8tBC+ThDue4l4FBjQodDVIJGcMNqDKyhrQqYtVmbcVGlwTsH2lLielO8pt2iIXKuC3FI73+s
2z0/QCko1OIQG0wMxjKseLXsAsT31rFCOT4GNg+hDTqdTl17XwA76NhwrxPnU4UDU74wdi+4/++D
a0MsB6QNuu9lA5GIgbkfwneMdFjq1AYWVO+skMCMOgEuJ1/2xxISt+XAz+zgvzw0seV4PYU+9dUq
xJqnqDRQHKVDoupXuczR0kuJdjGiGxlkpP6QkPipWOohvoj9iznvgEK3l8S0YBjRSM6x6RXbI036
4i2Eclhb+VAzwNL98Y5grl+o50SIZX+kUTSfnVJnc5We5zAVDtU8kcfVr+vJxnYIgTHxVkT0PNhW
vYZg3eZUIF0hbjE6/6jpJQwD9SaDbHPrwoOv42t04BTVWpRbuAScDygghjOClRi9ZJR6o4jSmPLj
BJ0dVssOwZa1iaW77kGnl28fC5ZeVb2J4QqF9xvvCEF3st1/Jkfi4frVAYrMNIArbFguo4p+3MaY
FSCGlDcXdj2fKpyPVxoVC54jtU/CNVmRBSHU0IsNXkPI9LQYb3+PzCVMRYioZMBG9k5WRinT8ElM
Jl0xZxPpcBdBuSD8ku7nxHHvONmZE3xPrnjJHZbja7ftFMz0XpzwZIv1i+DpDbs0rzfzkJ93HGn0
6Dm7YauW89NSCpFE/bTC8jWG/xuxf/SgPHBgihIwlj32GGSb2KcRWaxt2x9CtJ3nBwaL04plXJgL
Tp2X6SCpzV0d2C2RmpR+9aeQDbE7GVUm1xf6X4u/x/2MALfa4pAxtLRbHQ0MAsVry8IbkDCIHMPB
SpzX0iRL/++CQuugTD+MyjkRzltD+O9qC+RDfeG4Dy6/1CrIfrxPjIWdcjR3NMTEQJs2TOAW4ftV
BD9KJuBWOmOYO7CciH3OYrFphQ5N0/9rRjJKTf4pq1bcDYT0gPm+kAJN95XBjAkqmKpqDBaZGXOp
XAT5LbzciFlSlls9EWtjqFeVLW/iil7q+lMBLC0hbEcLu8kGvpgSlj2c9Hfa51sczsTjvza+FVEd
yy7Ysx2UvJgMj/MiOKWih7sRjNofhnozMDTGRl5Z1Ge64vPJ1IyI73Svn8bn7O6ixF3r+hjWMQCE
jyicM9wGsz58USCmG9IIse25jBL1rdbiUDHroqGGnzyxUvBsZyc3laSQPrksqi5SX/Css0MUZ+XF
PqnV05t06t22Y1cGYVk9Vrx+2rMnhTysNzp4KZ+w8oFMYt8Kqq+fpXmil6NrrUrMZYcrdkTM0nQ8
DUPEVN2Jal3dVAo5eQ5qz9KtvBBJ9sqyrt6O5iEK5IYpd86PifsSrkjlir1/5FZzMNhHvQLm7GQM
GmKL5Ckst+oTrNlmlsf78HaFuFHlflZmg+Q6GUw1+zojojfaAxLdfBEsR6Q+TAviFYAmCOwn+ECR
0FB46xuh0JZnlEWPFlCoZRpOmF+wCDMjjau8pe5wNdNMv1LwiQgJHJ62n/JUJwdEFhiEE528HvJZ
SAvB1NKWPIhcyf3I9x8JUoNkTqKmYgAOtnU8yi5uuJ8x+3vBNH4zg+KdHaHLxaiCBbmDUDoBpR+d
Vx27+6v9WftqCyjavBtzTbe/0XN40EeSc64+XnShBZLPXF+AzdG19joZDz7eg3WdWMTdYu6bnreI
0sK6LGBiTfoBelC9ecNeguaSmCRAHVEaR1po8FTZbjSDRB2vKn5eevZolsK7g6FR1OaXxfAxvOE5
SB1aD3nOlexinSQdoWiE8zKziuk4Yl3C93b0aZO6H9iD2K7k85DLo8mcmYfxAbmJFX38YC0+iIeP
14kmndlhg61v0cIumx4dFWzQ9C4QKkiszqA3wtP6cUOsfiIAg9veO0REaatPlfODR2sBjXAR7WZL
WqOvU9gXnHem8Aw+12Xb/SA7pQEzrYzOzA9cCra7QmxMnvheSwsulPCt9rRdBmJ6njbb46Enfe8o
xFw2hnUxgIrcE2jHeI0Wxqa+86ibxC0hw3noZpkOxx5sWKRIKqOSUs9Dj9qjXDBXoxA24Gm+EA5D
ICncgoOoIHf0cxh+Azk87iclGAap5FMAATr5iStbMJPOk1uXCqtRlzVbPlBhUZZ/vWjhOSUHdIy0
RWPHmkYMEOI6mbHE18G7WzkzkJPwdnOGTf7ndq/eCv3p/PBeVRG96D5GPnUQavCPRVC0A3k1LLPY
9BuihDiVS/issQvwwUWcXKTzMZD/QRnv/Wwr273Vfxo8wR5PLxerPW5WCYE295xB568+6GUOmVUw
gUG9Sovy1EN4pYeQjqwyD0i3oUF1diL04zq7C8o87fwlHkGbwP4Y0LVPBNALISsBmFpetV1LIum2
6YtyEIf+aaLTW9ig6Rc/ahVRTevEyfJGOVqomB5kvTJC2DYYyXeNgebSnp3vzRltcmLANWhcsaFT
hZ74/socFL2UFg8zv5JjeKRdpn6fu4aqu55zUYcm5jQuhmu2FuVQYEr0uFHi1Wk7mizUOWYGkTFV
xQNpZGuCDkPkuMiFVoemc5K6i595E5I10DLC/QVHrIBxN5J5ozkz+y8QQwLWAOy+8kU88lM8jirr
2yB4FM4RB+rTyfOpZoVyjxGZ8p2iO/3FSmitUtW+dviD+01bk2uknF8eKr3f8XSociks9a5nVyCV
BBKDRgPSb4diIGeut/kSdbyYvqhPfM4SX5qYWvBgKEAEkBGpP3Md2PoOIHPNMP21Cjl2fH/lXfYB
rOJuJ1/HeW7nQ9IPscjdrMRJj3ZHshMSp4D2CdjQkwhtTjC7B1REXqYY9cxuw5t4cxoJkwojaKMh
bPcK+qzJ5TTbLA8kcysKU5HGcwlsQ0RyIEoHpMzTmU8vcm66oAcUpQlRpD4rsZnqHPc+8AGB0cPV
4eRO8rLpmEQelfQFw9uTrLKnQuWaUSEFHWUWj8l14XNjXFGaVM/zpLX41H+jHtq1gXNn4MAIzGnw
y5sdPVWAWPfWuXsHLBfpAkgco7OoloxAntTy4vSVYuazbDKZtLzFdSFtvVXL8Uw4mDKO/ZsJbFg6
lFndVk/Cjt5mOsXEU7bJ4GG6BLWWuCK01CVQ/mjyHqBRqT362aXec56lcz6r5+vI+L/oFI7dXagG
gb/JleQdLU4gvs7LUEO/PV8FtZG4CDRB9EJ0FjD0cGeW40QJ+RJ+DXwX0SxqX91KHaZTyzn6W0PT
rsZumxKZdMm4vTftLfmY8Bc0AxecPRvRHL5ZKudeiokABoSfTyGqsEp9wMYdOA7c3EP3BbA1MOid
ObKQfD9qRwfUSuIKGcWjxxDBXDI9VEV+sTgGyAKqyBDLOebmCvN62NYXQqwNJVUvRn+9jGKXIuvm
J3h/My76rHjzI8xIoNO4zuXvNyRyEqRbRMjV+zhaXwvpUUT5RDSchpZ5S97ENhwcj8jUeq9lrq1Y
rc2SpeNHRV6nktqvIhsmylys/SY1xPQadyNydUNEyouK7I15OF8XUdkFV1wmeZqprXsFwqUlb1z3
+wpcEbRLTQ1tSw8F4whvZHyMdVj0xJiGL0vHYwYOCvALUhWUBxU79kCFsEo9gmWo5zK1/z9DEkV4
i6Yj6Xy6EtlISZ0QNkqk+s65A1VSnC22jVPkb8J/VMgp0x6M+x8x2k76bPNqQmIEtQSKYaTmxKMD
acLlbkeMkX2nfLbPtOl0pujZPcx9RejACcAWyh1KPxGDpdrUP/vQoza1tGTKlq7UrSGnIFVpWnob
lsVTW+FQtqpR7ZDmIUPqXuqOLidaFMmI8YslAk7AqXWSiXNvReKnJ70TNUDF4/6TWAzAfBpfAhRw
qAQncAKMl3q1FAe+wrTXpC+cDMdWb02NvwjSuMQu2gS/dRhtcX+JeIsadWhAdDNix85gnRee3Kut
hsRk8rHnHHX1vkue765+4AS6KwIH0mTNxdP9x+/iDdOG2ScZmsY+4GuVIBNZ7VFiClnwlMu56axl
2wu7PSK5jf8kcnP7Ecj5sL5Zc/X5dGwipA2gjWciWK/3f1/r2pPXyYaTObVDHKPF4eTS2Hlo7xd4
6PYgyRTRzss3rm3PSEa9sAnQm/qxZny3y7+S8mB5JKgO+U0q+zPoN00K8fJ7Ruj9KK8QDnTB2Sre
Hngqfzi1FkJUdKaziPe2tgvWCiwI5yyma59vx7YUgo6c5OqFx5W6NI8Te1mWcjudFbiqnZQiEtlN
QfEkkd/hHOHviTi6/dq++v7haQJ2jpAh/u0damn7w4iZuqas1mwa/fFlXDk/KTYIrpc9GpynxXGb
Vu0XN6fxHq4yDsak/MtBZn0Wv1oUjimVplg8Sl8d6rRhXOwwZ9C9LGuZsxw2A5psySFeZT5EL9RM
JrefuQW2bGHhOSeZreOLANHFHUwp89K+fgiiOtTH1TBtaOZBmIrZ5OrMZrjGsqieUkiHDdxnTpER
yIpdOcx/TTHai9a6yTLyTBYKkRng8rhS+MmfJxsJcKb2JLM/3oxgCpGgo0onAspaft/inMR/zFJB
JG8Y1dGrDoWxTmpd0OkLkAzxDkuh7Jc7vst/SJuemTastDTl8NdbfVYCyiu6L0scAgcyzoAH/arR
6TZDw9Lzp8f/gwtLVoA4aK5urRhAlgG8ekrCx+uQnsljMQd/2bbyIlQYushnxafsl1jMCvO6WpJ8
Hd9Ic5qcQKoVm+PmjFNaEPyMhb4cawqKpdPAaNAccdyFLU+OfWkxiV/VRdavSL728H2GWt51AefR
VwTk3V68cYkUPswSSzL9vpBaqFpFUjcz1scORTti1vg1TkTyepqvAHOhq41xwW9B/EzUuIVgxf8v
+oAB5RTZeStLVHZm3NIgoQMU1wLk0IOD9ZMEEPPX2KalrmFOo2n2/4BhvMk7zZ9K4VkLHNwPtMr+
9B8Q0NtlXEgwpTaPwWrwcRiOPkNBIpIjmR1nvEDDMmVXSWuHNZjGpgabGO5nvFWNTEQ/pBxfeQg+
6DwXUp3//E1jqs2LUz5mfMunc4EIRPC4MxIAACC6SSDxy3zG1D7zpAhVuIP2d6C8DmNEp/rEetbJ
IiDnOQlBgHImB0oHJWdZfqahkM52xhbqcBjXolJtXtAtzfKXPkEsg+xBvu/7DqvAjeupbXkRKYnv
TuiVqiY5mhvrdxa8PjFFRNMnjWqXNjH9AZzmV8wo13D+sie78N6/V6UaM0gpTFsfivcm38EZZBPr
ZqcFMjMpf2Y4H1zWe4HhR9Mpg7l7jfPLwY9eizW9ViTvqB5875OtJHCbul0jJxsIntmALeIhAbGn
+BmkI4fZStj/xNW6h9xc4yJ5AkDXMQqIgQvv8l40hg1Ep9KjodoRLW0j1HwYio2p7Uot/yDpKVeh
6fy+n2A95xRwsf52nDPjLXBjtwtr0LJejBoWxPeW8Kr6n7hCz2mKzIttJX8+Q7RBZpyPTyzRWUW0
Bj48j1ZzZxyxalY+6H6c/fMtKAEOkYS/tCM67Q6iAA7ry6AbXxwc+ghbn5hSWXXmOC+5PoLfxcxR
8FcjTL5qXNKnOLzEmKwk4y0T6K5H6siBnwaOaCUQlUHGfhu42FPdHmlpdeJZvntlpYSrehk4GOVx
TBIvRDA41RWXtspIqjsvWGnSuQb/NsrIEuRw99GgFECjyu8WkNSRPDb12TSzik3Z5QR3j9xgvX43
+py8rebUxLuYmYuqZ9NYYYwIvnm5CTE/RPnBcqLyGnnhS/WP7E0eRuQQWoiQzbw/2GNLYq6Qorr0
seYjMSGrEEcyOcs58tq+Mj99mPdFo3UJ6weWAs/TCMiTBWlk6rtCkpVZqWuY7WhFHXXhq6a/eoNI
deEqUZlQ0P0ZlMkFwu3oWrodhpZFHWHp3vX5MDbg+bBWqwOB4ZW1F4mPdz75ImQEtb5eeZSFrTPD
CSVLIo5EZB6gIv8LbHIizKCkW2gp08MW8EU2Tqw9QfzqKJvltMpvKro1qComJZqAH5x1XmkPx4NM
55xUqYZ7GADopdMPKR6Sb8lzFwGxVbtBRLcoN3GCcOJoDFYY+e49acjjyZ52GIy3DvBaEzab8UHK
wUz7NVh2wYmuAP6PjTppxlMxRJ6tjOrRey0Oy0F9SH6nvdw6fOvJqIqKxkeNI3IbTH4i+5xC3XpX
J5G65AXFZSv2dSnY9tgjioscDb1p6h1/hqUiWI+X6hQH7zyV8gsS8pCg4ru5Ktx0Q4GAfRp8cSDr
huTUlLzcOf5h6T3Z02fr0gwA1YGO/7QlAnG3EYAjiM8vwCXlalOTFgJSEkKJEe7o6McIA7HLdsHg
1UqZIap6TCfLrYJG+OLMSVfRh/0P0vHGTVbA0SvZbVXX5q857fI7V0ryNQHivEIGD3xzy0udIlJQ
vrtGvhNotftNsCiWGEOnPP4T1RQ5DkrayK6DNbcG55r9CTPuBBaRVAog3Z+6+B0bkQeVMBvhutd0
hGPJ8iHQLEL4yQaDl5DTjCYwidLBYBfDLWYc+1K4aCJmtjWagpx/558CH8WkiAUj6SDQ7OsYeose
DtEfGS+4p4OttbYNAUpdytILG29TDNh7vUiqMZDksn8cOg2RHkc3TcAzZ47Q92xVf4c6mPvBpdbh
VyUGf9A/LJ358W+FMuc2OucU6tOw7/0HNHFki1eDATRiKTfkU2jatAYGS6u7vvuIMPMLG97w3T1r
t5NKTz6CsHv11Fjh7vSwyy28HV2onuB3JqOHr34qcscaf6b7doxFuq0I/So5WHZlpAG0yU7coTwk
wcihd5QdwG0TUM5XS8Fu6PF0nz5RF+8fbYMvu6YtncBcXchvQRc2pCK1X46ln81XkFM8dodrtVqN
hAf9aelf6KeCYjHLAgoC1b3IUIMWhR/gjglYZ6Z7p5p7qnaBLVHCcniLMoDZpBFrKqmp5GPr5RtZ
3sqT6fYCEH80uRcd8CGEhN09qelCS/etHFUDJ+G6rUTfFP9IWXXeGO3IqaPwZtnL/OS3ui5jcxrb
+6Sxvfm0ZiJ5TmkiCsTlzAPyu3dgt8guIbdTzroTkxW0biZOU1WCP+LPLLRnMguWa8Qd5tf8tKJa
ae4HnmZVspNJdhR9mECvRllhsYO5dqNAiqBmyAWs+LbF3jBWMBlPhSpnEcWlV6yvudgOKLYO3Tx0
al9hr+Z3SlkmX1IgdIWp815IADOK60yeVwt3bqts5Kk7vcicBi6In5Ncc4n/suEbebjuHpLMlaL/
59tUxEwsnHAW+jhUCF9qMmAmR5jynwRRhqXXor+mE9z2iS8o8PeVjZva6Z2ZIiiQ8k3pQ6ZEXv+T
KVbPElhd+tb8JDF1/MDaKbz+xjQwMVABc2WbfzYlzXWuqmaBonFdSIJAcZiSk1YIiOzIYl4Soh1d
EoH4cmIZ/Xkdn8gfs9ICWoZ8GKLljWP4zS1Eu++E9gk2tPlmol4/A2d9n0MrkdXkDqlwXvZ/HF+V
I3bUdZ9fLJZcq5dhAGgmjxsdeWcByR6HT6szUoZEfQGOg29dA6V9ugTzB/B2uSktAMGaMJQ/6hxo
RXh+7mHv+4iTFVL+rtGngIoef1J7+K3/XmssYEIQXxHVglIbha9wZMdW5xWS+2wlTMXDhKkrkp2c
bP4j+9TOmTg1IZwQ8xU35TUWiS/pLC/6VuWEkEjM9GN4WahrOl+ZkoZmvmTlg2jLl8FggASuC4EL
ACzGOux8YEPV8WRkbFrPT1V6lTbV4spcSKYFTY1v6DvRDQH7MJsH+wkjseYj18kSY+EHI5QOvWKC
iCUX9ldfRGBNBf5fGk2ZGhz0BN9QURzwUe2nHGgAe4IFbbn47Qw3+wpTxyOnDj+pcpP/1puTvRQF
a27udu/tZKHG7Km8NOCcYdEZNa+j7pvkb96BjecHNZaeyDIGq80wOor3iNashR1R3psypuaK6E1I
SPkP9oqEPqtJK2NT84r0PIETGYfswU6Qcf8xfacl5hhscaZ9jka9TM96eXfaEopWfYisVdmmPkdS
HghO9VSFilx/5X4+RMCOK6GUrc4jz41O2IqslbKlrzh343iC5DH7zFBMxFSIaojcYyXSlt0e6RDS
swK6pOqLZArGCNaYQI3YndQGLli9fLQPFpptL6ISqlof/xXz/8DWQYGOKV6ZOxzUSgQvkhBproCj
rNpoEIYcFaYGm3kRDPbnjJf05/KE+ZvCEfvRM2/pCpKdeN4QKtXSTL70jJy4pAKSrqODbSLhRw7a
P5Lnl0Sh2veKmOAMzyIiQla8qPl17S5kahmewvMQOxVef00ngLnB+gYmoNzpdUNPJTOY1iivLd+M
aTOqNIIq1TuxvGLcAfRZzBwGUW3Su6ifrIfKRqPyIkqtC5zUYUga0nRz0ximwVg66744hhFMnyPq
Q178CfB2bMnUgiRws6Sth1irEUXgG91JlOumddoVmBNSe6x7D3f14Ssu5shLma/uwxslL5CWfUhg
R8BEyF+uJBpd+oA+I0yV1HUqmYVhd1J7ubv7WEMvoYaQF+4IAK1osEG629Z8Yuh6k+cJ9ny91oJq
Q8/tBqvORqgFJ6MiaTPjsqoyeu/waGM5NupFL2LyFIIhmuI/tMepURkF7ISMw4ODord35PugxrGC
KbkUNoZvbuBqmzjXHzcrwbYejkKbbB/XEr7o+881blZ39G4mCGZqZE8O4hbO189e+aC+Mam6m4Wz
IJNZWZqG1EaGtIFcjNjtNB4czgwpAUq6vKFzcyCe2nXeHevSJ5GPh/id3GqEX6WHVJKzNk/rZFCq
jY07Da7kyslGANoFvLFG/Wnmttv2rBt6wJQtMWEzHNJlBHKRD2kyAfsoxjvxSKLI8DBSl8mTU+is
SPC5RCPc2S+cX4OQ4Tbt3SO2CS1D3YuSzSIHIYionMqANJ5+vCgy2gfY2nkWNuTvoZ9l30hU8dW7
Npj6Ri6M8tS7K3AynuW9Gq9OmSeRTmIO7izeHwAY1zZyYHIqaGxpIVF/pJfcYqvtFFRN1vToPK5t
M5adf/OX3u6t9Mr6DSgtvm5VoHeZUpWBo+XhwAi7REk8ukq4wR7PAu5bxzIUhm05gfvYSisIiFwS
nlzZa6S44ZgDpfuWlhC3fjsEMRQxWuYb7WQHllp72vRawPkx78nFMdfrycqxml3nJ8jbwAIzpchW
olW6ujDloF7HOIWjIxJm4VbUbRwj6n3u5wJn204ti4aJ9mXQryEdk1OgMCsAp5oVmm3Co+LCeoLY
wwXTfH7sfDOEaIAv44NUnHth1YZLKBAqwuXYGdAChg9UShlHIHff0rhYs19FnGaraNohHJ0sye3y
4bJ9Q5TiLmXCGWANcF7NMOxAjsgZskqxjqRN8ETGQXgWRVJmi+x/SS05kJBAb6362VYjCgvUBaeQ
s3nKfQ0IVC8wB2doNqym7gIUSl4trovAeghVxSo4yf5xTqkTy+XKB/y7Mh3pBw4+3BNMp3Q6rLI0
pbjcT1VDUO2Y8VX3A4jX/VcBlY3HluVhejN074rxaAGZLe0EGeH58KNUezhs9O7kBtXsQAsredbU
8Gsiu81JCVpNa6LgKQODUWxppEwisH7CsvF43Ejk6y9db5RUQFdJlG2jwINw5P2riAitzWUm7VQl
sqpCNbRdziR7YtXkrB+g04CtBJiAwb0ifGC3vQjFSJ+f96g1VpZPe5MdSABumIX6CcMy8e0NMzMt
gKi1nugQoTS7fhf4b+I/iEN3Ivth5BIXRGMYHgNyaqADFhKisqyaCYWKRoujpGzX9zHejeKJymAu
gtiXp9sAsE+QbGUyQgWHWz/A5xqZG9QSbXXuudru6l/KEI9g/xDX1Ofg59DiX+XWGhvKUbqJ4eWY
xl1yTMMWOdi66Mji2ctN+JobW0hcvEJ0VsEQwzCaSxMUXavXI57rkPlOWjFz2xeKQk8an8/XdIs5
yF5Ul2Z5CLtRYGdJJ+n/Y8mWsyW2M0H+GBWA/6cI06TmzB9vgHR6eQcraURXJ9mFihVIykWKMt8E
DjT4TmCcehb7c8WOo9oFHXfOHaENkIQezVCsheJOmbwFuhkBjqIu0pOHgZnuTJ4k4XMYBTlELkgg
uS3qeWiu2C044bQqX5aqI5KqjMyJ1v/o6IefOCOq0ytWx/PdgRcJGrGgn+mRT5ZcVrY5Nhj0V4JK
u6gw6rcbrxUU9oXl0vIhsWJZit/LCrCe6hgeY+s5q91roPUipfM2EfIw0LpsljgxvzfOMxkOkjTo
auJ3aIKWZfeoV6IojZa4VNmLEekeuUAz9tfV+p73zfRTAyC/lkja3gYwiEMqPRZZ2oARhFjTdL9E
1bzfY9vLlEDWaNCl7tdKw2jBmleM1JmpLT8ojK3BgL0uNyqXnaq76NKEryXLJpASqpTOwjyWNKQH
YpLr/YpkHshrQ5jDfIPf7FfglSTafWQlwhvD+kVisHtRa5uYcoqMc+qqbu1Ococik/l6bAXNuiXZ
Y6h4PWBVMp2VDsIOBp9P/v7yILHWrcg4Y4mWS8a6TvncZDwiOpu6bqVKLgVBN49RcWSp6PInysfP
E3kEXcdifaoA+XcAIv0gkTXnbXjMoL0Q53+Q0a8k/HEMlHca3oOtZIlSBYr5pbWGwWm2Rmc+WuZj
aMYwhwdiF5fsfjTsB5ggyclWH0YY0KrYgkMPsHy/rFwDYegUXb+z5NrR59d6xy7zVR8clBrYmYch
LJsORf5wgF5KCMTjvZS2PlSkArAMy+Pjzpk5q3nXunzW0+nuDJSloYf5BmeAn2SIhL7Sf9hYgGue
CQhsXt/lD55epOArkaxEhJxkPJA9VciDj0lJMcFqDlzThgxLww7zgWftknX2IEJH325ihVtWW2Ux
ODZm5RDcfQkXCVs4VpX1PN/iCCmGc+GN6QUWgA3p7ktrGSBLdQ8LC88mjWdrzPZmUm12ZNMwBOPf
3o8gEi5S9EN/yyHku1dzt3oVWlMph/dzHTZ4tQGO9LBpByAh6mtQocIqeeaFV34je9ySAymDqxrD
exbsjC8tORkE0RdYlE1/3Vbenn4jOz6Iz8Z4TNj2KnXeGu0PSA8icVkjMy8TFWOIMQsO0ik8aTWt
EKliyMi95jN9Dq45tqZRyOjawLhHHc9LZaJtc/juuThyklKJQs46hWY4VHsjG2qHUi06vpDgCFOz
+BHU+URWO3Rl+4+Qu/HOTqhpTx8nzO68MjdkhZT1JHdFYPRhfGFfms0+er6ajGrVTcye08j2GVRo
yaDWa4qDu7hqWL5xTZHECln4MBt0f7gm9IWSkGdYl7vp9EVh21eRfysTx2GYwQuj1Wx2WsKQv3aU
u7OVTClFukwtyX369qdXn9lda7J8IxFcG8nMhk1x0Zdjy6hwXXgV1ADV5ujfgBdpr6OGSs0vDoF/
aw3l2O4UPg+GroDedH7pNmPm7BlgKOCbeYhT7f2TIUmj03/iMppIruDh5O/hFmwJuby4WznkTAlv
omKUJbUj10a1WMszztND8SIzgPmAXh0v42GNTkvEuxWCAAVIopAFHdQ1BleQHN1rJsKqQciu3tVM
NZew5huRrcIXwW4ruyat1yCswb5uvhOkRwdbk9Jlo+z4AF9QJVLWcplAxOef9ncMcSkLXda9HE2S
pT76vssj4dchkD+JHiPt/HKprayGKOskd3S1Pshy1NyNgX1SSqAaRz08PbLBRFI4Z6SENKRcg2rb
8xc1Qbo32/Q3IIR9EL+kUI7K0se0cl5bpKE+LSWo7vMR1j8m8PyRqwTDBO28MefjiwKycf5UviI9
DoEnmgUGS4B9tqKxg2TrVpVXoG6ackBVKDmfPuCSgOI/43jacMIVU7eX9jIWPTU5WgZj0zrDNMj3
gEAlWiF5buWJHnlOl8vsOHmdZLpbuVYQgmNyz20snUG0OYuVqA9VrOJdR7sEmo1vadSYbp+yx+x0
X7lKAnwvr7nemHA9oZqNg/lg9KjyTBINL4rPnyCLEmdhM1mEyk/25bEIr3wyWrM3Ck/WOOtainIF
/wspZynlfZq/51e/tbjMAXaH8uERlnj/2afOhPPHkyQ+WSQ/1H9DOW/+eyGfOidbFaY8XUioBiwu
6EbY/GkHESp4rXXu1lYdFmzYpcWVQhtNRNvajQ65wIlXSXX6nPr+VbdO3Gru2tV4GdiiblB1NrBG
LspJOLMahU3gAYPLCM1DJ6/SN2iLPgUX3a8/8PApc/Mkn+rWDI08A1aAm7LAh8rBWK30POM8jYZF
lBfHy7GcFa7Ou7ZF2yJuwOQBw11DwvYcgqsS7G0fGEkglMBdF5U2x2FkRbnpLg4hZAwtJ/6AwCf8
VLI/GTuQfsQ4p7OBwBzdDYs/n5a1yLzVG4B9QR+rZIiD0KRQ2dv53Rn74JvI3q1YmiIDA4msmAOi
JKtmz2UsjjAdhNsAIUTyW7kzVpze2b3RVvj4kjGzuulOx/CZ/qrhrlbFO/L4ggL5NeqISRZO+4mu
eadKGzhJh2lwFdR+GmrRSSr04vf3+99QPbDkMOlRHtmX1wnshFWVgaJ5JJr5ds/DYJr3VzwgbclN
lhsFOuDVn9BIMvf1CJrGZ1YsFVKCe5fv+Wr9ZMk2LV00DeED5Q9EjC671D2xO7eICEZRMMlXAPAC
Yz6xvlTVhmEB5jRDGh5xcdo8nLGYTAJiJkIOv6zlH7uFOLGTWkKnqBYBTYCz6w4q2IrmmxlNERYh
DibmsH3z2yK7hG1QPy+iMAFn2DlszD5IPZHSeNsavowSjGJuzKqs44vT+d5rph+i2LvpBPv6+4ok
L6tPPLaFvRkqpDPWmQJ0kb/zfaC8lkk2UStPskmsE/7uFwpMuXTQF0QyeYvlKkdL3flJKDi+3ZHk
B81aP9D6jnIxCk0CYvst7HlCfMeZ5IMs+sNPImCdBkwFt8dUPQiZ/740UzGLF/kpkNiE71Ru2sVe
g4QDUrumOWqeX69QZmuzRuQYQntpwH4DDHiIfVLuy+PgiwlDrR0wCwi5jnJuBVOb9EDizy75d7k9
+4MRyCZQQDb0fIZnTw3JIXJSqrASGRh3p7hxQdw1TS3gcuSADJQczPZelsBX5NR/5tHr+oDCB1Dx
LmxBdCaV3tmxW0Caha1WKbstGxPy+qhSvFYK5pKZRuk+hBP4fhLyswc21fF648zqc2gHu0EqjM26
dtBRhiX96N0sPrp5+lGLonKDaoH9MVWIgCfgI7EK36TZcS/IPccKLlNM+g8QRe5Hg6uGDI4wRRWg
048RHuZ+rhWvHKNMokMTbt46o2i24ajJ4Ob4mTHQDP7CX48PdAR7JuZyF+zPE7YV2+LZeTFi2W5O
x1XgQsKBhkrSLm33P8iODfU5FbWduVBAJrKfjmRFFS0owlQcHs24qLcuelAgp8Bz7Q8pAip4PQxg
rTxmotaZdW5W3c5HyEySQsUF3SOMzLdnRV2JZka0WKFWlri3oe/6Oc2Y6JeOfty4B1Msrdp+xjaY
CdKTNRtcyCbAbogap1tP+XyQ7d0NHNHDTyKBx//0e9lX9alsSeARMqls4E6KLvRg7WlBwAXqycWy
CBU3eki2DdJnr4QadQCdu9ie7GriRfUgHY3Xijt5bs0v7ggJAaSQe4HynAWbK5tdV/AdT+N2/vnu
23Q2Z4u4Wl4Lb2aHV+Wd+nAy3EDI9UQvS/JW6jxn0dUO0q5jpMs6LxZoi0kEy1BRusolqrs3RnRP
RbuiLfPAwPrec9tcvxTlqWXldgm+t6xA2wYaOaL62KWlAOSTZiAQ6uoPVwU79RUeZ4in7l8n+O2v
xK2OXl7TT5GWBOvutZJjjeFd1H8O3mdGY0H5eEYO2meGjHtxbmhtcKXORowIGCf0kucNg4SI/U1h
sFdV/xf6S4CVqavdoeWsSCSqRmzT/DFXGpm6Kld0353JxOrQGmM3DwuLV+DFcTpawSAjG6P5Ly/X
4IIh+fPYJdZuAGtHkNHSAq0MzuwLnuIQ986hmOG5aGundrpkxd1MIozxjI/klKwi6+Y2/0idTHUn
PkfNK98Ss3UHiChBSKbzKPU4ukiYXdvlsG4r4/s28Q0wO0VgeZVLIMb8b8rXd/PT7Cwmqd8rFjdm
Fts6h/oDJh0nfPOwOkayNX8s1ZZn3uf9+3jEGm5KB5IlZfRndnp6G0m3Tx63uW9O9HlLO64knm5a
eCn7IpeMxJQyB3Ttl0VDTZc9J3p8umeq9wgniUmmSbuyFzNPCtvAu2EfbBMg7fwrlAZ3kyIt/5VT
tbZDkYttRG0UuIwG3IQZ3nH66qgOrSqhvNlTXYtOcJAWY8NrF6yc0IDQOvlW7qiCK6hqtNT39t6Q
QcBbDlDFyChl46DDBXQ/r8mcHmEfHrcL4oTEIN1WK8IXMzv4etzeUzkVwNdU7jDCSVAWNZl8C0mU
+6faGgfG2Wlcgb9BIacn4ui5B+nHNpw/AFh9+bbenNzv94sOJmG1G6U8Iy6EOV44jvj/rbNipk2e
y8Zgzr0+zHrZgeG6QciCXkAZFIkbfLNj8Ionyxsw6CJ6E5KpaCBTJH7U5Q9Sj8l04maEBz7MaaPK
Qk/TXIkTJwhwwV8KCojn6Vq3kfbzoz+BQsST+ntCpj5nI5H0b0xwdFmxvbpsywG72aJoPSns+rzw
TNiV4R5TcS8/wE9ThyHJYtgu+k2J/pNNw6MyGWFJbxs3t1+GjthztHNynbomRwR6iQWZMgBrCohO
GBQmyscySK0gTXR0lHH+kbEKACXC2tAvbQjy43kZ9TKgolymPx0vJjJWyfwik2UKRFkyrmIn4E03
yw5UT/bCMk/JZ0JRjI6fxzdYvfS94NrLHEor2aQBoxamdealkhxG2L+cfX4Dyo1Jyf5OYIK/2e3p
V8gE2Cem2uSZ1aALktr7G6jqYm8/MOYWX2ryspNN+BHIGxVeHz+ryrzHzjCq4QUHZGwNW5QDa/6Q
1ie48uoqlJ4PvXc8FGCa3D1QeIYI9DpQtiYcBkgL1jlVafcBYbMuC791scnWLyxzybB7SBlLrf6Q
YgcOcTSKIkoYUOD/Z52L/BY+GQb2xSkOO9kXjp8ZTE23aWcSFtOBIDh0578dYpFXCBTP6f7VYSwC
P9707gCrcmkpf4vLeaDotdbX7WIkCeugVL7chXY9ZMkYDISDOxgU8k0ZkiM1lSFYz4pbhJOFvOti
thXaPayPmP/Nyy+xrfXTzIg3FENVX/W5aEgN25y1zEEUElVnOEaO2kyQ0WQguzcaZ2He8Te2teU1
+6T+DVs1aPfelUwrdwe01mXMSK4SS+V6NJRM209/WfzhF5u0aUScI2HmfkxjG4q6icysmDjlOD8m
V7LmcBz/glm1x2fd9hX65hXft8rerVK6hryutsc32r6QB/2k+QK84GIcv6PvDT4LdwJ73X9qvrfl
kv+b1vo7VfQYCpOG5ZtLxRkuNzAaEnk9aE4RbpPZp5uw0CKqG9Pzi5GoWKBI6Ao1MNLg4nOjJ9DC
++Z7WTO8T34oCQLmG/Gw0Quk48bK1sA2C1V26vAMjHby7CmEks2viRkygw8xZcZeNHiQRAPxQWe3
pceg7kjNg685sPO6vOeRieGKa3dHN9iyxcrTMEjgTWkOqizPOGFtA4AAGYxErM7SAErgI+bgt5xH
od9ibCUz3c38i+ZwlrdYc+cCZHPq9i0YbVQ8HSJ4BbrR3AA8HUeT7s1FSjtsh/dFcad7iJ9Fx7lF
O8g1tpSRyOBB+lpqpjnXxGKcr1kjHFMmsR0mOka0WtnVGIYIITVHkZzfRovJtSmP5Z6BxEvOXNC5
SSwZffzxXg8v2f+AKA7JyXT3U0LYdo3eM9gX5EqBLRNYtFDvqNEudBQCN/aHjmE4exebtf/iIwr/
/BcMNBQpka31R5NsM/3UvWXbRpZC/kMmBVBCBE8hvFxQmIxlpKqOs+zxpgPe/7qgR5qAky3wnGdq
rYcc9UOPBHigsMJdkjDVb5W9TfIKcM4dYHozeKKFE7rKsjBZwfKcjkP0NdZ3nTNP7tOr8JoAmvj1
5aBC48pptbdTW1o6ntqeSPlm9EgQ3G0NgofOoYAIlWzpi4y+69fxRiQ6R6WSxOtDVTICxy2gTQf/
ectV6i+F96w3egLlvetCLj08NknAWTzSyASxRR+ZucuxzQjDKgP9ektbFlgg2su/uW99fnEnXc+/
4VKsmeOrgFINs2QyJVvsI7zhiOJjthF9H5lQ3PNTteudx+pGAdNToLf0zfxM6GYCONPWa38iAcl+
huqxpXMCvOobiaHhsE2xzH6ZQHjm2aC9gcFFYeQ78SAnno+JUwBlSjvJKwmSf8ILczv+oOmnbGRM
gXVD/dxSBn0HmggEFzEj7GjkoRoro8+7HfRzvRp8HEEGOzPUWuKg/dU8X6GkOnKcyEP6/2bC3qlD
D+q69Zy3c/N+dCn0RHQwx3WM3EgVPxWuDyCmS1n84gE+xN56Xs6fLJxJJxwslYbLa+ImYDvYTG7D
/BwMdiTmfusqBIkS4Jcy/OA+vh3eO7QhvsErWUrTGqyoclYErZ/UI1Hybiv/8Xv7T41PCkbcpSVM
JaXr7U3HGBT+iNUdA99fqLo584dkG1BIYld/u/uC29zziZ/qeOEHjWGNRvKzyX83Tfr0OTPNj8kd
gkBCxGsmDnkjwPuq3cmFE9UNCuc2l44PJB/L6UkTZKiN9l8o7sED+7Uf0hTw2iG1A5FTRYhIhL13
wPkDGpkL9cIZkHLfbBMgfoh4Ahe3W0Vl3C/EnVy9+ruNSLTIk1OqqjCEZIClnhJdE185yaN/4qf4
tzlfs5zTf26yxCeX3orGbS38bdkdA9FvrCYOlkCPdWuP5yD6z/t+zm9EKHaB3fvNOz1Arrih1f5H
oqUSjtx1Tm9LPTuFKcLKiEhZpu297MOW/IbEuy4Vq54w9AEDdhAzIYL62Ai51f1RNBQ41TRX8YI9
anrhwQ5XEFpN+92mSQ0WwVTVjhQmwuQ//nvQCviNkNqyXYS+u7/3y9qgiddKq0USJe8DeCVbStYq
G5k4zHydqQ4mf+KS3yRgR+Y4wPuVV9zUTPEXjku83b3VDR8qiL4t3JNyws5WXw6j0BOGz7+ZXvwG
VOnrfj8skSAADUbEdNtPDE5uwDPbQrDjA8jFRbChxNGHPIlgxaG0ZzBRzePQrJEg3jZTCoizFKxH
SAiyXgq2AhgLI1dN1MD2U9tHsdYqtYA/KiV2KTZlE467V0/CKjOo7B3VHvW/NfSfOO6qS6HuOsJ6
Sf/6G9+wk4oWmd5GYYMEoQ7zk66seUlPxC0g5GVKchO4yxFGmY9KEbLf6knbdIQV0psn7VdJ6kbZ
kn+uVkE6NjTccwINtRfL0TZ47c9afSb+S+DT6+ww5W63SCi/abtYz84f7G5WScaxsW1yxeqdoZ3q
urtMUdBJRZuIhWrf8LDwqmLf+M01s6yhJp2Vfpg8mGFEca7wvskhvrFIx5yt6htFaWy3qZyscRJK
sasf0WdaoTpmlUZnGd73wItYXHAOjWmgaJMuTIsT3lTm2/IWYxZi1E7M3jwgauA9fAZB8DQHb2F5
EpRZiTjzn1nW3jMJ6Lvf4axxsxJpHwUWihUQCVoqim+iMDxcJPrhHde/82D5ob8xt+LV95E34ykV
NvmJmMUOt0GZRxfq29D65u4R6+CPqk11KZ0bU3OupA5b7BD1LaqHZM0STMlfXUWwD2XXrz2+SfJN
uw8sbYVVcOgSdIU27F/RAUi19BtEQpXBPOAYTkkGdGKfkobJZKM6uESZw7pwe8EkprJONwanWhIP
XWxTAsa8b5dsT59xzvSU2p9a+lrFSuYc4wNcrBR91NXLS9qIhvZh9e+kT6bPHwj2QPdb453gCX+9
Vt8QOdg+cCTYU69M8TZJYXObdTqQkAD6yqcGQauysSwG8caYO9qYwlvKbFfibR6iwwaSrdK2hvkM
h7Vv43NxROhiZ4irchNE+BtH8jLU5T2DIbqoOyIS2xRYzQKJSWHocSFrpmHVMBYNZW/hGKTcrE2I
p9WSJgU8hgBcEgKftZbDPOyrgxNpo92ws0VrBm/WOl92hRNKhA1rDYGT8DkjIWU1jyCpteZSedzf
iE9NO5Hm7ThECr6N78fm6cgE4tSEPm4+7FaIlD7/aTf+YII0Viy6rcm/QbBfepdAyMgtFC+KlHhe
8/b3cAxUhY8a8CaA/N3bV5xcp5B+GuQne8FmTjgPCaPnCDbkP9TbnesUd+ZWgFuecsgZNo1ttlOP
ZEyPjcKgtdg4aI0yNuKGntillGRhRt/cigTPVB8RKoMggO+1urSslCyKhT6u6ACWmoLuSh4+a7OV
WawdU+9J0hT2Z+h/s2zScuBBwEXsrPZtOLf1BqcFsLcS/YihAINWLhq+rd90f9GSamkBjvLAUXOl
74kzKLV7kTlDM2CJ34wikmJ2zhUFl8YYxn+fgyyXe8R1VVfJH4vUAX9cYccZ1NVYJUsd92iSApG4
vNeR5mqxH9f+NoyYW+KP2phai90iqHr9oNGR6IE1fXtkEl0yffsToA3V54rGo7lZR2igIW4eLztd
uGqq4pgQ2/gIJ4R5ZyRi76p/1YXSzs4RRsqP1ErGPjvXxUzCuodCjUpzWxCTk+BYasiEBSSIImb8
ZF1c5ftT2h9OeVCMaEc5f2TmgEngk159Zx8PVwoRzU2bFnpGs4g4fz+9xTCONrzIjtwxgWo7j4Gl
5a4kPH79S+aL4PBF+DwYwMqU7Bv0zRaDv3hWLGcC3UiApRLd1DeM61DBgnuyibvznC4nxaHr6bvO
rQ/2SUBvoG2wawJzxy0FxoPaHPd0itr9pbwzMfX9v7yNqRJ8d7lPOmQV00w2ab6nrdFvmyq3QKz+
DYp9OkBsWWmzLJyeNApJwjp7s/5Je7ezy0RF+Yg5MZj4hSHIyrclhY/sry3tIQvojyq3WLwDLaoP
LnY7IFgGMhH8b2GZzaXkI2cUx8GB7doBxqGAp6ECDX8FCojSL7RrwErlAfJNqf0uVLrCOgYoKVKk
AEEMSRgtBWr9neIi+G4uCvgd1EMqTzSS0JRvBb7ZE3k9EYOoj5H4wyJH0FZAn3t1Ql7VOywZp0WX
Jg9l+giIVicWBK+BnrqKaQAtY3eon8TGaYm56xxIwvR5QH3lFet0ZECXj29Mc9Ze7uLini6IaV2y
8xK0RUUttdKrXR0scgCakcmlaab1Zk2XcBFZ9FIIFbcHrZQRD1Nsgqajut9+V/6a3DYpOux4i7zk
8YlSE0++pUJv+80hGaRjoz0y2YYC535G2HadfZkVA4iVuvOnZf5ND5sm8mvk0Pb6iaZqog/ULPW4
V5WIl3nSXhS0lTg6sJF6sHpC6Skp4kbLiYxn2BslpSY+cq8uEjTPDSwQm2kV9dbvgghrL6lg6b+n
aLchLpnYqjC6jhapL+2dD+fbfcBvNwDMjbQGGzDjpKez2ag/3zjrd6+bsT3J7nmdU8p7Vhz2P4jj
zlAi02JIZzRSpF98B7JkmMB3M0CaC+RrAe4QXj2zv68ZolgYnwfJTAKzPYZ4anNpWSYbpnTqtZ//
LT6MMZ1BDzBynqrQk6S7fjSRoBeX4XLkFpD2jbjRiXIfJeEJsiHxkE3laXWIpd5MyPse6jEfIHFT
aMGduvwIWG4bZZ7Sg3EWHtPcxWtbUXWcgSxZGGVQoE8e5knCGnTP83a5hEoL49HIcgwFDsnmmm+o
/2OAdsEa2GDJUnX5P564c/hwt947ryA3GBfdlZoDr8b/s3OngFuM1Dsyb4OUCOBM2/MnkIRGLyIK
+PYYZRPFYGo8o8vVWqErZ7FeBVwoPYOHKxwsBzSohTzoiSfRXX/vHF5cpUyFxjg1+zt98q9yWTfn
fzj9cBHCVlSAzejpc0uzX6zHMr5DOIP8k3o/VGPEqg6aED02MAbttMrl4ZKNbqmrcrQz9XJrFfj+
zad7uC9rYoG3HA7sXE3rGNV8fEoyneN6VKanS3W6rbB/BfFnFQcVEMoVzgWtnWUmNbJvUBn105AP
G0dMgX+qTOxTgelysPba15bQZmCE72v/zpM0TWm0OYh9SrnSaXVE7YHFOSS9Jjf9rT7ocMjs/UIJ
DuLBm+EfQwN+Ql8lCC+LQEQGP200jAm8xe7E/bViGxsjlwU2TKEJxnmDeORzcfDicauir2yEbNHB
wQ/3aVZ9Kr59lvqhoECGSB0I9CMi/wuzKJjePfheMnkye8tafwHAv8oV1rHiV2iqPS6WgUaNADnQ
p7Sj8dGC5V+o5KJDS6IYp2AMhz5EDMllOD5sI/YlRAMeKRAtc1KEol13y73t8uW1RngqEh+uUsds
2Gh1Y+1R4QE1o0QV+L18LgZ2C+/GjBsoUSyojXI4T8YAg1RMkrPhm5VOchSnwapvy+CEA/MGjdU0
76ss+GxZYZBJNJ9VI4lqR7ZLCrkoGGAzNS66Kxkg6BQeO4Zn6H3XLyiy8lAsJrvWJZOZCcMaOslU
k3/RqSvc51X0YRvXIXVT8TlaeSuIkJLgwXsR5z6ekisoc2HuP5hT2bh8D8imbXDQGYSs0FlNL6g1
R+WAlMVUy/qoWljm1N0xxJOLVcoF0r4rvhveZD+eUXpW9HZLF6wJvLhDmickvLu8CetTWYwxsmuS
+/8IADNAzLyw9cnLEJ/6IgjSXarsS8QNOv6pREkFEFNOlhxE7ceN4G33O/gst9Q6lJZ6Vij8Dr2D
9u7mEfBImG+4kVOmWftb6dPviMzykI0xb5ZmYerHKHJeTMZ/v9LswH/a7/qgADeTn9qQYg3yXIXx
fPcWq01XY1m1D0EfeeBRBXb3XEIZwOYYdxpIkZkSUMkt6SfTuey17GbtbEzh2MpFcmjGKYQAY4vc
gfFKDruX+SSNiC8Oko+qhF1h9hJ2WyuFHbpwUXmZngbfjYx3BofE3/M8ot9DMSU5nmtzSNVM4qK8
+A81lJxk0JKa46XV0IZVo9LeNYpEjukXlN2yBf0tGTPP+xKqrch+bUsFgFFu4jRmQrhZ/HvXwp95
IOoqWGxiGrSv4vnYJDBhmxKHQXA8QLRmLqKtFnOoRZJiBy7rzwJibUpYKvJxrch00zjc0/u/qnnq
Zg4hKqQ6TjpMVOfQtd0rcZxeow9uxvASEBJZmcknnCD/Gy+R+fTEjUVYIIMyAyRa0nhhy35OlZJL
0YwojgFxFGqiTupq+xEZuc89TZtRQ2QhNT7Uo07Ot9o75yb1L/oFN32wRHFT+OzuzEiqeeZdo1m5
bEd+OjYaMIdpPmaQYghkoFE2r811JxMZgWKPzCzIyduO1SpzjRGsFc2PZqnn1WxsyXothYEXLTTm
eixUyNo29o3qXUt5/Oh9N7KmXcJR5S96oSaV4M9kV//vEDR7ZUymDwJvXWWY/DgVhYgwY+PgPrlB
z4ZVEqUjsuWJYEc+fSE9T3sBwXvZVsaNWxJgEg6lzhSd7k858EV9t5xK3H1lKs4OM9MCh32+t/7Q
tJYESI9CtR7N5rLFmMiR5SKH26OhwzJ/TUsn02SZS2tb5N8ZCzxSW6jKKhQzrCXNlNh5E4ZyfMnh
MAqoso07QnKmapTAMPmwaDQGdb/EImaefrJn5Lb9QmTv54D8/XQmhlodZTc6K3AkmXZnccnCCT0p
isgGDlIXW4LCmkYMKMqz/Dq1f2YC+Xnj5RWmTWHbLch9D8CKuxzRHt+cY515BuuyKVOY5sQlk7jf
OX/3YAgEvwQp6ttamPYoFnmmAhJjH9gF5+H1AeTNJlRpksPZsV0ZeE4gAyqLiEApLfeb8AqQ6gy8
zj6MsiS5LKiIAC4RNtrxuRwKDFrnX2tSZtdM+qvdPPyKFscjsMhUXxMzTjDh7eD2l6Oe6dQxY3lq
1atWFW07/EOchChDsO5Hh1ALhyOe3u5zPeBhFmuh31ht2CJXuVwNoNoiUeUfEYOUmlkAjgbKIF9I
ClSaUvYd88V9fXMEC+9d9nG8y26eodsUgJZKuOabxoXnic5G3DYxKcL9gCTiU2JRWr3J4hhXakEb
2+N0ql+HJvfp9btEl4ziAcUE0fmNL5N476t462bTRMBVwi5pkg9SDxp/CCmpUpi0gvb1vQNsr1si
8Y57iB/MTU12u99vI7LOo3HyCEN7oIWYeXTLl934IKDwRWvDHy1e2cRGD1ZjzhSY83/z+pMOjn+1
NCESwzSErWo6zi6VRAhi/QTGjex3WmdJhyIPeOSiTfom8xqpEW4Rz2pUfZf1lqTVrd3Ad7Fc6Oy1
+4izuHRrtX1e38XJJ1cbDxmpIeLcsW9kdqTOoSGHC/OGNSaHbhYImSFRU8pi3i/oPkr8wBTOiuOA
7FpVqgDbcmVVUTEc/3DkTAY8xAPzMQKN+JNQZ9jJBjExzp0pgulxDGW53wjDk1tPNEk88g0lvAyh
cd8KLIVq1EVFVBY0R0PsAG9HGYNTgvsiGDw/ezF/84zWnumlq9wbJ9QlNBk6Guq6/5ugg8oDyOlp
97X/tbu1ZsZSu4K9LQekX81qqOD9n0YQJLJmfsFL86e7ScfP2TJCM7EDSFZYapFvWrUvGjtGXMwF
WqiKTPcr5oYcqgbKRSNNiJhNsfXQceSTKCLTAAI27+WaLiAWWgN4urGil90w9EdtuICtVllHf6oH
QuM1u2Fgd4sa0gYOh+d9KU3HBZi+eBOSm750GLAxpDLVnPkYqDZT0Y6vHqrF825FoIj+zAx4oY9Z
WWdcCEB/bvfU1wF1n/fnQlwya2GLmzhU/idkXPatHXtlFKOM+Y7xnukIlheZmDtX5YVNHAYUT4wp
Oy3KvJaE2iMyVmxAthVoDyd4qLxUp0r7hS0HiacRwgcPzZ5rl1l3lZ9QQAMM4sGHPV0ScUT97TyW
jsvG8CRcg29hQkqclnJsm0YeOwfe8ebpVWV967WG2PqcIJb9dLbk47FgX2YRqr5/QPKV7Pw2J0Uo
glRuRab+8BsUOFK86aamPi/nmyq0tsLQShopXa9yWwv5/AkD7700y4OJNo6bZ8YzHRx28pBuKZf/
Ejl1oZ6ueQGmNg+Wt8Bg8hugx38v/BLhbNwXNljDHTAfbxHEFk0qum8UydD3ns7wSwMN1AVxf+Yi
oPskf+3hB14dhKoLUyzTNMK1++koCreEUugjeiai/oCFsIitzazPozUYgEYNap6CfickNTJznumh
/b+TuQQ8TGIbyCtvoYfFDfYjWB0ehXK27Bmq7x4XnF2kYiJ4+0rlZTLtNxCnwFU0JrgIg70eW83J
ScU+fCesPXIWOLhWNlIR+zRleCKlbMODkUViWDGy3ucx9UqyXhZ8i45ToE2WpfNg1+qCH+XmVvBC
LejyFkNjIJAs43jXAC1uZDrgzD1jtCFGK4H6BHc8yR/JSIBFwDf+VqXR7YQfZHNHFaltqaUK2asj
LeRKAKihT7TgJsXuXBK4d8dM3OkvTHrO2pHisXRVMshZC+Np9FkQFOV0bKipRO9cbAWLHSutgc91
0O7az/l5ObADJlfVFaUkaeAzU+Vl90AXERARnxUkQbMA5X2kkqJjCN+VoImEcTjfFeWGt5lYXtAA
pt/dXP20937y3HVgr6iXYgm2OZGUfR85Rk5QcJG3pgTQ2tDICJrVfT+lLFc/S3W416gLlyG2j5dJ
WhKHlj4i1Zw4PY/Hl6ig+ch7nIWXtwq3V9nG1OAX2hB93HaZ+P8Viyjg6PSNq6TBy+9Z0GlBc7pW
jY3rHjImkZKDDV1g/v8Z3OQEBAd2oSj+oQOgZeiaRUPB0Zovck5vUVTU2kO64ZbLbcj9UrPM+dYD
y6CyCcfbMYm5P0MRzzUXxpjoyW5GFJZxBXUu6/DwYFjuV3ZVLqlPVh6h/hMK0calF2wGSCy7uQzQ
Aj5DP5SekuFqj0+otVk1paREYqVw+2tuI+Hq+mxTnWpIvtDeN6g9I/iF5snEbTTsbkU3wCV+37XI
J091HeaVkE8xvzKwAn+u937iIkbiqGCbapaYc92jFGgQGRvxgo01AZq2sKm1ALJGYsz+bGGU+PBg
Pkk3pyHH8WPjUOraSf3omx3SKGduXqCV6MYH3W1EsbBqrgG9fYubss+SipQGVBOLsDzk+wgrtycE
0zFZ0jCHeuVvIWofoemETiNdvzDF61w2cf+cD4+usZIuzBrWbpo5F0Zdo1uZxkDSrhZRdg/hkM0V
EgzFXlFoKJPFtjAfbAZGdMoB8NTjMpM0v/hCvFShduQS5GzvI0HisJdVVs2b62gdIFxi3EYGpvAQ
Cw4pkOGwGuPYyuQ5FsS8hxJv3Qv+zZFLqRvGzturkoAFjoF7+Ht734EH9d8FV2bzwSv/xf+q3BYh
CDdgF9B8HrZsRMyjJd8nwt0CV4GAT2cmToUWxsuNb6TqBHUg48L/qXFaqiqS0JPL2TOUyARqynt6
O0Q6QzNRs2sSTIXgy86Mj8NFkIFMJQpQFEryhRQb2GepNDwjATXVOrgdUWConMoa1SNM1VBMqjBO
MgxbUKyURNzHgb20ChJ9H0cuxJLZGyfyrdQgn43m+uGONJ/kpOKiLzsPkDWIhP3MrZL1cStNC5TD
UgxDIckuna1XF6Ps//Nonc3ZHuvP9uLRcGWDJe2FsmWaSz2yXEZnlC0Qn5CA+uUmveE+fo4KO70P
GVKzicT12nLerB0PtvUaEJymHEyazG3WowFwhIivqkJJOI2pNtTnFCn5VmeuloYgL7UZwCRpS8E8
AVw5QQHSAXiPL1RMc0/oGN49h/n7wZQBsGQk89Vy3riegpg9SFLNw/MYVbUYUea4CK9g97kOrWtb
AZPMOvZ9HIUy94sAvqBLpNpTxUK1o33lnfCPlGHLMoAwbjI1xKtrs+D5Bld5DOxR2KJxwippPCUI
DMEzJMrjkQWPVqLZHMkSQ6LDyqWBKFD8K0ap5TYrW75CwuWyYac41BtRaWVNsZ0gZDld7DW/pH0Z
kWZPIMPXWUVirdHVmA7crfRY1E1SOFhuNErbTxUjzglm6hT9Pm2cqQgHhv1J0uFOX/XPs2bxP7BU
3IOOhhHcgJuif+HFa1UsIwXjNlWk91h7zwJ1X3qTGCw5HeUXWX3nLB8GVI3pUgbaUDCj1K5OzT4P
3wTCTOZGyEoVKlf5mBiLRQdIJA6o+6XO+VDKprqnnf895+S1Edb5umM8hCuKO0Z5VBK8a2ftRV60
Ab4dYK/TIf75Eo6bQmDgOiGtwvVmh2EhH+4sebv5WRfXibTwW8zAmxWr9qVIM4m2N7HKHwish7Hc
iewcrBJBkfLioQTOvMtjntJxCXLnzaDBKoSmX3h+RAkX5jIzhn0h+6g8pOsq4Yv44v2EuzWVb3PJ
Leuu1VOxqpkS2ePqqfMH54Yxrhd2OeMLqvlBQmRzkvQ9WFpadI8omnkd9oIclKMhKsvRiLZ6sNMb
6AKSS8jfNXvS6uOTMFYBxwoxueYGOrc+ueFnR26bjZRc5xMXV7sGBdli7etecrXB3QsKSyWBG0oR
xRa43H7ydG5JLJYt3J4Ago+caAjXzUeDUvfA3zBWfMCQ3pYgCnF0Tpm+Te+8ksd82sYIWSJliKXx
kTx3ss2yc7XWi6ct7w+5QGj6yCTOjR3qPfErRi2Dj5uIzSmSRnR6BzCsFW92nGy+JMKufgtThtGX
L2n3GLh6WyihtDKt6QxUh/68FiBcofwgi1KdgkMs6ULZ6d4HKmkHUEHK1RzUxAxoH4acoGwzjFj9
fM+fJczoC1hl9VJoVYLjzmei+hg2xKFqzC5+7NrVFC66ukRhdVeORmD9iR745G/7JUhXMcDmsooz
R5YKQHucbS8lSgJLJWakSMh/2k3nLPRzAYLIlGLgMu8KVPwatzceZqQaHt00gWYS3qBB+r/64QwH
niwGStyFtFeEEhLB5YbG9RY8wdFnixS5cVoRiakay4Q8LJPnF0Xik5MaBgd5C5bnJut2c8FnySHw
NaZbDzMUyslsrqY/BkpMW5cFRMyc8fPcHNkjkuayHBH9gVPLcW7socR0TcbpL1vPt+q1W7x5JS1v
i/Gd4tOq+CHYBZ9B4Oxyae4wmkqyab6fsfSbRmb7kj49ElgpNHWyMMis0I5ouys1LdNbdg5+tVhS
A6PPLJZXeWGreEHG+SIentF+mbBGRQ8v8nXfuSzmn6AJPBYuL7ZJubzHy5N/JAt9TwVetpN0G84o
cqhQG0j4CDICA29RrfybF2FUEVjhSBhaQdUusLnv0z2WE7tt/pY57FG/oR0Q3ufaYFMKbFrOzbXg
YR6SAAlVgCwa97eL7tAnY4HdDld7+wVMAhisrhDWWpsRMD8wC1J0vEDGnoOSwpqBWJr90eBkO4yl
9kvbkw+CMKAjNjpR9mgm6KcmfAncKO5wSmuhZiM14J8kbqcbkM7UjhMCmzCTqaGPL3sQCKActtOi
w1RWiu5s7JNl8Zt+HLt3h9Z/i4gGcy6U+iG6DZwRR0lwor0gyjRspRFPoO+ie/aMQjmBA7jNFE11
KqRLJJv7n463iYfbWseQzzHPWCdhk+Ez6CbF1Q1miVFaQZlxGd3feLr8Lu4Wkjs8+p08VDtPTyCq
xd1tezbO6/CAgXfZAztjIv9kKMFQ7Cbt4YCfWl9jZkYqISnLuP0WhsCMZxUFqjMuCD56+/FbPfwM
kfYYKImxg4NBWK5SZ8TsQTI5wWUbPZ6oyGw+pEgE0jt92JhUlwPnZZSGzwJo8CvkusaJYyi/6Kyi
ksqYRYTWWBO7hYvpVieFvo0ecglEdc06CKfRqtFygkO4WL/KALKX4mPqExwIwFYA1pAyfb/qYBSb
CHXzri5MWlq6Lr7Db2RbfZ9/vSESIb9cvFfBS8/izC+E+g9ffANA+rx8h+jHSVyQwxG0PdUm5F1s
SBrsp9sNhW0Od75YCDelYOsyULNBgJktERxDIoYp1WdBlejwoeYtBaTRMB2oOhO0ysCu5fHHS5Y0
50MkYvWq2e11nCPS39aO0MkNoa2yVDBulVrGtQm2tBk8DVRdODdTwZAXpH2ChQ0nJuCNdrlBS1zj
a7SekUcq5duvBOS8vRkGR+o9o+8ry9cfESvoNLoZeqABBttb/qFQSBg9fJrGiB+VkQmzZ1Nbk4U3
4yivxXO/LZtUXffYE6vIT/GP/w5X2xiHLnut5teR2YwgtEbp0EAxb8OXlFGvLAKEkdDoajFqy0Jx
zWATp6KVa/Xe6I9ImCXQKryp3glDh3ZoEWq0cbWUmuDpq9BZ/bwguaNCPOK5tB4HPnjOLX73rkiH
UWYv9kxXI7vY2dsZPI/98fOjui+o5zvHhKlmUAy6Pztl6BOW1W2vpGvi6cBr8AeVsYJUZc52n421
P5WCyEj287aTLNc/zR7wlqSSKM2cV6QML9YBMZvwsFFDGefR2sChbq9hntejDGehJxIf0p9QwahJ
+aCyKsDDSKla7Z6WsVXT1Mz5ltftSH5zAQbwcQPGwZEk28vAHWibZF2t0auJGvpYnyfwqaqZiEdN
yn03qMn7g3McNNKpzkFSBGQaIvb1eznNqXEUih6GNmr49RXCM77EX2sI6iZ1GqUUg/TY+/sZbI3r
OHe5cgE99VPz2FDoSfYB9BB6IKHkNGrBz/btRxO6T/5nwstMN1bJJu0jhAYpM3uMfPq8K1k/hoDl
5d1gOI2QYC8WPY7E2C/d15jwUilowpOmN0wRQSnXWHLrpta3CArczhPx2kxQINUjcH7JzGxIoWbP
GxvjhMAewqWL0wajk2GviOVoI1clbR/7GzCp9Q1B8rvZPGOmPvyD+ZmP19vOBSn6XEsG8WseC+Ep
uaq/h5cNbTkvJOFDM3C85Igj/B2Fda8OW+BfHgGu4FRgtYjo+azY7YciVXt3Qy0jguKLu5IHnyXy
DMGTiXfgbKIVx45MINqf8rjYR+GaUIXRkRX5+7uIFgVB1Z0JEsbDuoxPBDD8N8hP9+dp/ByVRQno
89wdYqBHkq2pCQ68phCZxWrr74GzuA4vzX53ii12ld+e+XsNBcNXYAQqLQZMozoFeLJcK4uq4tmt
+PiXf1GZsQdS9TfYh+WuG0HEBILFtp3jwS2SCg7yX4vlyVYeQeyY63nVs6J6xWhsUff3bSMY1QT4
DMpGg+SFx4CIHK1gX9J4KXhnfmlXT7fVwzHISC0Y9e8Olrkq3srasH5QECmSAhNDgIH8mQHPvlzK
XJlENiW1sS3WTLQVFnCQ7Wuo60hyixkwgFvVeb6uoh8BVKFxclMD5R9Fr0oHRbvV6Uwc7Wa6AUOn
e6RaqlRK66BTJJl7XtGBEROKq5j+tXvoESV+sgxtTmbYPNlG6vtHcF4y0tsfhAl05eMb5BxIlfLe
tjm3xk9TNOSprv6uVcUZgZNmlLHbzHSzMLo718XvpfG+9BwgkLPKm6bLUMwwFIUH9ie+uEEDyz6/
0yyc+Kp/k7SxuQQzs6elWVWPmzX7Dcb8hEn8KNkw2l3KWYtMJgvVf2Uj9SmQApkIq5xzudnHabVS
hVmsk8OloZ5usMqROyOycfuxTB5dXTijnxQCPmHMx23b2dIeKKz/pulbRgguBNCEYu1BrFWevPyp
5nda9RTQsCjokQ/2+S2W75jQ6ngJiSAftk552+EEOPtHsxWyrfO8qkDkW7q9IRSDw6/TRlZhlREG
ZamQxopk1wjB85mXVTNoV8JkuAgOaa8t7Mr58TuF0zKiHA0n6IdvaNCchTxwOpo9zTC0jjoiBLwD
04/IC+2Vt3SASvgz1GK05YqhcXuKRSiMdYGJ4Q2gzd7RVKCp9OBPkKY7a07N03W9Rbjnb+PiNHqo
wqpeNKXnDIiUyRdU+7MtjFhYsrrebXPExR5Z5ISSDdLln+FuLA8IQAOClPIk4ZQ5+v2JeZzNEgQp
X8qlxUTwawQm664JrneLjtl0YuDCWDU+dSh+x42fN1Xeoaa0qnw9AOmQmQceCT5WwZugAcu4j0xV
sxQ1qfob75U2KkHFQrFxUmoqLeUKqgHCLzghoMwNpEE9HcM+VbKa5ATBMSkjVFl36GWVw9p/Ualg
iB7B97DIYK5kxUe4pTbwl8pyVY4BGwFf9/vNXEzHU2FfiH/OQiR0YIGXZD1u3Ff1/ASCwjXmSMno
y5//B6B+64SkkE/0/mVQXevx4M6nBDYWN4SDtSDUsJfA9FNIDSrDQU5SnMD0aX2WE+M1vaWSOZxn
qOyW/Bh31H7ClbgKpmotbkIc3A4ElATbO4WSnkeYiLXheMMHlpW6hFdd9+6nPjVYfo2N2G90i8Ca
1PsRxPI8Dpvh2suLT7TSYVJ83MFYvgJ/+BMBZW45XDBv32PfQ79eqSaJrLUu0elltJYi8NsTCJv+
SPMBBpz7V+5v3Ejd2+6/XKY+coSbm4viugTVMVS8jlSVXkSsohYdndmdknkZCCwBr/epAvyRe8M5
J0FukuUWzFA1M4iX/ZtOdmcdrBNlqp+ux4Gofg6tFGpYYHB75OhEtTPiMHvPVsSaJpDbf6qcV49R
SU1aodXhvN/QJCDIfPBcT4JvLa5xknP80GpOEx7I/9NhUu8128Qw5YOPe4sk8ftVkM4bnsQwZbyL
CKSJlaRtkL2dd7Nd3nqZdRtkpxvQcu0v+9e8crC3dwLx2bylKLMcKl0HTyLAfD2eYbrE623sqV25
rwU35bmM0yskek4xR2szmDEv5q6CD15FRWQzp3aMG1vOa9yFyZRJdswXqC0211Xq9PuA8VZPW73Y
M7cePWukh1U7r5mnBsqdb0ioqDaIxhKzR23RtTft07qgEDECw5Kr9UYP7v8tjgh/vC1ohqgFB8+x
Bpnxl9hswSSTZua5TGuX2HcvwBRaINrKHyC6RCEwcjqm/96E9tPQPDYznFs/iw77eL30VxuO7Sak
KTjXU+lXc36ExkZ73KpywvBdFMr7szpVU25SvEz7ORlFgC04n/8fUf4IHveRwAAZYqf17rOAZOSC
OKgKzRIAu6BErYfpxllBvDkmCGPKp7Hj0dzkZ6GzJp18u0uAvb6bxRZLo6Jgm0vbQYhqwS/kU3vC
prXRtRCPES41Q9pgBtvJZET8XoZWejs5duF164z+i1C2JtDiP/90OeFNyuJXzlATMZxjRGrasnwx
nqLsqe9rQL3ztXwHQHhGqcdKccN3LRtEmDDBw9XmZAI3wBq6Bvnxf1Kym+Pxhg349j1GdVLS5S11
bt68xs4bEIcZHOht77Wtyu2Xaw5IDvthqn7dojOtcU+FsyvaqcZzbx4JaTOZWNmIOaqCwYdpaGqH
qOvsctq1Tqz5pcyrx4CId6Ld08RhVcc7xBYT6c5OX8r2JvmIJqkhqMEsugqAxOjDGZLoRIZIx7Jl
Rt9bXT82TCWvF6P4mPAfEII47eJiEyqhdW6b8mzXVBeKauEOLC7nSaNm56r2gQphnspmuPX1mYjl
nGPl5U6M6ZQJFKtViebCc8owxQIzWY0by9/ddJTxz1loCJMINJ3+ILMq2dP4MO7uaTBUjLv0+Gsm
JhDeX9n0grAWgrLWLznCHuTxGZA1rFqETv7uMxus3UmAo1VLQcXhpYMQsuD4VIzNad9rk4W1RiCC
272mEViTqI2ryIj3krizxalfvGOpnAOKTtUfQmyWWrUsgtKPDOAN1eok4FE+hMHsdX7suseAVpcU
L6Tt6S72k5YZwnvh7BbebZFQCvwqkVLdgc3m1e3NWnV/qVlq8ouTpfAoEZd9M5cm0hYmVZRY/2mJ
dtsXJbRqFENowSn4ZnLi9PkQw6w2c0bivIaPMYfIaVWJ/x6ruDDdmpCIQyZ5iLqfNP9T4ijAKyCN
+KI3RFWKp4NMbJjlYz7K3meDhIVFR9ChXaubdLB0Ka1kKRsGup5amClJQQ+p0KAFCT4sMVywe3AY
PW58+jWbr6iuE5yIjp575Vl+qnSNzWHBvHmIqa+X5//TCGBflQ4iLJKehQpjWS0zNJ3UnV+wPmGq
ZD7DnG7GiGuWzZG+9aSlBw4ucQcp2j1UcPrKL0UgKyHvtTLqnTmyk3WLBto3h3zlKbtNML++9C9o
/vOJIoSps5SApNGYdXPXBki5n/5N2fTgDgtuSgKZjnkXnHK9J54xRqCbaAmftX+9hYRe1J+fL0I9
cXDEi7CQC0r60GUIWHlS2qOUysyVsxD/rK4rvd4pALofq/hRtch9NBAEiByIGztCbNKaUr66VXii
BT2M44qQzhb1SXdSaO/52c/o7yNtTmdCB/2hGWloeRPIU9ggrbWGW7uTGpXfuPkUjHQGW76ez0SJ
xOwwI8/H7rrpDHKIBad/nncVAJmCBIYD62QEuu3NVoeEab2NU0xNdZcwX4tYnuIaERgPSIg8pBlp
ufJncF/lEkNq7DRtvxDu9SSK4sG31Qxg3V3hahTvMwqPGU1LvDSZPYORsFu1gbAq1M71vbDWE0tD
NcYL8WtmVEFk0OjXJ7ve4pD/RiAy/BO52J3Llip7pDN7GjlUAb5R+7l48qY/VPz1DIOMb2H68I+H
eiB8VZDyCczYqpn11AJRdw1q0GgJVSoHKK31bsq0iK7o1uhZBhfqRBUr/Rri8sVP7xGncE5WXMI1
02vswabWpYge6GnfkiFwd0Rb5XGmaDlgbUsUAqCUYEA6gzXTvlzTUPF6Yy6qzRUA5dJGuPjZ12j5
pvUeFoiU3liRSBnNcT1OPIpo4FL3L2cp0IAJBv99reP/ib/HClA0/Q7w2iJ5D2HbT9RDnRvIVeev
AFIDKD5vhpJfjiUytL1j98kkco68VCyHhhxy/d9NNeYp43Fw03fESAZF10BWBjBuxtI9QYBYV9DG
1e5POLV2KG/ESqEw57SedLV73kEpEvNIqWyqhK5ykjTr9P1md81F8roRb3MAKx71LSMzeqlk2qkF
fTtXv2Qt8S5HbAFwbgWEHVrKkVvmn11/Q5TXUPbMuVX1i9nSdWchxQqj30gXkd4yfSK630ODSDGm
PlPw9hKQun7f7Xd07uC0UdkNr7v1e5kumVkT0EAeZLAxKQ7pP17K8RPDI0Y0L6QtU4Jvw1Ng5XvV
8aa/GYl21xyCf5DJZsOmOTzNegU4sh4M5oX+Bn8l3aRSLZywsE44mR4z0zqqEGgxUfqHagzj7cmo
FwHQ1BW/Cim7/kHmnD3XNHYz4xSHXO/y+T8ONGEuEzQGJCBRvoXLWSRExMG143164sseFiVZP3p0
DfD1+O8a6ba0bL/zA6OzALZGYV65hVbP6KQ1JmuxQyDMj6klt5cmNTQEdGKXYiSgF6tlwX7zHyCt
0kS1k64bSH3BKUHgmaasBrLjyTkgKnH3OoavCuGF9ZVuiXBQs9MqdeeQm8nRxnfTX01P4L2lLOEv
Q5AJchPgvJowVssKiIk0KslzheBeAGWJjBI/CmGbZRbFLJa84dOvwdcUI1o4vgWOlvqJbswrzCoX
iFDi6C4AHbRqd+H6p5Jk0lsrMWCVhzVtLR1zMKWWjIxy65pwsVFXX1Jj+bpx7kG+qzjsOq4vpr5v
rQwGnDD1kLxH4gEAhvXjlnL4+KeHuG23yDZcFRTOYvSUawLo8eOO1JGa9xGUClyW1pIloG4gxny+
7m/6s6/xf8aq32ohLr1avLuxrf8N+DBmrJEFTQPNOv37wn14DmEGJWCi9H2lfX2d/e20dTMtREW2
erdpc9QMVWP8SffmHnG8WzDMRQe/rBPd8MOROgGWzOJMee6u0c0lJsX90qaXq0cncQJbI7DN4i9u
sB9J3g/31YPOtcXD2H/1VGvqewbTqtTw9EW5U9M+G+cjW+8V7cv4vMQ61iQwIxIfZJEQ89+iJW5U
EyNk8XrcV7dYSfSvXvF5pOkgYPBtJFDCvg69fPqf2lZ6EAFAlUybjQEsoHkSaq9nBkH60nfyxGE1
CzHdAFKMnz0wWJ14SzSRmOFWAZVt8+xTCOa8V60SU5oNk0BbNf2T+Yyurk+B7j8HhiLBqO4WPzva
zfHGR3Ajj9uiNgMkF9TZf+b50rMDcfGDcCmXWmgXY0/onWeOzLAy97COrQFmHgHYNrRzH2yCpjju
/Wg39T6ICTM22N7afHEDGroeeJVa4pFz3fZdgxbdQrOO+qpjRmSSzkJ4idTWEZVDKICJIundjkqF
kbtNLs+SN4OM6y1f3oSOvZei0ODHAmcJJzhF7YynskQHV4ZB2R6J/6mGU9cDRohVqJMdd/O9fGRT
zyi22e8z5fzwSg0hPwehe/Tao7Y1Y11STPBlc4MXn0SngvWa64TpmSy1CqeBUuTsh7wqEmfQAH1L
xVwCC1Zybodm6ab0nC/j6NsKXvVn7bi1RT7OtQKv20vuFDtT9G4rY/QaEgSJSlNCTGvXWFZuCSaR
k+ao/LNDqPhHPXfY0rFNDhJpfetpK5jZtP2d8iM+KXa4uvMdD9URAUF1G4o1oRDlWxn6bHvKocIP
YHIOXjaRQvi2z8E8BFFwapaXpjTK6thbmsBjJOWGfiMNHEUz3uMM3Y3v15MK8rTehKKbEuDhkwTM
F1eJlc0GGDcW20YFt7wLdi8mtDv6jGi4Xzb4ajjs1ZF5JKr0b3hZyX3i2FbkjwMtXVg3ApDkApuK
aoGjNT/62kuGgPrsuuo/kwZH2Gf+JexoBUk0pHHGrPj3votkFiAq2LW6QjNfD1h8zlKbvpT1CWRd
LQqkJAXrNhou8mKhpIhPesEeBSECwSF/J+GOVY73+acTfDSFT4We/DjxLsiiM1ZL1WWchZkC6PU1
t2cOdUPDeOdXY1cRdumuj5rMOgpZApzxCFypAS5K9D4ZN90RuDUpQvMQiImsDB3b9ei6yyKDMnlD
ULwaarcgVZ7M3i+Bcxd+3L5mI1cER+Jl3qX8nLPQe/sW2781kYgPZE8JRv55FXVnpfSWG+1klHrT
wXVxMouP0tukZhyaqP/61yd5kE4WlJ0Lp5CSU2EHslfNzjEZ3kL/FmTwRxbgQDYKnIx+VokWevm3
dC8AuMIL8Sv/EGKwfZSd3GPzxudZz8LDgl+yiU9qyQTQ96dXcMDTJZ96CqrXCbuQuLKMAKkR5Sde
/wEmwHV7gBsnQalQbbNpTNImaCvFDUpXQZzWq+CGGanW0RD56AUbkF70hO7g4ueDgDcoXAby2VIA
/g8xMYXlssIbu5scv+1nmRTbEenOClNYy3TyoFLffIv33oWqkEi+4FnjPVScEl32FufDnDfSnZEE
58jQhpwOhbwrnO5qMwfmuhGOZhFXMVsWEdpQCQJElyjXQLoQ39PtT3EH4zGH7ymGhGRRkzirN5hz
FVh9xYgXT6oxjmn7pEj6WRoQO1a4NLnsLxxp22cGZd4oEwhY+hpyAK+6WrVOhdGlkyIvA4SiPxcZ
FzdEMhlPn0Efrd/k4UayqM7dhJEEvHLu+RLCmMPsfm0FFa81Rw7axzgxe8WKNCyL/0oPpE2/dnCr
zWw9uMs2+CNNQXZXpdXveHsh2mphKpXRoXOaPhOdxtI/40gHUj7bL+S0v8ANh1kpf0Wzjrt1jrha
gL9XSdo7FXPi8ZEtF1WpCLaXvJCI7PrPmqNA+/+PP0KRmnptnvnDhvHBbOsZDYhDOn7p4DKq0LQn
7+/Qm/G1swE4tWISB0d1tY2UhBmkeQXskqdLKARUR2oKahi0xoII7im0XmUqh7h1dMN/6ITgL8Xv
JJILXZFJyFWDYBuzEL4IHNCNg2DZvSp/N7dVztRyjsI5G0HJzu5QGMwIyupvLyazl93lGb7siNKs
s93jIl98oE60KEeN3BitdRr5roONshYS4xP2I9WYRvpfPlKxrIvuw1Cim8WhSnhjnr6nUQLhL8Ej
YmufIH/M4K3XjE2yiXtvOESRioBvqLhkQoJrwVuvjANUhyAfURUBJreFWWr1J67wuvd01XAKiVoJ
CeT/2o3crL/BU89U5pewXe9GQkr+UQitrIoj3sR4My3k4i3ZBTfY+8ObhuKjYoQ9x4F5/QQsNE3e
a+LX5sGwOLLbdPqLEfqIR+XzbLziQwpSqo3idXbxaH38r7gjfOB3MqcnTXjh6Iee0uWQMa4FYPYv
+m0FM3y2bcOK24w1wQ1LohQgwLXd0FBfRi4abqjO43HvW2vjwPcy+R59pxrRnZSD01sQwjd/Q/JC
Eu9zHIx56M+vmLAEHeltNY0ZtDDaF692MPlJBFytV/vRI1sHwJ+eF33EJ8Vv/AYq0IRWxjATBbX7
YdyXb5mugOnx6s6BCVMj5nUXd1ARLYoLbvRoZHUqw+wKwtJzgYA0AJQSKkiWmzYDexjmg4Yjlgtt
RlpU7iRAine07OP2F7ip1AlKuUFmpwBkDB8K4qtzmOjjjOY1LshQwwbHalQztphYqobk2mvjjZfz
ESC9bkEN5Ncmo0MdSAAADUu3LJPdaFs/PqHP+zdtpGIL9y8rc6H+lKhcSTzx98S/x9J9yK8qZiEI
iOQgw0AhW0kDRoxvVAKm0GPs8FlcDXtjPHJTPgS71xicBCRJDAHbJnn6k2FPU/UWh5a48u7TTHij
zM097V6211Rl7c/HVYHx4bwlK+n0M5Nuw4ecByipd/ltrXN3RUTfPTBlTD+e5VFOBMoDkI455FFf
2c8qtfkQmlYjuYHItqmJZS6JrfJBHEttaR20aqvUX8l+Rm8RGWBC7H6czoD4ZIsidm/rct9fXBxS
iNCAdI/yp3KhYDUdvtigjlS+BSJ0Ak7IBCyK/aR6IFpq+C4q4RgSAKHDwSWwkw6AYr3Th0ylp7n4
dW3p87SOlPpAqlkLS7r260YydysC7eZgIEkgwZYwDwSmjtpRSSSOzd4onym1MKtvZS/cOx2bTFAh
GLy0atMetK36QlGu7PqE5xNuj5wf0sGDiYTKlak21a+9wjalShJ24TWel/VgMCEfOnq6UF5CzbCa
Hyi4uewW1qWrlhNWKQSSh6CA+QkpVQkS/o85KsB3aal1kolX0uLHwRCMSmr4RiyvNLyLGhidYJHI
NiZCvpYqHkXXyyZ1E/CwJnWMOyfD2Kqh82NuCWh8VFalvDFMPIroMMUhQiHs+6te6DcgU5uMULXE
rO955vmL9RgUq4khg6YnWriD0Nn583fYavphPWrqG8uF8+EHpjSgAVdh4zOxLfO1z/i9ABjDcPE+
ITS+e3I1ed2rQACHJZuXMEvWUDsK0QAya7UERwCnD+KxCbOq+9E7FB9k+vKawZYLv+3bA1d83LZJ
yGJsTIBuj0VmAWHNVoATTnhhx2OawiId/wcDq9bT8ipcUvyz8mlLkIERR92JyUlYPmaOorZScSTX
vKAm3Y7jpuApZW74mE3qYh+HOEIVN/fOncvCVAYtrBO3sbMYjcMxx3qccnTrHDAcLgEkkUx0aHQc
4b6JyuL1/z73D0bzfDekaVFlPL2rTmfdn4VBavtu+KCoVEPHqe4Yfln3djuILBawD/687luAoz4r
n8IINqYQEY9QHWAm0qSYjftyQLiFy66QrvCSPmJLE2WXuEgemZFByaIO80FpWqNnSWiCIBsVvz5J
trikps/VidVP/DUxqLqB1PXQcNnMnvYe3/Xa7pTXQ2vCVE5xAsFu63DPPih7VvQfSazqmP9ZcIq/
POH5MbDPUacmRxOxiSaWSSSyHtGJoy6vonfUf4/VJsi+o+KgHxCctQu9DZ7bFDeSEfxA5EOriRbp
DSDjpLaY5xXBx4GtqkiBVmTLeLMEeLdnmvfr7GFSs+uCWdZ/tE+OLe7WdP///rjSztRlKkBC4uZe
yfwrbcPgGBRI8CUigN7IOvdybOUtOzpA6cyrSHAHuzgV4bG2ysUwc//yQ9eqB78k1ql8Jun/T/c1
vGkHCRJAvM1mrzmP/IiHYbjVtmUKauPQc7hLHqI37v91PeJg/77XIofKD+KoDp5N8UpK8m6R0x5A
Qk4pNU8OwxAFfQ9Zinen2NHRMXttILUq1U+doTqwVgqc0Fr5xNVqi1OgqH+MeoGz3pYs799MWs5/
fl/LH53yGPo97thJcpF+j83zYvJQD6xGSTH3DiI0cszAzIX0uujhsXqi21bqloKsLg41/6Tj2hOZ
0YrbR1RQR8N9JyCaU3YbWYVQCUrNAWRHxpC8bpFZ47hX79PNDvtYZyF5TZT9SpPs3LtZzrJpEyb2
AqxuljPRoocwUbzmKB8sKZyBVGG8g4xZFEdeCxIT9qgaU7mfUFajeKk5lICreIIqQU1e5Sbw5jII
LQjWd2zPCbMz6dXSO48AhmcrIveEe5xTYnBfVp6zKbd+7zdEgxNA0BwbvIvJS4PS+t6a/ibj3Y/Q
Irpph0uJCXVQjtbc5F/dij1DxlTTnBPTh94JcDgdJb0OFCRQnTmR8xdZB6TAoFmiZdiWkibQ7uFG
zOq3NseHbFYz7s1ztXRYDeScIv8sobvrIsazTInjbrTy1pjMJsAm6MgKXekC8qFS2QWWSm4reS+K
qwmbaksIHEZvuOFdKbXRk1ObJKwKXqBBxt8wKk/7D7Fd2+3CyspV1/Qf1t1j0h/Am5DyKcR0LWQF
KumV+iPaYVQhZfS0AYLfZ4d7vcV4IdfbH4h1SWodACpSxvtBbLs1yNMo+Qa1J8zxrvwYHmoUM1Gu
xL1uA4xxnjQhFBuyuIxjsJE/MO8+x+ZDoLeJNpg5qmpN8NtZ8UFb2v/LCFQ6cbJiT4uSBSjWacFQ
t/EhYRoph6QPMNNBIY+qT4xcthPXzkTt7q4C2bgdRnALjPK5ke6Y8ORqhiIF0SCNepdHU63XB7tJ
cgd7+NonDVaDXYwTp5fukE1yApHKk07p6xfN/P1diseK7VkdwO6VjCRXjUE2H5HFEubgy0rHyZDj
A1mvdsTPxByRK5o2Ry35T0qbZCiB8UTJrHpVpzI2Tw0HtTIzORk1p9d/eWsI+ENBKCOdh6cYWQVG
S4qa9dEdp8DJ5VXOXfDcm+XmUH2F5FCrGCs6wMkrjJ3sGacysEGobQehNRpCKcKOxxg5swSdolcq
88FRNxsaecDWiiKCZMviT5w4f83SgPdng52bzVeCFi7w6f6APhQsPK1hjvtWduT3P99QmM8mwnNi
vKqU5YdUjRxrcFtNOfcZh23pMz/G31s1ZqESzgdjL5C70ALSWyTMn+Kd9jEPIBxpkIt1ICrnuw7s
Po3MFkhgFza70a94pJBAVg8+N/HTq9vXUaeDrmECb4Z8S9mij4FlDPN/I1x3O1qJfr/7T2+CKD+B
bwK3dNOwkMuwcaKI3P9qlQBUWPG64PROgon92RvdkWCv5VkMieave0KGc0I0z8c5hr3lasRm8E/x
0PqMIqLRUgV+ZOmFQWfy0OSIf8hwHsEu9diUE9dnttGbnsVzV2nzEMyRik1TYUhpbK2K3xHWfDBw
2bidC4boTga6orRMy4tg34dH6RQaibm+NSWHml/r6URgZANIvw1sR+AeYdzjabhQMGi/xGQhmySH
0zCD7Sv1Hnc4KA81MHDMAxGh3ajbS/ijsh7reqHS+voOBNFJvxytKNuXMI/QFhPwqRdoqPzTQx9h
CfSz+O+dRU6fPmLX8LPkVp5MTSBNHiD1XBsr//6b8rw/9rpC9uaE7GQ03DMqQtZUnseRV9zQZMNS
SCwwoRbj7YsDBG2HZ735BnDmwL0KN3mKYm0Z3ttg/j2v4pwSdWzZZGwzbOYjkMxF81FfP/kODfhT
QeLFVj1BOemfD7lalPZJ/wURkFXA+jSsVqSAu78NzzuuM7PJTri/D9hagNA0NWQtJuu5HWaIhiXq
fHQpOQ/6PWQsscq+Ecn8KvVEf6W9vVDAyysCV4qsFeRAIZJ4sktog8NcIJioxV21oS4PeD6Dv5f4
cM+xwvBX3CiS0fHuREDvRCY6K+Iwnsh5Qh5GwMkQE3FuHXsshlo9kXsAs0y1Lm2F2mvwcJ780r6b
xZlkxtpICqGz8xLfZkHdAAB4YKg0UyQsZiJrmExepTT2Dd/NPcajb+0GRgGIgRk9VSz1pqM1ywhp
xV6+wWm1Q7GVcE9EgYpe8dy8wTjCaZ7gi39VPlIn+6ub4//ZGwkgUkzgUfZqGDaLuuOmk/TAsL89
o8wEtsfxjrMV6+5aPgU3TqsOV/UbTDcLjitlhLkfsmAQ0HvhVI3VVf5YTmsnTge86FeZtA+Bcwo9
r6kMHT079xiM43KxuHAUjhBsa/v7bvatZOvcVk0n7PHs3Ngh+G8khxOBmZ5PA1NY7DPwmtfvDS4t
pVaGIfvfRyMtrCiyn9Ll0PCnAHJTo4+CYeGj8yB8Y3Gl21koplqQTVICpNDl6Miv8/IK9Jnn3INh
qA6c4oKeH2U3rSaF7vsJa6Qd7I/DYmUus28R+HXdn2wtiRSrkAu79HDpXPerwNDcqkrSytrGhHii
0+g1XKXvIjAFCFXOBzDoGXKRjVGdw021SLB8u4HqUSLclJzIJcjH8szavrzvaFXQUiwwN7q3WA/A
gZrbaOkuYKmz6VzWu34I0fEbxFTCp7SGeDSXWd56PEW4V6j1T3uAPzGxAcWmN5rGyzbE3R6FDsPX
PCtfiF5hejCtmzBITtYjgv9MRJ3tTlgfYHZSJkpqf7jm0SUzcd2NcrJM6DEh/JBVrZGFuTUMqLg6
OQdKTPJzcn+4pdqr7JBmSxvZDWPH0ee8RDr9rcc7hBL1BJur7K1N5wJVtfmIS2zHvyACZHfFnqnJ
ZsXjmQn5iiPZnzGeikIqTnzOTYGR1hcKdP2k7pBNZAWEFiWdMVbAae+K4XBCaLLPHdO/3iILKyxD
B+JkGQ7h32YbhlsOaSFK23GWxXXjnMCpWd+WkRkyjdxBV3UAFoKAD37N/4kmOaODX7ctVYtvwyiV
0fNzKqjaAdcPqfHuG+78IBmLX6OwMhEGBay27Yci93mT7r5f0IafOUQmKMFdW9BTim8Sx8c5sdVN
X3BpZpZrqzRnnUQUcn2y0F4koqls2H70bSjPaBMGN3KsC7+7ixkxkVLv01UkOMoFU3jZtrCuKORW
EQJMabGBSIHI/LoPhpuKgiHphZiCoG977VoSJXNNDzOQBN1CFv4h/DnSHJiTG7cWzw0ebAUTeShD
CTCIbxFgjvOBXgDRyhOGCLgaJFBnQem/clKwR2a70uWNwgqokYP0GAdHxh80GqpDlhPmG+joGbdW
slqabvtOoKdOuDnbIWuvTONOOT3KJk/JHg6rNIsfNSVBXkfP7nn9kV8037BXDzsDC1yYRcS+0TWh
dCvGaUb8OPTKe2qSzTRBmbsfdAKoFQd/k1q8QqCkJ0j+vt8gI501zLH0pvbsJNcTQduIdRUcGLNA
U2ddmSSjISRKS61UGBSVsw9ZQjydmykpoXtEKkNPoJyG6JVuLLGIKUl3NaNqElh4MeI2LuPFTyve
wWwRR3oapeT7w6OyQr27v3qEtG96Pv5fyyqgungK4vyZkjOv7DpS7td8d/TkO/8ywe6fucULmE0U
UlBeJ2DC8b8Czis7v75a6zayfIQ6Fr7Xpzc53biUEuyj8RSjKIUnQo/b2qa46rYTeRyGVa/M+P+j
xmM3o/aXgBHkI5mCNv+ryw5XBK16qMpTgc3PwEOD6vLgTTHubMnttsuKl7yBGOJr3nJnSw7+L3hk
hxaVECNn+mbI7PyplLJFaz/3760xlF+izh9qYJIjEnORILqBUf3zzAT0IAHT3+aekeC1kblPfWpe
MCAwK9Mj7nhg9PGbLywqxD2gy+v+pGcX8QsTmpJeXzcxH2S0Wp5Wd/PqppvtecWhnpZkCKq1MZEj
oQemoB1J9S+yawb56GDSqRjScM+hJl2Dx6DJcDlKj83ViDeOapEUHdo/BhMlGk/DYHEW57+AaJlj
EemxSEtl3nx+AEntzkjccMx3Vc0c67WIQRztu6ozosXGn9i/GZQYazdm7IGObmfJi/NfoQzY6Sr5
8bQzIVntUgzkZVEMjKFfBqADDyaqZN3URSFxp07QFNo4XsEHS2E3Fj1689y5get1hMuJ7XJUiVbZ
oEW7aUwVxGQZ8EV1a0Y+IosBqTBqVEATKaw+1BuctkA7k+CEvOZF5m5snOmm9KhQb71HMV2umJwi
5g38Mp8enhQH2HTIWC4tlxHQXRfVC9TtrEg9jxEjs7FAnQnXDHy5kIt/5VgLsY+aBrMQXGO/tJSV
fjY1h48jAD9RiHj6VoQJn1LMUHpiR47ZFl6BQbEmGAzBFPJT1M66SJu0T+iPNQSwRTd8kESycapu
I2KmRMgD4A90H88FAQZMlA9Yaz15bqhPnCa8a2CvrFYYPnRkvIgAhrJMnZ5phARFX9OWQja814q4
aQtBhYo/lVAJ2YtVbcezIpHH0OR1WahIH+HRL9zaQa/pSyUmlVwV2uOB2W0LPrFSUJYLjTHAmVmt
fe1IufrVvpg5Cb1cb8fEORTB4CN6/76CkenxoGV6e5ZN2NLsL+mep6EqnolCjoILKKfCdYnhrhU4
un9a+KRoczQgUCBNWNLmbWC0mjn8cjZHnYA3hl1nagRCQYUPdvtJdjkkF4lmMfzFWGBDjHoDXDbz
FGHPZZJdoH5LNW/+EXf54aHkRrU+Y1nBNfYS69jm5bXbU59ZBU20TPrsXLNh1QTQAeWDrahelFON
SOFqofqVqqnrT4phtXMpBrO+G14HsydNFqpI8q+EcMrv9tT0ud4Fk88FSOppi/fdm0Jhgko1iluI
9LCd+6RF1vPkLNHUVfI1Q2BB2SDlvrNGRo5cRcp5VcPNP6p9FW7RRB4ESN7PHp9GJ2j3D0QpAC/1
dwLTPkKLalFmQ3YjbYkTf0n/Wa68yD7LGSCaIbiTg93fDjlh4KzMbQnz4+bIedbVfEpIfWRGwVBf
S2kjR+eFTtkFj0SEbiO/oTFnIUuaL3RnCZzF2XbPRFdRc81rjvZCcwmX782q/pv2/vVwr5HrRZKX
QL3eJY1sGLyvUOYOcm28Zh/u3jZ5MLkcedtU+2e3wQDeb2iQQTLKshLxyTvyBpGUUlB3kthp8IJs
0odCmugLTQ1SBEJJ8OLoR3ZqgoDDWqo61ft1Z98cB9SFDH87GZ0tghwbF/1kTjsSxfr3wLQLoRaG
GF0fJzvxc/5LkARhwqToijjnnBjCqBORoSOxmCSr0BwnWkN2UN8eJU7jJQ0Aq/pgYMSuLmkWVEHm
9c7102V85OS9QLO4tBwLCoUPgedIkOWAOorGMtFU6wAYjcQ66eaV4PFMql7BBGDJ9v8GKcKwfdDg
O4djE25fDQWdQxUHNzBoyE/t/c3gwvoEB5IZWR3luw31YyDLCYnrBAmt56bPgKPdskkBla93P6N9
exCsorQlqMNUieXRY/wEHAMssVrcqxKUCi6OaHl7Qics0NEHcKK9YMuuLTLVPjVKI++eG0d326Qd
2NG3qonfYaM0FH0H0S3pbM6jhl9xrQbp/1JSGFS55J1qc1MvjpXQyn0XVzq02m7vOStcbinW9hit
b9inH/1im00dumXPR8gs0tlnrgNrxZCjSkY4lYP9W55DmBgK2SoBmuB9STS5lxUs9Cz3hC1fmmZN
VQrJejIzXklVT9UrmRPKzS7HaaxHkyylgDJkB3PSEuqodSQyN0+hDBLWSeDBqO8fTmu0UDpDKSIv
t+Nsa4983GIRBJphzsg707fjRXvQI5bsAgTsYbI3R0+R4YVNXK8wMoQ+P3DU5pmxpAEG4YsNjK51
ayA0ZfkaQmE8wTjOC+Bwrff61fa07oKi/sZ5wekQDBJxbR3Q9RozYjTRo6UDPyGhv89U49biAq+T
z4qkJAAg8G8QgQclrsNr4VDCRorWeYBJSXdcwxgpC4cAYibxTgW5khUHl2WkJ8kK32vOhDmJjL44
UKPJ7YKTo82ZiWMLmqhOxQOqN+eE4rr4KaZMlErai9D3fmM8mhOcSeb4kNvZxiYJWJ+Y14eoxeN2
mWDX+lC10KU1VUd6LKIAbTI2vP8r8C+TVLS58IzfGiSG3e2QlJ/DNh1UlHFugkEUCECvHddDxIjZ
XS0CUFDWXjOuuE+rdrPXJjL4dpLMUEdabpt0MktuHaC65w+xm03QXDQ5mC71d3rT5tShBDElU0bX
+oyvHnZUdKTivlA7lEhWZ/KrVFVa+71FYi9gqafq+b7FAnmkLDbJwKU1R5UekUqI47wxTruzukZv
ouwe9y8RsS9VJwDgRHC3H6FO5pzRBuUypVw+GvBu0jiX2161jdcTJE/1K1RQCJwz6m5TG2FXp392
9glOIyS2jzrSQTZk50yY9P4VNzyvXxzmeqLzW0HgZ6+N8BR6ark8CatFeq9cEkgnPNNHwoJZH0sS
ob59LbQFqWw0Q5YoG0rTIWhukvWT2oF8eoRXAMghbX7T3SpVXrdX2Pr22PPbFCqYzJHqvchT7Shr
pPwppSJcdAAmWviqjmScMJFOjZatDSlIgY2+QJFNaOLfpzMcrrUBeNGEIe29wkKbx8U5n405N7Nm
w/xRIFeiUro2WUIY/osDT/NsaE0HZOLBPSMO0GGFWNbERIWUL4m28OJlIg9hOzaQLs560iueM9XP
orchq9b+lHVYwlJVA253hS7YCXjMdEbZ1lYQcPuj+tRw+PFWo5br1cwkGvzAG8ctsr9YJ/3huSKz
J/9C722+/uYUoRmE3jgDOBY7V+ft/4/eVRzTVoSfMFQ6RVUcyQsc/zGoV35KfMRZNnt1T2OQ/Oq3
vBiy12cp84C/raggp9oKBepVUFtIsWg++pwcENStk8MMSSr8lrytjrcwLfSg4mtsi+viOgq7oDIm
nP4ac0Tgqjp5C5a4805e0oSJD+uhLSCRn+2SyaHJL7RD70AELfpm+RZmRCrulOc4opbNbJZGsSyn
KVgfeYOR5pTGkHSrbMJnF+/vw88L5CID43fNsNFLPUIXC5Y7mXiNc3vJ5j8a8bVd3WXG+eHG21fi
zFqwvxmQ2QOyUKngSmGIVjidN2btTgJQiYS3+gs2WJvkGJelotsZHKh5ZwAGAFKRdw89ImxxhZ8f
FmKqO/GsnBAXp/afV0nt5/Gbtey8VCC943TZDgt5hYHQkcd8b8YqEMLiQa8/A9PUnbWRL9sE1yTi
akIWnUaHL6hnrb3rhbLi1vpmF0i8ACkwKtBc11msrODxWU8SFLFvIuezFZ0FpQLNWx5I73eRV7fo
JqS/66qt4AmhBSkEugckTdBquyXociiy1EgUU9XEqBF3fQ5hW7uErbTHP41GIBMZfQzsvtSpv/06
Kwb1X9dH1ZmMSkGpgUxsBH+LncWBL/4NQ/e8Tq8iB7qOhUn7hMaozBxCXI11YhOLEH/3uzwyILEB
zUYCaCoMn6dT9iXLoTGRfntmxxAE4vTVTfxW3xErCMBfP5V09ltu2I6DnK0N5QSOz4/vHVbHffQ2
7J2/8C3I+Q+BCG0i7Ie6qSfANs6uJEDu/yF1kBoRHmEjzC+aQhz2dXFOIYbBNSvlc0TFFOdvFk+r
G7Dk+vRcPwv2yY7G9kxJtjnsFSTqXfJw+Q4RfZeJ5THGLfsWmA6sklZd/MTLHqnQ1dvo+vxntDhh
vjqG+2DrIniYGSe6NopbcpUjSfqZc9cck4Z1qYSa4vCSU2L6P997ZaqRplpcWy5TtrgsCB+KcSoG
Dq+B7F0vPIClCpJa3NtwHKEmvt1TyddSUv3By2AstPW/COAvxDL1a1D/e4HDQzpVABITruNoTf0c
G1kwcL2iZkTrL0MZLT0Ncz7YpilaBAqbcIFrb2ZDXsUpenAt8VsUihkNIR8tfbXf6se1nl6lAaTK
PUjRtRoO/XkUM6x9KHwhS59OUGq8II3VsMbRu5bq2YegiJWW2FP9OrQvR4A8J7cuZFqOJiePfdCI
LiqjOVu+kr9DWuMcKFbA7rqQaX7cGTDjz5oSxcHTFBYhFN2ioi8MswKb0oyjijqK1iZ2KfPXeEHv
PInOx+eHL47Uq1l/8gNRTj4IDLjkFQ0qsJOVyICzObSiFn5MaWAZXJ2V99RlQnUHGt0AF2UwptK5
rIIoB13M9viSR99hExijsMrTSUMqHtsRjYtfizsVoyTcUFUvDKQ5W6MPaac11jYRhnfsU0i4lzVo
xNt5RLAeWc9grDrFt0eBvvw6FWPyXPZk+XVzX8DZ1SR7HXsmJLzpxQu2l8licYC39HPvCkxtGNwM
OeuMFSdjXMIUQ9Tg2QaZOgDt8tfnzqGXh+EkKdlPJ+Zgw9uYAPRERm+8fPIyV+KMTfwzlb+UyVKU
caD0WXy83TXzDhW9IEtQuSXrBcWDQGO2lACyDPRD7EVUokuyTUE1khjxeuuVZgsHsyFfRc2uWOzR
cVLrQXhfFdooRabh+YmwMJCyStvH5TS/RGA/6NUslEzBPvGJeibXOchNqVQ/l147wcJmRocJyp9t
37TKxKjpVAI1JWEk6lirGzGm+EzNPlz82PlgQn/G07SlAyttYrMYCNZPSuLuJUUQvp/2T77mW7kx
5XSEWfpH0nsR852y5qTIOAUtRuRfSpuNplXNfQucxeuU9t9lfBda1JYzFCVktK4CILGnMwRUpL13
FWULAaa8cqUVK/3IYG4s2W6MK4I0BI+gDOeK3xjlNMaGfGMxdAnN2tOR3G0pUlnf1yaIgqRvmhKp
yvmds7KotKwZnD5LWez4pdOLE4cCQ5kGxVEkwxtUk1sWIENaEqdveKMG3BFH6gx1RRhiZyqy2cg0
/VpTMyz86M1RzWuaBL4C5L0TehUjqS3pu76lPZtzz97b2BBUn9LIPs1NEcXG7MP88VIc+oCZa6re
lbLHwGYaxSmmgRJel2mawMhGSoF/e07fFYg/GbR1zDWcIyUZ2PZuKHqugjwrqaR7AWUrm/XZVxOt
MqufPaTFiSK/VyFOJk8SU7VVGNzt15XjyuwEmgHwuf8nCDQH/qP77txPGmmofOrKY2wEHiA1jZnb
F/t6K6pIjs1nzQWlr9aacI+vI32PE1eONiaSiVcX62iQZUGpQeAU4ubzhvKdmo7+ZCmRyubQtFlJ
hyQdlZzgsAEPqgUTbhKk3gGK0ItfiW68uQZkrUip04fADNGkFImnTAxO531EpioOVY/k9OvRoIqn
c/sMqSYSsoUUGskRs+ajl4glpxdycCMkvjnMa3kqJU7qNNrow2x3cNYXXv8EkzoCRK/D+VOxF9Gy
Zq+doAXGW2VyRVxTSCRE8LHDVTfFMIhIwS2GrCa9GyIr4YEZyZsLjHkvo5q7dmppVFhIt+r3hw+F
PejP7gFCoXJ68FFC8bSU+U0m7T7bubjshTOe9P+JV6DOjAb/JNSNzQrWa5HyO95dwaPF+1PkO2vl
JyNHtlJZMxusA0Vbk3X8aDaSE4L7SjsPxn59ac37/wHYORHRo363IDJqYrDYODWte08eVru0ac1S
uCo3l9o8E5AEQPS6dNYZZ0cEdjReLZd3xN4JDIVy8HoMf9/mt7wGPSFiLrW5gd4uePMM50YfpKU/
4W/wXgADpJl6F3GmMBQrTa/HAeq/X61+X/i8+5nOnVggpaYvENUJinPnH1G40LZXCqsfdiE24wCw
azCy7DcHcSZWKS4ny7GM2NYpUFteUG+InHtrjQJYOu/vWSAoBWZWqNRkHx8H/+z1yj1Y4T/pMKS2
iAFyVcErbh2nipttRYBodaZUCMre/mnxnk6i69B70L9FAeIrgHh//PSHoZa5ONW+DOFe/LgjBt5+
TW2JxaiSpdY6r4Y5Gy8ml7jsG5oCqBTim8ivH4fkRXWuC9FQS5RsderAwQmeb2OGqXICV8IKmkTF
BG8bpVZiGG5VRwjKZB+n7oiceIab/mSiN4wGz6GF/olQLxl1biLFTm2q2sN2b5xj0I2YXLSgv6wj
KEhPAWunPdH4Ljkx0ADyQtjlHUQ23/+E/slrdKnSmhTp0ugkL7h8FK9VGPbEF2SIc2kP/6u3qzZo
FUVV9Ef4Po6ufEFC45WGOuDgFAaE5g6iz9thXDfFqYE8g2ztif3m1RgBl78QQje+LQnDRvBKUmzc
/T+YFaS9pJ85ZmyB4m7q8Awo0/6o/1EOHWNRvThIb1t7Ba9GGbZ9dn5mvu2Qeriz79FrsTdbBF+H
jEqI94wH/4VvqyzV8W2fZUWqHVqNrmKqa4N6hg77NAs+uuowCNvPpsNwPcpuZiP6Otlc043RJ03q
dqmAYkxbb0c/1Xqx3zpv7wNcCvDHWlCwnfrVtRit1D6FYTWN33F30M+vLEfsJovtz4xOVitzzkqI
t0XCu+nc5Z5V4qhvq1SBtMous4vGE3ZNF/A9vZjFy4o+UP2tCbWRjUJIlPBcM51r5+qVADtnB9sf
x4yeJfBthzL8SAgHEy2AqDMglASmsmPmdSdhemjY+82foY2wIY0DEUb1v/fziifWgROZAILEl6MG
SyF9/qHFQ1n4epsOs/r65xQNj80MV+tCwk3djoKwTrYmWQBHVyZOxQJQxbOn98tUw/scpfHoNyhu
9zkuNJUx0X3worZxKEJA0kT6T81EioyhNcv0RzfbC0DatCEQ5D5O0cOuBqld46emoRxZXUXP9atH
3JdvsCjocFwNyJieMRh6YidNUNtzBEKkK0Xxx2KnJDCTaFjsXM7L8ln7SC+IPP5cNhuUJMLSfHuz
rK/JZcP+iI/YVaRDgajhzge2TBbuXBHB8LVzwREZZQESSx3xAt+J6b1kT4hZUqVkT9hsnaghK5bq
5A/46OawXfkZwaEdE9WETXow1nkJ3z426UXb+A5ZhCd1vTKwpY2ZPgOSdgBZCVQZsUEyBsAgMc8U
Mff0akMf1Q5J9XB5V3FuMGKvtPSeSPFohJKAlZd/5y360cWrGDct2cOZBKU+8hwm2vrhSuWTEK5S
I6VJt00i+bVTKBN7sdlsY8kObLQDCdd154dY94VZjzVkHH0+nONPTOTM1ulHVGOKMyyt7DMWzzVy
kyHKkIqCgBgYrk6V+2i5oSv8bqafjtgrNnzZwTY1Gm8owNWGSKewOtpW00gw3Ijc3fL6lqdX27Z1
axbZESHJUoQzMzYg8QSX5vTLCzYUjtyz60cODqj9anWcHYs3NChsZU1Ud66P/wsRj0hZRm2T+Muf
kfKZgC3Vtos4MSPXGNFMh5ysak+u4blBTulr0gWb1OX7it9OKZvJPz/mL2dzsWgKfIP9pjaXCqh+
xf7X+m1NE6loJkMV0vxvOwsCTOVUncM+z8YTRh5QDGX5Mi2RnCCqipxHTXBfXxpO8kZvqI7mLIHc
qWFhsyinkm6ffNKN3pkY+1BZ+6h2uDaAltG2/lnWRhQ2O5M39IZotkzcjT0FQiE+K7NaxCOP5RU8
PdkaBbKeG/LYXkC6SS08kYHrLYs+ZjBeDVthVnA0kNFTgfaVOo6oayWyK4qIBySkbfqLdpR+1JMR
yr3iDtsIdWn/GyGOgwBOU8RWA7c7zDZdxxWlSRTMhPDfcCuL3HEWh3kDcRuLwSMTSz/PbunbKNMK
S6uYVbz70D2DGHKhT8kFdUQt3T9mhMfeG89ubA2X1zlQB0rwyp5r+PQTS9+IOsK4ufOfe2NpYaTO
Z3Yww+FCBLTxeB84R6iZQOSVvVPybTjgelaI+FOQFTUnoSwdSxe6B0V3ftHhrx8tQqce8j4L+qps
aoQOY1cA8zvTeAIeVzkByNqwliHFxYuZOIA7w6PaYCPyOp7NLu3PFFKy7dnQbWCRIuFj9VzRZ41L
W2F2Y0I0MAx3De2G/vy0axDmV97GjtmazUQB7TNGvpG2WFfQq9DZ38kBH6xSaT1vl+1G+C3XNwNY
jHnC72hJVB4uI1vf+4bS8I5R9oyronLckWup9O0VG3U6tmS3DHklXDkKRrzKCTN6pDr3rNNtuiiG
hvZn3YE1VkJyiH+CbTVnUcmayTqKqp7G04G4q5jkJVx04p1VMtC1xWIg7uv2G+1Jna2w7WQAiU/i
BIab6Kl4QTWm91rXlN4F+S/aKS4UMT0Yp8Iei6pWr8l1gm8my41pV8dBs47UVyOcLkWo/YwC2p13
1+whkkMH+i7jksc/5WFDCdY8LCpc4haw77Ch8eaSmLmApx6wpdfL+RqLY4UDUYNfWSO8YF0XH7aZ
REOnQqyNVlu1756+jmIRWiUp0WaaT27N/l6RlY4xISbFgCftbklkkzhmXS3HV2xXdMRGFaY5PS9X
aZtIHVa14dgtTXwJhf47cTMzu6rrx4ytTCiYvdlbmZcefKY54RW1vhrXdRGP/TYFXs8LkVyhdt8H
oOZkdKj3QwPhZkFAPMrH3fOgLhsqMUS7Guo2xUlsCQ0FZP6yAhY8IuP5Z4ZivPP0Ej0fG80gyP2t
bApQGhbJWE6gFmqWCT9KXh+IWuo/wh5oapMFR97HXaVczTXU7w3FaLrqB8CvhX8Asri0mNso4Bsi
aMj3xgR2hrj+sfL98025RHmU3Ce/ewwQF6aNWcdG1+VG9aWO0P7u9DQrmig8XB47b/vBYxJpv7pg
jrYu1ZyHD6+wO0xMqIZeJMeDflGjHegt4PU+2v2v6Kb5vcs5CpUxHOy2UnoQoPeSi6nPRrMlRTD/
eLiDkCxz6wLVT2CW+RWiyWaV+iNQ5lRmUfSThTYoO+TDK8DJD4g8NC0DcENMyjSspye4EfDtoSTt
5n5or7Jo0XIWlSeDK/0hDQ2iHcvJQhF4nnrEbrXTRNcS1HsLDBsKSCY8S1/oXruTsrmfxnwEEkYS
PTawc1TWOlPs0sA3Ii4ad4A/ZoKb90phDjtTJF7FvbBJxTDQ767ddJnPQZT8RBNlBS6aNC/2LxEM
8IDDNy2lCXUAVtMAh2UR5cBE74qc0Fj8xWae7szH+4ik2k77Lirf62YHWF0OJGfql92v4lAGJb2z
pjggn3hrPp6VnF2MZz/EKKNWDmHaKlleBPiFItQ5ZJ8M7ayVufE6ZZRvE2249ReI8IGCVNlEYB12
iCsYAN5SkrBcxrVQq3HnpKGxFJ7uFYHKN6cLo2t2L7l4SnKkaV/i4vVeYcvR9xnAJ7v+YHFjtukT
37iy4AJogVrV0aBDSXk9ZBINkXTRaMY6LtTVadkE/VAEvugc4DwVwHEvf2/a7m3KknqkhwuSmdZD
n6HdLpTDpuJ/stkksNapl9xOlePqgC2Y0TkPb09zkcQULfUZwa/+GGDYQBK17QVD/k50OU5oa75G
sIqcibPAcN7nQBBbUnkx/leytuWdBfcmGfkb6bOKbJ4ESDBWTzvLy2uGFL/M+uGlZScjZe9qMq+7
u+IkFHX4lQW4cCybEQPRcAUadP5a47RdKoq8uMcQq5uYwfCvq6Zou0I5nV72/yWI0Xgki+D2H+LG
0gNlMVTlD+S64VSiG4+PXt4I8yXxcjaYcCnz6uJjz0QQM8BCFlAHdlAbm5oFNdpX8B32hhHeVczk
DqcFHaunk4u0E7/70q6dVNKAfXry7ZIsSuqDBZJXd9el3dpSe946rBditzqSTmml58zL8EdEkiHi
S0yvd4JtU8n7FR7f9zRjVy80EntOmhnaCbc8a4uixfPmGzTgWZE1oeHx+uew6V77ZNNJjdJqNHCq
UBu7j9v/WknQhNM0Q2eGM2EmCHNwsThKk+AIOoCX1OqgUekP2BdmIj1ujIQ8bmnf6JSxNjcubYgF
3N58qcdwR4ZZkTUlJy0obCGCjXD4nPgk7KpYTs6FUINOPOuEvGlhP/wkOfri7ZXNmGhSHyvsSiXL
lCl6VLSZthS+GL+ZaUDnnJ8+G20DMZzovnasTmRirbetHhg7/JMUpzV8/wIZ/hOVrQs7UrBIAiNq
LLDSgl1OEYfVwKB9JtWN1ZI8pSid0oBM9HaA3U4xFqIf3cce+KN6jfVt4MULiZMIieHZVjb1RQLY
vvN6M/Y8XOM9jfWWSJkWNf5Eakqvaa7qhmAXrcc3wspV+tR4IVeccMYjr9LC49Mu7g+EAzbc7K2G
RVevVVmjhwFNfMeP/skPGizFaF4FRvomQVmpPUT8JNo6Mw9N1bnk7f+dxGl0BIp4wNAhQs0jB/CX
KAeDJWiT//7CcOrwu3i+Bd35z+zDxV0AOLI/jbMAvnB/srFgVKFY8TJLFDdaLVbaxW3/2Fwup1Nn
Q7m1hWK3iFGRbMfHTutWUR7atngv83J3jv9sgVDdNvs3LKiiZYFzkJMVDeadZRtNd7TYV1pcsMbc
xvr8PjJDyO9g6ied3mlZ4m1Y4FogMPRAx4xzp6EkDXf8qtPU4K1G+Q0/CTScs98dVnMXhetsEtVP
HawMairrT99wxzA1tJu+LlE0Drp3TrHA4UGS7h+ZKF8yWv7OJnPW65OvYTk0H7R/nImWuJYguiCk
3Wr851Tk1nMo5+9o1NeN1HqAmeM4sJt1hVUTGDMKrQJ+cANbGBMx5VCPumKSOVswmyI5UJ0N99Lc
GoYxjHsj8y9TpkC9zTIwwiocKNmiG6y+PHmOEFEcYCHET9cHvbQrCB+KinHIJf0ymjBHfzIrecrl
rf5jO9LwKKuTl8GFpf623IidR6LllUdTMqqcU9BdjD/1ALyO3Vv5p8SykumlGZyRAJn9doH21y4g
lG8iPQxHTovWlt17ksUfR/zPM/liqvvvMtsCBm2Zl98T15t0ji7pVnHgn12hAQ+9jusxv/SWa2VN
CNNR94htlQ26j//SEoTRIn/KtjJM9d7E0u3lEdF4pUNqY5hdZi4ULVZ98sIGUxiKD8sWjI8UfkE/
xIYFvZHpTPmKrO1xiwHKwi8jUfYcQo2PGzPTw1R8IPXn4tnNv5JADYICxThKi9uALGe/fe06QzVw
3D/QkMZMo65zs3qg26Ce8V0/JOll4WREba5wki4UB3fA5kX5oB/xDqUPRLkX6kAXOJ7L243WAjsC
FkvPS9rvhnOcs8MtPLGpFyBKWrlBSOTNO+61FBdIjkLhtW36rWljccchyKeGmoQkd6f04q4bMjKH
43y2fY8QgH3veOuCLqcT/NsNyxOJpXl2/HByCLcs0YoL2cUNxA6xFEL3XDqi05rTP7YqguGy/V5Y
iwyEsOGpuOmV01Z4j0rnT9rlr9DVj2pK07m/iuLhOT9lZuxIS8/xSti/LR4rvJgza2NfIwjC8JNY
KiRYFzZ1b93YFYz+c2A3/YUShjPoaKCLTFIRT2wDtn+i2l/lGMNkMfTkiC4+2rofg2aR88H1shx5
BuaavsXZlvXjdb2pbGvEBeybELOcE/iYkD2jXlLrOL7ZwmqCl2ox2Kg7BRnB6VT9h2pukhCKXnPm
a7tMe/PaGq+vntE8oq1krVSoirjqObkSx8atZwbkp2JARdKWTXO2u8xAkJn+hLZhQBL8XJZen+YJ
azCdi7pRnvYs7Upf1kUvMdKR0d84HH2rRMLkEF4i47olcmRz8EUiTBOJ28Xk3Zv5U0hNNDPCye9N
lhFTXWXK3XpLw6DjX3aW21o5spPrYocjvhHOYGtwN+xz4Oto1QWe1chK+/BrBDzNbawFfQPfRsu+
V5jVSQttazcb/n5Qo5ewFjUFfAomv801dPN+Dj2yWl4mLAiAVs+ZNgtas4QwykkgBbUl6mcZdjDk
Mr55A1RD/yI2Eh77afn7W6A8aFYt3Uad0bUNAEuxwmZWyRQf4jE/6nKBDnw14GmWlTkEdbSefSN1
CyMeFoApM9+brJa/TeJVVH92K3YqEIwXcFC2LPdvGDqfAMw/kTf+XgeVTq4LAdmQc1YcbKKDJqo0
t4fioVmGriFcJmC1gKjIp9bls/if8vJQYTMOLbhbxP6+kumrnGy1T5GD6cvb74zHMWLAbZwo7lPR
flNfjwqgmAs0GDlR4giLQHqyJZLTxM7MZZ0KL3XAy/KpCmSrFX6gkZ62Na4u90rZS5xr9y1QVrnU
1xT4Y1fjDFvR9nyUmKzAYoXWm1Nl7q44ukhuQBWwziXBRGTh2GobyfXlL+YtzT/4V+5FXSxrAglQ
qNAW3YZazrX6o5amho85n78Y2B3Z8gl/v9bvktihdbcEmc5lw9KQGliOxqCPxvMpIjkJ7g8IlkgH
YZJpUCF0UA83rSb+T9M4UOhtnlNa5catzdb8cJA7StCokHCGrLBwbqdmxocr3YYvc4GtT5Q51wd4
Hd3fjT7b/eSTGUVq7+fR0licxyj20VdIDWXTR4rgS/ily8K32NACKjb+4QEKUITHCTMJoTkLIAx/
SD0A/aQVbRo5rvU+e45DtzPFtd+B5o5bdqxnZTDfvYVRIRpEMIT7CAzX4twb3y3eznW09U5ERKny
G/v9ibTeQxYLqPyESELZuF7Zc7uUuzCq6yzYAsEDCTYDMgn3skfDJ0hqh4xz86kKUmEXLP1UtD7R
/phVukdjFy4Uw4KlWKnWB/WFZPlABxFIl4/A8qn5wHJxuhwN4Xj0NOTz8R8wAzBb8foLek3+amJo
rdB0JF/+hlCFCOACPc3LEDz61C/q6tTufT1EnGTQETYUXEGwHwk8Fi9l/AfCZmoYfFCiD224dwS6
Mcr3PseJQUV56zhVaedEED6GRql2mVjE1/aC7BrTm9t7oJprE8v6oHi0tPgBF2ZwngH/SuSJTIA9
EqKpuoDHeQXatEQQg9lReMFonWCF3Ivf8JEEhay3GpGWA/06Hz7i6AC0dz+RwNNCTaABubUQFIjN
O1zi/g4+MOVNXf930IevZ3TCwvavgQYxT24yiCJyC9x9GwaBxkXM8o1bJJrwJVRioMY80ASAjgUl
aTV8KGCm2HzjI6RGdWQ6p1iPT2SRcXkiuHFcAZpxzXsmKInRbj80Zx1PYAjRRnFo4qkDVoZiT9fi
y0/2t7MtpWu6l/Y17sbxjvy5SZaRksPR4SXXfdbJ2oBynBpaDVfnR8807JvpnSN2uVGCB0X8S6C1
AX7F9D5aSf2gB+8VKNEiTz23sKPm8CFYyC8TzAn1UNlvtd6N7cxQfAA1ierXh8ZxNKrTkoSSj8cJ
k006M7ClCHIQ8s6w+UxTc4taUCOz47+D10gpsS7q4G1LqIFAcWXUiFTokiRAZBdRGzCoKHM4WNTK
l1k4v4D4vv6XoeKBta0pgdN0Zv4Es8cHWRNkLXZ6Wmc+NnTDlUGBy/06kfyjaXxkxR243Pj7pO4e
ZuYtXiZvDwL1uCI2lBMXrT0f+pTTweQf32Okxt1wFsR9zfIXhXjRLgCuQuYCrIqxYqWLnBYdtSye
56HpSdjOvzOSX170+AaAs2UPCwWe81eqLAZrt1Yk2XlECJe8eMT9wJ8E+fyxl40OyjYQE2qwhJ7g
USVUyfzkTRH9pCwLD2aiFJbGB6e02BzEhKXvyeraW6q/L5m+73vvAWaLS68XApvlqPc3xJvFZbNO
SnkzjmBBrjeZgXKs30rBk5+Y9jq+BSHxZK3XAxzAQmrPLr8xrceyUk2IZbV0M4tKx7PffQigo3N0
+TXsSf/jxVyjv7lLVuH4wb+86K5uWqnSH2q2wafulKhaL9uCrHgzKTS1G6zaXrvttHOyGtA636uO
VHsYL5HVJvg3sg24BXctomAWATS9ImWGlrqbZ+P1SIpoK03M6TeHGwD28o9V0BImIJsp5IIhqAFw
5X5txVCRUg8EAeihYkRfzB9ZsuMYFnyNVhnvpYwBMll9PFd9V7Xyza6FtltWYbuG/QnNf1rsKAPP
50VFepSczVRW9UAJQNkZssGGQURTnpqcmBLBf1wprjjcgU8td4obgSkEwFHwT94RRtDZopPJ6qk1
9+nefx2UzxaeMT7H5Tlkt4fdiHCMbBXahO9bhcZmG2fWVT5QmiDjTJRPbczNwkMPbD4nlt2RbYDR
tCjL3KNpCxnYdjIDdetLu56epj31/iivruddixwLxXDZNF+aoIbcw8MbZPosV3EXhnvTJGh0FgbS
jH8nXoEA39H7NtLPqA3UWquULMLCkWI5G5NWt+6yB41dkJS1dd7ig+tmlYLllYGhmgibPK5ftbh8
a8dRolPKqY4gMyVglZ2DWPw2IJJ9pagkUdeKEAiiTMNqsCipLBBE2wDZAeZT0f7O1y9fa4YawdLk
B5QT4XDAUypViCcJFBjKs9lyIq28MUfDDcRCvxU/qVKHOZ4S0x24VpIRw9dEe6MvFxIatdnywI9B
dFYMLTc+IF802ERuP9YW+ylNaMZwXaAXg4gAlUDfCJDV3IKXGKO95ZEdEDv+4p92iYUHZUhtc7AT
r2TuxhXI1okDkMJ75BHpdpkVvf4MiZ2/0nMa88Kgjl3HWrBvJIUw8gDHsx2UkVumJx5js2Dtll0Q
SbMFohYpCB/kOOtwNV3QGKKpyArj9rtV3ua3VI+fUbOH/s/yESFqRTlkPMLBpH1GNfcZYkukJuN2
FFCPvJWX/FAkh8l2+X46Um0GuiLVcK8hxLaAUg389zJFR+j3Z0jDk9KlyZZ1wKac4zHgDHUULDbJ
T+HOttTjNbZV0OTE2g5Psyu1EVhmHy0XmtmUhlFkGHl8t45Ma+KKOfdTIW3px18EMAQqx9KpeoXc
r3IPu9yxcfMs6LjJLxJhHGmoVykCjyRvSW1VU4IT+tLoSpAZtRiTSYC2rn0cX1BsVJi7toqwCsQ6
dhn7upadztf+mQYXraKdu8YZSYoDRAjXiNjCdwlfskKNj03K/UsqkbxN0tZsGPdF39mkwP3nuFfz
11MjhMutX3SDx/qFoKQkEbrolQPg9BLY37lI/ekMFTrpecqDStFsNm4sat3+dGPC/Nau6LshyaA+
JpFRlZuOzwGcIAX9Wx1rdHe0Ugk7BR9tbdG2PQqLRrclYdn2T2bpV9lscLMvdce8gFkwEfMDWGpJ
d03zi+zJbzVdS0QedsxsIIYyJi3VTBH9Z57F85vEq6DR4OPZm0YwrZaX/TTi3Iy7rJDZgOs8l1MS
RS19OGKjeV0GewtV4fEdC1D7QW0/HJ/Nhu64SXPGUVJMOsdrF2Xz4lxkjF8cJTx3kbD3rai7ZIuS
TuHoSpCroECqKUT7m+jJDGXNZkEsMVINXuOXJRax47XWqxYfoXUTvgZfacVqOAPmQ7pb6wEi7Qvu
7fB3JHK0ImWSwlaJGZzPAXykReq0Ip9AswsSwPN0WeXp8s+92TFcEmQXa3o0Uia3yFC0MqK+wp61
O0eLDrW4hqjp3f6WnwvHolfifVo1kQfYkx//wLBCaJ92qelMW7gYM8Lrjn5klraWRN2okIkkSXLa
MHgi83AJA04LcCVFlnJgzCVHbBlBYBinLYx0Vm+bI9ScocIXCqZYi9dQeJtFFAcwcbYaKJCSrXWn
yZVyOqueOrUswGpwpymme/tdanJEEM/v/MXnV/Oo9EMetazcLPbaSLsDDm3yh9cp1GQW3SXYajEx
1eD82INWYWmtmAVfqu4ZvdiczxbbALqfiEqsT2sHwmoXqgyRYmSq3xVxk+QCbefQ+6zGvTnIsg5u
C7kNwdxXgHeU3G3PjAFbeENbqdq9Ky7si9YDMjwQr1A4Yv6lO8WnpTGzp/KdN1JHqwjduFtDiNbH
SgxnCbuU/ly+pdgTJHNjCsH7mke05F3zOhEi6t4HHZ65lpvDS90pDN+UPyZUFxAE+Piu83hXqFFT
lmtNZfBxmg3g5BaJO8n7T3gJUrexeZSRy6phhuBuODrtgkqkZPUxRHpVaJaRdY733aWg9k2EBpVH
JBjZvOovYpakrJ5oUk2hazXBNF/WqyX8FfQkM1eHQtGX0vx2HSp7VkbhGIGGtXFKuJhR2/OxkXaP
IWwAyiExxQlQzMILaguD7qHtcJ8/X7SIc2+RE7wyU+Raq0aWP/xnLv+qcINz5DZzKJ40Qy5H7+aN
o6KB585t61mAYeZL2wdpYVqh3JND5hweYy7TR6K7dmjOAc3svoJ6tiGwV6Jpd+2nxlQ4XjM1SfOn
nzCdcbb73vaOkNQTjpGDPZIND5VhVhToorI8V7PAFsbeao+VziEOBddd3V8UtBVA4czHb2DnY9s/
QQ+DM7L2EJfmzYraJvNa4/QeEDUPj4j0Aof1DQ2jPVufUQu3ZAwliJ3JnM7vg4R5kuufnnf/UHbW
ATCuaWE+p19yCVV86kaY/5DNN6z+AF1rBGXRMfM5I2NX5gqEyVK6K5XpdAXXWaE81ahG/OIks4ib
7AKL6VbvQR+Tv73PzTbaz3PnERa8cXMBnRfXu7o78gZEz7sobizmBvZRQpbX+aHetUsFD14HvUuG
FUGMvfGttnm0jy0TPUU82sARVj/kr+EJYbOvswTnhlaePVN7ZPidfFxWgPjvIkQNrc+qC6mHsh7y
PGlWw6lVbEJXcOvk5rQuT8wmbsJ1oIdRtm7q0tDERTW2A0cKGXfmqTugxygL3VkH9xXcQLoYc/sW
2qHqV3aH9egHwMKePsU12j/2krs6FYEUbByAF8TgBxVCQsCeqws1bfFFFv38oWitHJb5Fs1ILKxX
/Lv+nOlOBmVQrKURwmc1KKmnINGaMoZ0L6hkNc9Hk0KdGDGcWxsjxCwTxqxTNtCCdX77HqwFqCMF
qg2yiMrFl0XMkObnu8xML9IO7Q9SzPI0qDlSzU7fJ1savDbOmC0mvIYgP/meAhE0v/lPx5wbqqVJ
Te4L5bN2Jz4cxcxWTZ/4U+EiteDGuoex9RKPDZZ5s++Xn0u9vOTnwh7sUGmxTtzTBb7AzB1C30b0
Xx/jgrmD8L8Yrl3HAfPLAt1YyDOevprXF5MaNWDqlKiN6lj1em+Ulg5bMtAvMcNCdSSBlq3007Ce
9SSIOrq5hH8KnWHgbk8A57SHw75ZEwChOxGFHsESIhK+SYLABvqJgpTFwrQcj7pyWSi6Uja+TbKw
1flnTwiaKLuh10apuvHFaD+3JphBY7PQIQX1XWdXZYGVGzbG5RrEYRlSyaSPjPYKDUnQrTWrWmVY
gUTuqID6Q9U/asyvsKDGRszIlm8tNkBWp9DU42VVOSvdx45DTBt+O1JUTUhXq0+U2vwgHOHQLqGP
46L6IvF38u8CBP0k4k/Lb1+UPnJCOWdnLOdLqEWAyYsxaaA0lhFq76tAQevqhXKHBSYoQGfkrqDF
SBFrXglg2ZK/8+rXB8ws/an4p/nJoV/OE3xHmKSNmnmi6coxrpQ9395sSJC++H+qPDB0m+5TSArQ
sJhHaiKy1oi+RKAGCFyDYy+NJaEEwOalJzZG2UlFt7Qvk/2jGr/RUlaKixYHTSrHTsJ+YY3FqjQa
kppO8C081psEsfK7dPtsNJyyW4WrZr748b06QFs1TkJelR6AJvNqjZbsO4imN7MIsbF8CRPJT533
IbSxbISelc6q97mL0PQA1/tjafdbdfXSHdOmXEU3ZHO9s9Baaih8JYzs1XHVD5bgzYdVHN2aAsAM
STwe2wHiBl00k4j0/YLKBHuoAiJmjrwfTMXsD05uqf0qbj6ry+mGIoqIrDag1L4vDzgFrGWrhdn7
AvwOh+Uks7ywqgcc/t6cGrbEof2Biff0AOABBH3wqnCHya4nz/pRZIiFk58pKW4yElQLR05YTlfw
1zdsa1O+hxwcEZV+pzXYodL6vRq8spFwbkQPqKM3lQMaKoj3hOtYZbMAGcCGVllHiksJ/VQhEZRc
Tgz2J0WfXnHsln/eB/6hkYAAJKa1mXkLmrDCGXjlwE/IyTtsTZMt4/QbDAo2GWFj6rtZkMjyQFq3
wQPWos7J7sLEQhlpyT047rOPXmISsN+OeDSdyThHbTvyWrH8z2at4PK8D/HyoFWoZ8GC5+5u6E25
NwMe6T9NWmYH5ogAXpNaAwlDY/wv7/FE4Ei+9k62Wfgox5zKfgUiYRsifTeNrdFNkJKrslKpgOig
CUq5g7eyeaUdpAdWdx3oT6kE6kFd561+30ShRpA8K0qP07oXYMkcuEKeypNK8LjN/ngkqqzc3Khl
8GPWDdRJ8CjmM87hVnVf0gkVO/KmWwDbNazx0P3r6RnCNXBs4zRk3D+invnfJ53Nw1M3eOb2Wnt3
UzIbcoq5kCl0oa8fqsSxKTjS0i/4Z8rb9gDoQ4gwwijtRzlEKJTP4mGL+iW6phd9Rb4hLd1kW+y3
i1AlSj86IB8P3lyQJJ6VPWznRb2FaP36s6OCdkNkuFcLJzEWu68ElK5WUtIK1oIGvWGieW65kW4p
qCwtVEAOnxke52tvoZ7XzhvQEG1i4VXwMkBQw8JkzJfJuKe2skDvc/VSLdf+q0QZS61NK8oyqLUf
xYqSsfhvs3AbRIaQiTI9dZ3wwU//dfSTXQo8YvCO/Q3NhnTdp5jFXIYPET8Qw0EPZLRFA1ILxtWS
HBjffC080gCNEZ+i2748eEyTZlH1DRWzaF3v1jEapwzbXxQaXBk61kecoPbeQUBrB4bbcfqYX1AD
SuGwRYEA89QjFCZC/Cwa+kY4NKpgqG7Uc0f055EpPwRF+k4Voze/FN59Tqb9r7ahhyRQJcDa7eik
iuQwfdvwxIxbXIvv9JQDV105+T9bNIEIS+idyBT8IG4DlBLdLYVg3wC6YRDH5zpBaB5DhTRSPzTV
wqBx7/HaTUxqmjzWQIvq9/34g1U6UcYk87CClTGTT5RNDNV/y/IaFX26yw68KwoaBK1vVxQ4dYM0
k+Q001RF/pq2UkRuk0NDVF4zGzNL297/oWWfTcdnezx/in/JHIJdvWTxSP8EkBQwypbtDukHofzN
RzirjMh6TEyN4JGt/EREvoZxvYF4Y8O5kN4mOH7tbT5eBozbFY4pL6WJGtF5sGT+ZLhd2MIgUhFA
QOq4js3B6ts/fUCZ8VD6nWPiVCOh5rD44rFMqEcR3Tj3fsODPki70XawDayqV0btF7ryfiskphAV
Oi7cs0BlSI2Kt0CGTNSPkWUm00xhPLApDAoXZooyRjxn1ywBGmfFmhb+WFij62oWE9/7C0NgsUe6
MsF0tflDNjBv9JdNHZWGIqGJqq4ErdY0Br62l/YtGLmuhAgkJy3oYJaSWcTfQ0THMEWCpsD9JhWN
Xk8QEY9UPF6GKcxENeTBx/IaVhWJTgXvQxGrTxEspRK2AZNCNIhGggwhD/EGVxn83AafKH8L4O3c
szBiIpzlBoVpUUyIl2BImW4TK+CBdI4YcBfplAU4gl8Qs9ZkUS9n9tEg7qCgdNLUOMJMFFmJZIx+
oKHUjEGpspMR/T4Yp+uA9pEoVZELVHq4L0f6+7QyZWPkQqEmqX0pEUMTK2SHDM3TZlG5IxvbryKt
mddJoZQlo91omIyLdxoO1yI+7BcN2KEuPYMTkmPtrM2wzIu27ODZO2QeYeq5316JQQBK2ebw6eyK
DgYwpZOlAxoSpU+RoLcok8NffqDfafXTxX2itYBA3IYvflFSeW41u9HqTJwl6+l1TXQ83m0W5Mcn
YRElzGRzdK5430riYA7f2lRhEN8ckaSad9T2b4f/AfKV/SLdC3Ll8v6loOsJ2pb9ZaVwQ6XJJm6a
zTga6eJJa/71Bc+YTiogjp/RcU2kUDEt9XeBJsc2K1sCfWiJNAJtO2LCiDNBmWJMU+1oE6CRpTNy
RYmHo8TFS7J6PmO4ilhGIFVy50poNbRxHhz09q98Fd5gikX3dWGDAWfj0niZU83hr+vQamwcKvcc
b4lAPVTu7lB3eZajr6yT1LpM4elNnocKEbAOb7FOfiWOAS9Db2uiNuylKJEvWI1h6JbSpRF10pGL
ulbPMKlrF9xNS57RZIYP/z/BFCOX5AFaaCPjGhbYcrV5VOUy9WPLmJEqBOICEBi2DP3+Vlnjs9SD
TZq59ohdNkuUBHfZGC2kkwgMEegIKx+55sDLNIBOTbNU1h01rp6KRhi8ZZ7O5Ak2JO0wskEvl8oN
Ae6Zd8SN0E4zsBobsUw0hlOXzswNX5UBb5VPxwtuPtEh2Rca1z50I8ylcLUBHA7QyVq/ud8NbFpp
Y0Ydqyznkmu7bkDHnu95VV3h/Y/P6Bailazr9xUmiRtwpUDMhLRYLYz1bahaTN/doeG17Ci81jz/
wuB05b4ru/pSfOEhabl+D0CF4AIsd84kRPwgyqoZnD2BW5SM52oTpK8n4DW/hfei9hqdad7helwJ
GIi0qxqVEBG2oWN9MY/cjuru/GjSpEpa1INOkep4S3IUrSMZ4J7X/Y9vE1OUn6WyzepUTTFsj5es
3cIX98NrNHfQ87FEK893/RIsj5HAPFIuLe7DSeXmx/6uzuWqCweJmMNklYJnlQlbols4rLUsoUvv
wbtuiFAF5zevnP8yfayDgElabaU/XPXVDugV6/MLz1gNfC96waLdJDTbUQo7bhaTLBvlObtwZY3d
BbvPwBiXVyJyMOa/ArP8K5d62Pmv8A+IOanlWyTPQvRAH2v13i9wetsu/YdrhatAQMRXvFIJRSAh
FlDiOfLWvy17pJjIRU7PVSeckT5rHvdzzzB1k93pKwskpi2WeaGA8u7t+ExivbLH/i5Uls5mBl0s
KrBJf/hSqvO44XtVHAWrjQ9D6XipmAOnEnbnEZpEHZY1E0rEtYgwd3N+Y9ecd6cUUZTpQ10tXljK
3NBD1oa2E6V+itdxqs/bbbEp7ZkPp6zblFpxpzsVXvUlv5PeL7WxfR0O8KV5rINqOZWYMouIVpPK
4A68tSAlIjyxNJIU3hdjqfuwath/RwWsyiNBQnTw7eEqzTS33Fea785E6cUm9BzCPvNtq0UTqD7S
Nxc2fjXirumtdIQfz2XiVje6rIjLBlzshgb7isG6PMlDh512eZHvJmE7KhAhb9CgvQkv/QK/NmwA
W8DYPfiFkKf38gbp8O6llwOEjStlnSvSh3vH8lDMebAuUQiIiFAIx3ZwS2FrED4IiqtM/7BdMz3L
GXKQx3RP0kr5TUs3RA1nYV6xrN60EKNa3a47OLjsLB0QvY/IA2sHdBG7dVnKnR6S2XImauB2q40G
+UXeZuwKkNNbFvhlwMCHlXnazuhFByGvdc+/9juCkhl6TVTbj55JhMCzIzZWNxpVQI3QiLWQ4sC+
F3Jno58qAYULc6twuqGAsawlD9+5VvnZwZPW6J/t09m0QlheMvsdjGwSl1gu81Viw3u62M37polz
X2knsb5WOuMJiuuhoTWRnbsxNqaFANXv63Hm1RCShS5zMh4D0tzaLfAo3YA1mKkumQ6UiBB8VNvF
+7QeZbHfsIOi5dkvOX+yzLTfwmYFCM4pYPaM40YJMG8F2C3fyUCrDLX02RSmNXL6bm9ZV6bZLBmh
y26KG2SHmxTbFaN0p3dXt8/tqi7o6/+rFB6vfgVmnOXWOrrTyRtMXX7XwhaxTP8vumbXoKyQTJIs
BSh+q0NgKXuDnNCU6VEmtbTruhW1OZr5LmCguopMah5CEg4xXZacCSKop8hLoToiSRunSzOiYvWi
6g13zbHZqW75qYQu3fD0GWpj9FElVSs+X/Fxi6B0/VhCN/lUoSHA0gAixK2A/gIf6cZr/x+6PPu0
7Ljfp6yKNIalVAenowYdY0PnaJ9Dq1hhz2+ET9PMzE5JvuaSoZqcXW1nwruM4Ss8rEahbTGz8+89
c+kAWrZNHz29qQk0YpqnzSn1sSrk+js4fPkWm2h8dmIVy5CkCQXhZgrOw2Hbw5II7oT5MNCCVHEl
OM5ORp5xwvG5FSrUjUMwdLVoPsM8R0egIOVoPnwpOh5AGXVHDkn3Biflj567oAMSZFwk3ZihMZpJ
xrZyD5sVNsSkmMEstzbZ5V+uuYAZGyZazkNI3YVzEpGE4fv8HJW3QpTeA8eKykugTXNS4PcqaCFk
kZuqkHkwn+wFBg0PGZODQz5SvpL96CLV7dueeE0Pv5Vd6NEOIGFUW7sImh1m2qIFYqYBe6/AYzjE
pD59/+j5BSRFPqeGhVHOhS+xZn2jeQfFtpcwnTIlhkDoBEfCAtfU7qpVM1YI49OwDWhjTdqrFadO
ztavzKYsEadk6rdZM9jpu+YBNYUXFEy4f2AQfjmEG022wh1AZrMRtQYaEhmj2y9kFjvgyhEdAWnA
+9VNhKgvBUu7zsG/19LtKQA2XqPVcpV0C912vNTboEGj2VppLZReGtgYRDFafh8KDFgjk7vFWiyG
73z8TPuepV85HrwKprvfY74DYp4MKNmWJk0pDaHUj7pkSHMUICgBiyq+yfY0KMx8ba0IK+axeHlv
zxYYla0+yAdTCA0e42KuiPfptoS+QmPVIqUNTifHQhLjTagCiQdVoWDq19Uk3rXQAx7BGhKUo2Nj
Ahu8u0pfLlvRbVtPKjY1Kh8yOswjIUp4/OrrvV6lMt1x/KmZ1K+yyIZvjEuGT1iae8aioxkd40Mu
mRFURKEUaWluy7BdAcL4LrsMF3xWNpjWONedkKSsmjW90MXVDTcyoM60xN+U8lBj8XMgSkswTiTB
/PpXsCZ4OJ+cpJJPPiKa1vjKW3nk9BO8VgcJvPAXnLHHyr6bsxAJ6WUKMSfmVKl9m/Tc6Kgskk+i
BqwFDXRi+b9hhYuJbhCKtGqC7E2Cma3wbDnrwY24p87DslkVOcNAoaiJyXnoaL5d3XsSlrnxv9tY
CeGcUXwFlRwgyqr2wLNjijqjW1BvRHwhMLk0zGX4fGmhRxDVzzeisnt+0uMY/HiMysznbZ/mJrv0
F/ADXRss3YSILzQzdljmyP8hj+pAXSPo+pkEiYtA244DHEa2VdbL+3WIB5WBrVUCsHKeOCF9bZ/a
5Dj59gybriIVhcg4APBZ1PDiEjTKV1kaZbwAYwokDsjHWlMKQlwPoCQF8gIEYNibM9Xtmp5g1LUN
nmkmJuARJeM5sXvqp4FXhP9JUtjez+4x4xUW3S9lFcPDZab/RGKkW+n3rR048uoiBGDYxNVId2Pd
QADhWHXdBtfiftJO2lfeZDCj52ql9GKLGhesgDvyDgmQ8hUBcrEhEUNxcBrmPsiPIXZzLdInHt8m
6K7ag87oWo3IhHKncUbg2sTZxfIO47tSSYENnYsKdBt6VLQ25c0q1GG2wiiPL0Jc3TyJZVRfnu6o
IL6LCHxEUyRGGTI05TFJSaCgjRkREvsMWb92pqwKS7GIKWTayaOVNCjOwPl9HLbEkwJ1vQ24xI1e
RFQ4i/4JpZOI9mI9lhRlIxPuaR2zfoLmtv5qpG2Ui8iTrUXnjJ+lQEZaPRHqXkcM2dm8XWUv4y+x
y6XteNS+WVkNtM6XhnS8nYMs7u+plumGMOtBEHsjSC5+qTy8w+z4bAGFTEr2s+2cJiRxtOvOZZyP
SsYoCfG/n3D3hqUWz2JXbh+/H9EkdZrPU83CgekgW6ikJ2LedyZz5xExQFIuDUZ6/NRKu0VvoCih
gDvpSYWkYhY7VGRrfvxBqUJY+SDa5VrYQJjLLFKG25P/qgQx6McZU/h8xzaOx4OReFr6DuRMTSxV
c+H6IwCvietaCmQl4uP3PgMysKCsn2qLcxX/+q0GvAzD1yTu4TlxJsst6QZqnj3iGhBHapptOO6R
ALhlxBlPcV0HudPXv7+QjYfDN37H7B7XkJZTyzfQNhp6XYOBH4vjC4xe1SOKd0pkawjLUwj3KyUR
o6R5JV+Rt8RPQSWI+aqPtdx5eHuMlukJOVin1o+nqVZAaXsy6ha8zbq25IVWwgLFYViKooSORHIB
yfjntmI5yTTpofWo5ObpwA+07kPnySMDUJz+r/1od5wNn8CUbEE4qBU1L09rABDhelKvAr8VBuhD
fqbblTf2bwbn0HUBaqrAFFvq9iqIqIGTUe73Qa4mkjk6qJeVOgANUz3sXeZCyPpZLfZVE1yrrVxH
Vmz1I8EtUFl/TZSZz2I1z2Yijc+oPs5b5H6BnMTKDA0YX9i/iGOF7rX24xT/U31KpAp1wYazNKW9
5ELe9onnUAyqD8+mDPUDdB/bGj2mqGcpEuAbAcx4cWFmdrVNuIEVghRsyLZ2r/y3sY79teFBZbku
eWyY9clZSMAmW1F6aD7kBm7b243Yuy4NV9aBJ1JPSQSBJ0kyOVLL99614q0bg18tXw6DiHYsk8B4
j4AJeZxUZfcstd4n2hn5Bn2KeBOf2mkDvukLQAU0z8Nm8nrjX3tt+YzqSBrrDnlmr7RIVarFAr1p
1CPAXRSWSOjt5ExeYksqu3ZtvjKrQKOC9h32i1WlLrqeoGRF3sQMzcjUZP5GYiVD6aWar8QjB+Uj
qExUuSsJ+Bx1G+P/HiTDLGATHw2SxUSNpU8T1o80oS8n50hM9IFHwwFkssFwIZCd1PR3oYO4Vv4e
oFFr4JWsBObHDItWINJYRDjVGb41UoJcoes+ZJtsZNRRKdty0XjQDeGTfIMMF36a5KcIqqp8gD5m
Xj/Gsy6Oe+42p1F4tWiadRaTeYrGZXFMiQK31bj2AuiueMml3L4bdL7EjIUG6c6GRkOMFdb2oPBO
s2BqOhBZmkzdrGD8ijtK+VBKTf+mgBiTu23/tycE4V42CVJRuCx55W9GkALM4qYinzKsSd2wvF+A
/xFcgteLWPMBqU1RKI50pPvS9Nk1HhPjC91huOtD+os/coFuPsdBocGUbW266znzSIT8+ovx+TH3
NQa3mfvTi7wI/XzTranXjT0KSfTeLWUSmkARYcVV88cYexeZkYeYNrflcoH2mKiFBHD7LpHRhmdK
GXpbiHZuD/5JBpmxCttU52xFSIxeHui3HJHWLNKCfi1vLChHyhxnx7YVgUBAch36vowNNZFlXYEt
ay9MwtuLIAWNl+WeIgN9uWX/g+99Y/s2i42tkO2mHyjreoccjaHA/t7CdOe6pBoake8paUgtQRqp
Z7ejF2LB1J+rlCO7Wo08zMwMyuaxh5ThEgYo7n+a5BvJhfklP6evJpuScL8JlkGDmCdeSpiRbrMh
7gwJVk9egYKFo4Kw1aHZKCDYvR9W+nQLxDjHCFn/LPGPY85pgQPl9AKL7AgypxWeoV+WPrS3HLZT
lIZr9nVQ3JYnKAqZswMFmujrWQApOSxympmJZelz9nIVkQp2lLH8YByNfFMnKmcUE8XsRhID8crl
pgnf1OO75AFLm1X/YDquwj6dfGRgZLudHZlBdrDD6nDy98289WzXrOFzWIKJDDY31sHMkAici010
Prf0+VBH7ukqRQkR3IQvvMpl333Wug7VwEH6EdG904dDIO6KVePusKS1fSrn1VBhb0cSneu6qvTg
V1K2yBswsJ5huM2Bq7Rt4guuOfhWzf2UM0/Yc45vd8QxGVv97mKcaDUjIdfkhlEUVw6V6L2mu++H
5z0QUK2p04VzLSVEq85Y7OC0a+B+RedReIG5wexJW0hdl42tv0+JPAAObhNZ2gBYSr+f2a/58XC9
1EgAvsZ4K8ck8C8FbC9BchJ5YiquyNU/l5eIzQCaaq5NnKgY4O5divuNaWNMdSKz2arUCl8VDzBc
ukKk88uuYpOjcvXtK9dOdpmFPZOURMuGqaux+DG1zrAj1bzbQ0zisXQsBnkEcxg6ZDeWfQFnZvxY
Q47TjPQSOdC6Xc1Pe3jOUvRPE+vMruRalnBxFfG+V/8/+ihV1gFwWzMLcYf4EaCAS8o50IJS8yNs
cul9gjs/VVFvhfa8Jxh3+Bp6mwEUDQ2awF75hxSH8OrZHOvHfpMHhUZLYvGJKKVUttk8DSjGyth0
S8s2yY8K4LAqr0jgcGBCl62Lbda5pcAGrH2dUVx6JZxkilZ4uW8ubxmKIHLHWU9+l8e3Fx0TKBOX
0kIV/D/ygmC3E+j3Yqzs/mywYA0I8lLTBJZkD19A8z4Uey9/dNzdYkGC5DG71A5vgrMvPNZLy9xh
1RSu3bQihjJju5U0FhfuFjbEaDEyWp+w+hsMLKKuRwkO/J9VD5a+K1/3XlOjbRphVLZ52eC0MiDL
pLknWeWboZ/F7YwJ1upP1E//Jt0aWtraNLxbte/05HaYk34Nmt3htn9TfDwdnfGCZ1Y0Rz2TlZQO
HgM9tKPojWtS3wGi8s/+nazYekt8Plcwd45EQL0bC0M2EnWcLaFn977mh19sXbLqFwrwY3xEtXVO
UE3rEFJOUObhU7j0nN99S4JVMR1VPBUd2Za2jnmZ51hqefLMwGRpszmtHtiJ3M+h2B2gIG4v5Puz
uyOQhuRfPUtOCGbEXoLaKE3AXbuTl5OrKCUWoMP5I1Hnl/n/U8WYviBHvuhHyqZXYfSGgFZx6gB6
ACKTlAasrk8gcMa7VT+C4Tk1a/kwBRvZPnPpOj/pGkXChiPQIF8LTXmcE3i4YfVYElc8I+RiaFU3
A2bONFIu3WcXXbZtDEz4ivrLKrWJdRCHUj3DXn+3ldnjjEPevJfbeAKPj1jbgjCpAqD9Yi2EnVaD
wql0sbJrTQH9g1L0hYJWiLnoD/fKduVooT5oPmuuvI41znEIwxgmKFoC9riRaX22lnF6Vr1yIc9u
oy4L9STtcdvFJEo7O8sXHfao4OmrSH3DLagqX/+PmbOYOPJUK2rjGqn+rxSy9A4RlsTFzzYl7Gx9
gd6elV3HUYFZ6k2OTaPKAG7wDs/ZBn0aV9hg8lMtMkUtMj577Y026AvJTRFnjltofj/2m6fNu88R
HirpuIb7RlP1GWwW0UubXPi0ozmBKyQRj6dDEBpOhjEI+shMMPMUKUHFvSL/M4pbk+X6PEJSk610
owvwgtYQF9AvAW1Uqqy++Kl+9QHVKZM6IQ6DyUC1D8B+dr/HWyhLN6JVQoCt7RgRATc4BpRo0xMt
BdqeQxJZgt6x6T7fgEbtYMzIVEDkgYQSFZgqoW5+c/AAZdQZkst4sExmHav5J6Aq+yStUcVG9g3p
TWSRmWJ7BXgmAFx1S1xJCeqbsxxZ5n/SVE8M0SNy3ODEm+ynjiKixaW0vHLPqNQWQojuQtquNuJ+
4heZRDknS6scHZZcXd+RYR3jFxncVlDv6KOyQGDFiFi6lPzqvIck7oZdcuJKYgmXQAdA6GK1EMZ7
jL3lsofDwRCQD5+rtLZlyR8mbD9TjwNHy9qBzfEtBPqY7gzdfYTqD5jGnfSM+QGGAnAWd/sXY8BK
RI7wK6lHmoaSTR95RjC8Fqs4FK1emyom/x6LrfThg/QNudz+oDkUta67p2DwPWj2oTTanA6kFA9V
IRfJg/DaKJPRu9xD4yluXlFzke98PLgh4liWQCbtQ607N8ORkhnRydz3EMr3k9kOlbHaXuCiE+4l
kvHXkpiksDgX8cJO5QIZNICGAdatih0kjfMusSdRTVUyAgz1FHKVJ9NgqjTmsE4ZEMoYyPnXfxTk
tyCdJhlOJ0EPRRDZ5O6J90oPkqbfbGvdTIPh6vEX2WNr4JSyFHEva0Wa0Y0u9KzHStHbUWPBXZ7v
aAVCwrUCsBNKHusCQIb0bjYtQT0HwzrUj4KUEacTtH2D108L3HvKlzqPEkEzZohumWlr9m3BncPK
DEjzmnoaxXu5hWsMV4fgEDEOGYdP+fF0j6DOpi2y6H9wjzQvEqVYSd1tHKOD5UAxqjNHlLMbb8eg
oVd/dZfE6mUYcDKH7t57jGuEHGlKPJwnZxvR6ZsFt8weNfbXAcqOiGZFoqZv2y54b8Hzl+LF96ID
tY2oNfeMfre0n8RzLYXA52hoKhgBzs5ELy/nQHA4h3NDhXLa14Wvw55AiXV3jvpXy0XM7SInt2J9
oFABsMXlRNLJV+92YzWn874FXe8Q3a+hR2QrnZ4u78VHXXYKxBw7ahsbOeIbHbi+AGW4dQ7JX/L8
18BYrkEyyt0wtjmkalD3Je7MwqklT4XbSYi/BeM8CB33eJ+MnqGP+E1nR4Yza10J/R/5bUYz0LXO
TWtpQZXPrFsrSuudKA0hQWdhstaHWtm7cvHZ3QUOB4AN6wVZnY0CYZ8FRwG39w2pvE6BUTkcgyyn
UMs7NT18FFYvlO7BUFFZtXqY+AG5joT35u1OGyTc5wrSbX9Y0iMxG04a0CYMBIlvUK68Cw2ccU/A
eqob8vL4xoReEudIj/Adm30uThSusCN1jad4tK5thYqSzoRSBhvLgnuUQDnJYslAAMjAgzszzAUh
iGyJxFCc2lHsK+hNKpE64sa37PUqfmJLu/ckH19rDcwjAuP/9I7Fg60IcQqfJnERvPZlhZQdNacY
z455YohMusIaeZzxdLxX29Ym8+bV4gBF3nHTMa7+YG3OYF/p6cbe45fzga4SUd1mAV/VO9ds10Va
Vsj2d/gROm6wHverjSFKG2SoNRj4oAKbfs34ep346K9V6pscIufhACrMPutsrQSC2171EMf9WyHr
YxLfAaF7xkl9N9U2pRegmjUUXzbgXLkUwP0Z/5w442eVmtXgk5ISWccWMAzMlBUeH2xl5HhvSV/p
ZuJ8kvHaRZRj2mX+YSrVVKHrbahjbeF3Ck4sd1Tju5qq48zJdaz8NIiT1hGMiY4jaec5nZiJ9egJ
/Gf+RwApj1KFLe0dglqf/Rcewii5DPLeFr1/D5BR+xjEZWwmEwTHj9Vy7BXyPKN5do9CfzcUtjWS
XaduI8iIXW7J7N0GTwEe5N83MI7mq08ORMylla/nZ8X/hGRsVOTwvQS1ENiE6L/QkcwPzCqAxBQq
pv7RUpDL8dv5J8z1Zn8Jtx7+dCKrzUQQHOIPFVWiwYkXvu5umgg3CLxlMB4a8QdvcvxIw622HSLd
6QWrNSNXIXflxOzapr90naIM61W7BT3jOKeovy+tn9Q61zFm21gS5ZmkXrJe+RTIaX1QaD1lrSE4
c/Z5wX0GlLpluBRSyMEnDvYwdzmog5+iZcn+foXl/RoZ7G4BzAEa/H1ytQu7yhY2zLvEVj8zv2gc
ejc66OMtQS30il4Rd4F+p9NLI0YHbPNfDapfP5ZwkKP419BGdgLNvoptOyda47TrA5pYuB3YaLze
CSUjPS97dyvaFZSbgJ7Pb7iiW2Q9xxoU4md6X9S/hh4U/S/IVMG2ZHapyN0Y6pxHNOPrVPfUYFtQ
uccXYZvdCcMGWGneeXAUHw5KV5mg8jssipELZ8E/faxpYKxEUZMJHuRO+ne5R5jHz9tJC0YieWiA
mb3Iqn1slFYX90SICHiaB5F3X3q0K0vvw205Ud0rU1YIc4XWjk1Co7h2xbR27+3o6dYtut36d0pP
kOYWDPngfnkYE5eudeRFXZSohVlFZMYsAi9CL7IC0VfwcyP0aj203vmW919n2G607puE5MOAxHV0
xnxy6F/Dp0zP9sYqa7C49fMQ7bNXNvmR0Q7t8657xloK7kqYYF1c8BXhMaWC5XRFG8MpXtPe9vmY
Gqp/VOZJHoVwIh2nXnm4DAoMyyVWCmjy1Xv1YPTgMBYeLtx5vCxZhNQF+Q6T+jooMr2pasmFMfag
NChCOfDW4lFCB00HtYe97JEI5uqoODJjQTffyGrtYe8X+4sN8jaxMjwhzzFu//czWgV7RvpECzeH
lY6OZeWw7wwzCInES6G4nH337MDKHXBWloU3HTUSVsO9VPKI9GpKj6wd4UdFQ0Aba7RV5lNGtFIE
A8fqoHyRPbyUaTZpk6/HxCk5iPk4AXLuRvG6tkVSAiwS5MwLp/tOJ4xiDGaQOxh0eaAskKX8FQeG
QfKS+88PGMAWaQA25y4NXWPA9YhX4MMk21hlIggMZ4+x8Ug4xqlriy103xE/ns5ANsMseRlf4LX+
MB7i6vC0MgnoaClYBTPgZDnAwnYuSO/PY4ezkTvLhqU/HD85GFznxUVwrc86iAisXBa8eFOmb5z8
AqhZYcE9m4eUj+jTCDsSZZWGMn7jMwJn4+0zCEKMbNkGP+4RxlICvx7vvoSlBi33ua3bRaAm33C6
Ro7Aq6Dvtt7GYmT3GBtoThi/rNaWoXxTAh2d2pGaHSEoUI/bdjiS6/myoeglhxAO2eNQ1YRkHDmw
pQSBt5ZCRRROh3jm+Dj8+d+GxAxNATVvpKIUVItQQM+6kXjMiMjoSdTAe5Z6XuG0bFWovfSos0Tn
zmhAuRwXYhlODbG1ZQOItWqutMiU/FHCXf8cSlsTUvjubba7tBFeDFKTwhtnc0HziAybFNBjc5dB
LW1Rx3EPo8ijdYARPB8Vpk/qTs2W7tUorvjiz3QRiKrW0MuHlw69jVmlPRaVF/K1SJmmSTwmeMvS
TQ2IxDNJfeXD0ibbUIKnOfNICKhmS6NNEpPqwi9U0whf6UG/pnFq9Mdw72FsQAlo4j95Mr42Yixy
VtuDgWRajN0Ud5KonMTCz6iYiumKnj7Mi5DF0hO6s6ksYYGXRRYwHbkMpu2oY1At+6td9sb/GBq1
sTEJyLqWwCQHhkUdrGmXQbYvFhNGnO533ChjbUk+iMk9biyIrWFtrh7qRnRw2TpTDM8wlG15rdBR
DO5AlVAQdySNOoqC8GUlbdBJHCSc7GfUX3TJO432bQYpgp04XhZys1r90s1poCTKJjCadHCBSQlf
VpQKJ5iuAoWLULEjj5+dWBvavkRqGBdcystgGdKtxTjXHWesDnMAwNxVK8+sv65Do7Yq+iRJA1Fu
bhpP4UTr3k7F73UrSxIxLWScKVNCIAgo9gdM78+boEsEtFEVyQCUMroi2v+AIB2NC9wjX/leVRTg
fv6sLQZRmO+qP+80g2o+ShzA9YUAbxmNiD3TLz+7DbfA0LCuJ76PqXPM4BM9j/ytKZzeIFHbepzP
zbVwjsWnAFCw/87ahn9Jqdoal9+jSCBoUpecw6dWIiXgATz9dJhdBMGCS7iSjFybEhIwfyq4cDo9
Ezow0FUL48TSvbEBnMFNutDSwx2kBOnVgGVLGPiUSnnx8LASyqf2cKKNGpSkg1ZRJFIHvu5BlGXg
/31mWwN/PrVUTbooZPE2Ll037sKLo9gqxFu6vyOoYMCafmYesesWp7smxwP0ce0BdNngoDQdbjmu
FDYZuMwQUNVCRjhRxTXkjP7GlD8bu6xth1bJihnDeDEgDyBbulw+0GlWhfDJVhyiVZOjKGSgNtcG
KhTgrfB9RvixLZ+eeIoGyFp08mn7lOgGiVYh8V0PzFIwj+WvADoMkNopVGmF1qDy7kdxTadK3sex
Mdi/tPGB1UB96p2cBisFDzsoubvt29ILig/CF1jLEuhIVefmrBnVqR2O6OXM37mmk916DTsY7Fws
i2GT1q8YumtrpyoJpHoxD6XR2fDKj569gQBr+ClyMRKZpuF1nUI3YkpFwov6tU5JbncO8msgo3vW
j8kyGV62cZN5E5WMURRURApYZQOjNkta80fGjTkkegfXwRBVY/nfzhOHArlzf8n+95enmVCK6MnG
7VfasNdV5ghFA7zF3x4dYvSidb9HSQDWMathxdGyVuiZ65ESlbkIFL8xRtBfTh7NddPAhgOuNp/F
XnCrw67SYQPCZQBOdIIs7a4C7pjDp6tUuFg91uMl5gC/+Z9L+ceAedjkash24+/KEStn7V75oyre
NXkdHIkhooX9M4XTMupNA96lxNHJw5rkzEHj/kHLkI/wmGm1s/7NWtpvcTU37Q7NuMAVGFGuJz2w
1Sg3TB5PiSk2iUr8QWZzV7843h9LmmyItcTt/DZgY0THNv0BTvtnxgBof0AcmiB/J6cTPGoJsMeM
6ekp42iUSEejDq2wewC1j7o4eFzf/naGld9Am2SuBEN8WkMi+iKZOwBgr2emz1m+QqoP2zNd9p2q
zeBAMeEybWmK/PWYjValW7oJro2/wj0wF0rakJma3F1ukWZYePh1espsZcNSrSmnnvBAgvwdOGfU
SvxkdhVtsRv2MVGDR4wJ9baBvsbkZAVNGWRNzYEXwfMZMW8N9vvZX66ul9cIYrFmHRUbYHF2QfW4
LydSlFV9j5RsIYKS4XwlFrkC8lxzPv4Xz7J0B/Y3p2kbLGEKjtxI/+6BPmiI1cR6+UrYO20+XxUj
tfJdQ4ZUsmf5ixYJ9INbGYKNhRw2DsPq+T07cJ2M5qNjzRAjp1Sk9yb5AohJqMBANPoKPvsR2AMp
o+hbKC6xa1uTfYLvBNaci6TJ8vO/cZ7FvvGLBLbU9oyqAG2blxvht+Piv3imht0uzBLI8yrGJA2q
5wJcVkNExm6JXtiggNJf/jiEy0fBNoz7G+oGVTYuzFhtp8SwKtIPMD0TWC9m1xQvwzVMIOd07v1L
XrIqr/ssNRoXt1JMXeK2pDmBHmLpKb+279rOS0PodZtZPCvSWTLVZTjCCYRybFawQJui7qYTEaa/
Tdcoga5FSbe1Y70UIYYsFbbz1wq+6S0DN34Cg+PFvG4drk5DtOaFZPq/e/Pw/wAT2yFKYP1LH09W
jHl2+goGU2eBLcKhahp6JSoLZNFJApHqr2CSXZbIsrzLOUyrnbMcrYxRiM9N2+37ZRwcaOwwJ6Cc
MPnop1OStOVRlhsSno8UdrKAgY/3ViiwN75ZcA+PP1xQAhYc6BOd7fzq+nF7fgXTE5LhyqHj1/qU
0ibLy3cN25LUL/nTTMPjv/EmnAQaNrvHDKfsaod8tgJYM1P2II8xFSdeVlSMqeguTi8+9SvAI+7D
mTkXAZAB0q4GlWvL0ArgCmXjGkbUqfcX1RjMnI5FX5TW3qvIfJvctFmhda0quBwvyFrwopEubnJ4
4z9t/n7aSD5peXUa6WS5PG/BKNfW8sXoRV0iU3kk6uNlsQa2DDaiKMr5ibnsfPVLn6HUQvTweTXG
CHUleLczhFZrEBouvz0qEIN0llkN0f0Hf0iI+LRD8sjCK1vjmkBKN36lAHhXWCAvs6obpemyp4Vf
ASwfSnyvbkcnSQN1XLm9BoTYvZDd+a/bKq4Za/dDdF9ZXpSWC/f6JmPWsbakMAYcF991UASe5SmW
STe9L4Ky/KCDpc8+CQrgnjZPcHsxGZRcWlrnYDH0GjXCMJ5PaXei0G0dipcvxy1nzBmfMzXvlq1v
OWvkb3T25wpUji1GFgddW9F9j9kGT/sTtzdg8NMlO21HVUWnsu4xb+JaDRC89VsN9ntPTC1zSZgg
J7QCyTD3DP7byaE0tlSzHiqT2TebwFQg1dU5AuZ4U1zgzpSOwU4NKHROsQcwpGum9IDzjD1Qhtam
EtRrthJMYU711/ysN+RB9LiCu24o0UjRRpgKgE6oBod0NoYWF+ScXkPnz+2lnAwbHfwtzeaCXe9w
Y+GiYXJn4KVmAyXNM6jopRIeaPVJ9vgzjwnERVYNS1cHZ+4emHn2Xv0mEgQ2cguoPmk6UJ0zBr1F
ljiUmiAE38E5noJ3LltL9fV0+hmWulJwfxkiEWjmiuWooUE1X0bpAbTns2gg1hezxYn60994Dcgk
7wIQtn+UuMkERz0mFPM1RHqya2LJQjG3S6A+CpIb3Ky+MiWiWAEvEcfVG9u93OXgVVNCZ2VLidgC
BwkgE0GeiTM7mimE0m0ql6vPKcE7GSIyHJU6cAskc336M06GjdreHcQLJqNCBV3qZa/hAyd5o6Om
nEQtdESXstGIT9KbF3HseKdWBqzPBvQSGbxolOtyn8HujVsA8uDIDxdTr3atwHV5mr8McApkvP0h
x/sFEhjgAh4rhSrm+x07/aNBmgA+5Fsle10fYUw02dlSr/skeLBplZrQlQzPcLoqqFu33t3Ini9x
4SxkacoG5pM5gLTanKyzFqyQJWJR11UH5M2xx15ETc4tTwPXk1xuMvesKupKDd31cUw0f5yYE1XF
dUtpKV80YwRRT/yKrajqlSYCG7BRBRTakoVvKHBqOmVbdxTl4BD21dcKD0LZFBVuLI1m7mfQItZ+
vTJZj7IH8syEVfVmhbCWPsYErWk155+1C6mAwMZUPn03Dx3SaVYyPc++6mNEsjbYoileOt4H8VaC
FHa3J9rqpxoFgw4FsxH+IMNyTu8aVbiFvXXFgTmT7ykiTNFkNUhu6eWY5r/DQaH0qSlJn49TMFuV
+WpTPrqoNuEhFNT9SKFVLr04qw5Mu8E7EzTfCSbDEuFeH9JeUxnffaxqtEVGmzmMGMlr7J7K3WBp
wBcod3a+fgoYmU8afYg9z9+tXIG7QUe5kkL50iRUFb0QTON7wEaMi1xi+XAWeStgzU0dwCZ+ihFS
JY6Mb45WDQcuJSq2zzXJO6hb82SuhA5XZyZXJehrAFqrXYYtOh+xCtAAmaSZOBovy5BBBEoCWv0s
frb3gD+5wNJFU0zXrYBdudMbM/p89vk5VNCOax1QXHRmBir+4oSB70JJzRBIvrl1ERccW9YS7B2Z
Tnoei6BfVkySf4nHNA9CgaOl8MOOLLSUs5skMxBZN/oFn1sZvEAPZuI2cxL2pN55rTQUlC4gwnw0
Yp8aiWo66XOCYBA5aAVIW5I9KsJJGl0n5GlOO0ueO6u0vkIAij5LwmwuG19X3L+2Opu07vml5Q+n
ZAwZhe0/COG3sMfzMSt6t9YaPw1VGDNLDYUBzi6o09rAr1IJbY3XMMsi1URqFkeyIle1oTET18x1
mtvI9HKxSrZAmt6pXM3gEfxmJwmhcCQHKeALRIMU7eLOhRqhTLBX+YsxIkKWFltKXM75EmiDqmV9
wq870RLHKw7R8WrVDuBjpoxRrw9kpKGf/Uk2Qwnqd2txDVhaMY8WSbKuQA0YeGS3N6OK2Rb2S1Gj
9wfb0qBFk9r8jmmJzjLd05vj9bdhYWB9/6z6LjaVU4iHZ3t/tKrsxeQiK5MYG4dHn+Vw7lAxjF+d
qkTCYQzMjjuxiHN4wjDfqw3dO6qCUoGKkGKPcIf/I1mIZ8s86BN4eUG74+WLGCWxyOLkO5f9SPOA
QgcRcloctdoqUZtmkfwhyGgrdiK0uyTX66/C2mjhUyv+EY+IUb6QVaF5tczAfZU342ifUoVFtf3F
1POA3NjhFUS5M1wFUI+CBDbamoHFG8Y4P6wsMILDGkUhU8V+OAg1oXVzm2K/6/xec1pSIFk7QBYg
zPl7qlaaUBMRp3GGRxH8jb/IwvUPF9XPxg3/UD9Chil3OsBta97EeWpxcQPDhYr+Ckg/0zKeY1TA
RkfCxQvVnrvCImM/NHBX1MNFlv1lkGorVusqVUUs1NrFeN9270819F5AzuDXWoQ1UpoteaB4FQQE
88QNZqxx/6JLoAdMRq8KqOrbD4/LxGaQND1QH0wYkVN7kfReQNBbXY1ryTC6nwtm9UgG9G57T+SG
3dsQVPs66W9IjwAOFsQKKY4n3cEMjLb/qq1WNr4p9hOgGIxVMkE1+TpYJPfgIH7a79P0lu3PaicQ
9M61Q1NFvi415PiCUrPunXYOwpwPkb4XdoWP5EoNgCkG+eMEq5En1LyLEfsVYfmu+0PlqmxbVcvZ
YyHSxS2/wBB6tTLCSZm8gEbGa7eVBplAHsWVyTC2AuAIdqByrDyQckfnelwIQuHo+hKAjfFUn535
ReFa+YBbaQO0Lx2lHVb1VBUYy10dNBa5jKQ20Hm1FfvTZL1st8YHydHDfx/v9CVCPWW+6X8lY0W4
S8vR4IxROY7DiIGA2aVvnW3/PcT7jeZ/VmijLdKvZI7y1sHYWPc4X7MsrHOTCPOnVH3nxZX5I9ON
uU0xFv472td1mIbWEVrMc8Mdrz8ORJ3dijk4/okGkm7KfgXDe5aQAWLluTufs0pqu6rDwAbLgZnM
xvCtL2qM3R0EtTlGV8XZTH+geRjfkWLeHehsRBVZp3p0LAXNKdXyp6vhTlt3dEe/9GnRmq1ccBkV
fmoR78YPE9F6BCfzmJt1+6tv0FbjeQdYl94gOr9FfYzRHcBlO3jAtx5ooNnuiRp7BkGJiWSDwfxW
xO1oG2XgHRH9bs84vcsM5C72l5b2cmxq4/HkpzCpHYnyh3ui83c/kia+gI14WWiQAAnLA3NWOZe7
v7fBJLyG6jiH0Rr6eIkS4hsQLGb24PtWD5wz0GNGFm2VWm9W38GOqzhTz9Vm8ZK/grl2NscfK1iB
Fa3fdKTTGEhv2A8BJL6bLhSPxV6j3Jofx3aKTWk/5sZrZ46xeHs7p99jZE8ira/gpUVE2U3jdQ5h
RQXjtPsbh72Zk6ek5pVFTAY+mZp7p3ohr0Eaqz33XQceP88qkRJmC7BNesjtnvzt8sOLpXEcaqIJ
u8ZgcpQrwbnnJ/RNEUu1Dvdu5gFV+qZhKVvpGTyVF1D+wGVT5oC4B/rkXX/PqQZwZTNltGrddQG/
l0OcLcK0Q5RC2I4XoM/wP5TtLhpTC/csHZ/KILuIdnIG426jc8CdaUIGT3+SBJQH+fUlfP9DS66b
sBlAr17/Z79+GKVsNO/geRfwtH6Iii+sYknyMtag/HpBcVBKTCbhjp9DBpA9tDZyf5OWQqJbt3YA
EDUO+N4rLMP6ceQPewFs6NaCz8gdZNDdpVCSTXo8VES6I3M5SX6HNBnz6AOzabU+1zIPGpGdsCWR
lIc+ZEwEr6lmFga55J7W1ctHG1A4gW77GFUL1QpM66AYPiXx1Nkrt32+XJzOhzPrWq+YPEvb6BXQ
mLq/UESKrNJiEmfvInvjot7mUyNWyqGUeqLYPge0EF57iMnbIuK3eu3ECJtSGbtuAWBe9sPltd5N
RkI9L0v/OL2QxriCP8/j1rtwu5WYvCnNcn9QEgCqPVWfFh/FxUf6FBD0aUbTqDCaQDOM2fSH0krN
4giaTzr98NJVsVzYMADuDkRB6nJ5JIhjoLeZ8V8/DxvBll1kyYPl55AMT06i+1aMAa4HkhB1vkBz
CaK5Ea7Lw7IYblnyC73m4ayxlNoqLuEptuDQJnzYhZVNfvVO4IZKz1vinV9J+kHll7Yfjh6qVc6k
+yv8RhR16OO0aiFB2QB8R3hgXphNEn6oyP2PVOKvEYnQOw8xol2pxWdfjEeqd0LBSUlYHYyrHCuN
A/v0W3S9CbLsXt1uia81Qmzh2TKqhlngaUN1uvx7NBbEqN25Fy6hNlrfxUOGtAwBiul4aT/Kz7KB
d6OlYku751v6zf833lOnnkuYpApEg/gRs0kLxBjWq84pXcYTFf5/pOqJSzg4Gk3BJrEy1crXejvB
OHoBpn7iHTZ1LpNfaIsxfm5/GIMKZwYaUrsbN7W8tp8ddhtCdAXeM6/ffHOG38tmzPUxxWqpCLFg
cm//Oa7usywY3gfK1wMdCpLFGHzs8/tn4jroYXgLLhKdP9s4w2WZIhpa2RbKYvj0YN5p3EDDwyLm
3K82GEobfU8f7wUStGCDGorpetoZ7Hs4uLO/iuPu/np28plJCgpt+Z+jFIgtWSy4WXt1gbh6uZeg
eIskEfTWc/6rTQxEpkG4mxuMyownuVijWl4o9b/U/V8ByJPsIX8l+QC/BEczbA9bIFm35o1YaNDY
7ABD0P1ZD6n8q3s3niAAXgF6wNCP2/mfSadQxsge/X7u1i4GcrEd4wC0jZJv0wWtJZJaLJEvH2dz
g72xsFlIyTCp1gCBSKUslvAcZIVxwcLggJ0iP11gPYBw7emUWdTfVMSYfewPmQXxOlwKirUgapvD
AktnjIw5/NvCl55GXupDqgeRserbZTpatibGc1ElMHoZ8IGUuLKOvndiO5kGIhpBVcKe3qc7RVqL
XKVimhSpUb+qR+xp8s67ZbisA/b9UwBbQwM0sV5D5vzezuKSHuQysfY92zfMvA2DCfnujOgIggdA
LDOrfVi7Jn41l1dDyT+j7fpsI0OdQARrnJTZo8Px83L8gOvLBuLPug0yaar8+XZFf7uZUmMMFcCc
8VPIFHI4F21kspXaUJC2WWgFj0jTnNJNN09d0aML/ElYeH6971PNUqyCCVxzn1GYKwYoc2T9BC2s
KWkHzxpqfNM1EJsX02+cUPfzf+SjHh8M1n3WamRy1T49bB+veJ4yCUsnj4HqbdZIcodwylBJnqNN
oEP6NB3GDjBr+tB+1A6PMgdZu908LHX5ZZo3/RSF+f7+cWIwCrwJaArHwivpqojD+unJSanjMFpb
pH+USfmCkF3zn3ttKl764y5NdnU7RwgYCHgm/49wPswIiUX76gaodopOxI7/KCQO19F2f6O1sff7
j21BxtkidXiii7nuYb7T22hZfOuxx+SuvDClI4hC9pxWSNlcH61OBA53Txh3ErKtUd2oolCXEs3G
AizIZr+Mvu263Fo905ykSDLHf9SIcXADilCBoxK8i8YzQzPQwE0/A00JGH37VzfeT3fFV0dkz238
TnIuQKT4CUA36E9lMaMdHoW5LS9HOPQfmCjKhkezGIVdCrG3pUti838M4CVDPToZU3YOE6oIvpW5
JcFfi66jntPCPzZfabV21Q9f3pZ4Lc0ag4V1caMvQQXYZbsj+3Ej4wx4YrxTYAARF0j5Yxh9Um/C
Ppl1aEllYHGKOmHK9Q1e/RVSC5MW/OAIYae+hHIsdSqnFFphvD+76IoOaSFvNNHyNoimB8TZouRA
IT7POgIrU7mnXd0CzM79wCEZmCVq7j04NcsVmcM467dAcYZ1rkhGGZa8qvdNA4gu8Luqfa0NJtXe
ETMGZLwzixMdZqdx8VBBZuxShNYMDASIUFtZuYXKX1RUc/No3uw2kSssdr84OSFCMhNDGE9rxKDV
dYY4RMbs8qyTRBYLfmoaQJkB3u3eyIYQOyTSG/II368D8uTh6QInkr6GWVZJsXWsf3ss6vqQ8mlZ
UxdcCz+mxSr//TRYp/Q9XVBArazzz5sbL9/19PbvOg7Jn3BT6kBCkYCRCX0nkRbzQhkUECCcHdxI
whdIBNz+ENdOh5qLZITARS5kfcrlTdRWBimIt2L8k9QGuKjQpJoYO7IozZNED/SqTOalUQrIqq5f
GEsq/xuIleefCv9qT9Qc5rJDSNZEl1ThgSRgHa/heBOrZg7sByGZcWV0SeuS7SriJ4CcvV8VHFZP
QivVcxx/KsePxRR5J+AaZEGLiNzxteL3tN2jmWz7oS9PUtPDNAsV7TDtRTnvm0+7xXZ0bJF+T5lq
v2w5FnMADFD1gk6D9wTeW0TwwCs4seZgAtf5RKTdbj3y03+ZXvkUPISMb907JjKA8wUwrzQhvpsF
9wakdOizpRFjrBmyluT0Tu/iZu0DQbK9XVMbVQHpoyOHziClONQJL5dUqOHshcNhwAMJVLDkfwr4
X+pi8Q/ecIhY3oP/QYAMS9Kq9Icn1t8xsFoSzQUid5wEwCRGMt8o8IlnEesy2ljF0TQPP2uHN3s1
XZC/ZAyHd98uJEPUdFn8VwRZeosAbJl13IetAf8esvN09mGBK2JcGu+fPJsSwmJMoxNUtLK8bVw0
iGEKBNo50nypsOXjKuot0FmjsdGhjT4YMQuKID7LHG5Nz0us99goQb2CWI2z+e4zrBUZ2M+TZy5S
8+JnH/fz1WTWh0wmhBfz9tPip1qLgrlGVWoO/RKYGb9c5GVwMQKUoCEypv1P4XGcFRUPyR95kZJd
u10QZ/CGukuVXh6uVzL1xykcqLG6uR25j5us/m/F+N/I8A4LX3aAkbI62FcTbqt0KmZPCvtFBm9X
vzD+errERLR/IP5jJP7ySi1IUmbkRv8/PdqsTovp/NpzrwvRg/O0xEONpNjeuLmU7qRzGy6rF3DP
DZcRlmZlEZWWOgnsla1TxAbDxJlrZk42gAPSanTU8yKlaFoZOavYjaN8qV0h4mtr7MkcR1oy2n+3
L+td3L6VSrfVYPgqD2zwfzOP9LXsJsiO29pEOrR+ltK8DaYNtH5U63kjRG792Ex4DC7+jr7Y78pf
WYV1GHPsalK4Voo7coLCJIOO8bIhKzh+a1ujBAj/L6WACG3EYCbZpC7gUgARSY5nknoYdDYA3l0e
Kx40OcR6jPRubjzak4Acd9Ggg9LvZS5lM2oFQnPbNfk8wwFcUAoMaP57LPQtNYOZCLi3tG5tdAAZ
0olDbNQl4FJu4BRVkXhuROZ4Op65tFVRm3zCTRbKn4igQkrHmsAsFziTe9l6yufoWGeJNX1/3NjC
xaq8/aO2z1sAZTyPQuD7VBsS2yIsQfztF34jrypwvFdcberw9ZyKSU2Z+BYZeR0j0E5XgXfkYpxc
onNMh36MSMi2xAChKskEepRrj2U8OU8p5IRNn388nB8xFPu3nKr629ZvUfCuVLiPSQH0ReU7t1ci
zshKhJh66l+GVRfU3fEmZWFIESDeaKkt0diwPBiC+v5W1wZIx69s02fcxq2xqB2BlAcfSMG4K8Xt
YFBqbP6CEw8yXrqZe9U6vJiowZmn249+wzzV2yQplXbogFRHC706BxSq1CNatoS8BU6uVZeklezn
9OOrpEeZ6d35uzaEIMkeqtOeLIAl1M0F3GY3RTRFMloggMQkKfa8dAoOqbZSRdSBeq+mYdX+wwOI
+jixwUy2gWJmAuUzjU9Vmg5lQDR/Scoxn/q9SREjr1fk+QzGP7sUCOjCphysKlI2HNrlRS9cFxDU
edxOpJTdWvr7HvLWdFoFO8ASjgHegQc/3dOjMHvQJAxfPovZz0bF21aOpKO3jWi4JPxuwRzvVMlv
XYy8kS1KqQcKD2sGuxqEGp7eqz+LZRP7gUNycam5t/69qojYXnaCq+he36Q4Zeio5pY9aSE4ZSQo
e/BXj4hGGOp2JvSc4d18y3eoOuKzGhxBbmowbx3UhMxrxRMd8SDm4ggFd4G7qFHICeqmPXk93HKX
KBiUBO2v6wEjYf6vhcydUSTM8VsjLC8tGXecejj1Z5ZCKTt0ZgoCXqyHNUl/DZ0kW3VM8zKlrzzU
LK4xSoUtQkeuiqWuZ8aAzK4oKU/BTfFdp7hQBxM9sOzcIQoyuNkxT4gGOhvZed1SCkIBvXk1Vu/a
6xorLEQgoThnTU3EnUncDIpQC3YnErEjvWOab2Aqj4IweoDw73oHTS/I07h9Pt47Jnvyw+ld/8pD
rjOtkuoIManA2+qTqos8hv9Tqk6WHmkh1I4J+RVk4peB21jvxtOU4OVt7t4yLqAZzs7Hv4yzTpIU
DBzpMVwIgJhuSPvGR47WrG7zb2BD13gLOHzG1yA1/o+hTZJJq1GX1PlW1cga5jH9coOJPMwoJce1
3T8jBMyHDPp3tB+EIOcqWkYeZb1UHit4FCy8hgc945Ea7az4ElbuNY3ET1yKVrKzoLWeAGD0rCyF
cPaIhbFy55tIYUhlpyQHKHqAFaOeJIL1Py8/h76s44Fjav9zDox5ofrsxYK1RqmzZuwEztsq9yUX
a9DIePRGKQIXymPZRY5d2CE9/7rAjegfE11CI1lmV9rnAhTA322+tAImBotIqCR2/5RTErn/hbQ1
mEe4idUVtMhzWAHWF2qJorp52j8QdZCmZkYqVi/+1jWm/MhrL23foIPSCE4dYAryTxLd8OG3eFXM
IrwRGy75MQoIEb165qEsj4lHeKlTaRDvH3FyeK4+5sxtQoXU65mAClCwt2NClkpvdoec3q4pV9rZ
8U9QF9xLRkHrTAEUaaheOtmsK3c398e4Aw8IVp7dMeAX8FW6IDVOmH1bDyqbqPzRUxUP+P3HZ3uF
D2dQXoxSrNI96XNVkNABRGs8KmuEkNBnD+M46d88g5/ahAqabNgHTNzdtqGejucqzxygee9LjXL5
tj/ZVZeMrmXLbJdkv+E8wsKGs/nteUOH/yEB3E0caCuOne6V+FZHyoVLjRPIJJOR+HR3QEmGoJXi
oMJHHpO7+rMFxklA213PY+rmc+KdVK18fmWYCGt3jw5GUsfCwtBhiYfyyPp8AlOWeIkuZflZhWir
8IXp1oLiz7nGKU07phSzLOpBLr20crq7IKhOoiwrRhEwFJ8ZOMy+ItfhCGUj10WCB18kOjrw7Mn5
/wyr83wWUjIv+Qh5yf/3G3P9svrZsqf/GhYJOOe2aUt/PamWNIjcFmCJcp47cvJCBDO4bZESSg4/
1qdEHK54fkNh8rUyyU3iYO/Z7vPuKYIO7Lr7xcEZ8kul6Q/QBM7b3H/3sCsasmE2/R4X1HrbNz7P
FEbONowT2jv/oPNhA9Caf0kSjFpyOWwqZkUaTJrzOsHkb0GprVLiJc60OT+v7xuZrhQ4cDsABexs
Y8PCw121f46e3+kFOvo9ikgcKVRN3pic6eh01tPxaFW22/by8yrRAwEOUeuKX3yRvXB0LEdXOY3+
sTimHgBldvPxgkXkOXZCcAT12DaocrKN6dtzZXwxwsIxcDyHRlVAqNJTKOlkin3vmdkcXsmCyE+F
QI8lrbQLq+v2Pf9z1gybRWC43S8nFDaBV81FLhi5uQJH3Jn3HY62JMqF4Pp9gULon88N5HvlYLLL
searNYUs7KY6UY/5I3n6Vo9T5TSjdQYodZAB5mRfWwVs9oqfBwYEaC7NOOBBD407DaVTs0gav+ez
s51zekHEzV6DMajmAlxamelXIXxkgAuuQtzosfVQ3QpzCqdD+B9k09Oclbk3SQtuzEUzzFS7a61g
S/OpJFSTA9G+9mtZ0f4+4AVeoBMcbRoI5teZj36e5MoMVBJ3P0kIuTlY6SQRjPBXXUvS089Lix/U
FaVQlbUxIwjrFK0dDewOQJrjziEIZ8Nw8k54OvPSVZAq5rTUvXJCzFatBrWxMgKW7GR0wPm80GdI
HBvIqqG+rGTLX1+ZXsPkYzUmCDjPzdkQPzdCq75J+FHh7htidgJpykPY6y03nnvsc048cmDa2+rT
iYXUg7cIVjhVy5n9a+LNM8Hc1BwCY2zhqBO60HQD+FubMqbFppowsbQDtV2iqPxUOBJrvrV/u6/C
iY01gPRuqVduDFjBwrZI2OPi6bey6rzBmMBPgcWQv25wEGCFAWBtVyfawofYiC8Oia3YkN81QRwX
U0aXvNXYkjskp2LvRadBn35xJIYqV16BAbZutkS9CWpeAy3Y1LYyF9lp1/ZcqeoBYjMM+SGMkPwa
kLGPUv3WJuZ3lWuz0z+Fv4DD748w8sDXeEZBfkAm8pFyPtoYvcD9Vx3A1wP5bvwb/dilzyiAGYhP
UKH51MxJQWYtvUlamYsvn+AKqhOqCLJw33+UOYYCBS54vqMXwhGgFMDF07UiVwVSS45o0eTfjS1k
jvdeHzElQYQXfefLnyCeFY5/j3ZWWmXp7MtTIwyKg9A/C4TPXgJV6Ws9bAqkX9I6Csl5lXfOoaq0
Va+U+v1URQPp6/fN0nTgS5oCWSkC+9vK8Ern49gsY9HdVvtNFSn8b4gEkpsZRqrSkIQwp6UgGlgk
/coyPBkcBAMo/WNr+klSMuOZb+PtW0fszuh9Q5j4Sah/0WMKFzUuYXR08PHo/wq8ctpwBbzAbA2D
u9KhTfSWlO/ZJTGZ+VcUOWLCjpOpNeTavz3UWA5IEmoZwWH0PG/iQGq53qLRy7qkFHaD7aXmCA9F
CQAqekaBOIKuD9Ye5zVpcZrbH2v562fU0QtRtZoQXzjsTFgA6x5rEIUtCkyvsXiXGxvfoQ5gbA3J
rzJ+HDjL2RhCFq9Oa6qIBPl8kiHvydYEUlikbwkjBS8J6XW0SDfXzu23VsF06tpAp3qs1KMqJnZ6
Nl3jZ0fgvChA85lbt1cmBA9u3hIJQkC4UbzgcUzCHQcKano8zXdCfOesoNSLTDY/ecPzbsXCT0qv
MA+wwp5Dag0k8jiGcgvbnCAcWsxa6V1sCaJ8ZXsQj+ba8eueuKYZkCLN07jmwLLGK7EuP2D9fLpw
yr5W8SJ6Ke3FUT+h4iSIkwazKgIWcRi75Y7R8P2Q1FizyVXvI2orYItr545pUM23K4UAVptckrxV
gm5I63RezESqEJLEd18DLAaaF1QUc+I7mFzBP8wm6hjsmWNjYGl1i5WbiIr3vhRyENQpBEvAWoQv
IT1okxEbGj8sHVd8YLIn1sOl2hK6/yGg7AH8xyFSF1Fhf6Cc/Hf3ANPErynO3c06C0Y8RK64LYDq
E1Fezpc/F8PruaYBP8FmtaKLNkHT2UbaD1du2eebxg2DRjRXRQf8ThEnYAIMR7bh1rr47DuJAQbT
wrLT2u4EqBiq4aB+1ZPF9FM6Pp/UXACJtkV63YZZV2S1vCA7VdptbxvTM5PBmcPFH7IyfTCoCO6t
x8y4Em+p3Tq/pB2T8rAkdVtAtCQrxxTrWu5PvPkSoURlc5g1dIMz6ZxjdyF0kx0NuIu/D+NWItqD
UH7zf/34wH8l25waMjhOnZOuvk4VEIGFajjGqV8IL/dt6ctHXSXozMZCXrxwSuAgqVM16nkd4wg1
CU8GBXuaJ+KKXIepihzEmRr6CJes4zWjUnB690Lg2dMV8QS/GyF4yXoqpQkFzcY0AlweAXfj8s7e
frRGllcq8KHuvngj9z8IO4qncs3ApnXlTyKTzwc1f6fjQTTNgOZ4MEKMHYHiNhRUFqGUzGWIA7ya
dDhFA/PQyKu+4V7X7Y2tImBHDk+EE2a+X7jkzTZtVXAsFrJetBBMm+bMvhbJznHGM3jxv7nAZ8m2
i7nhpLnlcyGLSrziytWLvFgMCPdgzEaNH0FUHCYc8KS1fBQGeC13wiSsXNCmnLV5db+FshvNDafv
xCa8LaTr+SRFk7j7Myh5WJFoTur7UDIGm3ejxFsM8dZNcsVU+uyc77oSpiz/jz15frjLNOvPv7SI
b3L6hJw4Zmf6T8ARO71WVHU9D4tc5Y+/iWIbUHsurN02CvPj4cuaA8xG17LnS1/WqEGtF1h3RSXk
z11lAkS3iRGM0LYe0wzNPyes8/7N+RC3bIebsBwd45RwfBzKa6mx7TElrgnlR/207pSt6idHFaY6
Oa/ycVfFVUpexIa4Kja/eNM6iUBJ2xz2oTquKuBv4I35yl6Wuxi0um9yfMS4OV0sPNJO0a/BvEq1
GiJrW7aW/0RrmeFWq+VadhpvmMF3GDPB/enuWaS45WfVP0TiOsZA15P6znIAiuBX56jwbXePcuv/
fS2ISFPtyr1iKVSu4GeQUT25WgAMztXwBlKBdJM72C02imRwdLxIHeD1wjzEdys8mIEFIC2+m3dA
WP+S1FkeSLa2Gh0E5gvb5C9PDd//IBgnta8iPKyRhvSzgA2CYgGciKuce8TjqR1H8HVBYiWT+XG4
G/+x9nfOG1B5pjP0Zq0UuotQmOGzF0Rd+k9ihzA1xoqb8mCP8i8SlKEVd4Og8sEwYKcwoOrKaw22
U5beK7UJvslUN0ucn/lFA7gw2BEtJvhYDvUxCOzhkGgnhPbFCzG3xdR6j3cphZLWuzzAdDqtxf6I
3xMZie8defya1jkcpzzmH/dOiWhFPU4GpQ24aiXYvZu7UPpLc1QtCqKmaXDrGKehp9CXGEtypc+h
uiKiM60MIsB+XXa7ta6cjbm2ANdm2DCkhQ2uSHwR9rJJ9SZ3Nw/+HRfHtvcGrD72t6KxOdPiqr+8
dg9KSKir7T36wNuIoSAOBJ5/1nIhT9gJSc2CeagMWeYzC+wGSF1bn+1vg9HozZuC26XwomPVHBm8
mr5xE7tOPbK25JISZrEXJigBbuiiJ/wea646VF7q4wgT+1qy7m2upyhQvAHTGcC1bGHxpYDk4+ki
aEft/4hdasLhHjMKjhdSSlRN6HOEM4Buk2MJ5pQIvlV0qyUjOd+AejLHnspIWD/G8smH27XrUk91
01NwQxoktnd3x7dxfL3NTNZfz5iWr5RjF3t69Zu1claP3DogFc+pbBlLRBtYGdt02VYMgb/LWpv2
dJWEBj0njEzfAvtbAvjCBgxJQmNjPHqx6zIyvofNZd0OUr1fM9KjTDMmLYvi367958c4Yn8WOiX7
FYiaXedUZ94Sagg5HAZiV4FY8etkjQluWlVfSvHe4aiBAnZ14K3yXAV2EXj9Y73iE44P/o7EBWy8
y/S6WFQ2J7S/y/j0M4lUDTmdUIVJU0k7sFGy7pjKth7oAm1M35N9dDd4cP3STsZDJS3ak8H//pEy
W+dIeg/QUUCIwljrYNDnN/CIFmfEfK0RNqlO8LiaeGr7LHN0AHFknmh4lGUmE4hgPNRJ0EuGBD6f
sSjbmG0Ydx+0n4izH258y5ui2P6R43m/zVFqOK0aykMJj/EpED6UD3oMbRfYQ8f594ynKsuU8/Mr
hvYsRWqIrUx805f9lqDcGbUrjLmLvUK7MPrvYS5u7aPy5OnzyU75e7O3kpjpPqjZTpNpIIHOC1Ih
WbzLzCYWmYIwzHRg6+U0LMxyxyx3QppE+qFIeL/Xy+eVtlvOsgT0JVV+HthtgkadR+v+4cThoL8s
hYs6CR99lSQ0H2hhSdYFwaOaQu7ShKlDDRGwoWHMKC8meKvJTHW/cK6mSUM6cPFA1j0+RhK2G0pL
5m2wVh++SLDTSM/ALIQsiZdkKbArD6Xf5brZfwCki9fHRGCXb0+/dZdYQtZyT6Q1hTO5+faX0xx+
hWyfRE3gy5x1KOSCluE4oSb6fJdL3IjPzUy8HiYvEg0vlFM5gWteNKUqZYv6yVRyLefoFBQjXkpo
GNTMG88TAVi9d9cxYw5ampo+kCds381G6bpIoP1WwVADIkLkMc2X4qRXLOc6WUSMV1Wu1OWuSQrD
9+Mizz7qaMla6Xr/tPvQ4OdWUpUtn1qnov52TLwHy5CvnmP0nF+yxDaAZfVFLi8cT7rsQYUZPjNN
xF0JGNmX8nyhcdM7hzvFpAuhuUPSwrfk9LSliilPfn5xmJkLxyrsVDoKP5Zhm76eB79KF4XBlib9
wp0APC3zLOtgJYtr2arBO5EddXCkhbCNu16LmX6KrGQfL4yP67Sv8SGvepNUetjzrA/LOImP03Mb
D3A7F5jGlBQ8rdsgohZCSwvZrlVQx8SaDUO+GpedcKAQ0RkgaZKp8XL3G89M6MG/21LwDGtfxFL1
4aSampTHH+u88UcMUETqOziSRF9KkiFvc/GyNC79vMMlTcHvszWCm/MWiC7X2w9EadYKHno1HdCN
2mO2cXPK7iYQfW7tAiPG7QJnhbZHUrWPtzIwBhyQ+ND517w4ZbGT5vmEo9PVRQJwqLnbvsZ5I2UB
wv3ara+wn6pHdjiUpPLOx2U42j5yz6jdl41IYqCQMVaRajoy1kuRLZH7w24G3o7XPmY7igUMax9b
Lu6lA4nniXZqN3QkJaoVaQZyOZZkcAxjZw0nz1CWqKCdJve4bR7DHm037iVKgRw0OtK83WLYZw7D
z4sGF8ub/zcdF3zp8VcZzFqtS+kduurnaAkObnBTdv2XbWeuozqRXyWWkE77WZr4vzCOUOS5HA8F
/wxJu5GaHRBiKar9lqaUEcKxZtFlQFzS+haQhEPzgRBy5V7XFLStpcJYfcnEWXMsmuhWsChnVtbA
OTMzqmbegwPUm8P4flSz+9vfCEj51XwflkGVOqAoRtJmT1EthAB0RT89B33CG3wE+P4j+vpGB2FJ
5eq1FJLxbxGYPa0GFdDSaSbmBi+zS8yRq06kmWiL4NsE7SoaCfwU/KqZkCq6I91OIkdIn0cg10Pr
GSXVE7/Xf1hjx+DZKOML2fGlwzia7wEp5W8NTMZXCbfU6WImSSzj49waxkadPVs4YrR00HNp5ozI
HKnl38fQnKbHN2kuXvOTmMi2v2Loz3CzDo1Ko9Tk75QW3uaRFan9uPnDanQ8jKa5TUzhUjhJ+F9P
UElk/sDJPSK8N6+j3NTypgR2fzqGJ/Q6OhvakdRK4LvQYffZ9FIpETBGevhAnEAntq0o4MvqopIX
ZxnUlcTSBwJG6omxLPPR07tTM0GgNmqJYFF3tw6nME8AEAJ7+gs19lnLxlLTCZTyyGfudiyJ9d7M
C8mDZ26CE7PriU2TLPFoI6Joc9lH4GSVmHy3iVyG4qKnRp7VefUQ1dvcFPiFyymERqSe3XMTr6cC
O4JwwpoZxhlSwoJonhwQeG3ScJzQXbhUH8QNZOBYH/x+MaHu7e+pvAitUSPjnJkKhmPlkzPl+Z0q
tqKwpxso6V3l2Na2deBbmSANXX6DpzxKkSazNEz3ywY1ulMIZ2qHuoUeR5oRbt7X207W2+4yltM0
IsTUu7PW2DKh21vRuVcbgN24jXSueSG+PSNnkTmDJHQJmChPILjyDmJw2PWo9/f9DQnTIcb6xups
NSUkLKWnxdv3eZTTpr7nuRlqsDAyBftAQiavn0rsX515DltOjOrf1DHNYqT0ORq82J9XNePPdgHB
xf14LIcwuyVWBDQTitw1++bZ8ukHj6USFEIXuzJSjw9zLIkncDxemYUBAegsinhnawBs5xdEdhht
h8drrUPTck6qf1azCFKXsFw6BGFihy3EWwETkFcn0ett0+XN91R7/KULResZGbm3n6Ds1S7/H2n4
xVuk4CaLvSuXID1ewaJDOPvaCd+p3TUNP0IXgXi4m66YpFcYiJxDg8DBNvrI264kXsUo8JjGTb1J
JjgehBhFKh2zFEi8j4JU0oWrw59tVAQa5VSYHh4O564nC92k4ZtArWj5SRUMbqUSyruFqWcD1yTs
1THuTrcicfR/RC41RYt15qrFB4tR3Cy9w0QL7TEZYnJ94t0RMhcf74QGskoogeiew0/Q3qqoHONR
K86vnSxfO1lHzRGfXWHvySuy6f7o9YU6ak/YVG832PeEC9v8GZWA1dV6dzEtC5EmUW+yaujAr6ui
kryCTLKbohZH4vMfrtgks2uBJy8KKE/RJTjFNQEkG5Lrb668sVkiWtbHwWcWLsBiRWtzfgo4sZrH
JWk0GOXtNpny3gVCXJYSB//XTiRH0+j6ugBNPulDiTBl3BqEiMrKdL0WRB2gnYHT+NCv3he4IpDS
uF1d+Nvhyv+gs//Xs7C5CvFDY87+JwkppbzUrhu/EsHItxAz409OLZvqmeL8nOBOO6BfKiKghzF5
dRYaGU82aBMUjIzTfBmqlq7Ze/G5GK7nEdY+rR/1BnWP1bcYW3DA1/hA5g3HFhSpEVqqc+foHAdj
hKyNqdnJSvzgqi/9Yj3a5KjNcfQfa1sf6sWcw5K6Rvg027XmFdDIqiDYDYmyWbSVjPwCDdqLPPVl
UpdJ150WKut4NTsRveQKt51+GnIxDn9nttjV3oZx4YVXyL+3MdO83AZewP+bhzA64t3gI7p3oiUt
OIsdvBBp5Qw1UzPqN3zUS9uSzZ7+jAzkvORcjCrxWsS9O9w8RvbjKZ6q1+ax/E028N0JpB6PEBFq
hdOOxcl3Yl86G0NIw5g7ECNSCICtSPSu8FKD3kARqh7/SWFbSzPouTZX4oxVKqKyv2ASD6bDinLX
c+ukWD6dA95Q7luJSxeo7j0eroLnx/Su1xfoXW/tYyXHcOhrFbt3akfEX4+OfEpXg5Ul5BPWKFoj
qbruLJ0f2armIaYn7DSIQizKJKkTuCuiyrXBZFF/gJaLI9w0C20p2xxDCZIq9HttyOX/yN8zRi4A
Nz8fBveFpcAI0GT+QsP0YKlnA0dHQwONmaWm4WvDkX/7Xc/ezBj7usTyoD5HigoPzroObq+cGhmM
g5YzGwpTjL6HxpyABcn+mA4zYnwfpB7gavBVEOWjp4VHiIpEIewBysSuQIth8Myv37SkKDDgxfDl
FKENbTK9yljSIlUST5eYsZ7dIUs8/dMfyd5P9Fq3jdO0GmAOrDGLTzHKlFiwSNUNDNkXVYdSHGsD
6y/Ztf/SciLl7UcXOerjsIS2eMvEgQjNFHSMBfnMhwzx4NZkSO+CAs82Wq4G5J3Bmc+RBUBpjld3
qFu6Hv9HyoZzpwc/JJqX00ZcMJrTMYd/SOrSf/vE8VNGBUTSf7qtgzmXpQIgbuhyRBF9IZmIsOE2
6NZvuS/jbOkJzvTF/748x1V36RCz0OCr8EtYK0nJ1oArRafgX14d2+VYay/rRCFlg7xkb1DlNWx0
lVOJXUB+7Pmi3LA0/ByqUsuLDjFSbRh3QS3HWttG762XcySZHutWlvdfTi1W1fKUdLK8PkRht3DG
1WkMSNs8XY8kLihOM9JPetqKXSVW3KDPXO3z10DPNV6jkIMWZi8WzhidRoZHvOAAkR6sHgLP5ldn
9GiVZgSV6xOScz/qLfCwIkCVcd0rz892Qc3Vk3yMrDkWh7oCXEQpUwcvdup4KgmPT/ORwA711t5j
0MPZSztNNoubzoM2BH97VPJBt2iWHy7F6ESTmN8kIwXdJXrCsrKMTGCPiV3gXmDVX3Osbf2Q4dT1
YP2Iqa9L7wDdprzgr/YcM+72/yB8+83fbPJQNFvN8NebEF+2rMAkA+8Ds4oq7sXZeMvSxqNS15M8
iEF91JNJW+ZGvyll4zvBt6JkRskGq8Z4pMnC/m1qZv106tEJG9R50JEZyfY/JBzNIT/dVMhxBglO
q35un745iyDhOq7rDWlH12mjR9uO8naryXKu4C78eb01IGtfOTUSkvtYGf7eN+F5xi0DcYjWeXm7
5S5iIiEFgd5G7e2gyTnNkL+feUZTGK8HUXDfQYOCaiRNA8/80SvnVbjA94FFahWrKDq3UXZyem97
jW1543JQdzNUR8tNxmIgdt6BxPtQ7Hn6U6WUtdHpmk3RR/cPX6zxhIe+O6sh/c7np7gZ84C1ddAK
5W3KKhrPs9JOdy5d1ysnHlfn3rAvNRIJd4jquDTpvw2dGie83q4+IMxbkw7dqVh+7TZpXOomZQbf
9ZCm/6LLlygXMbCKRJT2dBAHpBBHztQexhCqLMqgekcLId1JInQDhiYkTuOl4tVlfVlstim2crTj
WosTGtBgrNZLQAqV2xFGbsn/2XJqcqP8zkRSplXONVaz62aXF6/pqMyJ58OivFoYdazW6yBK/2Zi
Vu8pDvo/xBZuuApHaKZm0QMrl8qtxRArmnFUawls0bmuEUvg0sUzCMT9QKqJ4skAEg6rWxrlhnER
EinQxp/KY2iqWFG6lFMUdTRlf+HPwbS08FbLay6cNTByP8A74mjXim1bl3XFyxmTytDN62DjJa8K
2hq2XBiN0xZ0aRz0+WtWirH38NLyfpfGHTpRHMIm+AZtQ8WhUUZw5RWHGSj2f6yKfaLJcUnEhxwK
KcRkSR+lsZnGPckofj6AjoCrBEQuF2uQMsQf9KcG0voaD/ALUxp8xqLMcMazn+eE7qPz8QRBDd6V
qfUmIYNgJKp8aEUZLO+DGEPWm7AnMq/3QDZYBSVMWm2fDI4+0asOG4z8KS0tK75pG/Afc2vy5P4z
TVWwlJsNa6kfcnpxtG7jM/hFDmbbhwk+T6XB4dmEBOFMbjjHbz5C/hQLnIGyxB/Ap2/LgVmA0XMM
gTwFW5y/4NFS0E2mY+YpEm07nMYUBPd5qjQRwc/C2rAFzg3FNX0ywn8wxZZr5NwSPxVPHtBZps5U
ogQRNGoaC8PMce82BxQi6YwwCpzj74I/8MK8cds2s3rZrPdSrTGdgSaq+p6kSTR11OZiVrdo6Ih8
orXH7iMZeLsDPjhmvJhZQbQ967Cgtr9dgyu44QjcACsn76dHqwPvr87lqnTTuEQfpgM9SvKu22d3
PsFm3y5P6druvHOEjYOrhb+WuWCXRQHMJzN2/yaMRbb7PfygDgBDMkdjcghAxSmK3eeE5jb+D2ck
qfz9wq15Dci2qaUfscjTQmT3Snjd61DXFTzDIM8HLyxDiSmpJalapIf5sag4eBMIpUfT+Vhdym46
fBVcqXOLtkUfu/2r4/MabPR3vCcQrQZueMhxDz4m9Ga0dHDplY45dYJV+8PbZwHJhwelOiPQsj9A
sW2i8MCgBuQuJGA3h4LfleM4CG4eqv5D24r9i33XIyksfBGyCDmvbU83wwgvlQ4OpvFiR5tziits
i6NupnSt2D/PFT8JQ22n/KJniOwOTL1TtRMUdGXDbFRNh/5hpGo8eoisrA2jabOYlK2VgwI7J6jr
WkCBcpiSqDam4JLlcX7Ch7BFf6EcQ0/0QNGhdUp0KwZUs0+j0TAa4mTPne346WDwR/McuGkqwyM6
Ibb/CakPhGJhVghg2z436zyvY5yzfydIO7scy+nfB+eCnu05oY+CD8l7sNFqlxcwse2AGBEW3ULm
1Kl+l9UJ8I173Ykokz2vjzs3UldulGNVXHnxbLcifsRwPpB7pglkF5r8jUKrFxqLfQ9k33e0rLgD
+wbGfA/Mo31CEYMldt3YoA31cZekpe9YrXqMr710/b4Ld68N5m4hfdBuXzzBESXrkorXJNBq7ion
qJxH/xXazlOZ/G7Z17kWwNdrKJB45ufbyTlCUX7dAayysRHTIo2arX1syL7c+/H/hT7k401/oiOs
G25PVtMf79cnh1PCW/OlfuCQ4xg4u5iP5w+4TUyPIqQOYsbrVhVAFbvuQUjR31IZMXWuXXKPLKru
l0D/ELUM2FzBMfoUJK4NQnS9HiuHRQhGBNZlx4B4oJEkPY2PdRH6eBCKTvplwQ8qME5FNDl5CW9H
etcVVmy5r0Rppypb00bYp28AnEWuIz0lenNaz7eVz2fhxkoiCaQwaUWwF1CLNFBaYy60QMIWJWbq
xhHSIqmwq29GKfzAtjvd3vcKPHfKrxK9JpzJsGsiWe3JAu/Na0QeGa8PzkN5oPY9Fimd9eRKUc2v
YdMghQyjTrwwSqNxkzlXFzdzZ0qbeSRpJjMmyBc2R/OVJHq7SMv6Gam/flv0mnCm5T/nfAqczg4P
HPGEvB9baKHbnE8PF7J9TpZTDrGvCgE5cpWfbaYtYtFvLK2kY5nnuf0gQQX6a9W8ocaMPBqzkp0Q
1HuEmLdavd0HXFec1lW3ZguLn9z6Lzz8hpGK4nW9PMVPFhCy+mNPs3jHWzI/SutPiPC4tb5iReod
WHGE1/DpMcKrOnfSSG4yJHUuZFQxCKv7FjeJfwBdjHpsJr/zzA03i8Iw8p9koE6K+GUYYNUCT/xs
p3tos6QzjRRUhnk7wFN1x6yc+9ef0q4+3CCnvwgvudzf1wWfglWEJLOdUXR/yh+YVOyOCl510PG0
jnV0PAf+4kWeKJcdE1BlDD3l3PT/6DPbU7uhoQK0Ph+eKHTyFUE9kA9K51kCVDetsLt0i9IY0ci6
/qCuFQ+wQ1R/O046hwk91EG42M3qJSPSuN0NlIgxwhyz8zPlf6oTkOnRyI7IPM3Hxh2Ek3CUq1JH
6fy8NpEr0GgXzBK9uu/ABB1BV3LTVuin2GKWr4zXXEJg16reGNbyknxupcLQ+P5l7dNV0HTuekUH
7oEYb8YVFysRn5hFcYhDLqtniCPIkl3ZkbKLOs7uK3TeiDq+s2Dho6A39F5JTQm3ahC+v7BbWsfu
7/1cnaZWwV7Tz0wAXlm2/jFSSzommb3tzocp6SuHeBUINQQgxCgQIZDGKyuKw02sVxZnNvzgwXme
m47Nyd+mRi3VKDlh+S8I/ajWLQ8MSAcKZqvwRpe27UNe+LlUBJAg2MJGQGcVqNKdg45Sn5sVI75p
LeTV5Zhl4GAFiPt4jtoRRU2YCZlOTWsOxrZsosTR3AfnftlzWB8u+SZxMLkc+JKkCC9SV6qyej86
tbJFHtLHLUrFL5siESeaUPwQ2+UNv3ikdpymSPkA6N9EEKT9K7mwWbWouX9ih8asTV6TEf14PjmE
+ZVl/iSdhYvu20HNstHNQ/Xdg2nJa0q4ZvCeeIlb1WGtqzuXLAVz30kKik0ZZGAVtHWoOyrvi3JI
ZXHnM12IBsiQ8K0qIF48f3BPNGiYSQZA2MWdkzYUeHvDtGXgwyl/odI4vp/EGNdNr2xCV69H3VA3
J4T8Sqx/LiJmhSPMhFae03TkJvEjhnAKtKxy/Io+UPbdLiM1BAPylEWjmeSWlT13N4wfBU9jhKeq
/nKXg9vaXdrlNfhDMRlzqEPS+5fTS5ssBq5QF6Mynie+/QMqrc9YegXnkX3+amRgguNIZnBZfUNO
qDqEgMGNk/llMGAa9bsjl1eVeaSy+AW0LN9nVbRd2AiCETCXbnVpAnTV4PJRg+gesOPo8wSipWeP
zGUvjrp3YXE9JySP6labs2fa6VIUI+k+hqYbZTBq+KjKpqbMl2z9vymYqM4KOmwNDm4qyWIZ7daR
5jNdZ0b9z63MDe1whmP2LD2bPSOYalaVYTrmH4INjpdTFZVNW4UUlmrRawQyo9HnY8x4xe948aN+
0MLEZ4KkmogJZs0o9h7l6leqTUef8I48ErlYk2zKYkWkReutcCec438+RPYqNYLKV9UWfgWpph/5
QWrXPynRo/aSHKHO0o0OK3PI+y1z3/mmgU5eIKNnWZrJeF8RmPnprPcivdbRHtzhdF4Ckl3BkJxB
JZo/kpujvJzzxuWmD1RPjfeltGCpHc5oTr8gtS4kJ3ZTtLq9VQR2as1ABPeQleOXRnZ0EKUjIuCv
7DAQfygQ57uysMLraJyI8SYZj5wzilWgAO87m2y5wsxS8X3p0UZXGFyjLrpEaGeabhHr+ZeDiHSz
/s/542yksB7K6mpyIbZ0ABYq5mYDUz7eeYoyoVACsEbJOP6nYIlghMfz3gT40POM2tmspnKE27a6
Nma788tYSUKD9YW3pGZ4gksCYOG3QTW9qDp494MVvg1AJBqG4sC8YHD5Joeii8UoeJZwQXjnHxE9
yUy7dVfIjf4LO4/nYFGMKjZ3jDBC3rHFqays/tgCcOgYoPnl2nA9gi89bTR39gQp0ZAPHirNDVbS
+kiNztjOlUfKyh+kmkgFQ67Mc1BU5cWbsyImHBABN3VVh5Ffu5l339M1u667Yu1v3QnGIMNhtVd8
BFgdtSMcFmrU7mF1ApGIDa7eQl523pgBdJEe5yIX8gW6mpQsnJBkVxtE0eaJbbtAFFINjE9E0ohZ
eZ0AUXhqk+kMVWFun325PpIb1sGYrHl2QbzSM1ATWOJByrH0VFTrED2+vf3UAX2TQ2RTDPNTpcPn
wyV6i+sEahmWpq/lZugi/nkvqoN+LppCCX+TdFQapa/ZU2FTZx4ZUKuAO2PkZFrMg7LqFmZIzacw
x7q6a7cNBmSJKXTvwg/nFR3QrH7h2AOnuKlkv2ej2ff8HTD6+CWRHxcFeBAPdZozlk9n5wss4Od0
vRp3mIlLvtJ+vFckRhGwOqP68NyhXSDY7OfY69yuJ5pZPELnIdd0El1jnw3wBLasTYqEkyXyhKBE
wIGYL2d/t/fZl8T+1jdsRDF7mllnIJbRQi6l7kgiM3rWnVrRLv7+XJOkw1GO7baAIfPYkX9gItxr
q7WpS47W00S+19Fl2tKDpbjF8m4y2P9jMe0X9YOiLnTVkgJLRj9rNohlZpIrzjFumOe1T6jMZXJl
i5MSN7QFuSQQIuTNYkDI/HQGleSdhFV1qRk6vT1vit5KDtk3/pszUj5eWM5RGXjGiqI0UZhQW84K
F0Y9QAm2k/UA/ZkEvjIKaGTdDad/CR39DhPg6emCJc4ATMgBzD8rEQMJUms7EH+4Em9gngcdfBbt
wZxpnIr+KAzJeJAzijMollUBifxVd12AHgVKO52g2BAfTvWwO9OdfnDARbQH+mT/AGZIpHfZT3C7
Srr0ilag+WcWtYtVEhao1Z4JZAIzBSPtCV/JSMf3HeqP4rnoLjKb4VlEgNAM3EmDd7xcDJZnXPeq
pHNoCoSi1sf5cYYsknWkOPGcYRYUzRFI+KKiuav3EOFwik+naPjGotq7VFEOe0CoUvo9n8hSYt8L
Py1r8MTv+Rg5Ixn5tiq5J6wxd+gfmcs/rJlDDaWdXs1cDQxL2B3Oj9wGWDm20JRNAbXKfMaQkk03
v/qfoBBDFjyrZnWC0nfEIuhft5KXdm/5dJ904a62rLH7SYIIOB9mPoC9JPVA3pciBlVuflBS6vX4
T26zzGT717zzKyMx4hvaOcg1/cfJ4ZnKyKx1wVuCPcAf30YiM6cSJ39soQlI7GQDXZkss9uOxScx
t4zlQHwweAb2QlIrgJCrrbYIj3qSDLkT5s8O3kFyrGz4VFozn8Q9DWLz/Pw7MIIDy9NEkzTAGkP3
nQnvzAj4rEZhxuGlp1dx1iOEwozBWroKNA5GewN9ZVV9Z6pZjjHI1pQBXNxPqJQ2bLbrs51qN2vF
o1zb3d2KVRsGZze4nk3l+D1mLJlqDUVIUkDgJk+gu8lazCzvU3gwGh6W18OG5U0eby5LfsVB7kMf
DeXgDqoFRYvE74t9kGPRvJxqy7dFwygDysbn10aB1jE29j4GkGpw7wIGB1MXbtSah/1nMqp04sc3
iqoSP4CrGhjrGBgY70o724Zt+046UZDMs1kmF9ZGVEkjb59l5wIqVnxq5b7pPVHCkVNeGq0JEYZ2
pKHrNo8rrkE2ZCsnvO6AKPjupUXTZHS3uM/27RL0a43pY8cA1ihNL0gx3xyuTFB6jTl2drH3YhC2
RQNGSpM3jtK5kGP72vt2woxfUnmpm8Y0b3l/A7ZkXs2hXi3cujSufWm2vfikuqdQBe8wWw9rGis1
QcQJfGjZvGImLse+9dhGDwijP+AJM3ayPZpcc/BGjj0ReBzk0MXRouM79a6y8sDqLHvx1L5dT+Py
nTKuQPYfxo9pdgVltmp6eyKzVpwQiXXaqtiTdXaPZ8DLyHzaMUXg/G41NVOK74pbN/UXIkJn2w8x
zXh9OVywdVy6ejGOhaUmAZfowfucKpcloTpY1Hj9Qytwh5iaG7d4eAoz5fgW8pZS/SKU0S7Bw4En
YwEJX6RGtCr4+jU89UtQFtBFPcM5iFKOR7eiWOkNDY6hyKEGrRvOUzrM387jctVJ83NkeVypOnTp
DkLdvxJhXBPlmZzNk35i+ERAdV8zj2rT4ZgD13jT5YDpLrSR7if2VZsvcw/uQQhekVQ6G6gYsWH0
wAQw9aPrX/r5WjZujHYsnhArnyCRSMmSn9MPCEKFsGaFlI1nMH2jQzr4wXEotXUISqChpgHGs0mx
N+al+0QWX6A4MmS5AeJtQhnoFg7Z0IFFSdDEbdn4yrI8p/iFu9/y+W6nHLtc467DdbOFotnmoW7h
m9e5Oroz26AmYzjJ7u3g8aRZDJwKkP0nWvrro7t3QANw93Z/y6Y76h5azHFf97I4oUV9xVrkKKX9
5b5aNbdpOyZBAawejqy/viXlWbhX+SZLAh9mCr/dBKScpoRMKSyEQhu7HrP9giJVMWrDfLSCxTgW
NlsAUS5q+f7miEwzKhlCTAStrDhAUMfd7BgQkrT5SIJOrIxJAMdmhbjmpde5yEKzJwwfMIKBxjR+
Q6EtZG91onChJhfdO3fpP0mF4WBAvgXLG2bmIPdi0xANV/Lv+MCv4uqtoCcq6Mz9QcPjg65AKdos
Ps7xywWxzR/oZ+Yewu8cyAsWCxMVoI23fJhZew7QrCdbhZR/ZSq9mAr3b552teFwzvGAB5G5+jZW
uIarVCPkVl37rmC9OWxoBsgg1xuMRpQmm6nco8UpCarhRDbwkKNNKRcw/7bjRsxwMvFdUFuANTJU
F0BOiDKYtPQOzDR5DUVREgrK2fcdO3hPzGi0CVBrMu2b7dKcf3VVi4cfTuAEuABNeO3FI6tVOFbR
v5vdIawow5oTJftXXG5N6lONCxyODSSaK1eipQupets7hc/B6he9YJQ/Gw9rqrUDSzQyVJ8w+UUL
eZ/RPGLYHGjW+QPVJ3xxb893bLDx5ph22mlHV7Pkj2/fAjlSHkUMmg0I2iV2g+CfXWZG+U10xhV2
fZuZuf0hxKlfl7VObxjlgy9Y3iel2uEgyuKWeL9O04ZeFbTxGzjDrwOdgM6mSP9/aXLnQRCuLBJ7
aKAoMzutfHXnOHvGa7qrTJPTzkholR/qrVEFxJhLa2Z0fdEy3zoQSVP+DjUNxIkkwfh+B87CKhpg
I4CBPEN2ZCYgcL1d45PH/xDMgdOAQ9ttHw0YsSRd26+j1iuqpYQ4Adtdgf4BEbVgXa+NuAKOzEgg
m460+4HR03uY8d2Gs4Ot1U3Crx519XOnFTbLXW3PYBVMkhHvDEkUjqv1POIk24sfDfm+RjQ64Yw8
Zk9siI/JKWrq9NYt+w1GSLNvw2csmwf4je4ueFGGUBVZT6j68gTsOG7rFCZhHSp1FJuJnBBAMl3k
oCx+061HH1xoKAXcAhOBVv8ZrafyBn6dNokwQpBIeND3LF2IqNbw49D02X5sUSMHzwx+HEF91Fo+
j8BxKE26tj4viKppu0uJSvis/2bsb7GvmOfunyysYN02mQiAwgURLtqbq2JfJp2vIUYy8oKsurSh
gwlHruZOAcflCorrIDNpiijVOrf83T3URg08HTfsYfYVmkB7iml3+KULQoW9yPbdTV/isSBXNC0T
rBB09pbhzZyM9CYRgmf0mOyIs/SMOdt0KWsH9ylLZ86Wb8LFvHpmNy+L/Jd9YY680RihVLXAPmBD
y7AIvBjApIrMT1nvgRbHlmhjHdzGO+RjVVzDr3+r9BjJJtT+XKdGbFOg8P4ZxvSVBV+01hBctMKO
xmqT51LtRqMtqnGavU/OhsgyT6SLL2BwrS1jtwDtc7z5NRvh+vw19dVWMM/994UvelveDTVbKv1B
XEZPhkseJMcOmUsEknerymoNKDJHYiCvvtKalIql9ILhX0q0/57pu6lD2p+bcflkhPJ1D7aLEKj3
ndq4hpUi9N2ImXDAl2v1OAA1+jqrTSw1zWVbe3qGYW6Oge9H9XavlGbKj4zXMxdT7UeYB1Sq5XvE
OflGkrQ6nP+r3FgDnsJCeVNX5paUAf3mAZOQRIjXzf3uL6J2MpVr5bDNEJhLu7opcy4o8ZcF0LlY
99U6SYGycJvJ7HKL2KIvLHdEbFeXxOCQiT/XiDFqiHcwBC0Fp/AVOuMmDn3pa89b4Ip0PbtkshI6
5eUhfQ2IlMxZVrKMQfzUbTn/BbddLjGlWwmt03DMqs2Xl3JxGgaBb3pJ9eF2Dk+w30Lu5TzlYx5S
6ncyoWyHgrcWBAZS3NrH1w5eiuyaGzgYHSI+Gh6klpEohBPUe2tzaztR52lHsD1+VMp3eyIlYCn3
BvUO9pxT61+ztEAaGWFUFTyZ9D4ckzqE5Gl4GEE2Ko9MG1b91rJV9roXk+67TeQRXQTCr7UCAcnU
ZcInx59P/yn6R85hpEGpjstBqZj/YoHdT+lWisjOScWCNtP83Iz8neDr5S3wq5/FQrMQKw4l+g2C
/0p3I0Uh0PohL8C/F5AlWbPcBygQmPqJoi/Zi7prAzXYUDB3Ybluz1rjHvQrLb7+CfANBH95AokI
EZORVZ3vLg4mYzIOV4NaEpO3SISb1TKu8TkTg4JxqgFaejQVwpL8XY7AAD3vzrH4W7eSXxLd2Boy
Fvzo9aLoz9oDa3R/5CrSOSIuTqDF/zpnb+WZSzqYdhef8meAAO8d+EYaaGE/rPcLI3F1kTAwP0uI
5A42brL1ekNZaGOwU/hPicMP6G01+3IaF6v2xnFizAbjSIhsw4Mzc78F+ReJZwJ79JW0VFLjPADA
gNVbYhYO8XCZAdcVtjHLOQEyUGZIXerdgN7oO7FPxjiOdrETpLix/kisJyWKb4jttT2rRHGT888g
+tRNXPwLKNeDFJ0AvzfYtl/S/9z9Tbj77L3qGLV9pIu8KQZTlyZBbP0mfRIHW1VtpuFoinbbd/4m
h0NPZrNKiRa2Fl2jcEe5onCEyQagkBa4IxRQIObDKbc/f2zV7nPfarbsJy4aFSofvErM88e7ND18
V9OSPX93deFrh3S7AeVSsJJ8+4SUS3Z+90HnkFZ5QL/K+dmcJ0bI/NH68VBM6najAQ9DbWUv2nzA
0/C7n854sVZ1/a17hE1oD/j6a1opnNDZl34KQCGFHA9j1P9ACdkGjV4QDe0Y/hUnwsr2CYGBlT00
t2psw9u3dUpGyEjZRbY6nKNo+5ErZr3RWI/pI2NWQzVQd/sfE0bS0Mei70AClAKSh+ZTMzDiXuwV
+yYw3iLqNZ/FTSqNaUdcsj8FYt2sszCn2j7a0AU0TFVJKXmbP0GYyOja/lqaPjIoIRgdHaE8o1l2
ANa1Urlodgh+0iulOQtwGv7J8BGnZkwNBQ4M5aJtcvwqF5OZZlwqzV/oAT0nAkuJort3yi9nfPpo
JxGaUUhNSGYQSVzU5TIhaVAROP2JFUteWkrhVw3JU7KUcCvRW3G9M/krY3sSaQr/TvmwPsnSHVln
KpvGur+hJH1CbsEkVysy7Era3f7bHZ63AZrQTGVomzKYDvnRtHqR9W+iKvE2w4eMfu7rBBGs6olN
Hm7tS16TnVH++oeu1K+FEq2ywhtf1lR8R+CTCQTZBkT/QAm1zM5kRm3Ab2O0cLjIh40sxNYbKC1n
nehr7+AnQrbVe/2pHFJ4OdY0PIoK8vYmaf2hy7zd4xHfB7Yg4gLILNWfeNaWz2js4m7J7c3s5lDU
sl9RAUeokF3WH6pmuFjXn6tfjJkr/cgzVyE5n76Cq21UYa3xbn+f08Fegg9uudenu73rzm8XJUsk
I4+OhWI62yOpzMw3nmneJ8eUAo2xCMOE12Rn+vnlQYTsyQ9MNUL9swDRTDKwarUOL+6ZUJiVGk0l
+GwNmCh61lKrrna2NiAQyqQhc6Vu9fkKkmYJzsGO5OTKB6/fRCrWQTRu6YCbBvz1/Zdx7Tep/63q
UZahDtjCq/KMfROUlOF9OwOmrTwH8KHQa/dfarzTTbsiPQXtYrBpw1WLkQPA/IbZ+mMySwUqLdiN
OxovTV5/orgvcdSbfShDfot5Xj/UUxC48CLV4o28YWt9M5lX+N4+2loagDTKkYuMfVY6Csh26aAL
2TwDADdLNMHsNEpf2KVLI8R9NkrUnHRnA10Fr5bmTgcbeLnoq02dFfA9MIFsOYWR9ZtMVrjmhd1H
9A3Sz5apTi9HfhlOIa72Cwz1E+hrUfYUG/+zqrPMODo7yDLodVDN4j78YeXhuhgU6rLQa+jWMEv5
I/Q5oBS6fVW2zuz75l2aaveRob/H+MPLRy5/+BEjybAja1f9vvasd/oVe/n6ndVHoyihQzKh63rq
sfs4uwbdY4lxBMwtuXchqXY3dY+ArccEm7Bu8Yx9DHt7Rt6RnKs0O/NezD4LCYwFgHxpVCkjSWsW
sES0dTcgi1nAD2F62XLxqmkbBGmEr9fFenYStejEowM/1ugDFIntlHU2duPV59+c48kIvH8s4xJG
rA5MMe/2vRhrd/slXZYVTh31fabZuIDNLM6H+esSaCz8nTC0FmqvMITK1QErAaMNU2oGfrpL57bp
dlPWtTRPTRkpYPJtPY3/TBp3TvF51cXPkdaKS+ZQlN9lOGQcSZFRQTmMHRKjc/AIAci60WllgAJF
lzZdm9FzA4fj7yhiZGGkQRCesUjNw3FubCRpevY4JLmAjeqYhAhsrUFfF/uX3Ssk7g5pr6kqu5ZQ
4YpGBfqTKMZOU+gVfu8MthR7WsxCOeZE0LiyZd8pDlWYLQehBzjGJph8G59Ben5fT/0teZ68wr/1
m2d0veV6W5iV4V+lLc/5IZtwzmYX1Rhdd5z1XfUhEvQ7qIFxTrEbZTGQjgZ6lHjtPiVhmpdrYFat
MaXl8KP8MX/Z1PmakDTjMoUSFwLqVR7io1NCrT1JZsY+ZAhR/2Hho0/PCHrFR2Q1W5eWAnbgjVa1
Ilzg73AxzsvjbNw4/QkmSxIlbwkGFbNTouhbDz+G0HUG7rDL/w9wfDEsHwmEI7It7o2FdgJGfQVw
By2eEdHk1OXWVkkfLX0cpCmUdmDBMpVzRZnxBsLs+GTr8NG/BLXKs06+bdsUNH7VsWI8aDmqqJE2
VGEA1RKMetCAzJjjQUT/XEvP2fgNnwUHyeaLP2Hf2N4AW2YVOLVs4n8iKLk3DE1T+uOdwKWQUUFL
SIC7eVqSS2Y+QpQZnZEMnnkc2JKNsKSgga9fhrxu6ymbgEp9X6toJOsBTQIRJHoYi1XFG+k7m8h4
zTfjfJeKVYlhHL37f3Ig3ZC0at6+2Tqg8Bb6wEAKO54DL5LvbQpBgHzjdVAjlLekMwB8wgVFzetJ
v97uc0+DLOKX8twkWHS7ZjQ4mrf5ECXwdZJdcFcvFw6Ic1/QCsWfJcizVH6bepZxPAXwL6ITB2++
3FyprSmTUJHJFtLQdTTfxQWEM46U3W2DvDyZIlDpb4j2lVMeWYRYQlYONGHxGB5U+LkIGhtCbLBN
5CQS76iLj/NymdySW20xzUz4Zo5OJfBOje9eTsViLYe/d/IC0ISMWwZ4/xUono1U+ffu9UiqGyT8
C4HvrC1GgxPlGlwT8Ulx0T7R2TODzgTxrifjc2z/jFzhwexOAylU3Hc9S1TIOKpdY1FcfIB7Wijm
rO8wIBdVYAIw6XSu5cpezieM8t0CLPmuZ0zAAlyToyfZM0w7roCHmwUT/EQ0cJj3A2p5TowLXeGi
1nVqCh4ANY0a9umyXuQWMv/qeFlioV+awCK6LcYiE6H4vcWIF1Q4emp4QW3jxyI4hmJ8Ch5HrpoH
dlkCpfZVOntc2YDdynwh3rWbrse14ciwtF1dSu/4NP0o5so87iJvRSZYxSEX6l0Hc883k7z+tukJ
VqyTzQe37wAsq4UgHhZJycCwOMTph9gTceM/Xo75fgel3WaZrk8lT+Mqtb1KL2Ge2YT5gED/t5qm
/6e6w7tBLVM20j8hAFU4XozUzm3orA5Hu9N6CC4sej93Y2Fn7Hg0Ah6HLq5ktvb9Kt0vLQ41Pfhb
4BDzgDoQ3N+HwtBVc1H9Ez+9paRTbSPPXRgYk6nHzL6ly2uXTXu7IEZroy3ktNWBrfvDfWhiOvIt
hxI4vYUH5qc9KzABWnYLsTzhmUpJuomE40s9WVnnylqmq0Jp6kRkphdIG1NEz/Sqd0tbd2D9J3vj
fzaxptuFLD0vDYpO3sFe+cvEZjXUu+avgoWcOLa/I2WBsvcuUeCF2rDSiM4LGaRzdaGYh5PZwduh
bVGJ1rS8TvkhSzOf1VZgopurX/67ucBx41lqZXRxH2vIyPfPUQXt5AtZZGF3bQxVEgKsjzIDqqin
Mc+3lPiAkgnLs+j2twln4BFOV8+4UVoPrdvz0+m86oG6NiGYM8TQmtz1H1sXnbW9FwzERdxceLLX
5Zx0P7uHGeBxXLuxYX8subeItT/4HWW2l081ULhm0orVBVEY/Eodq4u6A/TG4hfNIJkil3BB3Ffk
h5twUXYOGed5ikjI/sWMh18jOSru9gVq3vMq1FGGSyY2vYF6o3t1w8uYVQoPle3w4LKv4rCNezlG
5RR2Pzt7cJi/i8RU5roK/GOwecP449nPqFqV73MrzJLjzdW/1y4gtF4k7dwuDUf34ZVq7rjStY0I
pMVZa/zlWorODe2SoK+ut5GWnce7bTUUGjngzx3k8hvod8NVPZRWEW/znNqwblV6ygmdGn3sNPjN
rs7m7O+KNDVVIrYClS8hOeprZlRygKxT2cINyjbShGtB+vkLJJvEbqhsae3nLUmQtnQmzesw+9aJ
7//liS3Sl5bS0LX1Qp+JnsKg4D+5KFxWaSeLE43zCE5RKai3rpxZDa9ZzjPi8tmcgWFNeZLJ9Rcz
EFOryaXn3+Ut4CQwItL9Ht7gTeel5RCQ0/Bbc6k0EoUZ9Tb5RH9UJ0t9NvN/72mZyTapvtp+dsKI
kYOGs6Xy+ZhvI2LoY18ep++xgdYGQNdxaGTRN8/j5dCE/s7K6qatk2/dPTiAQi4C9BOnD6Pi83lj
WM5GoqM2uIn4Xl/Quk5nSRhLiCwIm7uDsiyB0cP5tuus3hqTo59BH1LpzRlHXwDweA3OYuTTVQbq
BPe99kul7CEm6IwZ5Li2IgBen5yx8xF+aYYkbAQgDOO8uZjH79DgKdlArseCX1X3NFl8/toZSrHi
AG0NQQU29S7+qo4OKTr28A43wegkIGhXi4TS7Y+kioW59vqeUbo7+7zhxLElwBsC+usVf0RUY17q
/sXt+QG1rGdjl7+FU+T3zr0MF/OoYowSiIFFVoOayJqY2TVoMF5tVkgJlnb98LwBAmTQV+kzNNZz
hRssBmTa1hWKolf7TytrygvpoGaGoLanM8Q6Uvs4D88mxkEw74HHsSxYis6jDUoYBzw64w2StURm
GbdGXpyCfo+E3A+QJMIoOstFOtQfZ92my1JBeGj5tLBfmBps7N4LVCpGZ01SQ49cBcA3fXgvxWvL
vkC2fxUMM4mptuhtTOjL8krlkFMGCxAoclkvXADih6Jgjp1jeJ2EFNO+0jE2q/iycIsM0CECcW51
8FDuSuXcgkhRCqFh6pBXRYkX9R334n+uiTGUGnBLf4fxGgarhAqKHPPgcYlBL7HeAWXz8h5V241s
pr7BieLMZZjHhsEwbBmFg1yUcavurRhy6IP+vp6fm4d/CUZ8p8Rmm//dVMR/ReNJTJQbTK1W5D9L
DvnCK2DxHy+x/emaZosh6E+aY9JjdlCKOeawUqZFQtgOa85ZF2ygcz3lkdpj/M8qp6U7MR8Tmf+2
rM07crjLue64oUU5cbs8fZu22zPWE6cAq5pFxB7CxHT4J6hfJCzPGiSoBSrnriVvsc/pBpqPgDbH
Ai8OHJJqr/BsX6KupokI9XH5G1LzI9kMZK8Nj5NsfAmpmxiqw4DlwbnV+AC4vLFXmRGzRPCU2fYe
s4Cx9SypHC/2PUy2cQ2efWbsyEdomq7P8CeiUcjo5OuTZ+do3+mUAL2/3mlMBho/aGk9YFXg1a0I
tmzM+9VTV3O9ADL9RDPg4ZAcb49j2Nb8AyZRDmU2N6XhswyvewKKjwJ7eKXbw0AfOAVW5sFGwUoT
ZH1KQb3fKsvtVDwmfz4tMdRNF21tsqsjsB0OERRMZQ9K0TBaPfwgpLNMLwvxiYk3TADynIEtBCId
7rwl4WefneP+FDDU4utETKOb2ryB8WzpMi0NIbAQU+jMd9eE2lSDPILe/l/D6zWGBe7b0EJvK2NS
aq4wgqj/AFFf7fagm8+oeOejuXR2Kz0oAcFnKgM70Ei+K+t0L6TIhRQPBIeJYNLc/Ai4h5Z74usy
3kMHqmQTJdFYjpJ4awrTaiRCldI7EnzIV8yAbOx8RjdIIzjiO3NqWwDfZWl9Za8nvI4+/pets6CX
8t5303moUjvo3GFV8sWEsCK7Xm3sCR81pwN4hM/CbXRr0Fk+Ibdve4ukV/SKqTG3crhaVf+AARDj
QBZr+bcB6oD9zxDvHWy6zlvIGacL6zVS1vw8EwjYh2QP5XloftqEIf675bAI2axkMLyhaSozwy1M
HU7cKp9GO0wqfoLEhczbjpmzrGkDWczV9vrsbqos8j7eg5p4uFIA5oAyOl73ZZ0HS1hFjnVqWZLn
8adxnFeTQ97PLrGjjmTxYoF/XtOzoKlicEWeNKBeadV23t2NZeqxBBm+JDVC+ndHxNCvh6qEc8Qx
VEYGLCL3D5RIzIvcFNeD17zXPdMQbm9c/bRG3Bgsq8Wx5MKZMs6uvdgfQnoQ+/gcH2UYWIvSJzGl
+BD9glpTPeoZo6y+iY5iBdHwlbJSJJmQU3KhR9M2uT9Nv54R7YWdVCP8KurfsMRw5DNpePxtsfCr
dTh0s+XzmzYWIbHfcN2vBJ1cqWvN//1eTS5V2imIP1gaks99iRi2AA1kM8/4/cisPi+vywbTcEVm
0/AmyPutS3+/dnigquGcgFlcG3rm9OZZIUJiwC7EwgITopVVpDOqvfiyNjdsY8bRaPmQmJ3PVRKn
kyh/FbymWSXmxmKLtn69nMVwg1rZ50YgeDXkBENVksEWNZ4zeWHYZy6BGKaToZND/1UrzD02EbdT
phXqxxQipxNyD4YDwDUVZrq6PAoJgA6uHW4yi2JIKun9rQSdHkSybT7nw6EDfydsVPNIrqnQHR1I
oFXKU9gNgpS+QrqRp1nn3tTMBTm8Va+18+w4hu3sXeoKYb0NjPbs2MD4Vb++0ZkjGiWunXkaQS9c
UYTXhrjsOMdjLCkLnuiEWRgrLTTRpxP9NKljCQQxF1J94P1UChvAaj38Tkx+1Q7zTKy3CksFDFH4
XpzBXW/o5WEt5QyBTWEAJC8HT+88PKXHiORrxi7ZO3Ptq6QNIwCt5POavu0TrJ7uzeAgBTADKfi1
pMbdzKe3AxENEnnVolWf5kjgAqoUEzxPg0HqhmN4Y1C74an9f6FPFPmURAe2gP5q08s+DS8KYFov
WKdQ820yg/EiaxkKjpwMKZvPGytoArGn+xuDm+zPQHUtjF+Jqq+jUJBcsBWwGK9jK7L3o4fzr7/J
WKo9TBtOJMQXSxgX5SdZJNsOu++EmmICpAHQKu5Dbr6gD/3y0jYlyjsDRVMIH+3ft6LU37TiaClm
pD9cPzGRRJhscch9NmiNPsHjeDTgU+A3ZsDRl/1jUwp+DfZQqIG3FeRy0rDATLkBTZGHkZ60u/hz
Ru6AO4THJdAxm3g99YB5XUsMPob6hIyLd561h0hm9YHiH04046iUY9IJ4ALJw/nULpSYD8DpfaWR
nil6oVQw1SjBl1HMwQLlev2AO8CkwYsaJF9pqnM1mdn60olHMcUj14vj4TvQpKlMb00czkGiFLdh
o0e6oM9WM6AmUYEqPzv8PbaiBda2oCTdhGaFKqPVFITFzth3aSjU3yWCQ9xBY1s/EnaxPGckEHkC
tCQ+WZbsJirurzRugr5INInN5GRR1LQ9i7to638y7WPwUr3RWmLKyZHXfToWEYsczUFgFSwEB+c4
i43fULyz4XvzGqIOyf6MxATIcdY6fuyLu0HHhAUreUSSQf2yvmJya672dfb/3EKuFPKYRLd2ra5p
rGLzPiOpxZI91eWEE4YK6+hNQLB0deEYoy0+3vHqtK91RLIz1scDukHzJjyAi8c0cDLGf8LIUJZ7
j0y4eagV9lc4wPcGO05ybOnB0PNzZU/CIxLJt//5a+xlELP8Wvic20+ztw3q6XL5uCgyOgqXum2O
1dyENpfht27A9BouCgx+GUaPSzEG7HFps7tDpqWgeO51cvU+ibZnnaZkzd+hlWvH27NUe7IDh6H1
O1gtUwOQizmB9VXJVhf7L+fTpWZX5SDOLRM/bBMhHDgE0b3qBKtbErMMx5hauSxtKe/M5nMK6N+t
DNpqMoqtqtKKlDZrvbbbHSVIXf3GWdCHI5P9hRThHKEGkS5NwvPMaZUFtKvf815DrpPWfrKYhsu/
GcyFu03AcM1E3YnCmJxjKhyAm8RN/ijhmElOxVFt0P1+gpGlukcKRpqV2rykZqu/SeOIyPsQpeGl
iOIKhOM6dTbcdB5HSKiIID9G6NFFtzzZr9yj4aty8o7KCqVSZfpylmvQ/ZjfwSmy1th+BGOTfVLI
4f1q9/X1I1uaJzN61pRwmXaxwf5XSEAZX9YtdbNbePbxoDOYz5433Eb5H60Abvl4hccP52g/84Np
0fC30rJjSiy15Nkb4v+J5ziDde+sWxtoIBti4U1+JwFTbaan+mAUv1aCRqldL/467GqrcoBuIdcj
pv/EDy3mNnhaVrCrNL/zY5BaUFDdBYoAoJdnG/E6syBN2m+0mrididxSFTh9qXb6DVYPZ3C3G3uA
wlT/RnmeHlBCXA8HSDwbts3h+WrOZJoKO6Mlds63g34b8hmK6URZwpPgA2OmGoy5x/qNoHviOqRr
SJ9/fASTaTwJNn0TWV5UIjF/03m8DjKIC0sD7KOmW20c+4IZo6ZVMWw36t/xg4gQqshOxL0FACtn
WvX/cPcxZnO+pVujbcaRe1a4SSev62eXk87AwIdXL3ghhYO7S6zLw+7jurUuyu8nii5r/QQNFtdK
tkXOw01twXwfa++yrtR7uqphtdX/7SfQkpLj3ag1LDFE67jJ6vrEbS/T+o9KOkhTM+M7imHaQCvs
NQ9z/pl09wUz0d7zWomT8m4SrX4172tzY6bVXrhIB9uLYQruA8B/RopaSDTgAI3hztFoRCngPtce
WUO23aoYCNzzTja5mEwjXO42PSsUHF38x2YrAbf9aW8QCt96y7SbxiBEja0DjqyrfcuucNnSad0H
itnFl9ZuD6RIGCR0Yr2QvlvnEzenrWJhRosTTpdiCoBa1Lg89ck3bzxRLzbdmqXxuo1e6xCjyQa5
0Y2s83pdj6a1Ma8VrHGv6mzLVjORA5eRZXGAjvVAm5ZSCFSY8DfPbOh5eN8CM2gWFy+tkK+KLCai
1Z63qqpd/TNxra98lQ9PayW/a/QHe4gkf4J5E47swB5Qs2t5Pcz3rbwEtsDAzN7/H2iq1LJaK26G
saP5V/t4+CGNSJ9OTdj7L+CvX70nA/aUvwVqe5iBbwd7jlfiJMkXOgDLvMuQW7X3fZMAdlrwffac
yZUMqZjLHnQH7bbldBDLG4F9Mo9uy/pH+/+vDPSju0zpjS+Hc+42YUc+8doPpTQPW8XV7Wlf66FO
biPSOAmwbbVoKpVH68Xw8ImriHYqUk8POlv7N+4BwXwads2IcwiQT2r2UyjSk8NsWHYdPVSpUNKg
QahMhFtz8PfQ3CWgTibAoke8nQw8jGeDbO9GcNsftlmAYk+BLZyYefGmZZf08gNYpBaFtFN/exzy
y0DiU4OpP2ID73KVkFEWzoa+rK8DiW1QP2IIcOEv9KB1bAu/QtUeoLeY9MT/2gfkZ4UhaNQu0K/X
9vF1T1NdDfodvmqNHSW/XJYjSz+P2xMxenGyzShnPXoRa0RgVV0ltr82Uoeg9cWLLvsSFdX4eVeP
udu1v9wZgi4WtIP6qaFTzHQeRKXLl0v+q9xIegbjtYwyC7aFm5pdEZdfBw8YY3uU2SxjLisV9rvh
MZiBTd6d8RYAHDj+EuY9L8R9QkOwveirrBd8nwsg1yb6sUt8+woVsBCZNTlml1lv3bjdjg+8zLnw
fObSIIJyiLAdeso1UEo6AVdd/Ks/N1mrDmvC6yMZLgllBiTMKp6eRR6do+8gmwj6c48NsLxtAF1b
XUeGRNwgr5WMtCKDQzABHMTkznfZ6/xfwrK+0eHSMAqGJ5EulofLVefbou9KpdRJmC7nrgPr80Cj
r/3HiBwQlMm5Y7x1aIjNMiu1/swQGdh7gdr1pef08XL8TUC35IhLEAQPdcpPoK1h/xstPb3c3p6r
54pSSFy8+ZIxbmy9ApT3JkWleUzFRrEr6S/rNz0sZ1Q9rESSF9uR30STKvfz088Cu6wba7/hZyGf
H6q00XlY6b2Im7LxCQX132sN4BvsGDV9gN8LbmiuW3KUIl+YrGq7NM60Wn9t6a0GWMbb3qcbiBbK
Q3WESO/RqnuOa5nJpX4MS7EJzQhbJ2vKNkqy0ELIhA9U+d7x3yBoI3z65cgQPCEhonLNis0dDmV3
c91MI7ppm8+RFYGmCW8rO4sp/yzpAvDLzw7fTxvh8SniNCqEzVni2ojldA88E/I52vgamZqfji9P
juO+xTk4sdE51ANSTw65I+FohmUwAPHd9fCwGV2k26+kdaEyu+YOfF+8pOWOaEkrfOetufGOthla
kZSb3iya47I3LtEEihWapIXX5lmfkLIiX58dwpR1x4F9djlt8fP6iHbaJ7arumV3ChTcm+iay8jm
8gjqdNL0KUHNFYRGiFgXbxuq65NGmi49clsAhBpjbgaklQwsV+U+cQIsLoBoHeSBPywdMA0THubq
JzaedMdbHsEKnvq/10X36B8WQjHXW7hkzr6b/nNTu0JBnF901bSuydiIxAyknWNzjDmQiSiEPajH
Eg3l9FIpq0Dz3yIqm589xk8fVia3Izogz0tr6Saq/fsX+TEotgACOcMljI8nkga6RAmZuec0JEQY
eWtE9gmVUKHTFIvcVnpD75HqcLLYABXW1G/7gmJ5WCw8e08F1sESsqnN35dBfhkkpr1IfAE9RAi8
2mFqnUXn+1ZLoIv1Q6ZH2Im3VDY7lnyOIwVE5t7089mVXAo8nYQezsicmwuNIXpfuyZagzqWvo6T
rKWGKn0MRmosI3Kx5McUjfNdFyHRtabpjaNozPAIw7CgyRRcMa8VgLJ93BYcK/Zku0Xo45XKGZMr
XKsWzyJbHCSedXAlxzcklBe1po8ntSzAoBl9ElFB4Wop0kXUKE+pim+vlBnM0f5lDgumIC7i/aUI
6jlDI2QK0mvo4Mc+sDdY6nDy3Gg4va10zWFAjBp5KUs7h9OGzYiMjvNH9quF5hEAmBWEdZlyoY7E
m55nZKxx99FBefVZ19Aqi8Skw0K6/Y5aTw3Pto37m3TSDok5bO/Vf2RekmbCxr86zb824QEfhpWM
YGTxS7vHIcyJ48qt0Ae/9tsApmsXKAf5ZWSZEa+lBi522SNL06sX1NXOfa2wu10+ONcA9PfHjkw0
2q9D2te1FRf4VNoJb7uvfvu/mr3wF2Nm5dDok9UIN5M6gOi1H+UIPlZNQPwW8x4i3NGYmlQqPl7R
r+FL3LqyadfewBkwePNlzFVHEWj11V5vkzoGYGFW+HUzAI0wzP6CLewx3w848SmHMi8artWAF8gN
oCzldaQQX4Zlj5wq4j2fk0XWCyk/6WGeu7Cihf02wtao6BHqVEcTPSs6X9dprCcdA/7SRjj6WVbS
UpRFthE7QSm5aUWk2MOr2ADBZl1ssxBe0EqAsd8404oAbwoGkcxAy4jfhgsOk1KidOHS5+9WaAhY
ik5CX9V9naGsHOT+1nCNxzydlt/k5C+P13sdCNdZvyvbWXW+KXDRkXRBvgd1mQ80WneeCAMdGNpX
PFOByrhsHgrZZOrIIoTUBf5Lp/W/8/NHJSW/3CefvTRIcIbW7I3xjNa7msLgUIR5go8c3jdJN/yA
YZy12A9LfI13mFbXWUtaVIZskDf0WC8LyFnX8//zo+1dNG2n1/6+uWuLGD7irTxVBhoYVfdcB2qn
n3P+zSQiriNvve84a78N78+h0x+4mXDLfSFw9NLws384wwyKbZWHjW8t2+5wAUhaw98DuYR+PUIr
jeENiaSse8de82Rfcl7tZNi9mU6GUyIhxLGO9ObK/128Ywr8o3ooqSRJ2Okrz/iSgPTyKmBKMBj8
6RN7GcRRppQPQTc5ISOdVS6AWm8/51ZKmsGQBFgFjzmsPpkFDYYahgCGR1uMV07hP9Ped40SedTu
YoFQLlB0/w65cjh2ShWqY9GZojIHghPQuBnwiCeKBVvEqQh+3bUlTJbnNnAWnhvaJQe5PtcNGfj2
QbnvfI/KMfThiXf7g4deoZhnGxyWGOZkeysea6kpjF46zjEIuRr4WdMxqKAvywcZMmT3XCvy1kbg
JIT9Y5notr15pwloAsrrkfyxxC6YilKKwwM/RSKJJ5B3kSn2cb8xVeloYOhbggXj4ImMrV2kwx/u
SjHZdv/2u2Af7Wv8onahA2ZR/ju8UDUhoPosY0SR9KoEqyiyppr6bVckrqqYd2ytt1nSeUIjUflv
6aYcx8oZ4jk+e7lnd6J3A4W+JxCPx8J/jkXctos51yY6R6i6TeSKMqtI5w0Dn3KXR8RGdoIOdO8t
21GMB4uHUeYJA1YNjtBt890X4OCx1LHp9iUr5h5zjlas++vsqa466PzuW/Rb37Dzhyvz+GmQ4DDi
3Hb5j1Ln4JRyri0eLM/29wPsSle27o1+1h+TYVpb7k75i6sV5A2KSMPqMU/Xtb+slw0K3jeL/46p
b2/xgsHmT08SN9TEsoeZCyQtIDvvkIhqYLwZlDtwUaBi2m0ZbHZJhlgwHFbZmn+hDoa8z7NM41xC
PZ+PNnvA7Y6hUfnCTjaCdRIVU9PzBKVnwRHF2h2Q5EXL/Fvq/1tgsN4vvQdHnNANv4UbNPYRIy0o
aAVoXcUIHZzO4MUHqToZcholcn7Koi9WVuL1own6MmfV4/bSDqnWoNkjcZGNbcfPLLk3REoKoqwO
l+SeOTTivjqup+UpzxoPCRqpZDkh1lG88kYFban8ynRkA0nCTexyOhr8xUnqWbkkoO8+G+WazwGS
DXeP/pAMVXtwiIuYSJVSZTxtUfBQsDt9SaVBIE1kZRGbVqwNRWLrr/GHaqBhjIGTOKHxVwi55nsk
6zJ7R5v0lo6ALzEuL1/0IHTNrURbHL3ntS0EWnDKVBmnlLD9ic013oNU+gnRIcW41W8gmWKqHezH
lDR9rscX7V8cuu8ysOHyNaznjQXyJFHQyvt1sJeylNkn+4XOtuXhkXuEFFxHi+L5yt7o9WdUVqJ1
zNcq3N3uNx5YJ7AbHVA0OlH88KaGAs8SeVyH1arO0CFDO/uLstaL7fkXgv9eYvWC7WIwEWCS+uJ3
QZeOpFu1AQOsEFtIUykleqU+suG1PSSZX9S7jz/Ch5k6lry6BfyKANbBAwQdQ/6cb4URz/RK2bxI
gYxDyxvAQ42AP1EE2DOWUV4n2KCHGshNAlV4nHIucbCrREluJfkX/7hAwzClv6DQhFgiziiHG7Dt
Qbn36B5RHE0+7V1+5WpHeBPHXZJGW8I5Jt2QuyM0lwfWfaBowMtyC9UOPiq7T+52AW2tEt3g0rsu
kAHVPUcfcMb+FYKkOXyAfq5ftzzyYm96jZAwXK9V53ofX43grmcjKHVixbA6JPUaoGDHuVh7PAVt
W3cw867156UXncrD5h6Ii6C6xcCMnw98Mj8Z/GvBVxzjt5BxRz2NZzU6Qxtpx6/SkfagxWb0qt1B
Kox/f2rY06cEEnxwRp4+0DYAy4ioQa4zaDz3JGsOZs56t9M0ZG6qR1QpFGOBLnptQGL+Y9fS7QMN
NDrO5QMJ74FeP2D6emJAngvPUMfJ3Z5542rxhdpbcqVHeYH+CBvkcDZvB4S202fBCg/7/DlvvfvN
NUbFRmlCwNFVzzospXgc9bAoUelDiX1kNq+o/65pNh6e7Vn4NKpo5kjDtdJUqzh3dLlD2rOfN7Dd
3s/pUJJeWgQSBuqUBdw0yxDjQbsxuhDevFfU0lnk8AklG7r53zWxsbKGeEDrA4trZALUPg5DWiT1
kzml0m9hej9s9n3CjqbJGu1u9gF8Nk0OLTgwtWx1MhV/D60INqzXxFsz2RNH2J0SgppLCmu0lKI+
fgg6h8c2yuBVyYrCMmAUDIUWonYUQXiZPq693Httdm7AQLBxpj7inOIryqOHAdSKO5JKVrjH4WHf
A6MWQ3t0ktGG5aBrny23iDKaHUCm00WNNGK2ItHS2CrAZ+VMe+V++A3nT0FrGXYrlrS4SE7ecU3d
V3Fw3kwic98lp/CUfIW6dC1zPVnxTANuV1HVYVlnT7oxcxS4et9IrO7v8lb3W9969HNuLmJT42uS
0w6esXIkQkC9m2dTuA6pzotj8HtWk7VeJKx3VA05lByfbF6HV/vIsNqXhcxI2LdYaZw6qfIX3KPf
s7JAbyYwn8IHJCvx9UF0tYlIGiic78YqPH2juif3vBTkHEC3OMx3JSzDEB4yfUEfWKeHeHc+ew9+
/zm667jUzwr2KO1vN+SrTZXMgfsuGbwexrnoHymFnMHKEzfcFL4IkJRVnNPgOReacBmuvuPu+C5u
XfJMUXxRouIqwGS6657+b7HLAwm5W34vZLpXShSeP9TOamORGEKbEvKzJhnLyhpOaJZoGPU/ItnY
xN+CgG869m0vpREvgaNbKldEzqul6IX3CWYyfAT3/pfiQyme6RPScdH3R+McBxIapFIsx6CX0r+R
K0cDy9hNsVWFcFK+8NdwRhuwTcYLgCmM+DFWe4Nrjw6uXfyha+9hAG0yMNrh74Jvp5VqyWyAwfo1
fRnlsH6o3cfETREgABqlpgzuMVUKc1pT/50g+v0kYYiN1yoPpxXRz3Q/Da1Ygnuhee3GA2l7SByI
Slbx1sU2pFk5epuVl81FvoCtqQZQSJAQImkP4NhuoBPK2L77LmD3A2saJxhrsD9gOhbvlbHIKLko
FXGksoMV0wVgRkls9Gh/fJXsbAfFlmWRIXBiYk6x3u35c5zloDFFw8nrZouvN86ZwbA8F8+tTEUD
cpFt/PqqZaxIacF0NL81FZIyf73kAalS+6ezdfc8PL++zPUGo1nz94BQ+M2NJ7cfPzb5w8dwDvKC
rjZRFBRpmXiei10u6EQJ4KY7Y67vNNGDdYNZNjvaIWHDx78tO/KGNE86aHewugBuXgAjONTDPdNW
gXJ/1LghIyEzf0u+uyq/PX4dv/PI/pQJLsLJVWaQ8MOtuCfT3zLFhmMYWQt29RIED5inQunw8Lhc
Jy/kBg078+SYwU8od6GDCVC2+wx3NiZ2YjZ+sqT4vICe0S2eQpKns2xlebkp+ShmC0AiiuUGL7p5
XUEVxGYUsL9FsLwE0qeI5bvd7AZ1dO3qkHIBGNVBlDMfKMoyN7ii1OTt4qBQVu4Gy26Wyi/vUNKp
0V3hr7sIVnRV+I3KJB4KFFu578pF/mLXC65WznY7vVH1ZgkbvXbNiNUGHHo5FvVNwzw7yJvKJDWa
WfMRGt+G0ZWoqWhDda6IPsSVo8hQkaxZqee+vjAzUDg3mPe7btfJtyvo9u1YusKeYvkhX02GQ2IX
PWle0HrykYmHtI/T44GaS85Amun1etsuih7QaYkLNcoOF0Qgt3UevWSqlr9k8V/XMVH3NKRTBltk
rvuFHOKO7NtMhPRI+b5uGyA6HZVXvB+rPnjW+CLuStmsGtfBSUyjBXnXxZ2JMGV4CEJfYb3q0rmv
L9LmO2Gk/whvBTKPcEcO8uSAiEC+Ir/N/aPQdUEuiltDkgFNUtULFbnHCGlnCl64ChW0BM8Hcg0p
nx5p6qe6eCID/UAWkodjgsip/SPrUNcpeGMjLPFmf8WAMszefRYSpCLMmsns08jl8rp6i+87ENuQ
/pdx8JumkWtK7kkohzSKsfAfW6MdGHIaM5E1cnSSAPJq7AaH8jGXkMfijnpyEzt995fQ2bGAw6WZ
2ehwAn5k8MEx4zZWfLPxBGNFci8zHcRwd9V/AnMBT52f7XxIPDbojkJE7Qbk7LMBoqF+obkbyAa7
BQgTj0TCUD2RIOhzpvuJOZUZutp8mOw+Puz+zZkcpjYIqPM3GXfSenHUA78c4dzv0HQrl7CGRGru
ODuSMhfbFs0x4vChgc/0p2tP8SoSAlSShRlNmp552IstYhyecXtvA/W/oU4x3SbRpwz/ihj6HicP
Uu3sCzQp8/eqP1LULwkrVQxclBHta9vBZHmym8v8J8i0w42YkUm6hpYQYHSn/Vu2fhvelSBxogYN
5q+cs2Co3L35uRdKjOOO5uT031kKp3tiZrDyO2F4WKcz2z20RrSVcXGbkaGz01dc2VFr+wwMVd2r
eYNnDb6J1LInxi+CwRyupzQ3jNcXElclYDIccjV16kUCH3IkiJa7Sz+LOtI/b/7cJVSUfTQHCI8h
2H7d9dFvP5fzSaSXWIFqOItvaZnaQGo/OshDDKDSfhpgIhQL476qt75zi65SyT8aFedaYPU/tT6L
JQns1tLQYUP6+kdcqyHF4DBmQCPTHKVGHbyQp0jY1+lxMNnXT6NcajID9lS12UTS3savyalEE6xR
VOVW0Lnz+O71iCJi12TN1Cg47RLG5DOPn3eDzPUXEP43VINnDuYuSMQDz5fDDmhonQ2xsmT37Hh2
kuq/ll+kjZXY+wcujgpFr9uzYwRTSodAGGULN79h98h7qc/wv1KOBpSFFNxS3A5gcmSt3S0CAyCi
uUQNAM4vVCxnwefU0c3NqXkCSVdueA6ptG2OdVsJU0Fv93WnzxdhHBAc3B3zDFQ6c/RB+JW/8hcv
mKRe64JHYcBuRkdCdkptfPjUSlcQUhblojCs0WGEhzeuYIzIw4rFOPhG4AGZdA2CitvYrJD1re1z
xxNDHD83cJJBfIFittFPceKm6xvAI9rXUoXFMk2aazBn/5j++gNmO+qCbkH8LMJfZd4xti7pN9Pd
Ph546YyvvZY5IScDhbuaYdnZq+kqmROdAMX98CvwyiyJs7xSqTPR7hUfPWMMj5yyv1UXkJpQHmo2
2QfTJvm09JJU2vBhFmDxYA68IahwU1+xyH6vVm2c1GOs86qL8WSNPfebtgU72TlFN1QCBibeoxZR
4Tb3smxLcAqkwf+xOmkN3+5wNPhi4/u2X6cX+SGBO3kg9eViKc4mD6j+znZ70uxVYpS0jWSWvWds
gPayIACAW6vy2wlM39GhrydpI4D9vbTUr4G6kD3CQbrqBOC7ujzXbsCL39JkKdO3FZ+zYC0LzS3w
SeVNjlSEh2mBwtjR83r8k7TVyNXq2494HK47O2GgcRCUo7YDGzBJBWVhqycT9Wwfi/TmNdue2Yld
XNhdpdKYvugxuY6SmKs9/WBl+NriidNhr1bVyTFhqaNwwpN9Dmf0MBMG6e+gdEO9kq5C7j46TZZj
gY8cBM+AaM4q8+E7ONmKr8mSFRoHy577onPLw5xSKwrSc/F6UbvXJGe47f9y5uunbhKne+JLTa52
1ZZz+VXAwgrbye+ZkM6pE9g3wil2iDWghSmShKIRqzEeujELfwxT5JKeHiM6lrf6Rk6lYSCBvsOk
0TECInTiXj74h9DWCsSrwakLe9bUoJ+4Vr+O1zwC9KZ5UAlKkR/Ux8414CxBRkaDjuTdfmM7zOec
3HouXLCuzvenfRSe5h6zmpnUv1scg/X6VSDLmfGxV31aG97JtCfyYuC+jOns3zPdAtTBTaGP1YEu
4KmG/varePDCc17YTuCzh6UM3vuewvn2/i8erftubKayZ5chtp4DEIE3zcEEM6j8O2PSXOxydg2s
mM88sXCjKrhu66R5+vAyE0khcT8xh6IQkYVwIp/crK4QLrvQZSO6N2waMVl93ZjyG8wIgVIAj70b
Tz5O6c/1Lnq+5ctUVfwUzyyZ4JYw3jTDDcGr/G82S5bveZ+PH72a6Q/r3/WFuwrIFrhqjtDvyxbZ
7t55Dl2zsbFkom2ICjKoNTYUgH6SsY2nw0l6FoY8O6wv1DY3g2SV/n2DsIgLdqFN4Z3yEwwCiYJg
w9a/qfC9a3SqaPya56aSi65KwDcsO2uUSymPNCNSHmM8Ard88d6rq50F3BgstMKmEEEi9dRKoOv8
Xr7K74G6vHmmBBWwwhcZSIvuEQYzF9NmFK+pgDkysBMo/+opTRQcsegc6vHOuCmr+xJoWlyGwa3d
e18i6eT4oEgDzVkQSoi3KgIS1M0vQN8TbbflpI8I3SfP9ukJS9SgG8pWbPdaf5HKg8hF9xycy5Dx
zVEM3cdt8U+XMyqg+7OC9D0axIITKWiTbnDmfscldrasssyY4ZrqwEj0/VZ+R/mSTHNVGgO2dheu
7cxjl5JruVI7Sb9vk8SMjisiyuwLn6A8uGN6Atn5cL8fzGj07VRhTW9ulRqffouYdhVzUlxbCDmp
NCfta+wrCvOdgr2M0cvw0PCUn5FhDx4MiaQK9Fk8/BqzjdB/vr17vFo/2d3YSbIuSYOVNqJhkxfP
aOIlodXmsM1OFt9xbp62pzfrAGhChBRPKRWOZE5R6lAgDNhirXfZHHknsvxK3d7v9xx/bOwdigKQ
Cpih2weDLcf7oGGRQ3KXWXDdjKaTR/KBYAN4MrM7e85+hc1kqjVCGqOZEjQLn05F4O8WKyi6taBB
kGcXPFrEC2hZJLBdu4iV2h6IDtv+5dtvSANlhoFjiAjyYNnpYuHhCFmk22g2ryUnEl7maFgVJokK
3owPMawWoFkcCs5TE8MxOz8obftJ1P1NuPEpVY3YCDBRIZm9sc8/T2YF6AjmJ97o1e7EOtBfFvPF
8wypiZ7kOcjt/80pWTUClSOKMpYkGWFBHTQqxa0qXEb+z78zOzwAPss5Tfp8INSLfpqRTuaJS58s
KTWPKRyEAdtpQui+le5fCQZfTW9H0XE7oAa9GWRm29MwCHcLj19wqKQ/tXmTuATm+EzG62A2jcdB
PwW0mxSxlmRnfo1THFDTFm/I94gMl26+an3aUN4cKRYw6x7glCU6HnbIeAGVAizq9GqK5KfJPZJ/
gaIXFRmUkF1NrkkL5YM5377uKDP+tA9IXUY9thaeeogB1v5YxneOi1JT6sD0xTXSf83muzCO5SgH
XDklxh2UlwipwR12KEkHxyQ5AljPrpAQwhP24N28np+fBrJmV/dVyEX8kljiec1mc6OMXtGVOngv
HPcubdYIEq5kLyzc/Og6pVkIbVkXXz55bK7jmRp4pqUu9aEPik7+1RqECZYZwvDwPIXq5OvJtusE
CLC5U6xKlZpok8LEw62Yj6vvb0sNctzXV2pIrExHLI1c8JE3MAGjjwxnC5AINmXHXgI4+2bINzCK
Y1dZe9igIrLK6i9Ry3CdkQjFTOsAlOIas5halc9W50iUFb5/sNeba0VKKK9HDVsY6UDVPO7XHDkj
aMVbqEv2g7eqwjiTZj/kD/QX4ouVkEZNOyTiSllLDoBy1bt1nL9FiQLHhlQUy+WISifeAtTwOWMK
qBayM3BeWKrvIsC/Yx6WhP8++FCjJaaBK70jCDiqn7IspxVx2VfqwUoEjVtj7IWqz0qRV6SpCgGQ
tgwwSSz4FJYxo0+b6It2APGs2Xbwd7Nk7k4upU6M8RL1JWdJ0iYiCj9n6+6eAs0A+O37JDubAkev
+GSR72eJVv0ODukdxN9mMljiVrbucVcQQJHLMIECKeA7rrAuX0j6R7268V8o7A65oq4pZIOWVm3E
OeVskIWAuS1Zdw6hBBejvz9EiqnjtT1DgreI8NWslvUoBCRSEmuxg6utFa7kXfxtxwbCDDLkrcvX
2f8YNgg8oUEcYsG8dUvKTaWQgSqjnxtTKdoPVqTzAlwtyJwsNkO9bkwqRkKkU1yEZLIHjYsxavTd
NLC563yj+iUkKaNmvMVzlwofBAbQ5EEK3vXEcmDsoHjSy3yPkMiftq2cyO4EgDbEQXBbGry5cf58
9tbDcOkbpbEzhfrZvGBf+bcg5NVpjwRB+i8b+wCkv04VQmXL+pKAEFSTgRZ4hOIFNaz9t3VjTyUz
jbZlBXKY8GBvsyvr+mFXGvbfFeuwoHKFa52q78e3Sd15ssomFnXfdxT4mgJFzu4q/P9VRHGM+f7/
61flkoxRiax+L0lZhMHYwRYdYjeZSGh6wnN6C/67kuDH9H7ynsoniUpWb7JyHuGgUqPYSDlBDNZA
Vb5BN6inzc4i4XixhjlTfB9rutAc1bjXNStepyMe5XkLA8Kelcpp+dn7hjpFKVFIa8RTutNdRTrH
iM35lnzJFO8zWDSBzDCAHtq4XqUuIM/c43VfRcFx7fg76KhgO/HLI+SET6RlM5KR5Za1t5k2SSTH
PPvYcDFTwukiMubaUEkrlN4qN4NOadwA3eGWARZdpfX+zB0xWjAmlZeq6MzC84f5MW2G43KqAvMc
p61DAg2cly9muJY7mea2oFgEn0ZWfvisp36RZKpH6Lj0yucHIfdtDO0KzrYe0My9gxiIR1gXoK9j
rShG4cIjmTkoTsIKMuGWok3oR0g6d96ub+Jf8lL9qtMP/Lzjui0TvWEnoeBvlPYKxUgL4K/2dhJ1
vLaW9/dzOcUORmeUcXvzj7Cu4PVGXEDNMNgTJWDqOXqsS6AKn0WFbvb4oIdCpgrpTn/nQp2r0m1h
+HtYsT9U97wfZv3OuzQtnFPssMYmPjK6Sqr0pcOGrDXeo2CDruAx8WjjfiCL8XfUxTb5K1701nbw
r1xKurkNRwQBlPTpjSpQHmA/1NI1mBzm9DLeIRK+CUNVlnvh5nmnLv/BLm3z7yq13Qd1wyEwrOiK
Gi7eztvls9tjAy2CkQCyIGxqsNHm4yC6G8qnn+DvwbvmKCr3tdSrFvYuZwqhBLnGWxE0CA2N4AQU
SmQ5JnC+xn2tAzsfK8NZx3nV+KIof61ysd5XA3b7o8AcbmAEB8cp5tj7hK0KHui6eFjlvhQYKaWH
oq72U6x7C8Iru7jv3oXjUe0X78Z9LLagKHr7uGV94RjKZKkfMlegBfiTAr8OpS6S/KXTEuKM5wsZ
QldCoSl013Uh1MmJdeIDf5ZPUxHy8EUJUgcqWAeRjRKun5K65kwv6iqRQJ20FL+gniCmzuqSVAhs
RjDKLEP13TS/ZhH981TCLdAbM8ogCoE7lQB6C0D5ztwp5RToKFhSTHkvLU9LETIfj+Q3ZyIDynQU
dSwoKcUEpX2TleZ1exElCdIABvw+dfkmfrtpoSoCer3Yxhlj3ep/e1elllP4eoJHTeFoM5NKaJOo
qAuD1MY+ChMT/5UlaCpgsgM9jG1OtVlYkO8hKrTMIwZOu6VSXL9faMzsq4gDry6bSgGnLWpZXjJB
QXF8LrGQQ7FVeWwVNBqEcAHmu7vqfxbQ+jPzbubfiMcJSqtOzPsCJtgBA1TAqkPqR4FG6dVhXuVJ
XPzKh2WYiocKwa3rNPEojsrd+PX3YMQBMrHiGKvWf8lvKvax3uPLwMQJZeywfLklkhAH38PA0+da
fx8mdG8pqP+dVXXI9XFyfGhxrZeJQtJqYGYFXRW3a40bruhbYu7LXD53GlfYveboPtqR9sxFwOfl
GkvS529wO1QgZru+VI9CJZ/J7rcH5tShm1gdlwCpqAq1BIiMtVHY+N1uOPMrRc+cWp2Ln4YKkguX
os82dUdsJSEokTk8yQ21DehOkcSxvcM6b6os35ajfmzpBJdgIUjqhjd/0ZtjZC30622ZkBetMuuT
5EW4euEsm8E1wFPDU5qjngYNNeNuWIerZ/psh2FDtwmNkJClLcujyqIfkPX09vn78drbrLQMKgZK
sOrh+gOhQwOjRsNLZ+waKaqYN1ZW/w2gxjC1c8lM7aLK8SzfBxX2z0ItoaqaS0TSPh5aS9dD4tjo
SyIAiJv+dOE8mcvwlKBiskOoH/6+NpF5MufU5n8vG11BfaZwSPqESqDc5gjW+gUazDXkXory1M4j
CmMbviGZ255nncOXPIQlfZnRKXvqzWccdcNpD9I1eKST0ZInPoRnevzcde7RMRGapJWIzRZ+5qyo
4dmaZa5fGcL0t31ng2MTzKeJz7t5wmPBHN0mOoMZ+9Lf/rviz4dtvX2l7+1BLNKxvN1mxbzz+bLO
EKAYntCLCQQ9XO6G6GP0BkFxprVWi9vEaHA1Bg8c2u9HMw3eSuB9uJtbI1CV+lUewEXdGvrF6h8+
pvCcnB2ImCL8+f1A9pqpzk9j24JVKvV3bfXeGG4r8zcNNCGn9hH6xqgXEd4HzMfgm3EmG2k2BZYA
1LBPoMddpvNlOFqZ5LO4zs28Ufr9qy0t+fd41VAlOga3K04eFdXlbMqstVi6BtmrdDcCUPnxp1gE
plLxS+3U/HKh9mOQ/Z+WJG0iX8DB5vD3k0Whz9Xu4eDFK96WBKDp3oNolhdp0HlFwiW37l9HFjsE
/wG9+vm3YJppdFZMTDCS8l6TScmVzkfKzVd3FkvxQhe9L8osCgvt4s4q8feetq++ZfL09y1Trxui
/FEX1rOTBb7wnKMkEYkM53iDdSWXgIF7Z+fH5uHhozbaK2DsukniUg9mk42Uqe2V0WrVVzC/2dF8
H/INCZCzezeXTnXtroZebnibZ387/cSXxy7wtjEJYCw352JPOa290whA7fFmkn26tT4dUZP95pAI
W7a6XiaqvWAfPs+gyFZMn++fS0wuDwigUH+xUBiYR+EKIKJSPQbzcGpPk31+0OOIaXEnpK/QyepS
PzQAWxM0zQ3kaR/UN68ZKu6F9/Baoj+GR1HJuZNJYTLVwJLdnBbG3nMohNT3RD0cwVxt1o1mwJhB
uxTiZKNlooEQUAGp6GXbhKOdrXdk9MvCdALHqu0TdbCQuEFdvmn/Ci3Tu7UD6Y/+ezgKYb/9snYx
oqwxNEE3RQDZaJa14o5sWqTuSjv24oSZgBEPjj87zsveGBEYBdM+1ibVEGwT9aNI31IlkKxx0y1h
3yUCGBaYTYFoK3zcUXw8lr/E/8g03UN3OgZGyoclv5iZLx9ZQcYKQBKnV8dhKEfG84y8Wn7Wf82h
ES0nTfa8ohuT1uNLp6Ndf2sAs9RTi1GbzA12KRn2sAHwH8nj8ZSNjmmujUDDUTLI9eqeNomi5hlG
i8uqrIGTb4TMenOBLJ2fi1mOFCv3cwkRVLtNHklHiM6XAuuzlHb4/rS5Co/YH1Q41OLL/EM7i32+
peiGedLnaPKWml8JfyDI1wW6tvDnrAxOEGPhC4ayiqRuz7w+3a+D+AI4/vv8c1ecRpD2sUqEC+uK
DYP985Krp8wQiRntjl5OXEGdIAJcyqP3aRN6BZwlF32ZjiOBzof6HQ+AI/5a4x9bEpdo1WvzHXZ2
2WNpnQn+Wv79/nRxjnxh1KtQXcVUhlji5ZQLRkFvBDIhhcuPrNtcfFKglO1hI43gUFEqla9M7R9t
W3lyFU6yLwtwHq7sgtTapW08avvvnqyR17oEH2ThlhUpup0ZApWE9teNNX4Pv84lrskD0fgNJE5G
g+lGVUVgEv/fVXhW1FzQqKpTMxEShcGs7C7gaSygG8v29U5DolinwfIazrFwbrO8rWGELOcDTcDL
/Xmnn2LMIr64628yRtedhIWVy7IPqWqJpFh0nSioWWtgnmVR5/pU9B5rqWi8zJkndJ4LONx+aG/P
qvpHFASrsMFqU96kGuonZJHzVE3GH4accROh3cmQ66hO5SUPoctkYSlKPxZoH0YDXpxa/KuWeC8L
SQfI/OKY+Fl4+FH/ayUviKxkXXa0BfkruQoNogtm1JrvpYHr+uYVMkHG9pCfNqwMRM7gxA/TZFAy
2tcovbyWLk+R33J/2BUSYvjNdjKPL1mKR+iVQKcHSbyjIQAr5Hv24PWW5VGxYGVzshco0xybLAWw
MKgAYIti2M9ohRrzlc5N5kOV6z95/6KwZc8huPCoNPcU0XdyBss5amsFeY2AHTCVXfTwVyt0n50n
Ih8mejph/+agZn1XQK4vx7mDgCdzsECJhgh+cyFE4xwPyrC0ALXVClCPVN2Sjs43PVoiLCREGZM0
SaWAQfr82QWQKR5GxTMz0Wq0BtKfNitKNDgacQ8W18K2hNnH1m2zNLIudsZRzvVy97edCvh6VlzP
mzVMnsiCKYdG+v+Rl5few695pMe//H6tN7gYKntfcElL2Rn4LwuUJIHggKZXS7Hhuh7CpFmPK/OX
F9Bgaanm3yeI2eB9T6I5iios8f1XlZpmAX2IfX+zJFUUgHd7HD3wOrGcN8YZwnn2CSYnqZH3GQOR
CXzmHsB4j52PFuaziMkszgMS6s0A6Qp3hZ8IX5L8C0oEA59KRBMxaof1HveNVzc5U0GW1j07E3dX
DXIiy0Ese8OUTPcEbc5dSqviSAB51WT63X5ivNLjCRzWyxWvWmiANH3rTwQW2+T7SzJROXJZFc+B
R79naC3TIC3DyebKI+kpQorTy04J88OVelAYgdp1H9wT01/VYeZlYSApuATllbOPZwqv3JhcODWu
4IxEpZnw560UMWmy0XaNJh1W5CAicfRfh3BAZEuUzUEJnDl8whrYTSwqWWApy+WJVN/GlfikNMQS
KXsBD6dEFfHazFa1AkU+6P6bDZXkiY5pxxqfRlvjHhqzOnz4cVwFhBKmpknNHWOIcvahI3tIXxZ9
WEUBDgAJssWpuBUdzSw176uHE9j7vfStrVEu6sSC4J2I4nNZqXyMSZtHFdBMvy86F071oM4sN0V1
gdaqD44cNx6laLfUqvRJn30TjxT/GiiXIZUsPsmZ7WiZpKN31JA3eQGdKRZfD+Mgq+kCfV0zhOSx
TjCbHJS0KPFJZHAj3FBGA7vwNT5CkYnpTt25tpUfYpiEMHlovz/m2rMIkZFfLmams64MT/LDBtHa
rpz/v9MMkMyNBH9IMiB5FdbN9r4GEoXPeu4zi9kJuD6hFXHC2Nq8IT8UrC4Wl0Tu1c/2s9qG6MKC
tKijv2ab8Uw8JNqc4odPlH3Mg3RHoKCXcSBl5JyFBwI4Br3xTmOAs6wUmJDuSd5CFglnsMSbwsG+
LQgxBIo/rPH92HvIsVumnFtoxG4gKQpl4pwb/XRDZ5wlSKBueMCE9pC4t4KJZNEMh+Bn+wyKX68j
MHCYTYKL4QCHhgecy1hxfFdBWDp61LjyKsc7Ewss9wMMDX0notG5syd1To+Uap5cQYPK0i9XjKiG
iq0ItT810QLG6HdL6PWZIJ6ycyCPAIpbitOcNWw3Pz0za0ydz88WzDu0Uj3TF1aeJlVYx/IljpCM
0DX/1KQ1cOegR0G0IE0Ndcw3YyNM9DndqOBRkP6su+X2hOk+NQACObd84Hintq5A/BTC8e6wjcgJ
nef2ZrRGpksJ/hoGxeh9s8HDEQyk49XSIGhQKI0Xn55dJQdNbIBAn6fLZKDW411VCKOtd4TAUi8C
guo3+7Z1gHrPucZuzMYkvC4TSlzsfBqAfRKbJthtjTc8qnyZFKXvuMg9b4NCZTicAl3Q+eucRyBn
aOTqBRV0ABAH7svorjoX+mpaGvJn19+icJ8gdO6+0MqMR/uY9TYQ4txwMrswuycVCicGpUqHxYHV
C5o5v2GMkEpXbc6QJTQgxYFIVmVXws2A+bsYFlpfAD5z7jBzCwybyzavKVoyJx4lS7aWFOak/9Dc
FT2Nl+e+VJLukb7E4cktEraVsRnOyqGxb2ATpCNuRkLSwY2jkQVST69YX9j8VqX3yY2ky5mfVX7l
g0c1dX4qfn59ETnghsMXonGdueDGiHpyMvbSUXa1piM3/PxOSOdrLyFfYkJx5ByfVel9erJn2R3R
a83Y4cNt86b2NBsPnoELi4T55OYvqIckKdzFezVNbhlkkrXoUnOSIHBogQLioBYojEnjMDssQL/p
/NGTua8AwPlnYUykZgm3RJVaHvlPfkrynBKtuw4C6trz+4S3kH52qrw0NiGriYDbbnNuvMCzQLVC
kxpp4NzIR767SPJcB8+JSipxPKwb4qcGxM/xoatB/DSu8nLlQfMKNGj3F3HDL6xir4MZz+pAgieB
5lO+k/4v0jn9c9HzjBvwEF8Fls3YgwmZRHGkPSd2+Gc/Lh/2Pn1sY1f2NIOW9Y9UZff2uPdghvsU
hMT2aY98zzTOmsfE31cpUEBEjlBhMWZg84oWFIyJaWkr85VmZBpyjvA/RG9WDETfds+e9xN83yRV
OoqHrvshqOsKfOIx2B1RwR+lmD6UgYqxxs6DiICAAs0RnEKMdC5Iy7SzNi/HBZSdSthcv3sGBBVF
WDusYaNKCLy14nt1FKQ1HXBBcjLGCUApyP2hM2iTjn/xgHLXCY3SE5NqIFfU4tFOpFzHhLOuWjW4
CSmmBKG0ebxMnoHkUMMmyC65GfCNLLvVbrhT/H9Ify9eGQTVc/DZz1DabUV6KaQRC+U2gyvHjgXM
nAFcO2RayJl1q4dXw9iRunvcB2mEc6lZIg8jcTu0Rz29rJVdkRTn2zBv3zdxRWvCi8+aUsDKzqT1
7MwjymSXg7w+RMsyhLWRz4CHDfKZa51QJMEWe52fPI6ce3L+FfC3LWOviolj4z4pRo83lwx0U+LH
19vlsTd7K5A9Qmc7bljrchx+GB9noxaJBumdjSa6sf4yQq0+2UkIuKMOoEHP8mfsSwsroWWGo1nX
k7sUn0u7FGUqv+an1tTE3PKTeIOPJsRpYNX0MKwiuCdJpDKHqRR6Z8V5Ix44H78cj4lkMpv8q20K
iQjwbCqhqMtegH/xjE87kgaur+FzcTexrS+roooGqTsUkjxEJ/VdzJc01JeYnwGPM9o3fW+gCtqf
CDLnmfz6DiNBtPovQMi/U4L+1cnzWHRBJJucOuuTHIXxcHeVM6Wvrm9fVIaK98uBIfhgXMaCdTwj
pwOXClzBADG6GxSVyzooNEw9GYGf8CGZuGUbf4miEFu6imwL/xv9cuZe9E1kQkPxG9hbGGrsbAAg
u3VK0iPqRy9vtuJ+C+YLl7Dy2J+1xfv4yc13/DrgdBMTsCn2Dr77Tyo7cCyr+8JIDUwyZcwvIrYw
kuWUGvnXRuFpRMBlWfRzAKHQQYD43cMLbMA03i0/3jXHGuxheiXRveS1hghBq+ALCktni/DWqUwC
+DUtM4Sy+Gea7y6D2Oam3fKz8BWmhnqxLQOrbhVBMdejALB/Cx4hHkUfDIEKUBUNxrUl20+K0ihZ
trjP681UVUREQx8jJUCQdsza/T1YvXSiibYK9sJTT7Q1sMqA67iv7kwavQ6QEJ7N2fs+sSBhfcOz
DP4uiXXqpx/w/IRddIt+mIxjVeCoSskpScSlwBuqxlBshUMyzkjzMLI11DYSq+L58vDAgjqiNnUe
a86+0FBbe73v858sEA4qq6KNHC72CcwctKcHexvpzO22Fw8dxyb8lMpHyKsbg1Uf8wxMwMJGhTTp
nfVBB+vetdNpWzlDf1kvZ+Rn7vCZVE67gglbtWokVSdVNwtceb0FOJhs0KNoZ2IEV5DR79JnCJjJ
zX3wD26hTSoQPlBQslYTpCk6KvITQIgZo5A3RVPvWvtTUZSfXcz/Twrc3e3039OD48WEh4NakJiA
3eCVAM7FjVMRQAJAt5HNdgsb1rWFviAfp9GV/ZkECrmR9/2E505bz7DQe+jdlW3cfL+R+pNwm6i2
5GUpxxwRsl0EkmAn7hfDCsP4NAwLvR+LS2PssKh6HqDccd8NrcfpZb/eqkSdc35LtcEWpnQcHGoR
Nc8hVUheCTC2eb0JNQNhHXS++jTnu1Jed3ETe8ScV4v6Wb3jVTyM0ihrD6azqXxMYHc6isgfsiYS
1zAetl2lYHDv9y70E93INo8Hjjz5ev3TIs0f9HogbEz//4ILL0XJS9uEFo+h+eiQ62mqwlIn2xbq
uL7rL1ViOYynb0HVtsU8+WIRrgOreP2wGpHU10FK2lLJOVgrembvh6rQZUjQdxfphClDXjLuAH4l
c6SxvWt2zXSd4XJE3nmK2VC5wUDh1j1f4xdik7T/ARtQuS2LLLtm6MLV2/ni8kOHyb80eBgTT2wG
1NvRnU6Bp0vLoJWl67XvbDyo6eFoIRTcHP8jTzzIHHteQjbg7y6VmYd6MPMhejNj7LezScIPpDU7
WjhHLWdNCOHvXYcbk/2+qTbRFtrxLNVhUY/V8l8J01Nmuhp1hKuaRDBh2YGHJWysVvJy9ssG0TIP
AmSKqJYoJhArGsNq84vCxpxoEyi6lNxU4puW828d4t7NlKKJ8dNry8rYnAAWdmMHCsCTiFIXm/hQ
Z01XHI+Y44O2/GhSgf2/h4cq34BLdSAVhhWwLXhIkJSkOzzZyY/j1cwvwc2mQQ8tnJw8cRdtODji
C/b3jBgyGVDJIuDK7b47j/VzIcDTUxKcnlePiBIi3fw1Ufay+XA3aJE68d9jzCLiSsaV8j7QkIo+
ldEB2mE2gH8dUk1QKVcn0E4So+sCTYPAp1lsUyaKbBMYlg1tsuvN/OLv/9uqNjvOD4wndhBSGbR+
EQWuprUHdfV9fWvfoCV57+0sAYXeo1+YrVcSo5MknrtCyyoHsLuOgqxjqIFs0PGbalN5yGomUWtF
7t2pMKP+5xNo3vmV15UYUfFhzAQGs21CvUzM92wx6DuO98nqUEmb3rQmUNUBu0F0LIV8tA9iwg9G
UtuRUINbvYKH/v/c+ShlZMAhm7ABltfJQxYgmeqRZH/V+j/UoW1cPn54uR3WhbGxEEm5RXVrDF6P
rBjhEH63DkLNeSaheinIfruIVt9rdZD3PcFXxbKfwanMclm25G3aQwGGDxbTi2BN4if/QBHcyWUY
NVebxiGD16E/3R980so9r+I2Q4ohBUYrF3dbxbsXDgFSIsyJpBNmo8rKdldLOgncDqBKKZUlhzgB
mrssEAcZFTpYd16QxLuwowuAwz1ZycRYlqgmK40HPc5GpzCRJ+/p5yL77ncBCDUzzrne0mnC6ZKj
oRlYyKfOgw7pSw8gTjnKlnRES+eE76u6+OFaSlZwfJtOO/AnXxiYEhCzXM4DsX1QTmMdxCWa5VaQ
DgX53esAOX74T86ddZeczoSJFljPeD9vHmq+Sv2DS89kMbyfb8QQe5UVxplvmHSFmv1wQYImX0VI
OgQB/CjWNMQHS53ze0dC3g4JmOEi21ZeOwMjk2KT5rDwIH0uaJCUGRXDw6md6wfQtaHTp1O+yGKY
xf8kTet1IGZRFk/z1gzOVI9U2EUwjnPpE8bomvqLXJGhHieZkMSRxQuxgozyUqsyfC/OK97T7Brv
gGdGPfE6DNpj0FWJWnefW3nzWMEaqCcrW56B3mi1LZVV6Q1+rlI0f+YFNrAxprNnfBwyk2T0FxX4
CGNQ1neJtLk9tM5njkRAPwMLR/dhKW7mdiqy0BkPqzfNp78nm7nJmPjRzK7Xr4zG6NhGdsFsIqm0
ddgSVRNF4Ytr67p7HtGbB9mkzuSh9ao+EwnxqWXHe7VeCd9pMZEhZm+DKHzxPBxY9Cud+mIKaPfc
Ncks6Yx7Kydv3KQDl+1PKYCs0ZXI77BRuiXftlBqa6R64U/fz/0PF73p9RvdD160bcME/xPOU3b6
MFNQckmFlWqvP0nM2XP/msJiY3j4KX87GECyk30ZPc8519Vy1B6iIw3XesUt6Mf0NjhWg4Hthbiv
/rARQu5GAdsugfJV1uCy9N/DSE7+psGVlScDZSWHL/X+d0PyfvGGbAhM6UQLJEwNZ7MkJi5OWrC3
5MoqK6wvvrgY9o8ROMUjUFkMsCrl2/Lars7shYZwEIqvAW6844113mye93Yt1SZoBJeV6baCk6lR
HaOMghU+erms5OQfKK+mrqZy/AXawgeOA61vZC/526+rl0jF9zPaWOzuL8QaL7b+FXO9zizBGZrk
ioYksce0jIhfNHC+rACBOsQd+bnQTIh1MgVlNL5fr6hXB8DuO6TRG7HgyN4n1HnrCmNsZ+kVa5K1
BWLfl0Sinre/3JNmTGddyAdkhgrgjsdCxq+H2f7hx9gX9QfH4EERROcm6Wiu5Is5V4rP+b2gVfh1
rfb/iBnOq/mZ9/qfE5Q+A/dZwAob47kZiZoRAajrlOe89Nydua585G2FaglRWp3e+cKm+eVISixP
QZCISsde24YM1qib8P4tpWA59d4SzIK2N2eum3HBeLXrPcHotie8m9iqRmPLOnKk/dDCLkGnDd9w
OCTHk7FZKakydy7rnZ9aGPJK12QJXe7xl9Lymc8Il7r9LDAqs/QQzI0G0vzaAzWC3HiX4wHTi8g2
MMWqmjm8I1tq9OXX4s+rlAXpgkFSamYbrbrEPR1WzzMvtsK8E+95bs9j+UV2doB1QL3Sp81UHDDK
KpAzh6oeEdaIXISNojGEJxQldGu+ePccz5v1vMMueAGFXpZoK6bIy+ahqZ5JPBmgu0lmmVikUP7k
uCBJtikFfwtM4qNw+d9Dk/72XTDJI0rJXRS5r7bSnSk1LMAOrqj1ClNYU5BPwT2f0JJHS23w14jA
olU+6fY3suHrO0AiRH541IeCnprI2sp9PELyo/M2Dk2ViPeEKSvzd1SvZ3tclGgDzbOz2YB+e6OJ
GBHa3hhN41GoPV3TM8qImjScoO9Q1AzRlF++8X4BqjJqpLcv6OXbixMoGP1E7SFsUOQyoOXARIuv
d/Hwn5qMkOk+IFEVp8cMOmoCMj1VAXIn6mQib5odb1VC0rlHopxaDIJefO0giaiTE5O5blVoq3bA
8X/gqOMbW4nhwBfcRhn1btUZhaAMivmTPVABZVRX/yvWh4dQlVwQGzJ1jLuLRdSyoh+uYx43VzXl
OR7Z9eoCH5BlZTy5NgNEcd+CYlsX3F0srA2QIl+a+SvBfLPG0En8gbS1cDSCdMQiJ+YgWSliOHaC
VrW6bgFRw02s2HMQy+OplARFYF12PbC4VGSBTTA5UbGP+dVKB19//e14xUrAwxvVCnH6gX5+EMKS
c01yIt4C4x3Z9sX/cWYhUuNM1GwLO8RKFHnqBcro4OvUG9F5vPjiCgGsVX2Th3XM3rAz3sraNHVE
hhIA9rXllY/+O/e0ZYJNLa0iJQ2RiVsnu5wrbucmbVnzUmaqxozeo1b1eURuu+4fUcVVnXKxDw/5
hBYreQwYgPhGlQ06EuUPKgHWNKlx0REMEfloxy+WHWBCoufSjIpaYGE87j9XKwfuPjf4qtfrl5yd
6Q2QlGX9soKtQGIHgIBDA3EQhQR1zWpqKSkNvM308MRmI0e1rYoxm5mb/a/eaN5J7wwiU/JPGHaf
EOL+MzJEzV7KJKF3DTZ5RVq2T0lu7+wjdAIdzLWnkIy/QFudXj3Pt8QjYksUuw9KMbyOlLfWf/eC
+UWxdr64YVdv7Wc+Ej0N9IHEr8Xk5oNMlOjCDG/IedTxrTFRP06LWN6W4iGsXGxdzeC3myi4UEGa
2R+qGpQcv3VKof5nOuULwG5wDutWFy6ER8bJsPbIj8IYN/4t4P9cqbrUSh0Zi+ngKujnp5xzgaCj
iDx0eR+RW2qdDh3Jj6+OuJK4MUEfErv50l8cb1l4hPbBRbZ3dxUd+0syBgh5+F/YaJCwwvAcKDs4
NJYSalr5MCQSAE2cfjwBlDb7g4oi432gymHwIr0dR6vwBVLJwqh8xvPIcEssJIeNamlFAR+uD3UA
UOdDvg6u9OIrIr7rFLskvikgZwVa37CcWJAo/OJn/Q4QOCchbpvm9bdkQQR3EcUDHhw+d/vBZWCH
oTaTjaZPYj5ctsnEoEOPkKGdkvaOzXgLKLnU5qJgDuRpBXuRnWFlqObAZad9LLCb9nxOfgoCokLz
BLP5McrOiCqH8dQxnkJAoEQEbUzgHrUYrGw3lHCLo4bJ5Pqo6KRTYOjxO+PpSINPvxdxh7KyhCs6
GBywTFYTNHNnX6Gm0BYcdWXmiyErX+NAx4RapSD7nJXBrHf66JcW7u3MZab2N1xUVwW6/S66GUOz
mx03s1/6wGzQF5PbzbGxx7OjDAklQp0kDvfRNxLMJ2SPGAe6nbmqv6GdVBS4lHwaef5QscLERVJf
yT1ni/ui1jG1BD+7k1i2woC0MHXdLZQebZTRzmoR/bwX8uw5RCSlO+NSr7x2h+uuLraaNuAT7kax
6GxTwcKX1LZBnbHkFghxGKKowyRk65rN/qyslGO9wMbIuMCh8NQ2QwqmRPnSjQu5dao+7LjB23Wb
EMZ+Hu9ghr7jd7C6Mw9oFFVtyfnm2B1wMMaGj3v3/ascUZ/jBmPDaIEG59tCU3cHkjj9tUqrIgst
FrZb6sbyZVAHFD/wBl5b2OXltDOTs6jC1lx4Ja00VedRM5lMVgqeoz6sl72Vf4D5WSWEyPMqrLb4
Nfmki9+gSWdqyGapMFkkXopnEWv+fvTGxBPfUxqYhyi6gZRhTzhXiG7hjs/fBPz02XuPQvSyLXVH
raciQvi1/EaWD9lYrN2QtdPJd0/ThyTPchx9HE6pXCbFfSz8DDKbUIUgO/NhJiMiyXNhrUjh0DHl
nEkFtgorhTZ8dXuS1Hk+28j373FyaJ4x86lS1XdZHYhGOJu4RtXZp658rMIbBuhF2qCh/RaOa2HH
S0FCPauBnie91Ey+ogXmC+TmJDdv031QQvAw0bAZsP/eCb7ogffcjI6Yva8P86BLsPZrwQr2Lb5D
pQ2NvgxhMVQdqlOHH/krmBX2nB75Vq9P974HIqHmGutkZu2fdf2ND/sFtWXW7R/izTOgZVV3x/Yp
1+K3bCY6OpakfBk9OFslfWsEQYQICTKMGE2EyFaRHXAfe32H4dN/YtPfYkKzCwchfnQQuSvspy3y
GNR48Khe7TyeewtCjNHlOQ7l8HkB0BTmon10Gtv2FgGSyawa6Pt08a/r44FulrnhKHTcovJONeb1
/tnel+NUlUlA4b4O5JYdsOvxP+/CqtWp2MdOHX++EEIvpMorSS+MpYrCtIa0xFZYy67qP2U0dd4V
iwGUZ7+TOLQSH4xVzwf1e2tHmfBIM7neKBuEnKiBnGpw1KaJYVpNU11Tqyh3amZPPB0FEvzH+b6e
n1qYvthx3HTpefe6iX/4t74Eja2Sdpw6dZz20/lMXxm8lmqTWDQO2oD8Uy8I3kZU5VD0Kpk5kRuQ
/FFDrtjx+gh8GI9kPQsF7HAFWq6ru3k8LsXjuNRhmyJjQngK9WfrGNFEEP4boDSCTy2UJJCiqlkx
s7GloG/z6rvx/c5R4ANqEMDKBNr0vbmROPXek6RHImM9Oa2BgffDKe2SA53XkkheoRnWp+WK7eMY
oPtXXTf7WqiSxt+Oj4Mt72hLzjaX/MdJ/wkFVyIfYShvPJASxiJdzdRcwrGBS7JpBtaia038Sbf0
1Tgkk6307IaixMEb9r3kQmlYTxL508dtCWLWyBcueXOSFe0t/P0sPvYqOeAM9BQYXU22stBB+Jk5
J3/Ivrng87kJLQnb7AdKoiSrjPm9t1ui6fypFUS69DICIZH3UlpRePTXu7CUzM4tKh9qyvLs+jwX
RYyEXHkNhGtrv/MqyKcbIugB69m1EZWvrw7jkLAl6t1XuJaSvwA+YLjtCwJBGn20yZ5kYiJzov27
mLZerpmgdqG30ayJ2JQDIJjaldjS4jn+JD58CnjBbiN5BUC/OGXP25O57AQeXj3GvARGdW75+qit
fDeSU2f2W2DppDEwb5PzPQYzPPgyFpRH7yakzycP19MX2KQsK5n7/0fABMb+2lwB/Efy1WFmTDdY
b50/pFTmZ2JEveCUwsqHajC/Fcv7zOEg3vekoAD+jdJsxMXP8o51/+XNtdLO5dwuXAxnnaleX0Yw
gehEDY2k+Knkfy5JTiSECjrGUDRbDM0gaRxDP20K359F2ECt+6opFTl7RFmixlJPheAcVESqpSFu
Af35GNi/Vk2noCdnSCxczs/qX0vkh5tVHOZ98Mx6x+KJeAqh79FpwJQ4KwA4lOHQ/H5bo+E8jCgm
7x2PSgw6ZIHX01GnlWUA5DLobM3gfxtdw8DBgKYwBuq5xSDTFPN6O2nFldpmT6lFTuYk5CLXvj3H
k4EdL1NLOlwjS4RirouTtuDwnrilYLR6dIjuHSsu19tjg8c5leTq9tI+VV1h/URWHV6muqTBiFz8
tRRgh9I1ubzdhMZ+av4mZDQTrpjQ3+v/bkW4VGu89oXuY7iCol+9PaabcveEy8FoIDUSru6CLiOI
CFTMg4msBuHAJbB0jCJd0CEUdgDGgm7RjjfCFok0gaPuZjARS0AC/scLLqTOKIUBzuk0XAGzIUfL
k+IvuVgGQQg73I+B826RqM3hj4Wc7Ah62ldviIqru+/KljpqMr72+rKTX1kKHoFSN8+IR5fX3gET
CGhSCoYQRXATNCORcj9xvxNJyjy8L//7hCRY73yVMm3qEBvvtiLk1yiDEr4ZUhwE3xdyP2OOXqFv
/ej3WXT8VvghN25EGKCTulmYAkigeIM7u2UDZa6nZ8eT9H9Dq529v9n4iJtUk6gfzMCvJzRA7MDx
ryFjEsSjb/GK58aC3tCscrmt9+eHTiY4l9IBrgLPXkk4+5DPFC/WW4cjme26YkE/TPz0MU6Um/d0
kAMWaLejf5/PUsYBFAV/lYW7l6bdRuOuVeiQn9pgr2BXPS+Ndsz6eg8CsKmlkW4o8s2FRfuD16pM
LE37hyBM1koU4Kr2hCdGyXy1TXqsUXgHyyiLGnHzMX7tDGLiNamXLsFMT92Bj+BT/MfcE+H92Qlc
F+TR9YyFR793m7PA9Iz2NjIfB52mlVlpTjH5sdMvdNzndEZ6EupraNbG7Jp+0QmBdhB5yI7LTICG
hmJQ81TwH7skOTrdhn5b3Dxh02y3X4fNoNgl0YerHUsLqrVkkuXLvU/P0ZHAtuQv+VpqpaQTGYdX
FhleH8PDFZ1Db59jhrQNGROfTxW/cifUnFaPxydiL6bWSr6RCPGWWoZ627NQahw07KyK4RRqMs4L
Ks3oqKtL302pfo+DPX1LoNQiAbtUcarAdr8nJO6DvVcpw/flHwcCtDHJkn7Y54/Xmge6A9Bq766C
aRos116WZeaWpgHupP2lts/DM6pJyAWlFCm9qIINpLU9owBQGSZJjmIR9AsOKMd9TTg6nmJ9qo8D
OPwyvEvep/5usgYazK7wbNZpQ9cryu2Zgmde7nq129M+lvFh9nGyEaBKWSU/3Wb2dsxXJW7VBtX8
RPeUxkAjgtzPz/lB6UMIzAOKZipNE1Kv9AqHTBld1IWFtPiOoqvI5LvFxN/nDPgbjoCHWWAdqHWY
jNlK6dzkQafQQfYnpfbd85fSBt3V3JIHJKsM6wkdiEIuw1CP1ZO5u8N9MKazH452k23m471BWNdU
IPPipTvFlWKXgpaqS8QQ7znU8bTZdKd879np5l8SpBPMdCxISwotGX/mqkKo+gGwnrqwt25xoxa4
htDrarBOScKiDan5s6y2EA/VIt4k7dRSr+Cs9MX6clxepm6vyMrNQH5jFmeVBZhrVperKHrLsAnD
80EBigHBaquEPLovzOGB5CgkZfyZ+5FKLAhjqgMEnOs9XVzNYyRMrMexxIAPcslr5friDfDgHyjJ
H9V4Lp1Q4ZVmhvMQ0tCV3MFvc9mLUbp8yRBAwH3TZ+SImRW/1da4zD6PZXfkrRgpx7UUG94TQDzc
shvOwelhJINalqweTKpP6ozLtypF5ofnJnQi4TJjXWx+03ugZg6zcqNqxR5DhUC6vhrjK+3hUb4t
HLxE5ot3UfuvqTR44rswX+C03Mth2/5UWnOznzN54qyR0mGmT2qnEXWnR9MYwoIuQSECcSygTrgS
j2CF3XtLkYMPnl5aP7jb6o7/7vOIEKw+cARxQy//GNo7wj5vLEyA3Dsj63ltR/Gm9dBfMSHcRuuP
8H5jZicFxZzgX8xa649yj51afBC8FBae2iMjNlahooI7ux9i9USF5mE86dePln+kzjnKYOMZHBpF
k3hagMGE3Ipg4Y4tMSqAXkzpiL46xRiPfN2rpglhB8fbPWtWBIA5ivLA5EwW8FnhCNcHF2/WvCx0
hquEJgmdTkKcn1/L9gO9rEVXz5IbVz81tb6mUSiID5jshSb8/xD4UFwHon04/QqDJrziACELuQh3
PAZpfJPAq1Kud5ibRClUH24ZFaGStpKMGAstYBKPuGhHZS9KzGtAz2zhC9pAtrIakKlslffSacku
N8fhaPpa2/OjwF3mZ37sCdAGVzhidGDxKqh5ym/RR/I9eCEbeLks/EfjcVB/UJxyJ3xoF9ec8Pmf
I5VbicITaPpavPNk1v/GBxTQtT+IjSqUzOeOpUpzwLTVHlKt0HjFU9V4QGN/SDfRlPJ9gvJVJooP
ibWeRevj/u0zE4gXTNRzCFkXDsQ+Lveo7yKcbJ4sLr97G3I18fbcU0eQf4luvsV5n7fSjHuKBPnx
HugvrCz+8oCM4jSQEeBXAz7nI9e06699UiaM+hhwatHlXY1yIC6byATHtsz5wR31xBtsC4Ne8TSr
OAjsunk0G12T1UOWWz648IDTX0RLGJTvDRms0kKwZ6wCZkGcIz/GwQFS96vcVMN+iDJnr+oUSJgS
dnSBWW7q0fSunSSoAvceD2gwMn3yWw1JMDCnZxdZg3nvnRtLbOm0NdOCmgb/EqxBqsAa4UkSvzI7
izqkWoxim6jWdy+OLW5oC0LMmzvlZzd+6X6ddATEzt5U4nzugYWMSDexUNhdsfktXBTh7YTfw5p2
jLJr2sgp80kohZANWpc9CDJGYNywIgDgbKuWR6PTV2BcRQUO6h+PheoF8dUIGO7IsyQZ2Hfnkd1A
VLztU/BZNPc4Kvl/ZVhbZp0imexvVCthIKjHnTaTdXAuge+JzQN7g/V+1ryt21inY4+DqzRSMk6e
+lk4IU6Gy/4dmy8c3ZoWO5ez8MndC0QN7UlBfzGYwJTovJzaw2nevHp/tyiW/M4ojJNPfEmE6z+T
OP5Pv1/uVuEvQpwnHNvixLD54MjS+yWdEwnQtzbHkHq/XhY/zWiVBbTt18CrB/xb5bxvrFjPrnWW
JQw4Wrg23sIo9sHo9HkPn2n0+budIy4aoV6gRGiZHJUmJqAAuw5NXW/mK9J84vVKeXbXQRyraFnm
9501+esjueS3F14uO5dToqHghADHxseHu+4VAMVCx6nCGawPIz4XItasWu0IE0QpOGlebHIFGJL/
Qk/+t23dXjNtbRhz1u2mdjqR7wIOcjzt8+OQkjtV5jRBeA1qEJOgp0tOO2DDe/ufeBE38WbDxzjI
9ZHoP1/6sgjUGr0rwBNA5x+al+1oKrjKL3Yj4tVEbzJrQ/miop29grBLsIrROwXW5G5Wf/GYhewd
+TsCIiUIf6YJtakJP6QHwKDrmHdYiCP04SCGfJ8HW5BHvSVvI0BltYfsbJxMhaL2X1YZCeJvJb9e
L88leHxjI8r3QmkdEoJvR4S64yQCCbSA8dZkmgJx9TvELV95I0bE/E2pr3M45TsS280fFO6Uvy6D
4EANuZpBUKZ2lg+jyqEU+T08pzLm74PDKQmYDUeJ9e5e5d+FN5QWv3tPMU4/z4jCKWR+bx/4B5Xe
xod4SO69rEhj4vApRnzXw/r96FkN4aUv0KYiVe6OX8gz7xeKqI3JtwMiugQvyMvkk+8WGTKLatXL
iikFi/vUopWd0SvWcXntebnSAlZTFO0fEReRo/ynP/lp/DtnSM+gQ42TpSJQaGdklragiWjLwpfw
7MPzba4swNkRAyl5rVT4wSnjjPMy6/cWcTG0E5Ji5x1qiEvAsHQrETjHWjd6RdDeuK9nsTjZs1oN
OAgGn5CUKJKaBK/k1rWiHhsSVISoqsmD3TaJG4yfD6b925yUm2Rz/uUxUHBQsPDayTY5vc2iN8rQ
SfwkSuGJvlg3yJv+2PvQJZ91xTW+CDcEfY/QSQV0RksF5OfIk/W6+kUECZSytL0RlnONkZS2v7Q8
Xjzh2nfiNw4WYRtHlML+pYLLqU9nHAYCC61JqREIcPNNLQ0CFPRhAqM4c7C1BIC2fAZUplTYlh7k
xCDueuMuCVRvuTiKmSjp/3FOLx91zvJzaDhgi1gxD7Ya3ZNajgGQ2fQZwBaiVxQffbn4pc9l40xA
NNW8fMgTg4+zjiSwv1oa3wSFX8OaIrUKgSrJb5KDUOBxxOMfRZfHUcWMkpYW+ijEkC1zL/JeK4qV
loTjwlYLWuVEjfwEyYMTmbznS4SJxjc/QCLKCEw39Odflk8Lrjd0GtWcm8DCGCNRUSM3VcZfUFBj
ldQY2V6KYYWDQGwrUYElZzD1h/QdeT1MO4w0Jn93315g1GXgi4hpeZHZoydMwRVqFDoKZOYIrGX5
vlZCPzk/FkZIXtvCgASqlcWOUPm9ZuIfy09Z78KWFvTe11eMlN7xSpWzR22EmLtjmW2XDesbRc/f
9O1fBd9UOJl4aN3Z6CxxePKFP5h0IVxD5X3RoXEWAVZW5y2KoQdhPKdR70fCKEKiwoFgyp9rKHII
KACjeykFGe8jxUb0n6/fIsnKOTn2pR3QFBry1FWBmuqQxG9WAXC0c5snX6Wurxp8rAJZvHkClD1R
Dc4l0GmP06GcRovkR7QRdWBgQd4QfADLfS3JLpi0Zh90ATgpcyBYAQQDugJiZ8Ed/WpxTRk5LduB
dqdcCXDpz6gbQ3f13lNTInDQpgDKZJcTgQ7Zy6NWZ9yvxGsYpV/wQKRB30gGFlLztt0TE+I82p1V
dvJkDp+GV3Uls664lK403DCm56teCA7EQehApAZSnlJ5Ora3p9rMtgb4ZeEpm7U+ggMC7yw/7Z0f
mb7KT+Ra7H9obaYJcsPHPWi3NZpnkShlyOZ4Hqh4IqglwnW+0M6eO5WjHCvjW8uLsjqdFgtHmkzs
iCfoNxdf0D3qtH/7i+NRfkrhMhUwDJ8bX+yyzZY8P3y8bnkSlnR3XFDFAVZWBHxFV+v8/Rf1a+hY
RQ7+thSoHUr5r1rmYAsGZMg9TecE4zgFAi5mLj7N0jBNrUR9HS3kpd4lj14bVlCtAQDCgnYCQFg6
bWrK1/TLeC4rxV6l3VvOfgjnybLcSGxkJ65y2DgYXSUV7giAL8Y6ejZEtm0oA8li0Gm6AKUyeAol
hSSOqORsDQizN/3h0tVTYb+toKGPKGjeLYVaWHv9oq4tmP100st9muJUeBcYGxeY2pyI1gmGdXJZ
Zoo1ut5uFdBhVWULsPA6juJIkD4MPRlTsbfzp9q3een3c6pxETv8APiMI/p1jdfeTa4RkarAX1uA
dobvjrQ45SzM5agftHLVGiqrcoifUJYnScuxOcsGDDbF8/CwH23YupFrlbvlsf/OdHkosl16Fv4g
0eGUgVtydBj9E8VkEMoE3NrlkqgvlVRi/Q6cdxH/mXrVlK4La9wes1jsE+gI9diHNDcU6zxFR0nb
OtMzqc5OnWiaxUlhWKYwfgrHTUHxDx44SE91zpLMsnXW5jK23xVH5kHB0CwdzLhPLT1icSJRUaWC
KC5pw+R42IubKPZpcDOs9JB+Gsdn3CzD1fAUE1i88E8vnLKqui/gccC4Lz1KYSKPjKaRFrbfT9pu
u8xh9GdmedUx+9JxjCWDlDc+PhbX9tJqt9iPTi6dHrB/WXNlJLPw5CwyUZ4t1gFVoPFj7dMSb9SS
toRHZ1VArWw1rrTb48rNX3OB1aD6wKpNfI78d/ALirCY+afQHSLDZZpsAWzurWdNq+UIFrYv1fgS
t4aSLV1C3MwjWFpD3z+tWOnPi9vPQiUsAOPB/KygmJ648EZXBeqEBqWGMXRQDJ37QGmPwG58ISYj
uw9+TTWKp2TfapzWVODrv1OF+gYct2DYNnVW1DOdTaCKga0IxqzGZvx4KbfCtoZY0Z2UduMgkfXn
FLk5xgEZHnGWJauMaB6w6Yxsz+pi1IgZ7uCfsmxKugGqcmtOYWu7Q/pIq90YU9zD173ov3AFyg4u
0L3f8KUrbPyeKe7Vxqo/NwUIV1gEh4j5KqpIOPWN3pOUcekgk/kM0VwzpYT3IGydhwgUgzNSIwz4
9eqaczuYyZ8XviSN78r7M7R1xS76/0jfB7clquxSN8PFrFrZVr27mlhIx5R1f8ep74YGLutea3/c
xXJv3kePWY6unlXz8NF51WissN60+Fv2oP1PbLu+woYk091qcM+JNVLDl4p7iYzdHqjDXJ7s3tCM
3cyBCbUmXjlP59QucwUVCjJc0g7qsPApgk1xadKkSkhPzaQurr7rGEgixHGvG2N0fpzgX5RgY3Fw
g+0PLNjDYuVXaaII47HqpnDL13I0hlQP02hHKWfxM+1saStq6H/XLBbUccCMhQa59CBrAh1ZD+5S
BcU20eY70fEZMpqWIcSgLVdKhCBTgvLFs3z7JfKfvSnMz5ANHDQnI45sKU7A1PY1eoIavtvanNAC
FPPD8zZyiT88sk3yXnCDN2H+DryWP5/ivU4Tyic0DXmIe44bFU5mIpEkgIcn6OsKLiinqPmSy6ZR
K634eZ5j0FrN/7ony5xy4uL3La0bTpd7+fZqPiPD3I7TSHkc87juloWmZOlFm5xqBBqf4/hclm3r
0QIcLZS/qzTJrS2Taf/+SlaKThRmZyWd5eZzv9sJSDqndZJaBeFwwx+P8rW/P5DFvrumSBLlxJp7
blmMCKQ3XujsaiKQvD3e309xHbWSFRaHfuy0SEN3ZuSaNFbZkCUDT7JtEnBkeC6/mUuluzbugkzR
LeATFUDlhg/FXR3LfqHWWW7SBdu6WtThR+/Bj99Kv8gbSu4h+7Q2TfB9aoB6ZbqengdL/kskkLKG
WxYnOQhDmmFV0IA2CXf5oApM4vk98PIIiU5QaaBSGR6vZBFNA+rL7Ix81rgjBikFuOuooqYwdOu3
qW40nHN7Ikvgz2qx2UcYJOrIbWdLxbKNXJXr57TA4uiwAmxyKFYQNHfJntaAC53fN3klzmZJZVzj
+TTfi6gVxcKeBiQau7D3+tYRMleNJn5JuL3MyLqOFDzbj5VcYOV8z9v97Uv1C2tWEA3zfF/iCPJk
GwVtl+5f7m+xCLWN76GaYKGN+SDeDWfbyj0MtvcwcuDgzfRQgrvwqWgx5I4NmDPkGwcKH8WJP0WO
vZsBI3apUYmSdb4MMXadOjyMf9FCCA+0a4qic9G4Z6JDne3nWcdEcGIbpa5AcxbsX2BNEAkYvcDk
dGAr3rSE6x6Sfq19MT2XUhx7dgzXmJpTK9au+fy2FoI4SeEyKKaNfmMafVjPYapPGNuzu/paUL6S
x2KEDORcAxVRpstOGiKYbiClfEFW+UTGWTapbTuuFiekCvVgsZQ8z9qrSQoaepyG5oL92o2g7abA
+KKenDSi/TbHNLYZgzxGxObd7QaCT9cZ8f5ORfpPA+v0+60VwzMccu2EWQJtebOUEXJOQajwEgSk
cd0er5uNPJt9bgbxf/CjOBG7qZnNO5i+RthyUmIURK8YgdW4+/XGw3NtcCh/6Hb2QeaTlb4+6iF6
8D9k6/1eO8Tv48aEDT4BdzckxYXfg4FhQ0gpNUkulVAd0nKvyuCoU45tsdvZNaOi6D9i5NCCTz1B
U7U1MGqGwsbhqUalYBIrlMjSRxW71MMw2pXqPjIsFSJXgO5PPRalILEyttY7zdH98Qk/VvaGhiYn
9gFDLGq7dUt63dywjT+HBxaeoy5bRj+IiRT8kfAnvDxuyWkNNh3rmSIOeS7VcEKD+5lADLctwccr
yvgtDSfaWcBgawV76XdrgmI4Oa9ZAsiksPdp6lHemQrQV+8V7T7hIhJmYbgYcIlSqqBp9tCDr4zC
71xT1wuej4qWS+hDCpuLNxAGx9qmUxLeSRb7cQq9SD2DPiY77nNUEMSIs2zACkd8b8p0dc+qAHJR
VtBGbsvBpYMDL7FQS3PprMIW1/opRM/2IobjAAu4i6IzwH3lgFs/zgugCmLmyq9VbIrr0Ov1MUDj
6/JpSwdmPAZsgyxmJB5KHb1Dl2EGbrQXl1uIgElHp8P0Gtw8EcuCyyU0KoIUsAP/CNJhtR63FHkc
8qfCUThdDA2b3EGHOGNCK9GmdS0x22MzN9tRlxONXnBiKtepyyOvRo85gnACadBsXytsm7U9g1D3
4RAVNfYfK29C12gG0ULenz/fe+vweDjGdxkDZCxYcvFgEdJ80k8L6XvbS8UhQe/tADh4IR+43Xoz
nbTUQkA1ZuSqPSU33EGmrUx8Zp0SR/5UIs5fi71+9I2n9X9LP23PqMt/CNciB78V0QwwTqERBZbi
gv2xlvYT51+h+tOvRExLJUNX42O5K5sL9BUG8FkGB1jSnkorbVabCuYHB5KiyUU+hSGCgJAYcNJa
B+qY7QpJQZEgayP/msoeKtEKmhhAGEx+OPgrkEKmLZSEz3dx7yeQvKFilYHYvNDNA3G5/9sSr5i/
E+zvyYvvcy/N4WuYtgwTs7Y3oAfroIdpUQRCupGf8sSLsLcE0t02Oc91ZZHA+HR2KEbE84WVLd1F
AnQ6+PW7Lyt1pOLAPsrZlzvn7xen67uFZqILQy7p/FSvjKoPkJnIv1JKeqWzPMlIkzd0xqKrpH1o
RlXY03gYqIaal/l06dINdy/iCrhZe/MQW+RsJzRLPKAFwAh+OwAwpSwS4eHgE+rXvPgHCJpvjPMP
AtT70UOvsJsCuEIa/j90RZ1TRNgksBThfLv8HbxBtn4gItE8D1RPauy7BOa3oFyTLv4lzS4OMRDf
RnIgIBiXRMKm174ykCoBx+hUP79OwvcMtAiNae24SzvOEPNlh5GggmThkwVGjb//1XQeJClTgMoi
W5kLJkJMluD0hzdEGDG2MD1jO9jBpqkNFTnxDC7I6ex1njpsxGdRRjX5d6N/iHlasu+HRNK3xWcN
uE7e5udSUrqjBV9hnj5IGZwdpe+0dSN3fOf6DdBKFpyhwkeNH2bZdIM9xX+9gt0kG9pTa07vTtC3
osBHFSPRRHWccpFlxSui/bOyhm8cTiDx8SRRHnbhmwYO8dHqi8yF3XAoajX+0wU4H9+LljQgHg1s
oV6k5l+812OmWgeI0gbYWoRao5DWK7rBulUWkLbUXx/wltCF8/Txg0WzwQetSzkXe2fsnTuUfnKg
bedlHBZikp9dy/ZU+Fhn3Fyul2xreYn7obaPJbFpH2vTnT0zgslxQcUMefwuCq2OTnFsQwjKAgw5
7jNxmGNsHVc05gp9ZNwieKE4IigC5kaEcD5whWWvmKFT/69kvnkSSj8J67Ey2REXS5FE3d9KBivZ
rgaW+gxA+d8/ZZBqUMwB7FYyhwgd1xnDwq/T5kM2Udg4L0IYJMAyLMeKEkD7KE8PRsGiyYntLzPm
qmTiXTj2+oQUEnMKo3SZxL3asNUFT+3qiGPdE4O448oCFJ74TiEU3v0dq2m0DYIAneQcxtTKIYdK
C0bv89Zvig1ArQ5F9m6s58SVWdqR5TgmI+CuXN4g+ujc3rSO7JRlJ1IbfuYxeUZ6KMe7i5fApZb9
J5ZxykbtP+DIfRyglte8/blAY3RG8gjRsfWTyLQWfxNbysl4kqwLiM8i5Pi016/y3FLpRXz0bTYY
SR5vrs8luUvyn47NfSbrgH7AFz+H2aGF38fVM1GkLIxwz1w7kCSWP38eez7MviBmH0yjLIcx4Td1
z5drwo3ayZuFZG1Ko8kE93/iixBn2VJtOfxtBxsUyPeh0NqAoM9x/V+HnyZaUCve7+X4K3qzRvq6
Df/j76xDR//iY0NO1c3rjN0hhd1TFMKXKipSOozKeYn1935FHS43kk2cd2DZ1vatnUKXzQ2ku8My
29ssGEO+HX0JbrSacLCLQ61T4Icx8geebwm9Rvs0TvM83k6VeJtqUPdQJUUE2NVEJvR2m+li3eSY
VeboBWQuuogOhDKDtdx8yUOdxns+8gOKWjD1CTt27m06/8iKcCm5zE+6Ug7GbGvC7d3/tjP/ivAE
ADqUi3apnSmWosDguw9+JK1L0errlNsjaIPSciVeLBkSZ6kCfJCLYM+ZvLLzIm+BynUtr2AmlH9d
rkYQN7o6n138JmKc1ma2LbQAPJfdZID25pdTBfwEdoFpU27GrGf7q2cpQxGeZdEiUfmJbQ/j+eYz
krS2P/UIW3p25Ym36OygZHp5THCAu9NiNDuHD2ShUdaCjYHPqlhbdE/2Klj7KdnRBWOT3Z9cChED
QOPPKGsNo7fcCvgILH3/d0zINtZXXItRJFZJvhxZoUQuKumOlx2r6npWBO6JsaGdrFkERHTRY+z6
dI84m8O2v+WwolNaLHeTe18WrjhSL4VpjmHP8ryYKnCzYTwIr+1S7JCcXgtdK/YVtiyJceH/mn9D
C5GcsuVPIb+TdPlhAN+3T980+34CpR3sHT3AuIl0H5lnVC3mNPnB+sEJW2HREac4l656qrZ0qXUz
Qia0CTAspz74GB0wFk5ieqUvrdtmD58Xo/yPKgWbMlrCaqtiOnBIjnxFLFcEanb5XSGHhKHJt1GR
hL8/l6vo8ngojAp5OMHjxSY5phXzfkHJbCHu5/hH3HDolIRlhOBB99zqTNBjS6PmJbF5rCAjJRG6
3W05Ed9vwgs7O9KZnLpl8qfvzAythC+6O72WyR5OO2i3v1jeFwJdPtWCJOYzkYFp1m7Cm8UKfuBT
YQTwOzHgszhFnC5CrFbTzEnoyfVUnhjRWJthcXTaWrWvjU1vDF/O1XO695rbvJgvAQhFxaKfauoK
J3LLmunq6QfpDp9vTOhiS+2b4KzwE6E4vR1eXK7M1gMNJkSDrG4dQOWLtp/39GLz/HxQJb3BEbQt
ByulARR1PwTqcmtJnNktObn4D6XQ8HuwWivKG2zc9e6ysQwdk7XX3W9Gb8HeEglLZ7VlA2Z935CK
GZs9wPZESobM+hJwnZvSNM3hL43GrtKLEVuIYJLNvNZDYvNp/GEpJ1hQWB5LPUIdkTiWBTRXyIoJ
oXaCMhzUYhCqkNDAnJRLlvGtbOiFv0Aje1/BuUNma6QCVJ6weF5/pBN0sH4RkqY4kJmnhDgorWan
WAeQePFj859NcyovBU0G0WRVdOcBAaqPL5SOwm59bluAek6CZkHnlSw+FEwSawtrilieaCn14WsR
oKN/XZb3u1VA9WMBLsUcTVDC/QoL87sH585aChsh9Kg1QijBPPP3sN3nK75OfwcGTHy0Fn3WpNKt
D/L6ToN0hR8LlmSotZoEhiCHRwukqOE5mX3zHoCh5HWsaN5NgOV9EIPgVd5MG02obi9SY0RtFmN2
DHXeo2YEBopa/0Yug/VVJIIj+G5uKPphSRGmLHqbKJxDVLuvMarOXGzkEAR7llqernnVDwoNyJfQ
5f3DEeTyvkcpYxMWaIUfpzIuOXmt0OktOI12TW2VxoJi2LNq0ZIg0d19Ri+GR+S6bR6THacmsriN
Gn8SYBBJf4FsiG6Xm9FOQZT2A5YABvFyRlIc+OW3IVotH+7xQAVhwnjBXS3NWNVOS3yr0yDoGJF+
0BBlY3k/jVCXzXoHKCoFrNmUBmF+HvypiSP7Xh5mEqdx2Krud1yyLslo5CRS6jPe5iPF/p4YVBFG
RAObNNmHVRVaHQyg3MK4QG0aaVweZfj5NrbwG/a1ddqTMU3TKBo0qgAxz0MSSWkMGGXrBXu9FPSr
+NDY8VBaJvpVjBQ7k68mDqjZNcNy/iMo2P3ZJvBkAUXCQd7mOaorCY/Hjaf1sw+lX0iQhgMzOi+0
SvCEFU45K2Iz5/1Ap0cjdE56KLqHvpJmD0ZO0vQLVYAVzVFcOnKL/hzGmlFb7kNAmeZQRcjI3erL
Gzj86nizG9wPeGmmIvTrYnTgxyANfh+V+AOywLnz4WrSinotW/DUtwCMgAQX114j7mpP7SNA4+Iw
d4fvKvlC8Qj+qkxO8mhaNGCX16K2VqPlxrBOBd/9so/xvsXy1NuRC0SD5QKvsLhfb9ebGpzMpxG9
migFRkt3rBOCXrYeslPicLkRHg+KnE2al3fAHM7Q8pm7JM3QohgVst3KbyRrPIRgLxV1RNbI/Xlh
Dkhc+P3KryF/ZhJWPGr0DUC2o8CRBqgeCv2G7anGMtAYJUJs/YtJA/lrk6hrUmIzC6MNtry3LKzc
MTNLs3UjftcdB2lhcW8mQsGQjkWBSqmvY0CojAN1ghokL/v0DHRExnDzhAtcq5lJaUrRJDl+5B/h
F3WkCEVw4T4dMaXpbYwdkPBqE9mBdI8yzkulJnLXS73pt2FQm9JjTDpxTSZ3jaMPjnd45PgxHcnF
4mFXBR7ayl7EJKy9gmaIZ17/s8M8MdNDADen1lBnINxyx6oxpPACm0SDQUDSm2oukYU8kypbTAsl
a+xwzMNwksJs+fPOapURAwJk2Y+KusrCCLdMiw2tRzNDbznz7OZqtuX17v6ypbVTf++WD6+d/eny
EjPuiSFWmSZaF2ihFEtQioKplvKuHJryJytxCUxuVmbdwTafpI6AzZDAfCpC6jng1KHd0QiESho8
iPVgMmMQi3NwZO7j7E/624ByxSF7uie9GlftSueHXhMbAVi5EdGSQ5pKJGOUSnKf4SwoTZnoLh26
pa4O7SMF7N+kamxQyKgkDRsa2Q0p0JtKIsBo6MdnkOWpvc6ecq5z4s+OucKmvky14uTLyQEaIeDK
twCMNeBoUqgpSDlGDO0G6C8kUG1nqB4ewm39ZxhBVCF5F7l/Go69+KOQkPDMdr8XfwVeTOKUWflv
MHghPnzZW5iXN9WsyVftPwOiBJBdyxZ9bMCTgjq/hPbfhPrcW38CHlByvuqhXM+KCynm3Z6e+y94
TqdVPeVi6T4kO1nhGOUtRhOsZNrYAcXNGvd/kgM56Wr52rBU5sI6zk78qnWMXNf31SZxM2cKT2/M
1o1HZ0Jn7WekwbArRgs86p+RvGLxJbd97prilrCwgOwTefixU64EThlcs3GsbpbP5UWlOu2S5/X2
qnD5NGuS9g7YFcnEvB3bsVCfS/Wk+hmce/02S658gzuYZ921QRip2CqBDMQk1lxlSTeoT0qIA2Ft
Cu/URakW7lQDlLbO25/I2WRMXVV/+1L3Gx9QXRH/KtSbvfaJxvN1On9m2uCl5xhchVFKRcH5pC42
aGcbNlIJNuQ6krCTUa0fi875Kl3n41RdLSd1PCD9CwIUJF/9vVtvi1LtPJDWFBA2DgN58KLXW8Xq
MoRUaFD1VpE3gVCNJTwnnvElUf2ZyqaPa8g7SovAoTeHD2vr7T1QxbCArsB9ULPpGT8i+q/Aymvb
q/7HDd+X6+P+mHZfTq6qs6XiCSvZEW/9psxLaVGt4R505k2eiZP2vDJb000mtO8jUotwhKm4Rl/6
2wJfoWBV7h3BHzy03qZcQ0l11LxzNDj+dBJHzX0bP9S1DNQOmYygJgt35d3/nNxh9czvtkA9TrUK
7aigXXZsmcbja3jhtr/J5zzrIl7GWRVrywaLcsxhoXUD32h6bWuWOpy0iLOFKzsYZD6QrXx8evF/
sWEWdcfv6MgT90VCHDO081lCDy6F214S7Z9Tc3+agHUBV8equSzIIYD5BNb/GhGkAbDh4MJgAl9i
RJiPTpHKYdlTdrniclJQcoUa4+dd8AW0bEtSF/lKlCQKKUD+g3TCkGcw9W4z38AuT43rlITKzF4e
p4tpqaAnEBUZSAHxg3aA+SVG/PMfVpK/Bksoea1jf0h+UxiaXLd2HDGfQc3x01Nho3FuW3vBiTFe
ejhLHXLuDE0KSVEA6634gz8NavcwYISNaydbYcwKxW0VS9OrCQ9zM8QZVihL9eYexfm3sgEvhOHG
m7L0jnZVOrHZJ56GtISCGNKET0qsote2+h3LtBaLpda7iI9Hyq3cMp+MZIyo8z1dOP2FoOHbF4Ou
38vFPBy+T9kw5/c+vLfQTVUY8PmT1loPyW99xgoFrS0kQuRzqKdqCYz7seLi2M3NC7gDz/AiDLZV
WpcvIdrnC2QRsAq7yMzfeGS+Wbn9ZL93crT+T/uvTvOIWmYdwd55gTO4qJkdpuxSDb8AjsmUKa/B
fin1gi0i0L56B+2A4QZtIsvJ95vp5QnLVsXOGIc0kU2PiknBI2VWgw9oDkh8OBlmT38O5SxtN2cY
xM1aBTemcyObpgHsm5Vsbzg8eX1Lh0d6Oh0u0YaIs990zjKVpKePbDYS+J2Qx24MXyETnlfkhtKM
uOa3EJgZoHEXXvoT1RiCDPpvgdd6jOk9OJCQcnvp+vbKysriEZFtVj8OM4Vb0q/7avXsOzWhxYZ/
FS3S1JwYr+q1tddZhbVej4qNUTioqzXQyoQXa179MDakxtU96kzfcmedZPpnam43pNMaaVZIbNQ/
sLeycncliIqUWWx7nPNXjVOh028GWddvwCV1LY/WmAY4yOX7NrGOW4213o95Tvq8F8Z+Jsz3XR/U
Dh7DR9oDMs66wcIEk4/hyvEro82BKJhHSJY2dRJs1GTIU0nFNGOr2VWawwQwTqAQxT7kfXXgYOgp
qqFo1RKNvk00GfUfirGsJ0Fi4A7vCTjSQ+IoP8r5ExIEziR6r9ihZC1naN0u0fZKbCMGDEcyxWQO
uAOQ5WwvCmMTvqsLMG3zHL4/oKD5BRPTiRRnHo3RSn6aT3NAelYpsNXTWzizxxqRk/AY0QDOejjI
fowLULjrBzCfylHS/nm6oQj+Gsda9Fh16LHRLPh00PohDR58NXRyEU9657S8Dlat57V0g1o+z6EA
GSDyQXfQKRQJmv8h1Y0eKk1fmzEQxIpwW7QNMXDhBQwtjg85+ivJAlZLjtuJPlVLTfRAwaBeGfIu
AS1fHQAqq1/diCoMV3X01sYP2f2TNXIrP+8vmS6JMe4cNbQnDTWt33gG8v+5OztLsGF65DPWWwab
341NUwU56jH2FJZWNunngaAKscKpfigSDrPSFzqN8PI4TdkFPYpV+561b7EInWRmRTPeM6wg6ipC
sHlilNT7Xy79J+nLVt+hDHkUAgzU0eY9DHCe+32vv40+Csi1IpOj/jA0kznLayvA1Eul1uw34IHW
J+2aOFIGQPXP+Pw8PEGwUMWNEUnXtSAzcdW8JslrMa7MbnIMmhvzzwDo9N1gB+FCWVVT5CIDRV+s
Jfphf68iTj461E7P7FxlB49K1ViD/F7SRwp0g5uUMyA+mYHB04OaPlTJxgWMxuw7s4AytNUcS8Zf
mn7XUbuEs1yxrti+hgAvMkZFKXk002pdVn/yQC4gXCWdHXdj9N5FhyL036GX+FLaNxPO/JFIZ1jJ
gVInq6SHTidEE+Fj3p/7DJzlHtP9q6BDjUsUPcjrsi41sJPNNOkYzHIF0G3pUQr3UWW/oXPo2+Zh
YO3MJJ0vXrJhCICdcL1SFM6cf8+vzEbIM9JuGSkF0xYNdHreQGBf2vcsCSfrF7SscX/D4JoPFKLd
cPFl3rY5nAJ83/NWROQmH6xK0qV2oartoYcz62+y/chaYj1fuBGotV1/0WEfWhyxCcj+khG8jxs2
C7mgzt6ya6VvFt0nNQKYD63TcIbFIVdh/Jno25RM6VZrFjhKJKjGpfHfNnD5hov5+g83d4LXAR8F
VMu359FZLgN4Xkzy2kZhgslHbkWdz+PJk01n9iURAkatVKJ0nNtHwfk65Haj+dZQkqhLKkTpd0sx
BFAHDp0EIwHXawZuYjNS/Hrw8SrVGp8pmjhIiCkCQ0q9E3Y8MJDb/B3IVMLJmua+GnpJ6D+pGxj9
UzT3ZINKZ9ue6Oo0whIcgsfR0+lB9YI4S8pZpbM3o29ueAs8SDHnVpb0vy54r9+BvpJ7D26nQ+SD
YPaTj7j+7opMXIhAKLvPZancyhsPAGaSjhTcnenz07lRgmjmLZ3AW24IaxOEmTouKWishui4FD9z
MvSuF9JR/vLn6B9sX5d01n2PQcaaae2pNFIsNh/tYMvSunNFksW349Zcd7pJdPlWiol673OLoEoe
gd+j7U7slMONe4ATbpZq2nZTmO7i0xTpJY4rhKHfDog3CKU0SIczskA7bjYrccGehw8ixlkK0X+0
ak6SgBK7Y1o/BBhoIKm/QP+xLr05ACuitVOi6cucnmGRVNT3ksanLbCJdMaskDGg0NoHQatgiNN8
7mI4ngJ4UpzeWkZFqVPiKDdW/xEuwPYskQgsGCqIJzTTBC81rzuME6oZ2YpB8rcEcvAtq+tE8hCn
7bnJK79VZkwZuTWl1MoSEYau9YYdJDtmi+7U8yyYHPXwN20FapbrMArGEimzeSqqMoJOiCUy4qVZ
2OcDwfTP6ysoHtr5PmFFDNJ4ISj6Jq0+2JQDXPuCz+Eoptq2lizEDT0ecHKc/HsMGdVn6n2Mjjzs
EgMtL2IuLzhkagRUxIbFUJa6nyjw12GeVUXOeF2Js3pcZh8A8cvH0rTeNhMogEmydqbpdhhLSFLm
+dzmmcKNyqFKFeFfn87YWpiKYcXRpSRmD6j2MLY6WI7aN0jFA0GnaTywzYelPr22olNR5hGhcy/u
xogSD8B2CNRQgl44LIuRzIZBOSmDWwNqBsHgCWPIgi17rclQXjWaiQFEB7/9UrN+dnQijqS4wYnG
VtDnnR8Ez5OXyxx3rKdESYFOVB3MJD1sfYzRNx2Ss0YHiIAxkys2HTFlb/dnTnPjUeRti/t455KK
2wHyONy1kNi3NES6nvbRhhzpsNny48yb2Qa9oM5Q5QaPiAYDFs+/1ptGZjrdbCBKQCCZ6zXFY97I
KV9U8ExnYtAbqwZc3bli3rLgtT5scLgm3nDmVx553fdkAz3qnQCKi79qacNpS6X5ogiVBjT/cC4R
Uwq0SC6RhRlIJFXxwqBgYFizR17oujJo7gF8k2rqLQlsG6LneeNcX2FoVs2GljbuUd+Nzt0rwCIp
YpGfSNbzIWktgE0RDRs94eBQX10lp42VhP6+ei7CVBETOR0GKF04A+j0HXQEQxq/EbMPgmb9QvH6
dTUO5AFXS+7X73pxfrHWw351/71dNBpyaEpEjYx83khLbUsVvlxRbfusV5GSmI0cdh270zVT6NBG
jx5+XKuRCGRWoMXOR6jmyw8NmpB8C0lpvbuAEAgemxZWLY95c2PXiFQc/BlL+La5z8UDGM6GOw3c
GbPhdi2YWaWqCw7UGj1cjrIyhlTxfNK79jc+r7T4AxLK2vQLPi6OkY12PNL0PihueP9hGxFv5Oo5
ZV2zAzrpCGa7uCae9XAh4+ywvUu8H9MJXqZaE/oxcdTaPakUv4x0cZwQh8NBEA/Waw+C87NuCvET
9bREVYf+mmOA+6UCdHXYitfhJZm4crCHcQ61TfPJYBtPa9ca+VPlPIEfKNNjRc9bGegC4m6zshK8
X+PR95w/KaXcRf6FFg24pwoYBDmkfIksmtWxZwsHdYNsSO+VU4bEampvynr1cuDoku4gx35T0WAL
Ie+wtFod3p6ZssbAI/Ix8YgsEZTC7ACJ5YW/R8SaPj78l9x24UCw1oPdMx7pcI2T+KZtOThsB1rv
Ggp3UhksHdFClMpAOoFyCTKKVmAkz8K7041DoS0krlqBsy8eWgGOG1SP99Wucj9m07fjXvbcBmen
BDCctEVS4RdNiNxFZ+OLKWs++mrDCQ6TtFbKDAw1vlmHcfnv49g//LrHpDoVgpMUOpcJpR9uEamI
fPlKjB/fmeyxmUqWTyVrBFY/YSOt/r8QTc3fNGKu+9zNSuV2bw6moQRDrwZYK+lZBVkKiRxXkMyD
Gm1nawY057ujLT9UbxICgjpkyOP1oJa2r7XCD9VFWvs0+pyfLJs2TzG3BHpyKdxiZbsP+bqGfkOE
EMA5q+L5cgDoE2KlrWdCLR7oETloQBssN9IXIeB5z2LsOkPaqj/KLWP1RBGFaIYRBxkZi0ardL7B
V6fDOBOT4ebxljoYZfFLxALC8/F1hE5pGTEg+VPLzUkKTY11EKEprRr/iqLufJR5heI8M3Qc2aNH
XON+ngUJQC6R6XFDUblCNi488/ruRInabqFqLDT62bbLtHcCbLyHYlh7Bg52Lxp0xn/JjhLBKtnl
f1c378Pt2MRvOeEZfMXqTMTCWn/JMhVzOcZA/5RIW4XcWvpnAZ+ykmUv16bpbntq1EbTlz2lprXV
VcSQHsEKW4zyR/M0eL9S+bFaDL9gMt48DVf4QTacqrIGl6ZEZE8eACBuvaW4BUqVRoBbzLSYtI/9
jI6vNAtxHT35FART2rP1B8k08a3ETGmVMAIjBjPYwf3MBlCkITRXAd/NX+aEd/WHOJsX4dq9RUH5
09WH3KpLhTBwOwRs9PhCcaufDCSZRbjNt7Z19+ItLfq0S51Mdq2UZveGh7mVTlX2NFDpW7GBxrku
gCl6jXHq6hURQBJ7nBaY0ZDBMUeJltbNWGnEf81aAMyc5fetRQ23JazEiQG+pJ562/QWchioow4r
HrZ1eXGMGr1fvzPCM1G3Buxc6YNTY8S61yMD7jdAHmKtCnhkLCCcQGzVP7NbRrfu9ak4Q51ZqXIu
CN0zMjXG+SXj3HhEETgHr9r7SGjLyFBPacN68uUQdIbmCdc3LcCw7pb91stL//CeysNU+wICV+U0
SxaIbI2IMfBrQgx9jKz2oQStF4IQTWW2yUewZK8R0kkH7eD/UX/xnn7Pmb37+D71/Vlf3nRA0IOC
Xj4ojSyYip3x0sp/5INUcUzxjLs4izyUag1bKbtnVDy47FwVMsRIXBGuu7vs5vMN38eI89vYrRa+
TtWWvXaskiv4Tjc6EmtP4N26PP5fdoaFY55l+hO1dWOgJ71hJ7FEfEQ7/HRsSxltBbshs+g9gW/t
/lBx80wkgl+++z6casP9gfwQJVeaU3hnaaeWtTtL4cKDleguvbaoI3TP3pQIqDQS83ZKXh/I1etW
4Rz1r0YHAWukMklL6xtpxR8iw0pnYebedZtmD02oBfvJ55yuDauc6qpifBuSHlOktHdHwM0scj7h
1duxeozNDrCrRtahdPVoOS2BehzeqlKglur3UHRIk7cyjZBzrY/JQz4a3hbuP/kuw/0dzd8whbkX
xlNwVY+7p0sgFAiTf9oJ4wLzTQfhag8DDfhsFd+ehhlUwUtxl5JDRgOYegWpAyRrqHFeIACRQX7b
UUGoYyQMTqWGHRxBeBSRMndSL69rsCFESI8ipDIEjXiztuyvRgqj7kdimpumv4kpSE2AeckbSVmY
BpGc2e17DAAe3e/lMQ19Lw1G+skzGJein1zOov5N7u4N6L7CWsZrqySU0G1MNdFH/2oX5TuPxLbm
cXo+6UW7E7wN3ZJgO3sohrLLRtAMQOJIqQe33+SYAnopcuBh1hEcjc8OFFc4UvbAHM7bt4CtM1Pt
SVnfRlVZyHRIKDOkE18Mcpp/vicG62S3k9liof6Q9ogVFn0nXk++3he+5yG3+nsgLjWs4wEmRR0B
AXDih4tiP+n4v4Qz/YXvOP7h0OekwlCShhyxcIakeMYd5EY4goeC9h/ZWZsmPVoFut/N63NW//4B
5gS2jam77zDc/89gA2tPksOfeuO3DVhSiH5Wx4fU3pX99lKcErLn48m+RLFSuNxRjsHP3wdm4rsC
g4LS/Td80auUTXswNNwwQTsbs/CN3uqdpPhMlRaHmMf3tEM5NodDDZ574HJ+/SyT2VSzpAyLSR1k
972FMs7jw35afPDu2288riY33DfZOwQWL8Nu5oL/m9lclgi2vy3502GpxUcMf3IAFwBf/RgX+Nnb
gDzQqJmeYbG1xzeAlSBA4EKFVdguBCRhqRQ4fbZ9n2oGDyg8LFPbZEeHMYTjhg69ubnIbSR2of4v
YEQknoCyZaq7WY/KESyoGkjl1gxGBNUUr1zdBevW+ZQk1TsiGlQlQLu4qQxzn57jA8YTLFzYKNNn
qZU5kIRZbK4p98ZX/5zTlQ+/oXPueufOpMKyxPcv5YU46Nz85ypidX4URo7x/wHa++MixP1HFxvX
qa7BaH3E0GImGqrlxLI+0ZpGUtUmJOZJ4wgmkdiMIXfBSDnImukobqKcj8lPLY2G2voJOJEKdJdc
LA3AbKDbaCHQVqAOYOD0J6QlgIkOwN4YTPIj4BusZjmqtg4JE/L+Z/rL+3LV5grqDytPGGAp3dFN
OYV5SOjqCgBdXM4abbn3yUNXRORS92DJpAeTA4IM5qyaxuSBfVMIs9peNNzVe4PpVOGJTVL/xyES
aoaPeYnC/QNTOv0PwUJvGOYwhlhyAqm4InOUgZDRE9ChERc5Y9PL+lN2I2BkPKhQwxgEvyhsdYld
VAzxXNzDQo432RK0/8kmRd1dZRsgP1j8GrtkOYbMgXcAf4GacxcH7OxZwvZR67zEwmgy5DaYn4O0
LTMrvnTrb86HuMffvzocjaeLB2srRIOEYtqjGE0tjoMy8+GbssEymrlDeD4mjEBSMOWPpX9Jz3hO
fabndCb3Nd8dYVRf5UvSUZhWvmaiAG3n+KNSEXQCVrsw772sH83cd2CfU5qkd2j2qfB4w2sZEPz8
Ie+nye3LftxfjJX4HU621bg7yHRRvmJ5LYY2xDKAfH91Gv0H7Mppbvkw4dRn1zAV/KMf0sqFaCwz
dgJpGlRWP2h8yE9snrbEfhWzA4XF2+Y4SY3L0pAX4262QkNk/OOX416SZ8cfIdcT8ulnTNhTgRr1
jMVFFanoO73hs6EKhhA/6QxO9sa/FEFDJeRdS7jAbXZbefSa1PalT/r8ZKgyQe6lm6+rMyGoxDqN
7EBrjtD+rTkS0q5XIRa+E8UkYhQOjyCdbhBMObcQEg4vTLp4a6Bx21x5HFUNMKeuvDKQrYzVbkFN
eZ0BcwAfDY8deNxps06xcUKg5ctF3qucZ/sWnIGTEbD7XAxeWfIWYx0O1bAprjmJYlXMUm5Inf9Y
f3lnRvCTifl/P0wbDmPLk/4RCP8yWS0/IG/AlqwWEOyLbgGwzaPx90PQ+yWTQUTvO4+fpp/ZClne
hB24qTf3jWhKP8kXRWVGMbKZsjpuv5zUR6CCZP/1K7tVpFfAuiGfWl1dPt7G+oQGG0RNd5eAYdtD
yz4QER/bLCCLQjG1tmNSyW9ktTJ75DVHTnozuFmD0ZszmF9qNjI/l935idLTGKHxFYHJIuCdHMLi
7CWEBcfNIx1ujZHJ1dzB7v7lmNJCDomLOiW3w0xWC5Y2yDtey0RUUQciEOXtPK3fKarR+Z+Q/l/O
nTDzIWtGrvAmAd5cMLToUzUFYfzxV8812AcsxfroX1A9y5x8lkhBt/J09VlaXfR42HGazjS/Dxfc
PRx657Wcl4ugaS9IGajcMLmWRyvjSYU4yRgOzy1WerWLFu4UTVs8X2fhCN3pz7sziTYYVzCjkiGz
eF3tnKAdoUu0sgsJSTsXZxgxn0gJaiixtxlO+BqvI0XnEV2C4Q6tmoMV7vGg8Qb6sfER1Dihczrz
yA/b8lPd3gS7/GvtyUEKM+rwGyeAyW2MNvAkkxsRDN8Wp80a99cFbdTLY3HkoaX58IDglK/jw4W9
OEko0+j+9bdKkaVH3NEB7K4HKbqsccJCj+YgLThLtv2Hw1U60MiyoY0X+1Vx8EO0u4zgo/jlfPaW
IVid3w73dJNrAHbbsb4fWLxgY5Ow2eRkEe98v9oFWTtooqbfBzW6zHSy5JjiTnursQWUxT0+fnXb
8+SDqNRQ9AZ9TiEyCLM8vwYOFfoYJZntYA8983+Qvg5B6bIoMSOUwLbNzjpeKpfhNmVTISmdUvfM
8yyRtNzGWXm+krIjs2OI4HI9Rq3iVh9j0SITvrgMgaEkYpPdNXrC9d2psK86cKQE5aNLoYLWIkb9
4Idxqhy0UuMC921wF/cIRo7nm/43riwwv80wpQJCPtMn2c7QWUutj7NAIbCCntAYz3o9mH2EqDHl
GgYFN+fD2xmagHe6m0oQeKsdl2hX9TrtgZX1HF/FPVBT0btO5WMwAzPUPvOsoDgIMkG2BmgDKTzT
S6+wlQfvW4dKbALG4GrZMT9gMxQZlBIyDrHnKvWl9Qur2pHeeepoQlwJZYbb/PnztggJ5O5wXfug
0ZAJ0Pzni7hMaVl6Qbszzl9qAKBzCnfTTJp/R3NusN6WMxZ43Ib8eUB+3elSxY5vkjTYScaMGPdn
T6gaAxz1wnUI3L+KlZpq45ovFLeLMbAKhxNQoatjWF156+J6dz0WkkXgFXfqoAFKB6Arqzfm0cEz
w3EYpIw2qF4x3LmR4jjfsFMIkjLRQPftCu8tXFsFIyg5rSqFi7GOkaTPovU3lGXukoTTiBt9K2mu
2HW4tKNA0TXONYmrWq5pt46Z0yqdWc/mcCX2HkbbAy5coRAjOZovs7TH7ZbzQa3AaNa+KuaWu6g/
86KV9vRJOXIgNBtJqsphM/JcBgLsRNUwI9iIUAGi8APeKCzr6EURnJq1k+gcwqkWYX76gCElI8k3
FR4v+XTWI4PLwi5WTZ/AvdDdgp74jrdDFv+GYRveQKQUHlBaiTrbiKTZKhYTVuvgxO6c+Ve2pI6U
qwbiwD1zb4x7Uj2ybYreWPIQYhx6sp4BOUTP6Ix7wm9G+zbYJXEKCCB5TmDHpqKLBmJ0pgZ8/Et2
4XFSZExGvS+Rz6VMzXt7ds0oR4rWpSRChbHMMhq6wNvwF2WbzkBVWT28eE4EIfvHGTtTOlq0N/8h
+IsPahCWzhzdmJa8xl4N8LwG/EmqD3mP3bdlB5VfK//cJOqMjtGug4EFqczRw0gH6VTKiDzeBVe4
zhFduQf3CZFRWM++zeVhlGZ3/Ap5iTjqb9AJGAUNjkOHdx1GPgsbmma2Zd7T9LzTaOVva0MWD6dw
dslOMiczXfReBnGcksphRv7gayJdTEMXOpjSFzbQptYHcyuLDrZ+sQI5W3l7hr2a6jZG8enIwexs
pfRFfW8+PKBRYPSB1ArvLngSfYQJSdz9kdXH4i9HFwAlvzSXOMj+4D62Z8z69bAZ4G46OKE41HNI
VFyAU1YdE+GX9QoZM+qxr86TTgSb/uwxFWBaJWCV6nc/jJUBHqomdOi2I5vmzddoFBNmhQI7Llin
zJCfSNY6hQrUW0v6tvM/xe6RqpNnifEs4schTeOaRo9PlYdVWhM10pOIwr651tl6bb18YcXfmB1p
FAGeEG4ZRRyeaMFAvO2P+b0RIQWGlG5JZXb67rz5JRlN4Jd23LtSBl7TfAo27CbjEBOkCXEMyifB
ooH5a54iMKTA5mY5Xqt2rh/HHd1Av2uhkNYFqTirSANEZ7NCqZ41MJWARVd6HmEDkFYw+iZb6iFh
kLtGLwOvZQRtPxQOBrN/P/GemUXyyEtFq6N2EqVyRjnKdZxCWmT8VM4muCXy6MKExWvDXWaiwnC0
1dEb7pPLMm6nAvLwOTuilKquBV8o1si3+Hm+yncyBwL3Ac17THS2ciaUIEG7d6trrCm1dmZHmwfN
MtxBpmlXYKNBtTXF4IBoY9cnoiQCFrPlyBJwzlacuG/bc7aMk9vNb17EeAxbaGHuhq06vhmosqv7
1k9eMefxrg5tLDhH6yqYrKNXnumCyJ5eAGUqSuk4RzrGzDHwhYZp2TODBuTdexYHn/Oe4pfr683l
w36bd6KRLn5weiQG8h5BU46SxFne93XtvUrVISk6h/dFq0fldsaPj5dHHlO4P+54nVyUt3+gCkqG
7mr73vVTqG7pDxl8iurvLdZSRrSDPqMwEmCeAwMtJLY3EwFX0OYfchLqgyOcwHGdjdoP1mhiuSH6
Aov9UnUYC+wbyDlr/AwA6HirkAeUp4yFtVPLQhGcvQTQyq78CjOEvK7Bl87UVz7K9oW2+2mX0igJ
WDoRLUissuO91UCrV9YjEpG2N4UI9imr+gMH9dCh42c+YwbAzXF00kmvMdUxzthu7EsH3yV3BKLo
Zc1fuxI4VvD5QyCYXgRldGNns9ScRhFrTBQcwR9HM7JUYEhqr6yq7r9bBMP1zGT9SB1cMzv5z8gg
zyAT1lsm0RWIEM7dqlJrJf7kC3EIKAQXaJCtpR0prInyRqL3WxZPCJZbZEGqN5t8P5I6TDWTRYem
56UeDi2E7szw27aJIBr9p9qZTvMI0YUkE9gj+g73tHYOAiwyVoAiafGkkUjt3uejKejyoDaxvqiI
O3ne7QfTiJtG8Ym7jc14+cLiM13pKdP21EfYhvdRndNs9AvQ46oBmJGyEv5449lxCADGiFAtgMDl
39YhTTr+7Uhd49ObSKYEVjUjt2rsfgGfeOeB5z3hT654HdvXFWKySvEtXVHEfYWcOjz4v7g7pQvW
O4d+rVZ4/2EV++0iD2oaMAXDAlilje38Kwztj7chnoF+f3/wM/yWDQwiIOg5jY75b1accVkm7Pj6
uoBfD+k3wu+y1va8HSoMXE3Ylqrgy56ff3i/lX6dffqDT0+FknyxeVIBGG1otwnh11vHRV11qEXE
nLfBJucAFJ3iSa6A8lT93UdsIlCXZcFMbCT8j3eUqbKgv1+JkWJ8RBcS1n6E+tljQJT/9ntVxFkA
0VXIw5CrnB4bT125iXArGxXNtEyyNiHFLVhP/3z1nx/bUQkFsXRGU4BgOU/tHI2OL76RDohbRxgJ
5KWSfn+vQMqUe+3L0YPH+FfC1y0e1J7vHJr1xFX/+Q6723LNbjym7im84dlOEGiZBjqPoL/Uwpw2
Pa+b6I6aSWIkC02EOSSTeabl+PnUjRDj0bNzszM2l5U1S4bMVbzbSl3NcmYpsRL93K5iKVkoIgdp
dOD25LkgLTiNlSBb7udJ5FZeUUSPM/KL4jHPnNC8AVohAAci4qF8Hpvg/LvkRvF/u8pmmyGu30Cg
IJOB7SynTgTAn5diivpH72YhcTaFBPe0KlQGJMeKrezx8uyu/Wg/SoRMATwdQOGUPlLkoqpXpqZ2
WKEdMQksBGXDRhXBujm+LgeS2WKbNCTagqmHsXKf66We8c6BO8finzmBCdWHJ/xL7P/woxKQBvz8
2H/V7r8flgkw4KjE597G8db4C2z+bZOsIsvk9nM3PFlRoqxmTK8fDg1AbExNIBQCqC2zT7YwwVDS
5b01tiM7hHd5o5GDYubPsA5seHjgVaFKKxjcv6MbS/fYDjFHjziqJRhQj+AaAZILxwBYEZ6aEeBc
a4kTFjh8ZtJE0JJDWW06BV1kKh6tEmK7Ds87SKdPjH5g6r9D4TqpAss6/2pOWUZmrcJdDOM5GU4h
zRi5Rcbvq7Bf5ITfMvTlGZ8ywUJQbwMDsspBz542qmIXa0ymIpujkccqHI4v+Yz613ppNZVFg9zZ
vVoagxYAY7QbtswFkF8vvk4j19CaFvffVa+2E0kusfmRdeZB3S3sDrS4W2CA34BBXSKHFSKtFvD6
rjoZ5mB8eknUKvInYz4poxV62Ysp3nUOaYsa16uACPN1AkNrDx05YS4lDmAsb+R1ovElnLvfBG6m
tkbaXjbCpdW2msuu2OfR4Th0vl5XavNPWgDrRq2C8vRgP2B1IL4HGsq2UMKdGTCdFBQY4IqNjCxw
EvGMpkdRV2XFnEhO5dDUdtzT31qafCeTC6Esdq1B3KYLuxnuJEDhQDLQcd3GtyVFEx5O3olgTMvC
83pf06edgn1HWVzhhCUnFhmfsD69EZ+Tf5tjDeEL5Kp+mtZvx/jX/bwhUIoR0T/Uujn/zeJ+8hL3
WiCkffWfbbReZ/gdaAhdqIl6/frWQ+HECYXrGR5hcpjtpY5IpDOz24Ui3J1NCwlbqarV8OdEGtz4
7QkjiNai1o4ujslQEud/S/o/3Dy67jvcfwSKC/aTn1HdnlETEwvqLn8WpgjNFcCX6MH9Fcdfa0G3
J+4Rwp47b6vpo9m4TBCVbi/PzzfL5I9GjDoPKMbpPZteoYnPHQMiYim54+/v+LIPi1Wm8Hq0aI3u
HPeb6xBPVDwBQ05DpyC8AnhI8SFi7UBcM68TNdFE31WSau3pog8lx5UOis6zkU6gitMiQzu/4ysH
j+zIGDUHrufLFvqnrn/qSTfmasrINUW6aNsvDW1vmVTjzr77jb3Cua7YXJwnPzW7pZJLi5+FhNZf
n53MrjLaOetytJb293zDVEtPyw8WHwZ239YWfa/tHL1D3yVF39TzmheXGIIw9fG1S2EpOZFEZ3Nz
hex1xMGhedD+v1R7HdZHlzVdajoBjnbzEDX6PtZ9c4JvF3xxlzi2fjYsGlTMtg8398Q3IFBSOA/O
nkq7XPZjj+m/++vKZ6YxBMGqkD4LbbUbbzx/tp7aXqVXhCzRzmTMevLXl/3YKTEB8FrFUnMRCMS2
QedyTCXy0LHlq2ta4wrk+1mwj0dWD07QNMoiX5uaJ7DtQOA8uCNZbMb7XAM6jKlNWjqwIDhGzmwg
j6pnHTzjkFNJZiFQdgFvGcPLwsMaPuegeDv5z+EgAVitwGX8M1gtRn9AAioUnDUA5Ll+zv4fGBq1
w9osT98Scu35cXCPFN3D9XqWTsVSex7Zz1NpwXWZiVDz1N/SM/ROn5VzB3V9yo9IItI0cXF5Gxnz
2ddvEG0/dcweMtxIeMgLB5+69dGnLk4pYkAc+AnIZDZfptYnfkF4z2SL70buslH2iMlcZaQwndkw
lyKlWC1EQXIwanM1o3I9YsQ90242YG7chk3g6z0mp85a6gK/LRMclv2HrXXdTmo9m6ycwsrA3GEW
TSZb804U20E6aSc0leu1nCvilPj9aJjpYgQplVTW5pH+n2ZohsK2aY0kM6eYsr3j8z/qGLrh5K43
Sh4VBfe1lPS1590fMnO7lgA/pZG2DZ+tD0tblDGHHvvnW9hAz4RI9pnKiSnpvzvpNuVMFZN6A1P8
wJWP0/3gzDRMVwELeqzmiLgZwumbiXx7YHVXCi7McGLlT6O2E7jYTd/q2PsWsHoDoFxt8vvFr+1R
UQLD8ixIwkSQfEc87P86K7QPINeyK6XZcuPjB/zoRkJ67B1oqCncS8RqH1PSJYsduL7Qy2ILpDYR
7LXpGvOmkP4pR8NbJb0f4TngUQcXxJL0/2IeTn8nagAOFH3gLHXOvtNLgQ3eOJAabN/F6Y902V1N
OfJTAMhdfZ669HcKXZ4VKnhcAqOuEjk2mekzD4QIWLHSN8P3BMyape93uChDeuXOHixqGzoOpHLp
b7YmqKq1ioomNJJkjpVlYRqmtnyPCMfvLK/vM6dwkh6iGIgC0o7eg96kmpO+cEd6qyXR2Kexaqvz
BtPyynyfDBaryb4U/GgNkjUYrBIxb3Sp9ZXW/kv9vMSpKu67+VhBjNdivy1gRFRBbP/sFKo8LbAi
rWKFftZUOZ9QVHaiNPmHKmaiaBhXEDd9PwC5EyzVvRUwwuBPub1SMH0y7hLfO3v1H2wQBHvRwWPX
tzOelzgatdwGMaA5lI76bIRxcnhb5HMuyzEaKQRAKCAcK9B5O2P97D+zjfjfIn/NMDSd58PfSYXI
cOxSF9FX8HrO0sAjTTPOQxK7Yshr1SgjXOGPgV7zYqUCy9WjyKXdV3l5K92xVYEjhGJ9Tbhdq+Qj
pc/Wycp6/rIpS9QA2QShvOU4cYoluX9aeD/LaS9n3Ak2lv1yAirSkaXJoMQKb/p3i1jndQSfcmgY
ELmFQ3RjG2dE/7de2Ap94kqG3vCT0aQhRIth+PEI6zHfPIuJsmx7/XEo9uVx0R01cIDt0Qfru53X
qo3E+RbJ7c0BACS7GQHmJ/Am0yYnEnGBzAFzm04A3SB/hy8D+xr3bDbI+y1tiHsy6ondVtImJKaI
dOMWLt8Q8O5wei7NcC/DXULDaySMEYxDTjt3MotmPyCn5mt1vAH8z8KLHuHul0h6c0TbQCxokrxf
+tPSz2R4dFlOvYkaJgttGlJMzPz8DXrNyXcruh2x1cyyGkNyV7LxmIymxyX2McsqF8TYtKm+z63S
+A3M0bCe707OcfTS+6uWkVVy4bhTmNZM/n5RPHkew6BPt3oGLYFZpLdc8mXFt1gWMo4/4zYxtcIj
5Z+OufDX/+mp8GuLr0co5RwkFLjZVDtnG8zSQkwMC0jePtgnY8RxvkTnmw3FAGkah91GmWKiHBAC
CSIIBEHGkn+Rwuz/5czD4CEtw2AX8z6aCNl5RL9kaMECj5BOM60RVt/z3ZyXqiwAEpD5wW+9rPRW
hqEzUHQBbvJ9PjDl/+nvuvob0yC9Ym0zL24L9KvpGsqJxQZv5z6DzxbYUvb3BBpAf9eXv/TsAWia
r4x5cNNPbzjlO7ZN0c04ygooks77mtPgimbn4rytMt8Xq3Z3ULHQuLMK32GNHM7SqwJSB2zEhBKG
qAWaE+FEhG2SczPcXLMQpyclEmVVneLmp1HZd6vWombmsxK2bm5hbG2a6eqW0IzHCTwcKkwz6C9L
UeWUecjaF+QxxorjE47W+vsWyFmOZowkcT5v13Q0A6f28dBgLOHePeBuvkHRs8RfNzbCnTpg2bnB
cuPrIu/y2puxq4r6/tU39qD8WI4WEwqOOqo8LGcUP0UOhs2GVHmWkrspxkVLHxXb4IqR/hNx0HV2
OYx4xHl9bp//IcjC0pD0FhCkN7s1CdB6/udODpNAiaEtx1emcVI0HUJucpGzeLL8eOOEu/SsKb3M
N8/FX45oeJRt8Xu37OJtCFE6iFNNoo7q42hDBhA1FS5ulSp2LhE4vM/ISxyPONr62clnj49giQCu
b8BWUlGX48uqCt3bO724rGBqTVPXAC86IMeOakdoEKz4SNm6eJeg2nyfPPXbPFng1kiMpeZpYmr5
J1Ei6y/mZeNJqwBn6xU8h4RL/9IN2+cxeGoxgcVHQiG4gpJkjAcI9zdvx9pSo943XbCBHidbH8eY
o8z6yA60wM2HP4gFj+7fpp7ctrFXYnjEKLT+QgaL+yAedWzV1UvMsb2fLbHWAJ1o2AqLFtgL78qG
vlH/Qss7B+Ykv1jdKRWokkyWM1WdlQXtTsX7P4C3gXF/xvnurw8pSQas5bnQMH/qZ3YFGB5xXDnf
laamAS4xAcbostK57SUBEDbg4nXDvj0FOW64dwZo8m7KSwxgzaDTifC0ty+0Lm4qqN+ZkRGrt6cP
CyHk7zSpVTKqmagLdPn9PiVEbDoAGZmUKklnT1+Em92Teq8kFMus7yYcwtHxvV8zb0irzaEDeZP+
qNnlbp1GyHWuNI3nsjSGv9OyPhYZtrYQHxh5otRfxOC72E8VVtcP+IQusCSn51WkFqIa6BVlx6Je
0W9OPdEkcA6cCnPBkn8dNMnIoP8uBUJGAloMkc4VeiM9QoIrHUSZhGhbtDqletQDqcV2GLCxo00L
EO7ko8Q5qFqNVrlEkVnW2iFAz9QJFTq1cft8cj+nSGy15N3/2SosqOUxTbmFrJ4NLbjPHTU8SsLU
QsfEuIVP4GOYicPK+bBqCUiWcqy2nN/Y5WYl9SbGCM+aoj/9pryNN4D2+FCY8vKvgiYn2SHyp4YD
4K2uz6Hwe6Qqgj1TF2rOIyw1KClY38KHSUIQkKkAZ621xIicCMhw7UF3g2a2dRF3IywD7fiV4rP+
43IOH0O0KMPuYn/Jt+3zd19VEeo4WklbFxoiTZac7A8ZvKU5M1A9P/BiVqP/jGHRR4DGNUmygsWR
CxLHMVQddhN3P6J/cIj3ZJeVCXq1f9tSYCqKRZdY0RFUqaL8Ge6PRP12g8jSgqmcYHodhaA6zEcG
wey2l7GuPnUdt58/Mb66gkNSk9vBFjPuF5slMdY9MXz+dRobW87se0PbOcRCb1j7B0VlFHwarxBw
2/B4e95glak++7UJL0e7vhqXBKuxH7L/4mkRp/AcVwDZOoK8U8uvzxLCfNwRAiM4h/jv2/TvYUJZ
gPUruCl5RLnWABNE2kTqQ5XrJwv1L0pxW5zg+CgIFPRFkIVMRfoVk5Nk4f6hKK9qJ4DjPuoSsK9r
kexbv7vZgpzNwnlP5APJJY1peHVEi1hCQfTxRRb4dTllq9o9tQIg7tSLfX1IG0EaS3c0RACtyiHL
LvL7DzyDSjVojZtTneaIteOTJCAkabdVfHlDG+Y9q1JlF0bUQ+6YTForlZ19HFIaSPMk5DMS44LY
jCrJvrj1UlCvgFvM0eZIPLVT1E4WpM4YlSp+GKY8fdFZ8sbiBnnHvUGIAGU4yHm4xuVNbtY4P36f
cMnXJ/0Ayjd5z4zsqCSeOz9pQaCxUgdE/Zp4Ab/UcuWXLmuShfkE8tQs4na2VmUck3KNBK0tcafk
19fnflLShNL7EGWDYuVdlZMxU6qaaXvbo0gSZ9SMh3ZZm4xhRX+glWESFL75qH1frstBKgj8ZOvI
eeXCBenpSm5OgdJnSm59X8Kl2YTtbWva3KQ+ce3M9v8L/lB/ZAVd47N6NSb5zJszeUGmi8OG4+kg
kATRS1h2Jf5ItPnpyVNqlyrwjRQQiyw9ZYurEzBd8HdCbmFo4mUzZW29ceZnzDfOGYT3CFGeMTG6
Z6ZRuIqUkCoUTky5lPo5xmPy+Eqq7n4QMCygMURW/CaAhY8TFSEJ6IhqWJ+nANbD9vj1L8VOnsUq
OWEYiNEjJqsXgCpfSEua8S0033SczCvuHN3Wb7sMcDjVhxKO1ff07vAKNHxAhH8uf2h8E0Ge5qI3
mUW8nFhA27XoC0do8DXq3cd+j4pG+XE16IWyvpT3o60id2TsOT6FZME5FCEI4cNCka1avDMGCkuO
yNgIuRkOux77qeZ+yVL4t31J99hZqyohrGGjW6vAivlZaKrJo8huAibqxpfLxXRaA40qMqPQG6OO
aqmEotte90xbZDNMm6Ep4Bo3pCj6fznVdKNnmWBUFZOq8qdf30yLng8643LNwHXeNjdpjJ200pdu
mlc6TaW59w3xlvBOHGC1PT1c0nWabHZvrunknrFJ9aeI6uZD4sM27rH8g9LJ/u5p/iVSmGkJtc8p
I4YeiL8NCMaFTW2vJOBKi+DiY4ER+w87HIh8keVXWQPhjVzNqjknyhbHz/DnQ4vPkk4d72NLocXu
1/e1W5k/EM1hFt4XcFKc60jwpVibmtfFZGuvYBT5P55QkbCIW8cgJPjfIvURw+sk/0ghhv9qmbAv
INTRyfisQecEy61fbCelNptzwiNxB8VSyb+544ngCsVcyWEp6sWGYETa2S7OAX/E9pshaavsdDYz
FF+Oe7OsenVZHU306EyW3hGXyU7IxllJeLvb/lSYxYGU90WVkFIcqhMbRu4nvhbmHGBEDKPKGSWi
GsE7ArRGVYJvKlAOGWm7O5HiiE96RCURulqORe5krnoR84Q1xYOKZh5uZ05s8l25gnhgwDbplreu
5FeiGWIQ17t0z84OYi5PCxtdQ/c1azRwPMKULqcjM3g1xioEsUvoN+guJzCEcC1rpsY5E3+fcWEZ
/WlETmGebOruPnBzJiGb0vAG60atauqzqM8ErBkqpCjawWUnZq+EspwIWnVBCyI/A0+48iZW9bgj
oXghcVVqcGbd+kni2pHuB7WGkCRbUZ4sLrbbrVwmpkQQXLsjcP78kY6tBBd7+xo8l4XWQr4sLT0F
CfJIbZ8PtkfaCUHomtxw+pgBtvpu+iRWSk5V95sl0VSrXPzMbwFC4/up7M2jsZGToGul36U5tidq
1PyTM6O0ut9MpAxMAjyzksspVlsSWhh/F0HpTIhWkeruJ9VwSxbHSQNiuv/9CldIfy9EvbIJuKYH
SBsUE/M1JmBkh8KIvlufdxrKe6gkAar8gSiWgNjgqYuew+M/OG7ukeTxmi9d/2v53Pb/CDVf3pyO
2I+n3mcE/InP6OEdqTT3rnk85YVDqxS3C7QrkPi/CEiJPi0iN5nICPi+yhMthU5Kx8dCCW0tQyH4
+HWLtjurUSz3rUI/zhTIq0A5se1AUb52JI0iaolXs9XfvHNJJnwUJ4w5VJ4c40zbXZgYKCAcvalR
O+k/8wHtqXEIfEsDMSxQH+lsLewcrqzaHFJrDZoGOdrx5Rk4P8N3n0RVwAwzgKeh/gpwCd5b2azQ
HbEo7wMNn4zBh2fP7Thl7KbHHpGFBdANpiwQHcSviCE7e3I8X1+W3JH2dn7Dek14GlhVJeZLCirC
QlPhW5sJHm1jmRIH9jjzk77JyzWCgpjbbNlgXJq84Bivnn3Qd8NxP9nFyB9Uq2Q7ttx7LdgAgBSR
uIu01CqG/iq5+65qjy9gUahEV9IP0ljwYv9T+/q4XOzEUD0OdufrbtilXdogwU1LwDrdjcRK5wHO
F+yUYezi1XQC13jrQ8hh+IQLwGqLaRUx1Ts/cHlRGe99TLAJsGIV5en0QnHs0q/sL3uaAlHXH+dr
mZOs0rHvlXgqEUWHhm1aPu9rw4RLy5FmWdt+BKkBGo7FDr9hRetknWYNXdzGNHaNHuSMzDlP9awe
vzP8NXIHElJa7E1ogbr0xGFfSOGqH51z+t92Nc7PTA148n+8scZV1w29j7pQ4bp84Ky9sQXhcUYk
aJpcF+DnYbc0kGrH38GUrDmy1a0vpS+cSGLwxc8usZjfbXxumdTIejVZoWPeIE9ast1SIordulPP
7Yvc3Hlnrwo6+PEDAEu0PxUo/ikNs6fvLUBhQo+1h18bjfbrJOuVoBnl9YutJf2s5dzsVNiR4Etg
tahPH3QWLax810IAxHSYRu/NheAbf7BYk3EA39hdcjoYTC7g7iXCU04ls7QGE7G+Po0r2zOv4UQt
I5JcFQNqJyxT1G/OpgBHpQTm+5+oxoLKZbnBfKU2bBAQKme3AIsfMZ0mJvkoUVTcBs4dxVKObaVn
41RDlGZHR2DMxMxHR4IW0ezoyKD+a9tFMDfBSww8BAOEyF0ANaDrxRFNrPxnea7kFJfd0sbqgERQ
cZHQaB4yiE/B9grHiVCWNAl4oMQnsbez2i3IH+O3/bTLt9LIBp4MFi/cGek91Bb4dtAY2AbMDQu5
Y3N7FXL4tnl9aOwsQLxOBcFxn3S8RRdLGI9kF+qMK57xu1lTaLKrygIUktLxjONI2xKyLLnwI98s
3aajGaaipTSqGbex28ZYgpsSg1XexKWwI1WWusGTeCcFArwtuNNe/jJ1+mtzHDkkxtMINbKUzhIU
Qg1cXlCl78EL4D/eiKRRfTTeDIUwWaZ66W24lY4isWzoNKkPjgk/L4e2NGc1wqldj76rczH21wKV
Q2fK2ezgXMBgWY/5ECYGLYMz9dFjoRZK2G9klW0uMvC0qIDJCVCLoW02wbm6GZCW9Qu/PuwYnZxf
k6J3GVff5A092ChfPtwAqJqJm/93+2Hr2MjKr8dK7gJjeJ9tjvbeqPJ35vF9ienLOJ9gme1xNOVj
D1zh7ZftuysFTELLghyuqV7TRhCuacYILTOfB5bO/gH3UoFaFdNajoOYCKh5KEd5CDUwTC0J3sXH
atrqv2BA1Stbat/HKTR3Aabn/4xrqImdBlrLp9Aix91t7MlafP94XoiL44u6RZZdFtzvufHMNuVt
grzU1kalmmoZIjDf2In1MEdv3tSgNiGwyzcw5hLEs88Jpz9PqIZTQk0wzkCBkr0FGP27laGR1LQG
hvnawMUnCgojrG58WsnGs8VtORqDao/QVEZGg8+pzBUs6CZImpD6lj8WV+IlYHUCTca21YC/hth8
n/B0Dt++CNEcKHlGUPEh9K2FJKAK/nlSHBeV7CSWaJeHRhKQJcXkqDbuhNkNAjFxK5zcZDrq9hUe
qAhMZuJ5hs43OlLKWjC4BZ6Lu5Vx7KvXH8R89eJ/JecqpjgZmcb3udXMZWh2l0vLtd/Ok2K40sKo
113tNWTEEfR+aSZpdchC+UpE0I3xURp5G7WWtlBRbN7KM31Ru2ahicfEaoC+coxuvvX4ZaQgZcm2
4DjRTU0ZZ9Am8s3aHJ+SLMElqoLLKpJjkGYEDktjku5iPJ6btH0IuDJ9GH9ttbvaHhflOfOwWTew
kMwSAoNKcXKltjFyNBWiIq3d2RP3xOAmyTQNVF5qd+3rC74mshlqJZNFbLdZvY/i0zEJU8N97nqk
BwL+UwWulojwicbuhHvU4I8/Wy+RJ8Q2PZG97CC+bKkjCgXZvG5Kmf9dEWEpmld7EfI9+EUxMl9L
oGE1ps7RqKzGHRM48C8mOkT31FwXcXsKuhzMfX0nbu8A1IKcOY5JXlzgRk9cnKlR1/VnTg0RzZy9
XQsXZP8z4W2j84exx20PHzX5PgfIc2okyvIgqUh0zlOfQBKvNPPUJgWd/fQouH9xBtswp0SEgzsF
6LdjbNA9kwIzJHqob+n8XIsb+ecZ3ZjAzu7oTHzUIRRrJkhYFl7trg87cYJyT7yM0uqJGjTOOe3f
eQZsmDwljOQcOBBwoJygVfRgTt7BKSJkzrbQf1pgHEjjSQ1GBBEmOwf2iISTqln7KVWZQ31r/7uL
LZnhcW9gyhcbgxIwYbZ8MMSz8ZAq1sXTdbW506tYAM2JefcU+461kTbg5ZjhhJcfS/stT8okGomI
Gx/QZAJ/oalrgyXpZDfI7ZcqFE92zHxEfYcvT0EtanHh8jbd6h7VEOmYbhnJk7c3JlIV6rhYoRmp
L9Liik9c3ofhCP9RF2h75HeGc83zMtalxIQ+4rIkTWFbnT+YLzyAprNFhqGrHJkUHxEkdbZ3fJZy
P6Grxs+Yq30SQrfPMv75xTZWEVR6ocr8tJgUaEmk87bVMrZNOKHIN2TWQ2KTOSRLqxWodvTgutnr
FmnPy9v3qAwDTM2fuKTAx6HiM9iYcmzbQFbfZNFp8p6jP6Ascz4gPpU5JNUIZZY3G1hXgRV/6XwD
E+uD8SsX8exxj+cI9wrRHt8YQCSzDn3VqgFQoAi9nDYgvH9D1xFHo1HeSdr8QHx3vkC5l5YLjuFy
z8OYnavgo88DZZ2fo+Cgncp6KEHIK0oC++Ru5Iw0zviPHmyDv8QQeeuv5xbjiPsg1YddA1s31Djk
uOcEa9MKhW6hckDI+BI8Ken6wfNxnAbfl9aBOhtL2omE+Oh0LaEyD+AqUSBLogaQg6JiqPqsd+Sk
alJCy4Lwiufn/C2K25Y+nPJSJ35s6FMsrtWRVFdeXYQEdYV0SG7FTAwhOzCy/VVReoz0VqE1dfVX
9HhQgQVvd+1Q1jijcvCzbKpYQ5HwNHFN2FtRNxLxDCYtd8/sw8fqJbGlbX2afryIVODZrCuyTO4Q
OuFasZSytXeVPgsO8nx8yox7hefdNea2/FChyX7vXaSAxDj5O9m3evPofhw3jK/Wq4Du//L4KndP
78Ryqe3mZaA9xb8i8ZkgGeBFGAqNX51TNBTXqmdb2Je8TEn1EC1zHGAW891Bnl9AHLibSZ+zfmSQ
+YSWx/nFauMlTRsLdM0Q+CXG4dgy4aayzeBsSBmJKsagC5TGmDgAmhv0wQHa8Ei97h4GGfP0V1n0
/9dqvr87pb0RZdEzyXexhSbfvS2dXy5sgQbDpf7CeYkqRx+AJ1mHUE9dzsQb/wXGuNHP48hg0Iji
pr6VVBIo8M70GA0so55Q6mgUCZBcN3gFcLysEVeI2UarP+axzlXucqjGKFVqRNpBRnR3RWIQCMFM
Bqr/z8Fx4HTqY9d0njtg/viSPIktJUS+quei67XWo8W/YQwbx+43JVmDs3gcRBUXO3vEYWtjHLLE
DL7fI2Q8KLLmx+y+IV5RYsJmiN6Vs0FI43XXXA+9rkPjMFgRdKLylGn5KodYqEqVEyss5vS/BjYG
XszUcCLFHpFIMo2KPH+r+VGzjZ2t7cFV26RzDWLWBtKd0G2/0D6oAsKHF2lasyeFQ5IsCBCp6Ltd
E5wN87S3bGlN8vAtx4hx7veMWAfelA8KXFpJYIkabIdr9n9NzsmE4xpjLrI+TK4PxpV8DAkNo8sj
iBt2YYJ6l6+H1kGokX7j1FewP3ru09kUQVxRfHS+X2MoeQVhZMToPuUSoHZxsJynnTtx2fvAgujt
52C8j4vKrInA58q3Mrsk8yBAF6egkQpGLcNI1O2boEAGgroVOM5tAVpo9D31HSriRs2wZLTGSUE/
/qYyNIfmzW+p0mM+RZnV1X0ZKWC9sJ7qDBxkTMwZzUn6ZYTdnH2kKMDjB1d/KJ+1qU0dhFKoZk/U
mehCwq7aA6wzw4B2urpLbuzvaAutXHSItRbZN9K5U3/4jt/JRPLsyq85gctXn1cFnxSH0gtEkB4U
ryQmaEMujUO+OiUiEf4s4FCtbKqKpT53/z+iehv3xFHlO8Zys6VP/wSHdgLUWvVtUVzXIWtODIJ5
6d2yutPMWKd9zsfJ/mutCRwCTxbNmsr7OBNkI1mHD24ordTWQJJl9x+4p0VDTKREHSkqEQY+icz6
B8U5HiLMUqlZ9NJ/NiIynev7ULx20pvBtEx6vxGItmobpzXHOTYXA8Mz9wVdGwJHO3AOH+l3eFIM
bLJA75oJptqXkimFiv/qBas9eGD7WxqdxYoqpKZw3oB8aNr4grTlnJb4psAvFzvfZ4PnnJCEr4ib
3l2XSmeux14/J5TYs+Exlojjhp1bcyymasMZGCI2LP2JvquqRlASq20ols4lt5b0q4qjUuvExI+8
Sn/HyvR6z/TCYtfxmuqldEL1P6DVp33BjxMTPzpjAwZGY0YrKteoSfyDI3MAs3O0Wo2zRV/6PaQW
Xiw6YJ887e6FdUi2evSiVPCDMQ0RVIBkO75Fud0lH4IUsYlRDle4d9V79/b9vKIRmVi+QBgJOGWR
vZ6tOEqei+aRtx7cdg3ozYZns8FoXxwwn1S3NCXPwXEGKhBgcr2x0LILrMLUfcJBM6YZ5lQHzqQA
3wv6fSHKQ8r7dnXer8KXuuEk8SfboHOauEUdyELfSEHwjNRlMDbnObJCxQZtFSx7kg30me7xEZWu
1h3c1yjzZJAZ1E1jiS87IEm8cLjpo9/UVmVFe542DbAE2Ev4RzBbkKIEi3CoA4Mb8y8kFrTmZiLx
tw5pXTcDv2RX/PoG/qvaMTiCUJ/h1dIxSKeJgDVxjs8aM8ONFxapv5A6yNSYqvjO/AD+8sWqF0Cd
EZqkD1X7LCct7rulpfsivez6+/oDBmP5Hdw/1+G7wPsIUvVaIn9VRzAD5+fXhr0zCwcJmNBBkYuU
nNFMJT9raTf64dUUPXO1eFLShU7qHGu1N/2gaPV49YyMhhQJAyQph0+E7uTH+6CpVVf7CLnASjt7
Q2zQTtcP8DMGaxSvMw7/mR//G9w/guqrEm//JMoaHnXvGcNIKn4SFxg+3AlWxfgB7uDwX/fberNO
62HTFHuG4gTCEySyr273uSDG70cssBQ9BqOzh+cx3ikDYLy4gDuTC4ALLpaEXtkegACKFL35e8uy
8PDV+aFgL28qMDLHBd2vNJPlsMXTvHctFdOI7ioRtT5qA1q+Qg2BjtbwlGoIbm8tbV19ZZJcskW6
Q4nXwHbYnJ21Uaye0vTdSiFRiZOpUgQQwAiDreqKU/enzMhhUp4ZZ6TABhb7cjT5+AN8+5EZTNWx
OCO9n8Jg4ky0SER7HMtFMxHnIYYc+3Da5ZEfKXSn4vyO69JZUebchKnhh9jaVMAIMjp+fn8oNVV9
DIDNbO0bBzcKrZyKdazw2zRmlZZYx2QiQ++CK9fV8E+le4+Un8WcblRp79WJ7BZ1v25ZmWtwU8OS
rhkwQ72In9rasnuNJOvr9uZepcYAw6JixhLGJlqeSzmjhudgyaf6zqqmRg+5o5adtr6sGCrLNroo
EeQvT8ufztr2bVOC28js7b4RdXJ/1mZfLEOfdC5PKs56BSZUGi5zu8m/IMsL0lUC/tD/6v8tpeZt
WGe8UgcDu2ANnVnvUocQuKmjDGrK9YM5VtF1yO2/hBjdvkn94JlAzT2K+m5fyodlI0zWZhe8gFZx
g48jxXn22IwEI1Ly3ypUSkdJpFO+EbuFH3Z3TKmlji5NnXvsA5uBrWalBTFt4LVNj/FmShTZ9ENj
A55WnmlWJ2hK1DNlucyhWUdyXBE+9QH2Txk2Zj1dHHs+36YqffvNvz0FIe/G2vELreyyN9QrqCQF
+m12ikZeMcVdbOzPHFUl5pRHNIWN+BUj01l1n6uHrFVqb3IGSFU1aYGi93ioDWeBn0VI4G36jMB+
p9VRshH53SCUfyHOjLAozY3bEbjf2kJVtqEubh4J+j+LKFvjnHMkbYX9W8PiDoGqQHv/dt61qAuv
XZcPF8KBHicbr6IyQFTVVgGq8Geg/U+CFkOW6UgZxVN7srts5SGInJ2TmFeWcouvwSAyfGKJMGIX
k9tAr5oBXAnNH1QVB9Z2n7GP66eGXJNVHz8ZZlcBSLaf/TH7+DI25+Rijbl1cJkUrzETn93xn/jI
HjeDxHZcWqNRMgpd2GoVn+g+vF43iy1P1DAMFOa3lgR2xyxgKdudpYLevxTOv3rwDFXa0+EG9ZcC
EIJkJFJtO4jE+whfyPLB2U09tDh642BfHuJtF55pnd33MLAICDi82Y0O6ORXliZ3LuKGOmryiF2w
rnZ+qsa1NC8jn92DSIia37LT5XcHq5YcFInyOqwY16KjkIMbN2VgQ+z6e4jWmZp48YVWs24BXhyQ
ARdJlRu8CpkLCZ9S8snkvwLl3u3l8nPIuWAKK5AaWNBJ27qjuDmCiQ0DkXtdgbHvQzTj128oxYz3
z1nvCgjjJfsZF0hRqY/5aqlzg+RzQn+SeH7A/CiRWa839PSsa7wBtjJdhUeZuc7VhG+V4zd1P7PU
x6Xs5VIjovg6NYJeFBSB+p+WbUCfdRwXojA6Au5j6JX5w3YhPZqS87wvj4OkcTF9K2ANQfoaiREw
lVORCKRRRY+yDlInNtE0dcQEl4aH5VQ58iZCCAMQyA42A6ffnkakqf8WwKo24sRbD4gSB0nDo/ZV
FUbKlKQtb3m9UHEtpcFUzDzQ2XMjI4qh/ezdxNEaEbNTvehkW90LKFGgNFxJeQpL5w1CjhQfsMzf
Qr6YKRzPXGCekByii2J/NAb4C8IdpqS6w2Mkqmq+05YfnC6BUHvXRXI+KZLbY7nFBgjrxPn5UKKj
U07XQ02KzP52EzuCR5lRKv6aSbXsR3GorH7bbmZCkyCkKH7nIqwm6Yo922maG4PMFNa9urxZVn8Q
3Y3L3GtoQZFYaihUIliY4ZbuwzJNcyRFby5P4zJXAbY7wqcjxy5dr9TiUAt5lc6Pxgzi2sPVkFH7
HwL9GpLsX1gTSvn0iBnHgEomWOaUzx+Wmx90nlxHyAZ/gxdwyZ1iO1fStj0n2Y7Xsrm/lFVz8O6q
B8bI8SHmM9aTzxLSbMQ8DxwKfxxWwkLVuLuLq56/+Y/QcKu44oeHIp8AS32uQ+y+9vRCnFN2sowZ
/fA+0jSAwpAAIAyw29ZkUdEf09pdArisHcoPqxNykVSED+eOyGHYkH0LuoioJy9ARV8dEDTogJ6l
gLa+hWavDV2aYbwJF1gowiZrO1rdym3zxnQ7fKTLFU0gqUpam8z0ivNItNOwoSdEYObUrjC7id8f
+iHODHb3MhHlfGDTm0MNjgUVYPLq9H1Fa0RDOWsvFSDACMRechWCTcd+WdPOojb/8ONod7hSqR3C
4jNp3D56dddy9B45dXrRhc9fXYoc5CxOtHHVwCcmP+yLD33QZX6ed/sBAGlQQtZ2l+OB8l3b5GoO
342DZelzcqpX/tc378TdutUCLnnCQfUIkzSkuLRU3vOJO50M0C9vcxEva8F2jMTQi+HDBQ8A1Lb7
mAbobeXe04gEDCG2ZHqp3aRvemUclnpfhEVDlcH69lVhwm1mqU9Hu0TbDCuW19wMEMTAaSMBRzod
1U05OZ/0vzW17PuihT9DZkaeUWW0+xU5E+DllbaTnZm2bhttAXl0dpLEXvTBLQIHiAjgEIY/GHCZ
9eOsgSgHrXuCVsaksXSaZ6Rxr+pTivu7H6kY0J24YFHhyCjmDcw9nAvnId7oFjDZstUOQZ6BAKMe
bF//zmVnE3rhNHykhODIXlQhB/budfo1WkGX76NbCklHM84Alh89e/fWloagqkwh/Xc3Cpk+o60a
jPv3miab3EeHe3Nmr2x3D74h3QLHlrvxgLCFqSwlHK0u0Zt7vAZPmxmHDX2kAbauLj/RhvCVVcta
aDXQR4HNx9ZmZF5bxWSxp3wu/i928YZKYv1qFWcC4sZEVc0qie1TdRDF6hqITAsIcL/qg6+LTjdb
nWIlLB6iDZkfsHOohvgvfHN39fffpcU2YObmahdJUqzTgeD6X17+ZYK8yqbT/2vae6WMF17AJLWw
hythDYoCTAUnDuV678X0H/Gshnu1gbFnoErcdH4eJzOF9l5vfk/P2rQAJ4nER4hghHsOfmcvtdHB
NF4b3PiuaMx2yuK0iQg3NzhKdIjjH6chIH2MT2SP2UmdCYdVeucO0bfWwlaE1ihLbCL4oa4Obrg3
VOc8gXqALs5KBCisEyXZpZim380Tr/UrJz8thuPwbwB5RWsU8uNTLRjlvoJq3/yPfgBUQfHQGTmk
t0tE4UUnuFj2PK0LS+GxdvhdMJBwCCYumOycYWFvaJE5XXkyVa3P+5Lq2ptJ6ahQaybmFW5acPnc
HXajQ778NtfwSJT4RShyNFCJWqyd2vbVrwUhhRCt0piVoBItCz3tdCzGgq9LSR2/v2MRiz8nxBkt
8Cg5fxMB+zTdw2+H830Vi4mKIRHei8gZe/L0eIZf4wC/NM/HS4zYQk4t0TuORA0/Ge6nC6Vox2w3
P887r7VFBrH25ZM9SR3CRzDPKW3rtTj98yYne5RNA374xcRkdg1SSnZoL5WSIkd5UajHqqWuaae1
47W/gp+N9aeKLYpGydZtsvjRDCPRZwbQs+rqjNQiGib75FjEGP7vAStJ2eq/AZJuA3ysacy4X3c2
RXg6MfP3XfUvLkWo7J5MDHXTeX0/Lp1Aqi7bvSrVMcI5CFWDB2Fvp28JkE603THzREm28seVGx4i
fLaJ7ibW4W3TS9lESNfu/O9uAJ7jtZW+M/BXjrv8+OE3Q4gRQyZcYnm1X/idD851MGBm5stMD1Eq
PJ4oeVw4QTmawbgDtYZmW8ehskUI1TfXPYc7GwC75zEFFTNsNoXphY9uhucvmQiNXhEDDxhXYFo+
Vx+SohBW1QHRWoPmEp4Rnj3MYt99BPRf3WWUUTvUnQ+RBJeKqzBlMEvzNXLPnKI1n72Dhn8T4DDh
2snM22M9IANPDSoSvLdzCdmDhoCahwQtwfrk3abEEGNztS0lvMtmZm8hK4otWSSzp3/kS2Zq0Gsv
YVMUGI8lJmZBSLDLCDS924YrIvVv3E1f8jrZXhfCrGI8dLSV5FcVbC04zLxxI5D6szSA9Yj6TPfW
mbrcc7sAnj8kHxpM59zKx8b+S7bCeaZmyWBLhFB8YgMdb/ex28PXCf8A8PJaMzVedqqX0TCwpRtk
tz9PR5XgKfpPynu6hy54fyMXK66TjPgrRILTQIntCWdUPnypOmU8ka+DNAZBvS+ZgpN58HhbP9E0
6Fa+/9SYcURjQSH4BBfxyQUjcXj+njndJop0dKSbRE/DNrqam1RSDuBCFMb1q3eoWD5s+VhR5VH+
XLw7asB6BzIbBJm6/zDcBRCs0ZcXxyWjTIIfrYMB4SZclCV2yeTWROAeL/R3dUJQbeY2qm8jogwQ
ktrBA1Tz01m5Ivlup8jKoE8YVbBeK/nHETJKYC+2/s9U08QNSkY9N8TQuyoMCl9JRZDNMm7RBbD4
a8xlKlpsZFXYFnLztackKoYJXGxxluWr+OC67fbZCqeTH2kyB4pE3nLu30mDSJibvDYd72UZFD1+
TsqIiJGNpbXDbSP3B5w+dJqDPQ0GpH/ry7SOW7k8um1Rl6aL5gcOZ7PXJyorqC8fV0LK2g5l8nkj
N6COJfKEXJxoEZf2ygjIO7KGAz6warbdIhMiyVoSP+E4gExwJg2IHEmbwslATvWlKrZZZIi0CA+4
5NMiAsshjrfk4Jf1hhyj/VNsSPv3XWe0/S1zIv/TYHFJ2vwfwalDSE1AwTJO4pv8x0eDzqHhTo+I
iZ1aiZH1FggBz7KIZ+8Mk+kLMvYVJTRWaTAxoTRrxx1dd8yopDSW0kZbFbQNOI+fQBY7gowoOUB6
vXEVcn2b39zhCtXI69PwEHmdwIIwS5JlspLfsJrRAqd+4dy39NJEB9QAq+trOBEsV6ovZ3xjyRJE
+KcDdvDj3uePR9lGjEnGeyDOL9GcrUwBpIJJptNvTgf8AXE+wVWlCs2UZyLIAP4TWOduMlr5Ut40
Pjf7z6nMo8X0y/DUvT+5do69eRVfSiBFZ/Fy2cjgZ0FAaFYM/PWPt4POrQ5HwwrIO/aRllVJnwiy
ZOSLU0Z0GLdlrDv2gdgMUMLfH5z0wVf5604yVucbsOZehXhZqPBWzfE+BdHOqdRxZZFrWcT2/r5F
4ZbB8L6NBFoaAMfFQDY6VdcQPvIYP90wnaxu9ohqSkSh912drQwmmR9RJaliokhoHp4AfZ6HVO2a
MzNG0PSx0vfL5uT4C5YISxGJthNYtZpNIFgcmQGfsmPJK0UE0pwPoZm95kQDLqrWXogmFalLB0mO
mrr7/mY9aV6cVAZMilXwuTN/QA5J6/j0K6ZSREVwla5vNNqdExIsPNXmaOJCr7TzadCGW7x9Knaa
BiPqkf+wmLdKyVplHoHa+agu9kIPxL+hDc+Xklcz0KDd2yqcDPzSoAFJJSIfsxKMlYPY4BOMc++J
6lO3FBNnTgV/LdgDv27Gs5wc2NoyGdBrhpgdZL0G9dlwhQB9V6M4Y9aXNgptXnHg/uI34AK1md+B
26pPs9DwV6SE6GPLa6QfynJ/9uf6bxxTWSHKodhm6RIedds0AvJPANXLSDwmyRqiypueBQzIEZws
3aFaPn9VAQ/c0fPAgY5hJXcvDz36TJKn1kzEluApiS1PPfTE2F0DPrmPpJrr+UBw469duCKXAbs0
k04TOoo9O2VJ0gybaUx0NtsyA9rIHLxiRGG23e9crdlHualAR2XuyXY1oVLEECt6KaH4riryylNl
A2Ero5JD1HijChIX4HutWdvyyk4Vrq5s7r0nh1q+aoQsy5I9dShEoRMWXaAuPIHf3PBbfAWry89W
H5GsCp5MSVIGdbVJ3F4OcxX9xCYhZmveE2rA45ZqcDteJAEjPVOSBgnH9Ootd8p3XnnATT4N726N
vP1DfBuSq9ZyQs57W9ddpqeIsEcareT7Ri2gPUHUCHFeaAcGFE4tFYIKMegIutktv9OrDazNDB4J
XYkUsKRyjHV2WhrYvrid6N2dnMUx2so3VC+zUnIcDvVA2IwpB5xQ1WjAim5THYVMrgD6UnahePDi
lbrH0rOogStRGWBvXeImxIlnDO0ayfZi8HF4z0DoRJ7Drmxb5shNwYArfJkQIjeju2SLY8/xn5Ct
kE7/YW5Oo5ys5rPqoKK0uMvQbKue4GxXsHAVZm3RLldTmgoTcLjIl3TE4MimR+RUdElHt7HwTtvK
QvERzQGZhmhFSr9jYIu8Dyspfnn5/+YxfXQhU+tMRPUeC8E3IqEo3kOqJ2ueZp0BJ97XzZWa2Trc
CYAJsRSPrn53y7UkLtdFLqDdwldoOVMjhdkMpgAyBGAoP3nWC/jFAEHQ46MbsF8VgBZqnyAlxLLT
QMwpbqzK7hA7Btuj6PXvzsOHIR3bwM7LCaqQ5NZ1zQnn7ZKoBqO4XZiAJS9+izbb4OckVBxQAfMU
AgjVxKKbvtHIGwQwnz7T9147a5AdhuVPBHOFklZaDTYnSCe0SLqz0vrgUFZOwAnUYR8P4xbH/qc3
JpibDirTEyQBIepAD9qTTiWU/3Bk2WsSu7cCik7XtAEx23Ed8yH4oVapoXjhgsHhFGH+a7f1A2Vr
nGYb5XIDdGnpFlWUi/NZ5K2p6Ln9GTfS8iUhiZH/6ZRfa1MsNrpWvXFYAoTA03Cc1yLJ8cWlfq4H
42hSbqJX3t/TpSng5Bu28NcNe3zlLh3xF0c0PuSEIJ8GCs3+u5bR6RROPrj7hk5YQ+cqDHXOF355
nAbYzHb7AdKsaNXk54bCngRRZowEFg6o3iqkwz5nk7qNEHP9b1pIXjJAc+TZFJz3l7emVp9ShWpr
Fb+DerGAfH8QbZIaMYN/kZy7XluG1b/79Gsxqkm4EBiRpaG4Lumf/plPVvVzDkOvCx2phjRbAX4n
3Ze0hFMi2WhaUJwxoP6Aya7vNwnK34/WYlHb0uwWIFKDWypKbin9+L11Jx6byfebmXF3t5QlOf+O
d1QbhHbe2ri3cX/TU1rfnBxJudwU7HsSjKBPBHTZZofH1uLAzd23hcZiXi9eV67Sji2t6NSvTp/s
12+Fu4w9Y9qWZY+ts1jnYmdRhOYt+FanxX2n+yKc7kZ6vUeZqXeatMGNFi06lfaqQuceiR8Xc6OB
RJS2ZVdpqk45AAwrp1hw/bl4A5qtnHEqC8ZDMZEVxNkcst8kSoELgs8QfCQ6F2mMwRoGEUHHTquM
DthMERk1TUhANMSOfOXYBgprAGxPXGHb/Jo5SiAxn+vEuFTE5NB/kvX47UDkzAOpe7Qsp+JBnXm2
087a/lAMbZ56YIkiSrftEJEhIT6IO1e30fqrTX9EcgcHcg9jv/ZlbbrNsy+pDQBvPxT8o2+hcZ7Y
Pgpib4iSyzvR73MLCM2nHqk7A40Omcki6PmxGk6uLvTUZnAyvrBPIrlF7nH3vIveWcJbcrQRV0l8
MJYUoncKh9NaUtbqWEPF+988rErYZm5/yD3JfT+xaFgzs9XxOeATYTwEaGkF6Z+PTph4qocKcDWb
BDV5a3I95vsNEpVASiRO7s4JjJwcSGTLXHliaDz1o0r4lWALrvl6vnyRhjU5PWmYyoRh3lpiRgS1
mT35TJBRX7qVGp7u44gM1dkjuWsD2npN6LUJA4md/sviUs1Ai7RWB+XI7m2b/JLZiLEpy5FYLp2v
k9YjZLYrVTQ5sdT48x4OhEhj7WOQjG9dlQUt0ohedkVPoxC4XiyqSLV19yu8cT4gT4HkdVIb01vS
YFhN3p4bRnMVYMdMNjKMQHhBekg5Yc5Vl6YC1XOtcagjKm3+4Yiob3GGew7NIkBFj6jPcaTa/0OV
y080/DuMC6B0qQik+gxVbftXV+xCMGz8fM9i/nxFDekZbR7zJKplIoXuJJHTxx5LRhwxtdpGiln0
86xM7w4gmODPvcuaKdiJF1LGWRnerSeUgA2SX50gBSx/rc2HAkVCw0aKavyntD62SOI7yK/wGuZ6
PihCE1RlsfxRVKn1m88nb6Y4+rhzU8OMVkVhsZNihtIudY6QO5Se5eTskz1hI+IlKfWW1iGy3f1c
FnBYmSIowzg9ZUTMorryKQVmlQ5Xy1m4G9WQkBI685D418oXbpgvog1fFVOiwV80NJHMG59hPfgn
hBm6+pEflVJSc4S5yWT5ogsefhQEOsjgb2MViJSCDPbrkXE40qsnEgx6TWIwe6nizQH/Uy2NG6kh
AswRnusiPheQIqfXCj9infnYZi4ylovWMjlneN6xhLG4EHkOp46h09HusPsTx+ulhIDxnsbtcUcc
FR/0NoqI6fcuPr2rwIKN1XCx7u5IItR/jcKo0D5UiCjzdDUYL2R4J3kJ4hGVY1NQUV+6Eo9WbseM
0iesmBCkc9PWV0UoKmnhNjEBWl7nhzfK+4yb/fp1ek6062GTUT1hVMZeS8ooY/N3WpoQXP5EKmwK
nt8A8Yn0kyeyr5Co3khGgmW1TtMmQJHgZs9JNi3QaYzzFrXo03uC73WzZF1Mxhs0eckk+KxkgMes
zmpldCtE/jddPM11XeY6r2873T9Mrhw/keP87K2mRViqWnbwJ/RMHZ1QVyHm8tw1HUmKrtguhR2i
GBE97c80r21L8L2cg61mNulJ+UnzkJtWiwa9D21fp8bo8hAHHDu7uVr7Q1ZKTtJbHlbDWLkUO0bU
FeRR6/LT4wKTNkaCAlfUQdGkvi6TDOPx8pwMPo8T16ZQPc75UILaQNzQ1g2jPndS8ohd+VM5Yckc
/ko8+KX/SgI443PwSKvJVycXE7OTtayLE5aWy+Hi6LocNdVud6JcOl7u75YMkSEAT0vMA5zP29sf
oadSXsE1XTSS686co9e/VAOsKh1wcylYy5J2QZoD9HeYrHsSRWbfz/Bm3CaNhaKoB86vQxdPr8+I
HJ9ltF7ldtyJjtuLpttuU4eVjaMa8VyJzw9oPsjw0TKIO7E1C6INXNsOSIlXyrq2aXsf6HeL3BcY
f39fn3vOKPk78igLyJxtEMAfIqr1ZbLiAXESx2m0abNhEWDEQZUaagRlspSKVwgU44gDIGnLQDIA
lN069+DvedRX+wdzCUktsR1S3is1eujushCszDC2J8eIU1OhvsSGnwvqyQqd5WNVzWjeIopjbbBS
oTkAnP7uJAH7RURchCQm5tjkaMwxlXl3BdrvrOGi/U53HGviOws6O8SSIvcKF1XS5uFL0J2FWEA1
ANWySjKwhAwzfc1Q47ATmCqPt8xZ0H7POn1Dn9dZivZHOguPvchBAyyqZkoBEb/Uugj03YFfjft0
1CQkj/lCvjVBLmjrmm+3tLpr5bAo2FSc3HJyvr9V/Cui6DCowHUI1u2+tnF1Opg4lDfaXnfhXCmN
o/t2xbls6nWiAX68S7SWHoOdQFhFf/gvoEGzvd/kmwZlEl9y0uDQBoDItxHyodXgheAxtREDw8MX
QeaPNWo3UGYPEGM7W0YFwtxFHrMuWFAZTKAzIEJ2/uXi0Z30L8Oz2T9fDT5Mrj5fJJX6KbrB+J4t
ZwpsAnSnrWq1Z7xIGGV6WkLzONOWbZWb3ZjqyF4qR4pIr0XRv6fyX4wJucb9/mnouBY+SPj9B9Ss
gW27SIjbiVoEN1xD7uCTUJ8B1jI8NWila/B/7/en7eE9IY5leHLiW3IKArzDwsX73P5GXlPNYqYd
v0Jb2nkfAomsthlt2wE06UYyW+sTUtD6O10htLTlvdAmJCXFDmT3p8R4AbQ+6hO22co1JsdKFqnO
165V28Iqj/5aY3hC1S6LssoMo3fC4ilCizO1WL59VbRcW6RQ5VJqiBg+maI4IldSgy7/2P8WSgYM
WZNM9XQrUWAYuBbHVYhCQ60U0rAHaoh2w3hsJDdKTGSZe1Qz8OV61DanaAiwQm4ymSkxm5a0Qzlz
KnA9bdCd6XcWGvvK0xtZDXXp/x6wHanhDoZpdTrfxCphTgS5mr1qtMGPsYcyrc2llZnjmG6FdELx
3AGyBoEsWhVGNxhnMsmuwWvH9tEWQidOUJQUdYoHYDqoszqKnMiDtrvc2b/Go7V0v/m+HTdbZs0C
yll9yVeyBPKUXIq0nqzCaeD0AH8FZvzvZcEj5Ad4GP4y9jPdm+maSIwu7QQEsLWwyRABftpcFLbJ
VcxmOcyXiEu15QQtqEZUbCFCvKbTCEh2MLfiP/ibm8pXeYHtqiBHCx/cbWXQ5wXUnyYwDHfVg1Yj
mhQo4DBY7qpWQcH0OtMYi/t1olJ8r2t3Zrp5iiF9hQlpEZ2bUxrF+HAufqK9PJpD4XP+59Y6HX56
v2DY+pyA1w/mnlyJp2lx4/UoJj+ORqCny9eERGRKEWhp2KJcjLey03ST/sXyPSawwimYHTf2NvPR
ESuRYOjPwvfNrjCujGXe40ie7ma7KeWaGnzzpYmzkregvk/0JO9MAdqNxCkxGQ6iQGz4aZaLqSDu
X44PPWrMc03ClrDpNhbeU/l9iHaLIU1LOSpNYAisRp3lWhF9AwpJKZgnnR6Zh3fmcoNGjXlyof3k
GSMjLIwm77DXJYwpUHUfAOFw+WLp7iyI1B19NrgW97mdG/8jGKzJbQZuDSaQyhBtfnaR3bPHxHd3
cGeGWKAQMoKCLzH8YMKVNfPtBSLCJhR9igJy/tUpE/La/X4M4+sVFJjbFnml34ONdu0/mS10Z+9Y
fL0TJF9QRXiWHs026n/GCh4KDhBxFK2oIzbE3v35BtEmJ6Jjs/NXSy81h1/7djzxU59xEn7HVS7r
9kjob+2Vp8W7V5/l13sLsLtLz6k8tcTR3p7qbmN4b4DOd9H3WUaJYNTUxGCk1Rlfw+nPzvMAAS5a
AmuMmnBRigzOdk+r4u0uKzo2n8JRAng3XOROvw2sqwEou8DMRa7lzFRriia8H49A2lkUhr5Rsfs3
Q+YauurIiU6hsyHDbJLJ6LcpNnFXBUADOTU0oy4LX49hYfMGdKXyCy6iVqz06ZdBF57I0ZRanwAp
sb+GLwdhXQomIn7IczFx5i6ouwqEezdJV7JQbPxcEjZfO4XH/tV2k05Y6KkQ95H8pNmGb8l4BXJ+
BoluAZNDE6AncFxQ3obiFMFTHnn7mluNdLzng8QKwjI/hfzENTYt45YTfBzTIxUifLwABK3cjCAP
qxm5Xmq822HVKkScGHpUfZDHA0Rm9937f2G1KayO8fn/LOFYFQHpxc6QyNcjcqgyGBWy5Fn7UbHY
eyk/oOA0IOHQC7RXmO3qBLvBm5CKbRozvAz9/BGYCV2BLdfz77d+0qLChc0FmK3mWhpbpZJEE8kv
Levt5a67joau0hbue5xoXu5LYtRKf8zcdhKTzg+CfidP6FnJC673opIsAvRXa2jN4SBlm8qnoo14
PeUfU/Hwv/g96VBDKldU2Wak2i641LMSbMlsIzyjSUTVMXtgoRKkwdzvV0v/wJcywTyLmN+RQ87f
RRG9Mev04bL9g+7pOYX2eCPvjzfrLdZ9oOCWGlD2e1SOuBKOxShNN6EAeSiL682BQADMEi3jV10C
nIw80YNbkTNCrJyzQ+mNU0YeqFekV/PBFsxcBfAHKLgE7ehUGP/m3AUdIwEHMnWFLKajCzMTCzKM
dsBmVGx3uu9hWZ8bUf+WMMuumyNqbrUDuXLtDbiskl7tnVQk1Z022or+BsXpmP3O27TPjxREyzCn
UWbMGLqJry3rYJuYY8ml8teTh10+S9IR8KCweRJdCQh+RrQGiRnNoNJ6bZADq7vWcdYeCnP93zYk
T+wrxZhNsQvcbW0Cw5nDcutdNDvkt/qdaAQU37889TkqHEq/CoVOBwgOgu/vKAwOeYbUHPtEuj9p
jWUNG9+9hw6waoJ5UJWHKCTik8hJUPDm2WwsDdE98qCxlgvQ+/OIpvqXzb1/etEQU1x7bMqpo6fC
zc6RezbzY3FJKjHMN1n9XYqPRPeI/veq4KgaSqQEnWHTHmU8VH7OeYzbAKh32XLQEOIwVnE3BW3b
ZnyPpTqw0XqS8cuaz7lycS8rCaW2JEASXToz6jFYQDVPw3vXW83+jIIzl808soLDpYUAQ5711QSM
Fv1XQa/1Am36HLff3ilcsTVa65i5jSK3PzV9NJgzCsIu5XBHMv2qNEh3vs+tBy5dryok3J3SaX3G
kJ+n6Z23GjIWYy23YVOlXUBwYweHRKMd/HjoS4iur+ethEMmsrKc5kXkmJIjriHSJDtEAIRYtKDU
M+OyFOfsk/fLq5pMMwIxu8dFXOcfqG6WK5869Jqm3ozMn/hdkmp1tYdf2vL88yU6nOYDzOYsU9hE
AGgapDaJmVxdLXNTvTFE12pZ800hdskNm469JtkavFR8z5tu5zs0oMD7N4V6EB6fiUgE6QDKI1ph
Q6z89LKu41+0y1gMYfwnKS+2q3cqEqj4EKnBeydWwitt2IS26A0D67viarUXO897D8jmLpV106TF
W7lgRVsSFynVG7Zd4IDWllootecszSwQyr3Qk/mqgaaQWwW5hYdUt3ZzDjggkj7756DTc0ybMLd9
1FeBHjKxPTtozxPAP+ZMVHVwQ7Kgraxzi5qrS3AXO95I1vwZ5osWF0IuOylPHa9N+qjXYJ0/MpWu
yrSAQ1k/9Gnu2VwQKVMN8cwJH3jYSfz5qbvQDcSbGazygPyG44ojbgNKaXYyATBlOnPmWSJmeHXd
B9KcWg3sstgtlFlipyB5XvJrpjDebH9e43oNN0hITAvZLuc/I1COTxGHKLRKt6gvpAfiBQuvLqEf
Nn6onrFgG5PejeQ+dChQJaCl8bKzfZ2PL7DZtjPztirTzlkBcyJ1CZL4Fa/VhbpucY0tLZ9Y1kTS
CdW/ORRXoZWhDBjbJs0uhNZXEKXzUhEjDbOEFcCNzrN5wwHbYB6KH9CkzoYyvV+fOx2Dq8EFq/9b
4Bgs/GkFq55oy3yv09pZovQiDHDECcJgeBaa0xfcq7y/9SicKSbUI8mBlZi88tf8BUkcgXLz5Nty
e5Fr4aOkBrt3JKW2LVIuNAG4AiyR4q/hsB92RjOgjxRK6g4GKscCozdrpeovsJOLugmuHbGTOo0l
pRsSEwM6f4OmGqF1aWywnQZY8hTq9mFomvzv1+TRKeKc8wV/INJ4MuaYqdVVIPtmH34yUFelF6Re
zR0kzDLi4s8nbukkLtUW6e5+sgidwfTzAFdkEKPtPOrR9efvmdw56HMbwx9stRLii/SqdUK4TsKt
d9CcVXyWvzkC9mfTNuYmRhlVoGCfre2cq7X8TS91Gd63KiD1wRpfh+PxI7PKllAhmTMsiOFZQ8ep
DfIhWQy809zDCZ+5YBcKjX8vcvTG8zYxGfUBq/VvY18fUsPE49A8xoAtTgcti0qVSQlNmeqnaJ+5
seSH8hnPO73Qw/FGBMKP36KcSN4fFpELXoPJ4rofEukECnClsuvLuhGqmvtOL8+M7GOBtKiSNdH9
VCsA1zC4Bz+QgK454Ll+pJZIRTZrBF55lwV3CmIAbH8Jtxh1ZeUCJAlapHhSNn80eFpfGfprVMGy
OsjQaJIxni+qO3a+RsZhEeVsq3wOAngdc+eB08dqJJ1uus6cncE3WDX6z5eWatEZQzXk2comp0P7
P29ulrU2DTHHLWC8pv8kf5PZumBthkOtk25rsDDKz0cBiQ6WVpH/29/Ovme3wtrdk50m1oDBV403
RGG/Cyaj7twZnoYfnjdPEnaKvs2UQYDdNMZoI42Ygr4Pa0+iMo3CT1mUvk2fGC/rcW1aTMgnDjmA
fCNhMtt7IVHqdyMjOYK9Pcgw33HE5Ht1jWLGdeKmfv3hsqSvVakB7yjGZo8rTLKcjjgJvVBwmunZ
xWUpmqAargl6GxGgV5ClRZT9dBtWmG4fhn2lKPTAOhJndy7XFcfV2Gb4SMTusUiLZZfudr13BV1Y
TYrgaB3vUJ/J0lLJBDgbYviuOjDUwlRgv/b4qjkM/l8iAdSCi7gwyiPxmCqGDQpU6f71fd+iAhRt
0sdqEyycLnyKMVWIS8dCZnYpT8htgEcBDsOLhAFsE4P2yI7m0iw+a05mCZQfhZuAGzIoElFA+N8r
6cOnLX32mYNBZZ1E6lt31XwCgM55LzL2mEVwi0i3NLGFKLmAvVv+MfJFRcgRP8NAbSr8/ptZmbIp
5uFkFfbXPPTQp4591Mwem1QZFLSqSxSpx4+/1pfzxCxVUOGTkZxQu0SdHg6hwpDokJPpuLJMVP62
0eAXMmW0mPGVS7UMmGU+tXLKcnjuOYhlxHXnZnzm/wYzhkQLwnzGYumySHL6j5kV9Kho3WiLkzSv
yzFSCr1yr3QFKDrFujzwoNxW17P7QH7skIpal7Ov9dt7fvU8HnB1jbE/tFzNrRn+mD/Tdn6ewMU7
YusURZZDJbFV9dDVmwBdYwJWGtqdLsadtR0QTWX5Ef9Aurf3V84ew6mid+W5t9D+VK1REMcuhFKF
jOUoBZnuuUQ2b93krL8W6Ci4Y9ep9gqeGNdQafyZirJOe+Ot+yCHFMUAqN1fYEdXmnMXGBPeneB2
GQ12qlPzf2B1Iz4bbRfBhTz2AdHxrrEbNJmKjaGXjSoFBBxZEqPe8aqyjrH18gC35AOlWMbtFWjO
+ggd1ZNMr/B8TnxKJmUL3n9pd2AagfAs3itzTlbbZPB+vL98MFVSI9RnlyNto0/G94GLjhLMg2Ke
EsiOGtzuQzm+p40pZB/3vHxoL63pQymcftsXk5lUrG7lOGpTLr8KnU1p+TAWYDAXCo8c3T3/94xT
lMcJZ4hqTRnu283qpWx+EtR2AUOmUL9unA++vyTdImCYvvlxJhNnpHciHGr0IopfoeM35aogHF+9
5loJPmisNy+Dicab9M+U9s/cMumW0ezS+6O0IDIvzlOfNqXwL7ZXq/wudeD8FaalutrDdLBr1pPL
7tgooWdOz/76splTErxuoXdjX8vfhzCIIxXsmGLjObiF/ihUDd1kAnuGZpbL0X0RCMv+QxYx9ne1
Q+gWZm3DjZvNE3e7j86k9LkGCiMGbIXEqOLcKES3nd7Y37xztjS891TLLj7VHkZg9oHqmf5pyPv7
yOTNCWWd7P+/zLOplfdHkMNtFGjyPaMfQw/09Ckb9DZATXnUFlqByb5MpN6AoADvfDVBdFDyO/l2
a9t01prs8UzoODbUwsivRvXIALQ5DbYz/Xd4C4XPsA8Q2aXCM8Px2GgfH9z3Zaxo1cmU12JqW8pr
GeijhaPsmATwDssjn0+CKk7/l3EomX7PM94tiSIO28z9yquqJzLaXeYejUJcib+HrQYPDeAfrjGR
Bs2tusx33ZliOuYQZ22IbiNx00ExncUIno/vsgcSJ//QJKngBG5rptzi7GRiIDIhDl7Cd75Ohx0j
r4j9MRARSFubzqq/mbkpg0l7WPQnjI0lZ9BcNdYDbp0GbfY3SSJjyUuPINpWDO/9e7j/YB4belom
NSF11jl+af2rS8cgv1MwyK2rGjseNTJwuHYs6gjuizcTttdNPm0sUqkqfVusSDgaxVfs0GjoKDVo
HqxntL+8b6xEqflLbeyDVBrKVocwWtWygIjoD9I4Ch7/3VmVffmIayuZKqnwcjt9NHJ67HYIlilo
LHiCzBvfT5laaxdvNXIvnkoR7yDzuWF3cLa1RBrv03kVKA2m1tGVoj6rTybza3joOoqOPGNRe5Jw
hAf4YgZleHznqtlGPhhDA+Zn5dUOVaP2y7fu0NUGfc3WmaBTijA7eHBR6L1GAgHV89VDvkdo+02G
lh2Dz+tYzzcJf1N3IeENyFGnm5UZKLcSpEaoCdYSkGeNtTZYNXQp/VBClFkE+0lH7Bn9VewhzDjZ
IMBGuDxuTBPGvW15rlI3/SJVey8VWlaeKFc3qjVzOztZSJnYwUCHrZGqj4ihHF53KNI5IY/c2gGY
K9YYyyYjf8yEke5sZpGGJNG8GIZhosJ+I3nFFBorlaAjqFF7msVcMUs1JM3ono01PClQqsycbypm
UcISMe9YQEacYxszLbcwZO97ZNjLJW7lyuxrdKLfQ8ICMq2oXjcbw+rb3x2Ql6dxW3tNLbvDLgAr
DMhdrHbbZ49gLER/uTBgq7DIYWBF8GHqOT64eHMD0Qv6ovNU81uKpgGQRRAqukf/nui7iwp3JfSn
ogNBKhwBiWAuKgEa7efT41EZwM44MA/GUKxUmQgKcu9M78C3AzKiIuNiBHdx5b+Jhb82XBl0hO8q
XpOd89MUnhm7dL5afY8PwTpkHSxkMDpd6B1Pk0BCMsLyCW5zEbav7aFfA9dI51R8wWXJ+cgq4LuY
k7BSaKWmyX0YVlW5t7OFFCDSSgWcuF33BEEx7xL0ECydmQ/mC5I8wGWWyGx98eqgez5md5MC3tow
lJ9dhuXDm9wpXBxUgtl4YCJfaC7T4Jp2Jc4yO0J5pO0efjZsUIej/fkPa78qjjktbQi6ZckF5xuM
nxky6jTfxymvk/oNcbWOhSZDGljNbILGW9A8qTIbbcg11vWZkN58DNYh6rNdd6DlmHEtnYb5+TCY
OS8260fd2vp9P21uyhy/mJJTydxo0Z/9XPhj3yijBlxgZjenzqdLaI6oSGFMltTRq0fuPGcLPCho
O+tay8eaeji4XQ6ZM6/W9OImM7vt2ichHFMuJ/6WBAB0K0W63rWaAnF2Z+HT/Q21VUofRsYTZMyW
FYr8XRI9RKrlzRb84nsnJKVhRuC+6PiR7xnKp1v0NBWRXYvKqkqZ4gCJx9kackZ7L42ohUF2ikXk
5SW+Mz1LsYl/b+PlK559ZgyGSiFzM2NT40NcAQhaGRc2mFLctSmTS5gVPG7OFdMd8i0a6l8qyi8a
DhG2pxVN5LPZEDT84IOCjrXGvomY4yLfKIrFduWdrSFHzq5jwXrjlf/otFsh0I0NrLKyj1EQDsHl
RcoHU5/BfBATR9FE5rFS9zUcd+gxpJ0LAl+IpRwVweaSq72ZWq0UP3BBCNF5u+bLTlAEK+/Ys4pg
aLvyM85u6WUiVE1n688nn7nzu1CcSWxvHdYwrJouXkpSclOB9JKg/ShMSfpeKfvKZDYrJFimhSNc
VLm/f0BVGnNjDPcKMllomiKG0MlzzGwtLDv/NUP6YxOgM6TVFD03xU/n0CnMDz5RD7GszpSBre6Q
N5g5YkDYADkUd6y8Uq2PZuq44M70zg1D8rgywuKqGs6YnNJnxvNJoySz68gbnuvgDNfxerHotLdN
S0ZIrfm4If34FOgMT9udwvF4v67hCAxGAhNDEJ71WHQxRCUDMDmGC1Y7qaSE6T9cFZKFDRoCDJu+
UvJYYfuMKU8yOd3DgBh0t2CMOYv7e2fg9IYsLcZTEsnR8sHfcmvuqJHubj34QYSqH8wVc47zULqg
HsS/IfulFgPO2G79r1YIAEiJqBpSx/cC/g3UTUNRmdgbRNtuXkskzQKSKVKFL/aA2POeo/XJxfli
CDe2Y2yZT+HdDlzna3HB3DWo7daNgEg+MrM1vUzQtt4kWlvLql2E1CZ9BFL+mj6+4PP3s9WS83L3
StknbVxA/EmZu2HRRJ3OIwaPbZVNxyTlpVxBGJRPlwtf/KJpAxuTVIq5y/uKMzR+ZiI+bVNrraVD
k4Xj7XjI+CfsCKMc2o1OVffr8b5p8bKSUA/sE8N3JXXAekmw6p7Oma1gcooEPfE1Kvm5vQZvEUBq
6QFel/2zzQGkIrRmW7AxrBIZh0I38OAeoY4dCGxJRhZDTxBv3s1AoKph+djd43uHZtWKTvSD1WSE
5InIsPkpVQpcpafJ9ihm4mm2EXBD5xdPo0x91qtFx4zKBu9YaVQOm/fs3uWp9ZzFcUsAyg0rOH/U
/upQnN/EKKZKCwWXZNpU9Q2hjLScIg0swTg5uxN91Vm2sL4GqChF6/AunF0CUE+u/ptMQ3k00QgJ
TWM6FoAhsuZDNpxzLn8RBKhYKgyC187VuxAcgajcWUa0IurWv8lAeerqAA48aGKqBlaxzPQZUr4m
DBMZRHejzoLMp2pe8c550RXgV2+GHJTCuUwaimjOmHEMvGzFUn3pcoVwoGbyWCzm6KaRaGsT5yWx
t6J2CbdPJAtA0zFMkT7Qp2xxMHt0BaDby/JmiSSFuWit1MUNJivGNmB/IY4VYgjqkzDXebSeZxKV
TwZs4enbO2KXefGO6lnE8VjgdREM0r+5RKMZvi9rtGNus5QP+2sx+RLDY2LV955gjpXJNFG57IeD
UXOhgKq5XxAGSBqerYWmmyisBLbLxwUIVlqRmPSbHkWhCzuFC3bCDcXFkfj46qxime4rya0WOtjX
0L+X9FnREpn9t5uR58o5xmu9/hArRWJ6S5k5t4gw5NPROcAvLb0wNAN1WPVEhvhResr9CbG7gPED
7aJoSCrefRhWByGLe/6/jq5tIqNsFf2JsytVkaNucfFSgCDtnNa95kT3NVuVdsAfw0r3Xkdi4e71
tYbAjcgWrxSKfcN6C5SWvF7BlgBq8nS69V6V4NvGmCJ8Z0ecGnDEAyQb1nsyZzZeWQ1PRhy0QxzV
70iKEAD6/+GyXcTQQWmd+KvTh1WjvXXF1Fziz3mMSvvEKmd7lfiTzXeDdDuIcR2ylSUP1+DvZjLd
fhmjyLa+ymCrsvGDK5f0c3g86jcbfyhT/HSvkWgJXfGTYixKYKaFX6eWnIezqyT0/uz2Sh//pyxY
GtiJgWorNtZ81pzivdjfrJks/n/BUzpYwWbI1pph2f72+IkPK2kqt7yp2AmvKL+hUHJo+ezDPwPw
Zxgfe8AhKtouEGvBf3XQAgrYHA/G/DWKKeBeoiWAWxWVvmsOFkoe3QrJtBpcNDfdkqhnWRVPm/X5
8JizUaTXg9wXg+o6FrjvZTClveimJDz0z8r9gzJXtKVkBAoBM5ELiacpAzu0u5dfvsaHexGH22FJ
WDBg17icsJykRIdUnzC1kFnj+gEmaaERuSUd6SASSdoJI1/2oQCErCWoiMCQ+3I2hxfX2gGPKx0V
Ut6R7XHylsYr7HCUtC6cLayK5M4cQgn70X2/r3lzrZ4deMwTZjulmkbFO3bI0PbzPk/olaeHGhU3
hkmd+UUBZb0nM7N0+ISPCww4ctRHSbFVyG63WdjW8aVa0FXqYMIam7IoZNNuR8gCTF3s2aM/ZfEh
s1YEN0ByWfPy+3wJ39ROSHjVb54z10WKYQAnHr+BSYsifyuTtr/WwmwqVjWmvDx9eP8HNxgP19cY
x5SWWROYGfsPs9vVgEU86BrEvohYm7Vh6546ScQ1cz/5WNRxchG8A72c0ozYk7OV0UBwwkHmlUYF
U7DA/3amtRT+7nreNfITMeYONthU3KQrc4YO5TapZgtOFPVeN4kVDecTnp9r4HNpCU3O+sxf04dh
+gan5uZEBA68lLSmILxWvRuSf1fOBAq1Rm0PYdWHIiKnyIrKcmWwuWtZAGkBvdLebYSGbFtzwMBF
uce5NU9//+n9hEv7YHsJD0hgcwGKHJTFIx7FnATGzvXKsaGtDMb/ghhKXfZGB6jNtr5OqR8+3lUv
GnDtClEpy/mOfywvZ5HuKKxm/iD8EFrwVhk1e0FayNgKrde6CIzFIE6OmgvGD+6J8GE6QP8e2GTi
JkeWpUGQuaH81oC99rUi/mcsndf2mrI8/zK0GJgDxgutc6y1RlCHlkwUKS/GbG7qqxV0JSMfvCwS
MNeTfk0DqbBJCI/Z/V+Pi+zVILTMsZ02H8FQHMoPWtmT25zPVgU3VpetvTb2zIXIOBVjIiFB0xSI
4LD9L2CJRFIRx7OX9aVa+t8YjP0q0fKIvd0CFpcD1iX26E1FTS7qI5uHu3b/dm/2z4GT/eGYQUoj
HIurMoSh3JH8BFVSf+JBZ12faeCLHgnLUIuCaK02on3ag+UNe0RBtus2T5ncdyvy4lq2715IkFLI
7GNLRuohNeHHiXjAPcyPhK6R1eLuQvfUlos7944ba9rj45FwgibjYfrSRY4FSm/FAEa7/Wk3L4x/
EVaPMSFvOJlFIQxQR7aosan6iu8V46G/MgBoXs+mZ32BOPsH2WbuJBJhOOvQE33kBngLazEMVu2t
NZ10dx/ZDtpVpAFYF8ft3m0Z1GUyrIxgBYfH43WkTYkb8itZ1PzyJMhWIkCenuvS1fVocelCAlOA
I/dPJlaAqWEmUu6Pdej5xGLbKhAw73wVs3BDw1VHJE8gvZlXTSZ3yNXFjFvHQlc7igPe+qIdibgz
9jo28bITuUEBVZZ8Q6bzlIuyG21XhrkxR1bVN6Q5MmJuKeCY2Zm+eaT1k/kL+HgqDAQrwnHKBLoa
6F/swlg31Io49P6G4eIYpGQ7Fke+rs9d0aoyczwA/fai32R73o5n1jERU3qW0Qzov5Zl+4sNUgBM
dwhxfTutg5JYBoQW1H/uKVhmcdSyTW5MpuwmrVjp+VtcQwMzoVCpKKNI7X7+3lJGHUR2SM5JSIMv
nc0hgUQqy9ecJE6JbY1XzGqB4IW37O8gjg2xwofnMfQ/pvmnzHDP6zkpr9NHHLj2o6hfhGNt53YF
+kY1AxmRV1aYcMreZQMjXwA8/dOdJqWo4sUN0q3a7hOfzz5iLbkZKFYMBNU0UDfDRzgDcMiNzxYP
MAAMhQJ1nsUWptj56vimmnNSuhmQfir6KDAJ2ywMx6eybwjzOXwamiF1rz+nz+SDnhPGfpUh5+3e
ipvMZDOcbDGS2hDtzzbR0ZapM6TONJSUTgT+GTcH9QvKZ/Y84XAtGf/o9NO66yJzm4eXncBodl4e
1piOpllyCOFWnKBhN7IwtYyJsgaE2vJSW8O86Q+ZHA+fBkDwTqB6sU6Jo1XVTccFwFsj7Joe3P1B
bAGguoohVwot7JSbWeFUsVh6YPM9597mH0775m5VNKf9CJFSQHMiLzrq9TKJUYbz8kvRt89JgP+E
wYDRcAaLiKOcM7QTGZQX5q0gWVXc7Z+SFUST0q/ZenZVOfvcSXc2Z5de94SmLDNqHACdDra5u/Cr
OvJFwzJQnyt4nw65ZBDnLQ9XZE2LPWyk3LS+GOATs8MTOj5qI1LCtuuqAVh+B8j/osRPeFaLNkSW
LJNEMQE4p+Tf+CB+eXIX7iyS4eLtKnVrlUz8eZR5K8K/wGB3uyh9jsniUOz1BeZL2vNNWS7w0+DM
+vzheZ0VAH3ochsIBv8VFxDf9pZIRK0xCcZMMxxfickTh9/HUa6/+oE4O78fCNFLKE/tBx7ltGfK
mM8AMWBtBsg3aDdpkW7lVEGSGf9T6w65iV2WcqwRht3tMu3CdT/8u3BOicafN6JMxU8fnTqe7aEv
GPbJNKHhtnp1DykvsOmY858zDcfR1WejI79nf80aIwI8BOnBXE9n+HeCn9q2+aaCX7/LREXw2yrl
0OEEF3pxbZ8h3A/IiP8E1qVfn78Ot5aBIHt+0ngAtl9ba7PZjX1JI/OmuxeaYxIcsd52eeZ2xDSP
cwqjIzcmc1CEqAD/APLS36nBi9f20+ejH1GkA5VoZvjnBtiJPOUBAq0SUkSayypUVhqswqSwjgSG
LI5otZJgBwu2CunveUUVLJK2kCMgohyPbRQXCydlcurDKv1a6GekjwBXP8TJcNOM4RkVgoSZ13eC
Po/9iQp0+s3bnzSCA89v4SvIkpNlTBjGz2sYP1nwQMGIVsYUNsfKKpZorxAUrmUzS58IuFYS1IUO
IHIT1F9qc1KXlDvR32F+G2XUVlvSowhXo/14XkDvVJtw1fE1W3mPjwce2+gdmbreD0GIyPJmJoLd
/RcI2iQVICHvdrjLq/w3K8Ado/7b7f9VDM32w25AtRGLws2Ndy15e/b+rtWB9ZJ9u4Sw+sxII3MN
XXDmmhcjhx1K/Ke1KfbgdxZNJ0ST2QyIa71W7VWR+s533zsczyh9h8v3O5nCnPn7SBbKjk0Pz4sT
9/101u6thc1C+oUwGpEgdaI9jOdqdcWN7H26cRc3EoDAfAoArA5UEhBXKOjJ479srZg40fW8w96t
CAE0/uiMUA7OYGjk4mDbrY5K01TiR1nSQl/u+oZFEYhG65IQKeffTetK3pLhcnnsPbSR29Y3PjAP
48ARSMhKLCfavHYc7EWq4Uz8ZHMqQ57rKvL20nw73AGm8wYAZClEixT3yVbXHfokQkMljPEexp44
KnW1rTp/5hsBBHI8O9ntqauZrMQrn/9ExJ3TXDpoVG3oACkJmKxTGEjiAZEwCHnT7mXy7FdSRERp
qOIC/eYdGSC65YidHHp2GxxHhA6TzTD5rP9z70vMpLS29zGqIC/nkS5CZ22iT3CB3j+FbbI5Y3A4
JnwRWxccGfQRBT4+SZJTcv0j/U3Js5Es+qKIrPyMos8zpnJzhrkCmzdeFj3Soa48erGUFGlY2HaD
fXNgqnYDlAUw2Hoxl07A693VdrXMnjc5M5P6cQfmieNamhMRwKbagUBeg8tbBtVo66T+l7eCKGZy
lGcGeFZ4htIAShJtJqgh37EV6U05y+mvIImXam9uL/9FMI1t9x6F9ZPOCutm2l0KNrje3EsC7Gz6
wdU+AbQP8Cj+NLFa1lgyLcH3DMq5VYFiDvFAixdJhIDc5bZyHWD9Fuv8gtxodMQ1E/wY2T4J+Fi9
dR3Yjt9taaQLO4ZFDLPjUHwJr/bExlhxWJYCJGQ7PLRgSKg9M+zJdEIDwLWcyMMe7Fszu+u6OUuy
7gEsNc5IZnjsxLvlPu72niCM+zeoW4Uhy+GIv47RImgj7N9shXtEyVK49dddGz/mFxx7bzHm7ota
fcuG1v311SrtA2NTDXb0LRV84p722JdVToAS8nfnaV0ETCadIGveRuu4nZaXRSXEmpmQwBmu+vGw
VGVaLt8m2KwXD1LcSzLNGi1YiI0xTG43nCALhciL5YY5QeuoZ9fBHVZafNHJIGPo2jn3/znr6c5A
Ih6zYE/X9m/xnaKz/+JxbbBCbQK5e7Ahq0HoRAjzvrZEBrvPgyU6EOwdGeVbrpfsC/Fz3QyiCHm6
m1MHJUSkg9Z9oR8AcblhbfUBraWnOUNfaA30rLgnStmKLYRSi6QmNFj/OcBmKrUnR7RULmBlfvv+
rOQWajjz39L5jMuaPJvxUvLtZFAY0NqasGmeVqF6kznAOUCf6h/wIkwaSD9DjE1Nn5OSLsf4eGiy
g3CkVhonzsGFHvCBZcdi47Fdx//GRKFjz5zr/tfQDlnvUOeJeT9WcgXmzUAZbJZA30T8DQ3C1jyo
4mPRm426bSmsEL5Cfp0hRn/6UaeKFY1bhzBXZ+NAvwHiUQ9UxPxn+gF/hU8VdS9vi9MuAxKkx/7x
YHIQSymCDkeEJarzBqqt+E1zy/SQBMkhbqer0Zk512SfGkO1bS1Kv9nsDzRomYVYQronc76GlkT3
QoAHi4ULop/pt48+qzhL/Q2s08S+Ur+f5JgXt/LNDu/AfbogXJ1R2VoCsS8ZPsqQrTj3KNicUJCD
gEhcFuJA3urjS5iEgSu/uayoAyMz5dEG/Va3PQkvWWCCZevW/iKhABWCQl4R9lH0Ro2NnNyrk7Uu
pmWHSP/nFSBu7fSW+7vrCMwQ8XV24nqvAmwdQaThmMKD3EtwTfN6uEOQSVTXjPjbANWfhtTW7N5E
tIv9Qi8Kt6FzC2Z+xFSYxpnjZtdHDFRl7M3zbsl5NotsfY1wb9gTgSKKmaIhfNzPKfGE0BcutCpp
UpUbxfCnPyaLvfjNnfiDgsTf41ogG847XKyhuUlcj2Le2qck9AZCjkG6JztQ4+5GTNAgHPgK6UyX
sK3OJVwxCt5YMMNytFIjZ1nJo/AR14ltwnJU01SQL5y/ifmMXri0m2YMokipLnIxqAieTGoTLTGq
7glJyJ7fCko7Urhw0vo3ga5R/a7DI/jGk+2Zeo2OdySafMTuN4DHYC2CLOxtbPGpq1r8RxS7TshK
fL6Ou/9/zCZw3UfKpx1BA4EUfU3Nin6EfYThdOHTiOPzAcgYkh/RT+lyN8yyZzeIddk3hnekvt72
SHrWedf7bg8pU54LuE3KHneOp7CFTtHJbYrlG1puNhDFUhPbGf77v5cC+DbvQL+t2rEXqBhwLrvC
Bh8bL69wIpv+PXMFAyCLU/lEfqIvjlBTfXnjBQZmlAbLg7prludjXTW+1+ZWCTRjXSO1JQ76NkiW
Uo6mp4hu/z73rKubhhJ1rZ+eievPK4PCLVH5Yy8XerMvQdLeFdaL8vxAtDjDqZz9sT782xRvp/vU
V0IRYXi8K78ka9c9KdxSYSsn2GKSnwfmg+LLS+qAGuVoZMWNq6cEglo4xyD+qbfHrcXSXq5izlnx
ZWERgF/ubMhyCGFLdhvTiTfJRaY9tECwUyfAXVjLTXhrb27ORFeBaj7Kf3p5+Bz7cH6kDUrm59ry
maxZqctASMwu3r754u0Rq8eLwpKdgi6hBBKORHFuNHnnxhoWJ1/7X9A1q/iwnxNGjXW65ZOh//Vx
AMoTnw6G9W3lvjy6pNMv2oJw8UucUmzjSb9q3JQJQgYvN7FhNhe3Aag8aNoM+IRkftNRgJIJlo1e
+GVQB23Cug6No+nApWURVmhEI9FmH/J4n7Yqto7MvLg+dpm+BvMGTAPd8xc5OBa877h6Q/vHc86x
rF9i/uSn0OubGg9Ui1g/Me+yyWwGRicvrcBYcJWgQIj6oCrm1nhXv2EW7MO5MmCL9MYuenCXk6K9
RPbN8Q8g8MOS/3c+nNpPlXqxFZ92Fgja6dRYl/4wZaJqZ4ajpT2XLGtBiFsJhWsfGaLenyFweWHZ
xfvqn1XuQuPL5zP5Xce7RliRdAEVHH5lc2DnpOAV8k/LnGwkj40mCLl0er9lr3DnJdl5uOTasOxx
IfuQ8uvRslKwndNL80mLftMHV8/ANqci979VvBNMQFOVlTDZdsDXkHYnwNWmjoIYmaGPvjJEjc2e
Cvn0OE5Whb18O91DkJpxiD+OBKNW8BMxrKBKvwPjlHXtrk6rBtXqAwJA90w8F2tQe4vryKk4FlVp
hB2qBIoZzZ2dSMas2Vp/vvJI58lWgsslLjBvJr2xTBnsnFxUsQUZI/aOniNCuwkPoMqAfNcuMYvP
XYIghyE5meQdrCoB+qFzIeVZ+IWPZh6scxOcXj2LcdQNFoFpJ/KKB+4hhpVHKl8k+HgGHsC6YeIm
xWzAsDa2StlIKUSvit7ww8/EwIeXAjNX7xzLLh83mCvYOENpsBlEXsFvtW6pqZ/UWVfNYiiVu4dY
ccbCTVXXFZp9cXjYEmWIBA8PP+xAnMdfGyIVVF922s87JJLQ/PfYru8laDQTNIHZsloy0U/3ccPI
74LTtvhPu33utup35MwksNV5RGC2JxjuKYBAVKsd7m8RTQGDbMBo5o4J6luJWX3N+kaFcEqgDbjO
3aRhHtGIZGFCvKa4xSiX28XjXEtqqkSmsNy571+DbQ39XyBgSqzIvEWBG/N7GON0GvImvMGrAToq
DsFYyr6Q9TA8AhiLt49RfQS66NZ4/m7bcGlgezV4qu05YdVYxkvFZa60YdcV3O/pnQFutubHkahr
TVMiPSegU3Bnnld51QmUgZrNFGbxGbHZwKsX0q18twExAE/tTeQe+6haZ3Q12vafTAIjlD0AMkHk
yK/eS3A3rjqjfSO70t+4CCFu4j5V5nEsfI9l9valoGErW3AO/+FN0EHgz5SraF5M87ZAMGSZRakp
U7QpwuJLX967oYLuioDG5Tin8lr/4RSP6DrIKIyBEsyNsLcnxUSyL39o9HgeybCCkM8bSw9IXwAT
LWSNtVtPghKuae+TcMTyP2vYdq8PEn1T9klAAjbOXnN1nSb0fswuLkvHlgWcHHgQMnilkp3LrDal
kVla+KB56+YaRlX6Uud7SLrlNMgfkj2MKhQEYLCUT/H3haes4GXSoJy++QGJFvuApjZO5dt99ioB
gg1qtZKHNO1aFJpERx39nCgYpjx77ggUppyuM2pLB45NFwlPczgYsbPxTR6cvThPx0kSKk9qZrEQ
xYGYfr7WfshVQvoD/OORBRQjrPGAWxNM4X8nKpufQl+vRCIDbb5Fmnij4D/3pu7+MlusuhRcXoFZ
E/LkOCsrpc8swcQB9abiTYHADi57cr8V0TqLOyodXKs4OUFlvN1I8F7wSSUCFEnLnABM2udNvvZ+
ljmO1FJfN67HzjuKun1kyQgYBLuiq7jAKBcU/PDrcMUaaKrD4IP+SM6C00Xt94EvvpSBxXN+xPOG
xRSq/dWKZ3BkPTLDymg8zffKfvAKrF8t5zVWs+BfAnsCSxOoIlUwHm9fSR6Bfr1UPCOizhaMUCPN
C3V0PIPkN2AxqkFDpsLKQ5if8c4qoVTuJTONgMY/V0c8iCB3+cmx4k/gSloHtDDowqFsvUYhemyq
7DyEi5TCAOd59RqPyueTXpQc/G7JwosytH65x+0ernwNIk1GrYmA+QaDcxaWpi1QGmubUc6jSXwN
ElTW+C+/BtGViRpSz4VHP0bruxzkaUUSw5qZ7izJyl+Q0zKA/VPFb8FzbWj/nVJTur/dIuCki/AL
eKJ4QuyuYFPT1MnL6lCDeokZ8wGFavUfTwWezIS9zOdcVs/LsmIYLFoQOe4grsP2owykVNyq5L0e
oJInrwwmiui+RgVYnDaI+Xj6Q5I090vZxzXUkOYm9wp6o+d6YACBgDq0wZ0dSEA1r0UaZKAxTb6Z
KRTjiB3gy8iSmb5WlDaL2dMEZJCztqw0L6aTaMMRu737n9Knh0JbRv5zubRVxYKwxu9P3ulFtKbX
xpztIqGjp/ot4GsYi8ZBFocdHnCyMlQX1Yadvipi5+X8l/eBlTKKudsR1w4hWqIiKqsjmVtxy/2T
y8kFh344Wyjj8CWD04OBqrbMfppELo5twUVaZRPOLiMOptExFu3+O5APHaaDSG6uIMkgewuWNqOD
QZ7VyjYiUvEkuT1SFJw6Mut0YP0mFJvigD7mgZtvC9QuCN3Pyn7++9AO4Sq646z2+OzJBPPNvpmp
x0eYBBmdfaeuc6xkN2C30zna8cDce3wtlRc055v2Nh+A5R89Jy0naJgZdXwUP4bLdiyohyf24cWs
V926aBXR8VDrkJEdraHsnzn0LZOJRiPIRjApPMRPz7WViJoJ17WLiCcggwHNBcRVAG+ERIg8AUQS
dZeoT5+ql4GnfhO/Tb86Qm9rT1Wi/ZV5AZzEyjJ1MATM4wxwIH9ogo47x9l7nV1a5T6YLcQuLAE5
1f41wwAqvd/PFzFJ9U2hoYt1JxJG0uqWlNT6irAsbu+NPBzo56fRmlWDOxs7icSyNdBOjm6YAO/q
VtrVfJqn9gQVc0Oy+SZww0BagS3RBEiLpGhRPNeksSCKsUole4tIwNbaSx3zUX2K5GtwwCeAj5So
0lJKgPu4vi9WjrN2UnwjUBZrXrZLuOWEE4297oCeLLeapfqyEM50J59P8rjXzf0wrJCLV7EgFyy3
Z3e/pYtXpvyCiWkJ1p/swcLJ3G6H/lFCaHm4pK/b1CAL5j68BKYmLBfPU2Wehp/aFZpVY2T1WNfJ
muEAAoYkWWfqmMAlbeDNrN0Ur5pPdZXgAKv57tj7knUhBoXxW3vb9hykG6oaUbNyc6bzeLAOIOn5
WXtHtRDHZZWPKq4I7jUTs+koHCArgBm5KyOhoAubtAHKV51bMIormqMtnbYzXeCl2t7ZX0mlfKkH
QNtkIQtXDWSba8o4WGwL3Cqa0FYIThJOQA3CaZ2HxdrQbVStIw3ZuP+MuW6wrr0WFEeQaJdcGLN7
uVsCcTlm9cB+RFdTnozkhLzWIe5aG/l3mtVTO8y0IoaVnPjl7hmXdny8t/6RB7uj/Z5X5vRmSb7c
7rKh6+03Di+2VoSC9hxqV2Ii7uMZ/jbpFp/G4HOVcdP47wmhc95c2Flm7oFdrbJ7OIiGgxGnCTNH
jBjemtsYf4zWsDtmk+D8aTlEKewlVMpSSijTZsSJsZGfhPRF7SiRtB+pWz1HzC/qSzxggEeDr72N
1UO6ruS4dbtnthN4+nmDh0H52RpF8GspcKch04O10YHP0nX1MBj6zTP9xlxhEEKS/24I9AcOa5Zr
jtK/w5gniE7XZYBG2FfwtT918g0m90d7bAlIywR5pk4Zyb5MlbzeYdUNv4vQMshI7WJfGlTCklIR
FPJRx/RXmzUMrEWMiP+1Z4VXdYvUREYU0DrGWZFbulDmn08n16R9Gl828kUSmY10XWRMl6HlALGO
Si+8gg8Y2TA8/eoVZco8nUArkgFAsJsfTaIctXge+DQvnGatTQZqgzKT6JZjJQU1pdl556JE1AYO
HScg7LuFT4Ark7GgsMvCwHGnhPBWQMvWq2yFgLEnT5USGq8BkU0L2dWsDTTM5L/xxnsbyUmUy5lr
dYlyMzb4WHfHzze8iae22w8BAre15zK0vNDs76hE3VbCWTqHm3H9NAPVaO8YMz4mGeCwxKzn/ZeL
8OkADEc6h7nQCh382nUANF4MxJMj8U1PcoBu7GtIXS8i/UiWIAT3PBG4TZlhOVzsDDxMuqOV3MSY
bSE5OfTodHyclO9DmIqrO1xBLwXqLAwvxoFL/oa9qCmcyqYd9lFRcaGH9GLdVqoOMAGObzTk9EVK
kAd/LeiOJEQf3zfL+k/+oojLcOTX1Xgx8UCXJFlnDVnhNqPwPjDf2oJg4vF3DlzlPreU9Kwt/7SY
0Og4cTREVhP/1MfBGzZTLzoOjWXHD5Mx3DjegML+iigWHyi5mE0YkFurx6RLxqY0vfwN7LRCNHbK
VTBXkfd+cVLbZnM8X5dMy/JGMyvhVT4++CXCLYylc9reOhHzopAfnV6klM6HpNiczNOf2yBG+i7P
6u7tXie07Jsf366OkU3qA1Raypy3TRp4HOy57GeM4JENzAFZ9/HI2DoOn1DVwXeaA9muDBcc+3H+
RZzYyx0EHui0V2Zefr0jAYapJ5/Wp8zKMxUCrJi1mK7+/iHISlZeltbomoB6JM8TIuzauyXA1oxv
ftC5ZmYkwQTN7fAno4cAmINsah+dIDuo1sO1FMnz1P7njK2s58UzQ23vmrxTcOFTGeYAAvTElYN3
er84ZpkpQT/ujmM8DQ5C3xJC8sCWDatUY4JSbeVYeFcZYQLafCXZY8JKedVR/w4I6yf6Yzj57Dpm
w0R8kpje2UYxb8Y2asTZ0JVETE2R06PFjQvAEkQIuCxIaJoUpyia9nAgwP4sAP8ruHkk9Gr6EhOk
FcDsIaMB+Cy2/j8OZwviC+ux6NMKHBRwjfb3UVoVfW00x9idsBgkoNKcHA5PN257+3qfQaqYjbCP
Dd4OQQMwk9e5MfE2oKo7WlEjS/eu/GNwzcjRhBtyjc/nb9gAOKz25Rth9Jepthk0XUlQWGuW4gqz
+ZXWuB/l42qhOqeciGjCLwvzTT5krwtKYMA1/48HEfXFEAR37KK68x1+lnF9ycC31ky88dd6PaXT
3in47GCQgguKqfbjdHKkib4aRfpoGVsoYLUgwooqOfhikvXNbn7tnkvV47AjOVlSZAc6p0FWasml
0UOTY3dvGPjN8wnvKgAcIz/ueQ9yS+AhPO5Xtm/7IUsG3tbYj0QkMyI+/8/M1qJd4TzaX7YgKtlk
EBcBogjbGakV7oqJjLo3nJ7Z03e1gibFQ1oPjaNPx5kapguz//r4eIjEp7TAcvji5DKZsJPLG6p5
S6lBksB4ED7KffsmUgZy9PEc3NeJmJIRvIe0sGVj+QNGbIMaJoIKLjHMsXVFjKznmwICpc6RELqA
DXRic/wyUlDaUTRstQMySktOI+gkzleUh5Tb/uSJ8y6om22wh3xo2tGRpf6fpfNF0Uto6qCtortw
ozlxkRIb0K/ryN0Yk9htS2N5aTsDz0vRjcGAy/EnIb+PqywctPybAYxbwATDy9i9+D7T5fJ2rbon
m5O3vb6vxfeFlK6ZFEV0fwhQSoeExTIVWXmhRIFRr5S0laqnjtvr6l4h1Vm44t8tDSyHE4PR7hUd
PRA5HBx6Ukp5JhpGp1nm8A5b4AfRuRCza2H9QCBNRH8eg6fmPhs86D83Kcv6gENk64bn38oZu0QJ
Rzt81on/pBZLFre39zACeXfqWI2GQv+FRtv6Z8qjcrQLx4gvfI1JubtHeAk9K+FN3q8frXKL79D4
vUslohUaVRPHRIkzRx062ymqRNWLeVD3m0slXRAT2lRB+HHdndOG5Cq9hp0rGzvyydu6KmvaLyBY
/KaP9og5FNRbRtJ1E8JH55PkjnVZBf4k7nGlAEXpCacGdLXVQGQsSFB0BTOZEIAE1OKyQ+OhNpdf
N1XcKMcax16WQ5ds3T59HplukiAPxlMPZLkFvrjzdeOyS8A2DIf/2MkNUUWXzUJe0SrSIdUlUoOp
xxgWxHwYVbj1v1xk3ZRD9bynZkrV754xYpU+BKtxp4YgsZVyIPsAKD37vcHYLAf89Hn1hQfKK9Kb
DHN+R0WzJqOgXBYv3nxM5XZAHvlCP98EUwIoXylfRRkrNGmBfiTl/d+gzsGQqw4DAF5FpdtZk+eJ
v9QTSglUgDaFPu2kA76JkMEA/qGmOojGeuLXyCvfujbXCYNXlDBshHjGTZzrnpEsFpXJGU7sJGXP
Nx2lIRJmTXh9zSfmpjjtD/3wN7LmCqYKLFgJaZCmfSuOXzMuG19Kk+W7eGJdo7nlGYneNFuAHnDe
xzeB0HK7hDlGfetHXWzQO0PH/+FjvPY27EaKpMJpf2YkvJH0YaN5OPKbEmMcaVucyWFYa9rrDY65
rMgJPekNUQrNFDxmAUHhMATbPdkUR5vULLHZcGNZ3unDKAmMYjmngK5oC9px6itP7NEHrU6R52nF
gyDLbcMIABs73NGIY0XWDsxnSsMK6raAZztuvOuFIK+33GTiz0PgjEJd4wbe0lM0UKZCeQL86NvY
ekDbynYDAhdiQ6PYuQtOyJI8DnWqrrgbyTcDlEBZOlKdSPJdxzvmm1KiieRVwKO/1M9dpaXZUDIx
uvmfAXdW2ynbrlTdEKDyTx5ryrxSFDBKe1upSbys0p+JGvA5b9MqKEyH0j68y1Lv+tGEaAapLG8Y
+bJLP3GBaGchp9RVoflkbGoOnupCnS01R/bzwhRYQv2HGhhMTKRfvxJZVho9OYXyv1COxwXK8rQn
yFlieK3mPacojrhb0UYToxn9fMiZKVnXdsDV/swFe8XA0dfvtyllRCQFSIjO14i9c5bEyXZZJgny
Hf9d6xwrwdkEcXSgeOLpNGYgq2AWsE/r2JELWfX44UK7FKHYGTlCU5dumKJSArfsqM/aJebEX2e8
GqQSKsId10mcO6rPKxpJdYV80WEfcNe13BqObQ8PAIcr399zKi+y5l5i+nGgNUmDdqpPqJpUw7TI
jl/d1sbv+Cwcsa5F9pHi6pfnrMkP5PO+UKh3i1EaJxgEYAaJzqnRb4X9uQhzlpFzejFmipF49VV+
mbImzB5eVfCtVxbipTxKswkYq1j9/HB8PoUhjJ9h3WyD+m9qK/uBCOPr2De/wZHgJbuqH2HzaF7m
iVXf5i5+RkGaUPgRgQ7Y/s+V+w3xaVqHmsomhP4YSoFU/OE1H8eAfQ9oNM78MMJoUCV/LWBc6clk
U3O99Vbbo6lVl8Avkgd+7MGRR+dgIY5+8RH5rxQecAL8L0UZCiiUEpi2t4zGUbEQQfvQUE5LSNxR
bUuKjR2Y9a2DyuhAv31XukF15f29sTg7p6WDEDc0XBQigA0y9Ap9qWEijyjT9xB9FSYr5Frj/wx3
MTWDf30bOUZA+y73rwfKkLLdvR+FycJEGrmizY9/EPq48R8yEXW/c4KnmZCN+u/TZaTJ8X3Nv1g4
lc5QdkmGjhswSV+Bp2SwlWKf+iTbwzZQUwb4Sf6TOlLBAbo5Ze7Ng+RuxSsRJPkb38JkaEDcny/N
RHxgmDlK/BWWMOnK2/Vt7xy/swecCVYu6Du81FBLBcKRN7zGdYk0tSbdrgHVm3+dpYig9yuB06JD
6LgLJKGuhaYvSF29I56l0pqbxJ7Q+LgyLDQaHXICYqtGef4/wjD3Pi7DEDPoFdNf9dXSuSZZF3Jb
kWXkC5t6kEFhb0F+gb0GzlufnXGTD1pDwJHCV5gCWIYJLdlEWYUtsdYQtHNG/4VrCfH8gzJKxRjs
tHerZXr0DdaS5iqflarvDIXkmIFAMDDB0/bJzLePlhfZHi22GtnAzSE7qLoVgsdBDOMaY9DmqPmH
FB6LtGdhIeBTZJafI/WB9m3VyJuAnT0zbNU0DQSLjsaeZ4mrGsKpzySMYPgO+lsh+3iM/W8jlEdK
sHWf4t7Jy9VX1V+tShzZ3MWgHZt81FuNYKy8qSboTnavVFaqBg+Rfoaarf8BlEFqDwVerapQDNcZ
sV4uik0LIan6FcjMqAAc+ucbuEHSQ/jWtB5rTSwo/SqUCGd48QigVrOGQcI+NKAdPA7SnwDP83L5
JzVf76JwejN0M7ZntP/332GUy3mmbWWD57c66Pdh1FR77GzoTjzwFUJRh+h5nsUilTxoX3jaUnAZ
bz5eXXBT3o72tD/YcIXu5TdzUg7KNixmp3WPUuHMxzpnWlvtST6AULGYprvLSjqjNVmTXAc67k5z
ga753tDPgHJDVbjtl0Q8rEst1GvM1s5KCFFWLNpa0S9G78uoa9jYQPgIRI2zjCMmcQhEKbdqyu5K
GnOYdA32cNS1nB6A9JHsXWsici3J1dECbb3zLNZ8yG2As638GDHBeBP9Z6BD/EJ0N6/wBKLqha2K
omLI5nkA+uzosgNdWzyQ6z++KHm/UD8XxZ1DtdT7Qk856ZNTHDP3RJwf4ubR+o8nSK0/kPvW4PUc
8ADA78ac6UwFie1Q8HBomR9gEJUBvxks8MDICjGIVnxpMD8LO4xhR+zhXkaPAYPmtCgoLDk+hgq0
jEyVh7puRJ1zsDgqop08XqyIIRr/rUK8ULx9a7xdx83s6mW/FVrUJdKmVDk7l1WQLulEQ0QlQ0ux
t2NusXeGalv2svw+Azgdm6hKhAA3x5kmsznN+nwXZ57j2vA3G+k1R5ehvGBk0Q4p/NSjCcArYEAD
gI7cNunkyPBPOy2v5i7zk6OQx2HKTzfiNFQnfJTX+rFMkYDILRrWytb4DnDNrhWgBAYwV7rrk5Ew
0ra+eHkhTMOJ5axK1wfWar8WfLPM5JPBsLzM3zgX4M6PcaFmGhu19rzwO3cFOL2/TMcjkM5a2J8N
oPVrrXrsAAKKxg3V9vUPAZstImKChHGnBVTjLt3wxgblsAwzj3lT9aMc1FzMHkPz4C453s/432k5
0Q2bCm2v4S2USNurVP/tIn/8tiDU4c41BQnDe1VKK8aLv1c3XcMBnh3jT0WEL+HmeNRWHktJuxwu
zQpUMOenWBqJykA7em12iB1uuyFUOvOg0TU8fRS/VpVdyH72xCn+nUJEU2VXhsvi0Frm/X8MHYrY
AO77QYE7dsJZCZCB9CBRYkHGn5ODOWL79ztJJLGS2SPdYFKVnvVd4mlnk4yA0yu9c7pB99Aykm1L
MZd1BNB7zR61SwKDQdwST9CyWPO2q/g6oeNvVfwXukN1m9q/0OC8RWPdc84gKEYFdD0XQ00z9SkM
sPy0DR1p+Doj3g/Y+Hv9LSfJm/S6kredYAMFWL99driNxT8Ram+lfbpaZSNTHAMDmH0YOEXtVbzf
9LSgmrF2pC3S2Jq/wu/1Kv1GmQAnTfKElahoP84pL08E0CguBAYzmGS1oW05mdolH4TuEFpAaeIt
V/uZgGlKXSqEYbi6FF104Pmm82Aad+Zk0DZDhqheXEHSWL1Nks4XU8p/wIqmFrVFxw2RQp5tGyZ9
Yz1SCunAhyh/gpPf7Q9mDtiH3/wYuAJ8CDFEPWhIlPLJECQ1mon4a2vmBpPyWaJs95EQo+ioro9x
7NxBmx4hvx+2jmiuD8gBaZyDreAZF425eLWd0JvimFYDhz7REiipM/cOEdj2Cy3MQQMgqVBqnkz8
xJi6SswITJCASHajWW0k0X10+LmDbMsMHeV2euzjH21DCpEK63GS77sKQEhvgxyjo9IMz0q3cZsV
cRBZIxHkGYAGa0yLPWHCYEI88TGA8F+OeYdJsl8ecpcM/NWmrN238A07BXIznWnwczIISgdXDg7E
CXNarEeua1Smwb3p3TQal9fFiXDjaVqVk88rJtWwccioh9LrYkMrc+CDFskjZQuKlo0Uty9T8Hhs
7pnOHpgz/fejmNzjB6HFa32Q2YLIQtLBxBrkJQ00HXL+j3Je1gbXuoWdOK08uZ6MwhKMCCsVKVAY
Zqu0lAuBjF82JzJDclDlrbezjllqmSehCRyNuRJYI2XIaoMVxwVqdMI2vLpKucAIfesX2i81vx+j
i/7bay1o/x2RwKe1UguXPqlpT7xYHKv3poZEi2XHxZdtt0ZKOYy2Pu2vM0MIJVeIDUOv4mnpLdX2
w/AfQ75f2MDWIEFQU5it0PAsTHV/GaPhSTLd+Lu6ihJ0vWk7uHuAcGPwXNNKS+nURp/DdBbCEIDn
5lOJPwHN5yCaH4P0KDwF2oY/Wc6nNJcFnTrQ03vVvnHlhTyihhICDfw4WNuGa3OZezzTU46C3a1J
9DtO0uCYzaZNVyx+dMcBVspVsZTL5pzzb5GNOLmErPzI/JQXYXjHy/Bq6G7EN01y9SAqXSGrMyP7
y766H9jWJWzExl9l3Wn3ONwZolM5LV715kGqGSJIGFR+E9hqIerSm81h4UhbF268WZYw7BvZRsu9
8ESjsuc1icbFYNdrgQ7g0xulPpjTIWUgzPZJsrNCadP/y+g7faZ0v6TWe1scz4nA62rzz1f/dO4r
Sl3cnirqGoqDAj4iiomGlj2dJozVxy7taxCyulFe+QpXczPUrmgHab/0DZOjcubtmb1mtCcedDs/
ECKAL4Unxtj8EQg1I8mBorfYPHV6QQAdQM76Rx2rO+7JqmcV13Wr0Y1HVVtf4PTPEVZgTyA658N2
mxN5C6oRunUjmpHv6xN+AxktZAWO85jmVoPxHLZGCMA+Ea1BdtV+xHhinwq4gIDQIf1KFItP8zsm
9/t9yEeugAYJrS/KWQeTY183WJ5a36gsJUmPsoKnyCV4wt1JfrgZBjX99pXX9cAa42f+Qb7M7nti
3YAoottbcyDkGDgLttYT0GuuapJ73W1YrzsL3NPJJkRBC9VeD4C2JVpWV4xCrLK9xNPHbITBQSLy
CiLm7gQ7dq93AlI16YasLumG4iuDExHTHK1q8mcnKqgZTna0ZMn02jLiPaKzbWwJrrVkI4uXEvJB
2fJEekq+HEyYHJPLpSk6XaBZ7CVx5Yjy/FWYOZ6Ij894QYL74v9k4bi+30fF4xOF2ipqQL3U+oiD
ni6lUx3lL8zy4UeIvGrVlEV/M2Odqaf7ydZCSsaLhHSTyHCUIZCt8UikL/V6OTPz3u6km5JrPL+j
8NqXT9GH/8na4sDI6RGk1m/0SGkQ/rJcF8TJV56fY7DHmdZhfrldi72udVz0Sntd2+L1yx6cewCN
p+TcCDUNWbjS0DgSWcKw6b5AUkYN3vjDfFh3C+cMIE1d3ZZQNF3TFQyJ8r4PzS/CceJR4VXbwqVw
1p2ufq6dJoMQizCUhDVsn0JJSGaHFeDp3H6zgzaQcn7PZxot6SUt5k89VWPIjvFo/cCXalC4uQfj
SLzupG0sNkarqEjw+/k6ZXJG4iES159wyQiucowZtO8BDVbgUNvbLRGoiZ7MXwH1YCyD7l3gnifR
Zodeue4c01XjCrjZbOiWUFG2UgWKZENA6TGBdkazCfTQmmkngNqhSByBHsjud3iAesk7eMOQYN8n
rrpNSTQSB79gq9CRCgTuFDMKpLlRUJ+0sAR3BRLWoPncEyCAZs6bFh+NukEncB5l2eSjkwRAMIqb
MMqvJxkeIvxG5bjkFVyt57Ra9EWnp/DCdoaFZGO2HHTa4VhJALwcchwCl9ocms1HKzc4AX7EXv7C
H6odR719yEzxoSmMdJ+plg27c10lZ7vbCSoBcWivrJxAFE4tnMnrm8wZ8BswdK/ZCOz83nPNor5u
H4OBCHtwpIdslH7oTfHiHrI2yVLHz+0agc2TQWbh/nL4LnUVOYXLDcmstNL6ACQOukbySjgNvc4R
X0OysNeCw+Vv044r0aWz+bWeu2qO8V5Il6s6HqZ20VJ04lWyrwNzh4QxON7Umgh8O/ioyvmqRrJ1
dtG0sP+rvkMXqVVFjtoVMUwAViRHdTMS1ePvJkz2oby0Pa/hTa3bfc0nuRlQp3+kSzruZh5SfaU1
vjrBEMGQ3cAm3kSTf8d0pU2oelIFWY0kJkCUZ6n+Gwx3TJqu7lLiKIFBwddDGMlmEaXsuBT66l64
msAPptJNttpaGdfevMrshAjMF3L1qS/fogdZDwe9j2gHIaUNfIpsN18eQfe1W+rHJp1AUkR8ArV+
28D0nGGAODcS0MWG7SvT5UuAcVoE2cOAttISiyw4XUzeMN5LkneTw+srvzjMKkavuzvpsy3XN8ko
nniczEDgpZUOut4j78fKeQrSqjHRr8r5ihv/nf787qxqec4aCU+bX0IZxfPjCJUZtnlmVVtEiL0f
NBA8gp8pAXRYpxmdGvL/uz5TpzpufLXEEoivBzsHdvPgIijgs4+M0ZsU9NPEZooheHcmDDPK2KL8
ep1RBDfy44SYM8Iwg1UpBVj6IvNrrS11RCxi3yyHKFP8ZyLz3K0L0fRn6Lkz5xJjWwrLgY6/UT+k
+MiCQgFaO5a6OtPlRQzwgXChoio/WjBT8a8bGSWjDJ1/ygbhzT86uFssAnUByCiIg5TURpp5T9/k
w4/8/N5eq6yy1bGAiJOohvufPZ+jrvMWXGtqKBXQlNYxNIhwi8dsIfQZgsPuQ5SlklH1hQBBdUtv
IF2WgS8jxUbDmc2cvOwGYODNqGZOZ2UsH8GsL5gW0HAVgDUVqRX2U4xMGmvF4X/nGqflPVyWFejS
fRq8n9zR71uYbaeZtN7UUMFYxdbQxidTq29+jbYcTN5tR4/XFgSZ1RCW9Mwczl/rDDoKAUWtIuaH
SE748hFlfmmgiIAGcuW3V3TkwZAjfIHF9Mbw5rXvPxiwNToXRBrifUpBWcr0AAw1rnwVgCW8akg5
O96vUnzoJLiFZ/VbYvXWErjqQLc4oWjbsgjeFyDuerIqfaSmVnQ3oCamHa6sMxQDfw1mLZXYMgp0
+0LBr+YGGA3eMyBaF+a82aowDNkB97YxTcz7IjX9xcnIruNCCMDxVB5gGXwMIp8aKnynQvK7Sw8E
kbyCOKYOQzeuuaVWrSs1Dp6vbBOgNVlvPquJVB98TGcGCrqpGFm/9dTyMqHeEPG6ob9JAxKvfXap
EBk6q9syhFFYZLzYbqfjFYbsVzRogDXVo1QgtDon0L77W9xzUXkuRjqPP5xNMBb7JjFIYo1m+p4K
qxiwB+6k9QFYN9B3+oPkoRRM01Zznv9aV4ms8eVY63b5wIPymnBxr64fqsWSz48w+l/vVRaPCS9a
zWd8xi3MyBZzIrC1lzI6l55nHFeI9ryr7XKW7pzYKd0+qy06EM5qIC729yXpwFqgmT9Onx++U0Y4
g6xJ0RudOVyjR5ZjlGJ+B54LXYWreP44r+RXsJjPBVN85eSLnERn4D18BXc8lNv+990jIvEv5+Xf
v92uxKOP82DIij75WgyAeVZ5G7xzzF9MC7y9ZObqQ76OC50jJYAIZJpQETWEnMI9Ap8jjdW+K5lR
IAbIzWKQovvCUfYTKshNhLAK9PF0MvQJjIDYd4uWGVYAsWZ+AaGUjM902Ln2VVuysgKAqr486MY2
8nS7ttQhioEoPqnno6K2FpwAhDKeb/YMMntFXJRLTR8M5OMh56DpbjbHokubE3KfSZ9OeshnLOys
Ggg9R+tbbGGDtLzEXYalhuhPxX8u/+0j34vMXXyRRqBnkXxyzY2Bf+TzvBfDNgYcvkkjmLaILWJS
kxOYpfV9TrpWwpzba6yscbAOhXOhzF6jet+09B+fD2RbYSkKsrU/HCt5Lx704nY/xiBmjMPbq9ss
gG6w3j1L7RMMTjOkXAmbYRpkr3t/iI+sOaoCL35TqwGN3iD8hGFxIEf66GhwiQ6Pt3CICXjFiGel
D4jOHerBePBiLM5OLbTmAOuG1fqa/WGYVJC3ld0TqS8nka151Fjub6ESn8UG8ki8NB96/0V/zWV3
npQpE9/SCq96EddL+0yXgT/BuofxLU+ctdMNcbNwG6Wh8mX2Bp0cyVejTlLTqV7LZgvsFwY8AoH6
/zobrzQjy5v6FmONJ9by1j+XN0vY+faete0wVgH3PF7mJnDC+pYA4LTd/O6M2gZc1KABrmymM7j5
lx+P3o6hO32c0LmKwt4xsSofKU7Ep7azaSZj8oaIEo8r7jECVOIKJOinDl/x/mVpAftDPYaDyN1s
xWO8aTiRdmU7G12bFWxvQKoxsFPyeAJec5H9OpduhXtj1BHDB5oPsYuy0Y7p2Iw8OxdyxP+ngK0m
1lvX8ETZEmn+JhYf+53/j5E8EIvJ06gecB2Q6qPfZiSdbQTnL3ExRuoYHA5BHsEiPRtVoGo+ivtt
1fU9CkwRUgTTxngoQ3jq6v4Xt92K+WykcgGCCPkkF6yI3KeISukOoGX2zdxxm1A9yjGH639KH2ce
XaqrNJz7N/fRbg6o2mGcNYegKODFKvlS+xVx7ELEUAT9t+N9VwuVwsKe/cUguTgShdKroFnnU7xX
3Ipfv7vN5JOPnsl/VlqP9Oj6Z7hX7I4IziJJ6ZHs9y189B02LPcFYPHrzHaGgAyubqw+jAeNkySU
+noXgZH/og0DF4ODQqtXF37iP1OuYhEpczJrVr2u2iQixOBb7jIik3bzNbJYDHLBj0NHkuBkBkp9
oZKzq4WCEgIB50skkP2QttZqnpTToWma90XpcgnHUY+WoJkB3KxzfDznpgMnjcnrXrMYitSG96Mr
LLL5eoefU/LF2F5kgiGryuJwodaWl+s1QlpNZzFeY2xW+WEoejxE9w2iRju7CTSw0lzJO/HylILm
WEeS4qusTwt3Ajv55414977hBvu4fb9oY6K2ARYNSzHgXP7zUUrG+YeXKVLSIbVUfxf2pr5cKKs7
xS254P3SSMOW8/nAGR+B0tW7TzTV5MtCBu5cV0wkM6JW+ge8AYk/UiizkO14MRiynCfgLcuFrd++
WDtZdbynkrFUMznyiYcGRg+xqB40zzlNmVsGfZzmDiO1K9+rV9Lxu5pFS/lz7MGB9KKwqxhDK17J
gYZWiuqUCfiujMXOmjCYU9vpuDjRdeNSkES3pkhVDx5dyNv+JIr9BhycLMUTiFIM/RyB/VIUyLpv
wME8jWaUoyD0rzIYhXNxfvs4SgKuwB+F96N4Gq06VhJSEjRrdoNUG3tLd8Ec67KTxfUW0lJh71dl
9BGC7VsbwbtGmmiBSLJhV+yabcAawZGc/YEAC0X3jU5eoA19rpEKjVYdsK2e3YxTDRfyoCd9HzUu
AjtPxMHzCs4/RZgRTjSoCCVCnLD3yb2TBOy00dI05HyocHoC3Z+VRdwOUik62QX2l/ooITDphQFN
ju4e71oYXDVMeiHQzA53kXt8bljp+JPQY2+qChvKZ7VO19ZYt+upQ6O0++VXD+GVjcEcU7DiOkw9
JnkpAFCv7R2cB4JOWgjxul4PUIC5W5kpR+57INig0nQv4SRqw9O2epGJWz+ZhQkcNp5juAuKGgrT
gXCOzY9dHEMu/6tj13mz+zZQpq1XxPKJ6VFHwQ7tz4YfnzHSdN0b1nmZVSyxzC+fMpSw50QVzoSf
/AdAXstXBKoGDW3CUemaiQMWRl+skAf0S9ipagSQliK7MrZteawJGfdp+hIAvpq8prh5LO8UAlGe
tmuHs9T9F/F6ZRfFxfVZE7bu6+YweWC/OF/yChYPFmaEfjDEJcCx7xzRh1wSpQj8eN4agRJi6Vt5
OEaES4QRsBhtlSeuEpgykbi3D8LQ6r5dX8MNgkKMUm2Ol0MIAEddFyuWpO2nMXVlE2FzJ1eR8Inf
0dKvZWUc8xk9b+PZK4Ls2cuPeHZkFRO3liSIe+cty6p/q4ZJezsgHLiEb2KEnuB2LNzetAUNCzyg
aPYznVYEzsjO2EsMyCitIKlJhajyKbUE1syHnJbDMYt0fI0iUeUH4tVTf5AcszErVzJQAH/c58q4
TvxvPiwsc8YK3VI5YvMNri4kjtCzixEIEnIWuI2ouyAEKKpRf8VBdcp181+po3l7bf2PnW5uhWDc
s5mk6AQuXA55NMoC2PmlLwX2ZaCL9fOwyD9bz1V1V7WKUsbY2UpWKhOWK8WMGfI67F4utvQGG3hy
ELPUY6aQ0wP6P5SPZi8W/MDOjNlGcqS63Y4gX9Jojo3qmFHgD+mMFwrN1edIcLMuCYhKjcm4TGLx
nT2vZSz7N2SOAVZYBSDziDNhXFkgsYNo0PyeTz7oNTQPAfB9VzlcR+80hFtZJ9WRYGcfi0LvNAho
JexN/N/8HBuNHsmXPa2UDQhWxR5xDv3DRHzBCFEeS7E+D8xMk6ftjuMQAAqKFOP5W4GHxZFmIpzc
IwEenv46IK/x0Mja4ZX91fGZ/JDZY2HY/4N+D1ygzit06uINhevg8KMdTlp2I03hB+6aMNDxjUJs
c/tQpVNFtUz/MZqqOWrrlgWlF26t9JOwtvWuzT8Ym9nnd4EmCOVVFjTHrMiqT8h4SfeAj1WARb5/
XOKm81GDt04yIkia+nLgpI+3pEW8DGubg9PfudkLa1qFDK6PGG4y/Vi1/DLQqNAZSKTswa/qPa8j
bhU4kvRpx9+o/CwQzpMya4YdFwMj10d3NXCT0JGQEJ5vyusEdeZOhuvlGHyQVMGqZWJW87RiuYvF
5pU7oqhvqNUYAeInfMvdisflzQ3TKxM92G2f6NCJtGshsGmWhvr7ayd8cHaPz30XRrTubcfTZuBC
7X4Wx86nDodm4L7q4zGyhh0ijI/uFklt3ynk/jyv8s9VoEBfEuKOZ0zKH+VCIMxI3/zCb8cRiQV4
CUHLD1qi9W5Oh7vEIehsvxSzdsVF/+mm66IoQ0cm998LNNgXta74U1UwuOY3uKaA69TKOk6Pk9Pp
IamAV+z+PpSAgTzep38V8DrPWKZgEHVRxeWtfB8aPhlg5rAU0eXPnOsPs6JhP6mxDE7x80mmbZlA
WV8JD/Gz/rqPqYqdaZ0HeHU9FR1yZsCH5+af+tpF+eRxoHxtn2Que6nkiEcL9VgCJiQ3rsSAOhOi
AlGPzFYwurL+7aK7kjOUGTuCYjlRI31iBs2Z+SLtKBt05kRvsan6xeC6P+v5h+5zcNxMJ4Aa3G3J
9Sk3+sUwkfW9E0C2XUS+EP8v3fNr5j/TA/Ujrijv5/YdxsnDxtpLk7sBBVW0wqOlGPJ8z9IPcizn
QHcdGokY69KS4g0sCwQLDGJhEuU3Ix+7u5e8LaYQhZi0S37NJCLsss+N1uTSuRjzyMwWLNJ9TDPy
MGxpPmM18SXw6gcjjWTzap75s4JocbNMQTsUTeGs9+ba9oeawJSjSucYOnPPWgZB48VDoARLb7cT
jAECr0JdATpwspd9qQVMO3NNkd2A3t8DozbgKKL7F59xofpssGlDmQXxj91Dw7tiaID3djXeH0ho
9x7+rWDIes84UU+lpdX4gZu/P+apL7SxH1ZdxangSikjCCEnUo9/2gsCaOqS2J/AF4y1e0IL4biV
NJvXd6e0ChF+Jsv86J1+S/8Ztk6mNRvsli4jjcuO2SPV8mYnTRadzOWceVpkIEO9omY5mSkRNFzC
kVetRRCow8FmvN/O1DO7W+Ri6QQWAJh28KBCDeTxCj+9wgJO8XxDQFaTYEhOx/RZfp7VHAGqHepG
7A5fAqCRIcwSTIkfpRHp3OFv8eOBtFfypwBZmJs+bmA1jePpAjZS8EiQAt6Jpczp9fpUZkme4VRp
8jBxFamZlITc11TDJA+hn147mzCDVR0ePt6y0wUg7VvD3FO8mqplBbupJJPftZVCmhoL3F1qWg66
Kn5uvkTlIpTqJcqkUw9wo5Q342YfwypApuOFpUKyJiPj0UUasOpX+zFHuW6258oJs+/U5/0tMuSI
OOIFL2+j9WbRlmtNkMZY3HutasqKcemSBpvDKlrD47yKwBlxENpcrK7HmaydAVjZzJKE74pvXZwt
9p8LAPqH2z6E4HWaouhMF0oUcfP/Eq86rsdWAu9EK3O1Mabk7KMVYVmoQIl7VAgZ/Q01oNVmtHE9
Q+wFN4c0OjowO6aQ7icZPwd/ST46DCRBEsjv5cczDM/kfAooF9LxAULqQ76kF474rTZ7mjSTwvIS
SCFcGFQbyIDrKYq46jxbRx8zWwJyTvyia8zhwNpraeH5GwuAj3/QjORHvxRDg6OZyTcVijKrDi6V
Rgxt/9DwLa2VwO9BakqqRaJg98otLIH+FJdQueWqxkETTBnszvWrEHdV1vvbabeHHGIiOcllDnvx
SX2WISZL7laW3LPh7I+E0t6GJZ6w3T5x3gC/P7FimAV166mpTF/ncPRZ2n0Nueom+mfVm2TsE4JK
1Jhz1FKxBueuN9EeSNNoBxI6QA8rITTbbdRT7EP4I16nsur9u3IPMWGb/Q3nan8GEWVZ1lDoY+cX
KWCgh9/rTaG7mJR7PbVqpBsjPf+AtzCPRW+HnLxKtSPTQLYdqmviMY7hPOiNTrLlQBQxO3fBul9Q
/BQYosF9bCAKEkmzBaBoIma7j+NAfErQFRDmsktMaDIvjnDjDJaNn4pSLF912j1gPulVIbI69L3w
dZblVuyAblx88jLLODg+ROuIes2JbsbydNUsXrnJ17oHl5BNLGFPL4xUyqkO/sojCBKQHdtmlRPy
aPtAfj4e3h6m4fiaU/sHFThhs+58HFEsScr5R2Wm3iv4Dworg0gtphpF4NTec7YKLg/9jxEofdId
6aXvHUOI4v46mqn+pSApm13wZl0RkyAGkIf+8LqrNvjqqpIwjSRpvH6RQdDN8ZaRh+gFnj7iZPx2
hrL+RSyu807FoqBQ6vim5guEbswAK0QOf8UHjOh9Ji9ab0c3rzjxkOJT8UHTENyEvjZEfJsaf6DR
0B5agNK0oUWM5caRbjlK05Q/a6OdP6KuIDIC29krvD9+a+sRUyVtBxqksAFZVxSuNDX7MIlIDyl4
b7DSx9eucLgVfvg3G0kGReiaApy1EXlffa123vWeJ95zlLUbd0K35cXlKn26t2u3Dh8BYatSkObz
i628OniBPolwaO4AdICXnGeAoDQGDxPFS2qS6iW1ERrjUICj+KUrSKFPJKX81TYAmRM3yhYcdPS1
TV1/U0TdFfZlIYOk54vGemqCsnpB8mH/1bl/obrujpLpuJVRxauev6mDEBUZmtZk7aatnFu191xa
z2Cw1+a8UGgrWX4E6rsZ+EyzuoJOsCXzca+GD1mgKu2iif6hE1TVcbrfNp2I8KgbDO7bjB6pex04
DfaIy10AlVqWd0DK2PnybIh+hD/pHRvU/mHIHIc4USRKnoq+33ANVY/xPyB3m9fINMd4AggrJ71M
2DYbBvT25M1nYsWXh4LTPPX8u/nVYa0zsWlHJK3QusoVnC3qEszvMpsrKl8cBDz20OF9GpwHnfD4
B8Oe1DOGsBKTUH4FGvbZGe2DpfoVv03k3UcE/WRF6gExMrI7fBCh6RVBuGNYhyBOg1nAUFQKvbOs
3Jy5zsI3yvVmmiBclYVA8y4HT0bYzviz8V0zoYHeqywqzjZXOYamw/5WO9UwdD3BnyWIoYYoJYqQ
sRceIFfBLn8Dz0WC8r5HKKsi2DrVDkWsmVOu3/IRqTumMsMftDeZ4SJ60glH2eapz3MMm3YUvZFX
ssQdwKE2oN+HWLnx+RKwkrMd5ukh8xmTNf4XWpxcID0s84KZpUS5R5pRxmxdgcUS7ACNenL09eXo
OTw5ndaRrw9cMj3aHZZh7+csVZEFYoC8scofzow8rl6erEtq1+qJWJal21W4TIeGCe6uQEcYZMJp
zTxK9gei7lTTCVObOZQt7eZJLFhSNidLaDYVZpXdemknyTiSypmqy8vUb3qbZz1oeTLo2vHftaeL
mBDCbrErlDcgyqTYa8nMPnH5BxylgQxyQsZfFZkwJb8kIJX7682YRwknlhkfrEQ0lpVDHL054aMj
tmg1b2VWc7mfjfG7HswK5PvvUZFPeJn9D4aVBRGFQBXyqroZPHGeLb6wuL1pG4dehEafuvc2cUSF
V2MqnHmCtno6oBI5H0/iibJA+VYrnC4iCJAcM0iAt/Xui83GROnw+fFIuT7AwymdLFeipIbeeb5w
geMJnjtfGsP+rrX+IgxbftWsddsFqYt+VMnipoGayUZYVzRj/3ea2hVYlbLkW87k0rbTFXylVc/U
0z1J9vMhIwfzcOlYqfvi784Bv1TZUc3HjmbD6vUpaqy8n0OO3/ruEUC7utODMb8uFey40yHN/LtI
RBHHU5orK4nAzco4+X53kfaCoo4U9RGJzj6FBmk7dRBOt8Pjzs9kEtPMlIR5cmhEq7JhXl8LpXWX
yiag32g/Az1SmmswulJfS7jx0HLzdtMoAsKnJAvmB+QDDUHNnrY+BTCjm3Tp9cZ8bgBHb//9f+u9
97FvPDph2ai1oeHWtaH953r95VgfTX+jnSZOdclmb8kBdJnBpy0XPiq9+HaBurDXf5v6qcf2ahNd
sAY/jMv/6oVbQwBLT+FT0/2IAF2MoAf/VIOCgszUjK9IpAJcEWzcQm2/cxwT8oXUXiQbCgc/vkj2
u2ACTvFTpu0cyLa3WPww5dsb5kjshKPX65Th3p9AWapBTGVR4PIhsyjclcXSbYm4hWVsXKEHfhaW
Tqgv9nqt9Unre/lz20Wm0t4EbGxiUZUx68JG9F3PXo0elk8J1IAJwPCur2GKUFRi7JBEkkuoUpbr
AWQCKk+qvQVdBaUkUE3VGXfUrTyK0iNJ1dTeT1SLn6jUGiCcc05KCtm2QZau9xzBTQpQ0t1IPkoM
2FH26uoCNShv1a6YO9UV4bPXhJToZvc7dHIcY8YiHbQmXsLLVDk3di2ieieeETMeLpmWU8Y175K6
M2yWvwdwjuOPXRcp5RJChJxIGpVbouWaqSOXya3xKGPsAX4U9Hw2+eWAzWoPDIkZAXpTc5nIP/Bl
HBgSYnwFhF2M6PM2BlnW1hB33mAEuyXNiCDqkD5Ko2xzQAxJ2jpxB3CIs1tl0EyepilNiY1U+6tu
QKiX0XJMjIYrij/tl0siWrehDBNjzRXOXorVCXtFGU1RTIX+PrU/Mi4FXdvHT3htD7Yrs2W9BeWL
Jn36x8WoSm+EVJcOZO00PsRxY71j3Y5djw2eQ34Cwtmryd2OecTObit+iITuKu1NzxCkfxe4GJhX
TW2UYGjPOETIZa0/jKEnyg8N0nTOJCce12+VM0ra8QEgwjZclE3JaNnU5Hk33Kh50O/C9RjWYavX
bnMUiD688W7909L/XOET0W+WhsRa6pynt2csPv1lz5pOdkq3No9zez6kWKBNNtIMxW+OryFb/bn0
qF1MMZefuBU4bP8AVvVXnXH4sJIMVJWnP9KOiTJ7G1A6d5AnlDURsWnd13hqhPX4hLJGkdEOSv/l
bAt5UHJC2SHXeIiAOSUlPuxu4+dOoSffQqKmUnCbE7zytvo/xeiQCdaY7/CSJgDmbBeYMhhvrBkt
fO2r5DAJnmkXHrq9H+iKdj/seHN5lmxYHItSOeKJVCnPrDcRJtXNmegckVk9ne9gZJNj+Z8aqZqe
96yb5XdtiM/zaR+sqVDQvCGSoYvvnhWpqT0EiRAxATClzZgzPHrkV+Q8uznVOiDLi4DGZCZaWCuz
fQGAz6/J3dAzgEgf02lJlR7ZLfz4j5oZz89VR1VFrUuM4U2snJgQAD9mCWvAibM+yhTAaF+FDRaI
KB/iw62p3OfFIUNpTiQH9MJVFYc1+h6wM1BEz5Tn93kMxjI40oQEPujnRoHlK8ZAW/fi6iuxrRy+
f58BTVLM8Q/4VgM/lN3IDGugVXl6Lt7OL2cJS4auRffepvKEJpfypfbgTZdLxlreS8ngVQxrmwtx
JwFJ8+24frPiYwj25s3J/lNXNy4nZlyKfPZflw0kRrfMt91RgALj7TVnNAtVSQugl5Hy8Zz4l+hE
qTxeF1dIup0Q/sLsf5BecRG+NIth15svNE5gaR0VlAqMz8WhNOfoMBoKeIjmb5eiD8ciHbs2HaT7
XIs4kcqyRSfqTzGgTsHI1Ll6K6H1fOI3DoUGaFagKHUQrgBridIDi73Xgv169fv5Yg9GRVJpdpJL
sYWASg9150jHS/yyvzhZBJmW/SY3NWlxBADKczexD9RSLoQya9wtb/qk7slkdUoppIJnoxbhblbq
UzBRksSvnZVN2y6LwCSHUOTSmuJgHTNYRH7ZRdnqP+OsSJD6R8BYzsbbQmxUi3a6yEq9r0W4hB5b
gJkkuP6YpGuB/g6spxYiyg+xKJuebLHC5IyiR3ZGMafpjq+/uwRaKoRRZm5pIjSQA6Ip5aP09Bs8
y5nZOATA/SAxR8FfdoHxhN7QNR0nfa3fM52+7bpJ0gRSpTbvhTsXUhUjqAWdF8WAuGpmOAuq7CHh
R38G0S+DheIyNQFxKhuxSZdKKY66XBrhlolIwRU1wK2dQOJMpkvl0Xr4GXMxDC2wjrXPzfgwFAcZ
bBu71qRDTRgVp9j6pnTMfWoXChKPoHHNSMvW1lUDuKI4vk45NtzHFum77XAe/oOEexwwVbsXZxBy
sMZ6nLuD+tEiXpwNHkT4J/dXd/PPrCd1FPrmGJTX/5aU+20WfnQGeXpApA1pUXfUSFgkmd43ocIp
cUAY823B6yHn3/FVxV6jeFx7UqAO+TqEOBfOwYwQzdzcxPsGBL0rhDdRzG854Jbxse9KaxGO0uJP
qb1CE6YIeiJqvgNDrFPwZpz4f8vMjXuhEMyFAP0v/QrJHlVS9oDs2BXmI/SBjf9SnahlMP2ZPqHj
gjuhQwF8bVkXkglIBQQN/ZtlHx2m1t7oJi6DqNAEwCj6xNj+uAO8MAIgCsu+Fdb5WduazszeM/Kg
vTGvjhmjZuEZ+ADywNHTHAdA0yEelqps1OANn8nM13g02+Ul4PSr8sD/2/EvXfi5QQUZtZj7hGKO
8qpjDvBAg9KK/Gx5AlYu91EQZQMIU1cmjp7g+OJHuVOazPFPU/io+8fyNRlUsD9KLZ1TSSI33pOG
ZSrKlQCwveNsfGtzDBcJlWVQmIOAljDyymK2jyPdiszfBZkK2USi25EbtFL8FYfLAt1P4XdSwBpn
y20DGXR3pGjcT4bEbv4nc9ziGXzrMvaed+Ea6AwAtT+Kkm9ER0g1s/LTQ9I9UO1TtpWfpZbGRevX
32eVvf10gSvD9VpDI4xMER2jR1SQZWsOqt+HT+n5eQl7wCxIy5gEQv+F3Irfl/0yitsvSleRoxWu
j8rK2FbfDfjwi7xx/Gz5O7BU1w1NCFeBs9UF7qLTEyArpU2p0uc3M71WHk/2hLzEGosMXLiTIgWf
HcGKizgUWN9EYJQnw6YRylAG0GnarvAwjwTAkkGh/ddZEGKDbBZWHtXJGBeXGeH+3Or7Wl2o9beb
AKHQTUJGL6vQwyPBPuO4tCxjkrezz+uEPg0GPmoWtnV9pDI5Pu6X4b1xaK0Z9gPdqpfd6JixZPjE
W/99Q96ZJIaMMJnb4D/C8g3ICUi4fRdjv3ApwSAV5vW8Pw6JpTtmDI+Uh21vBLKfxRUcfw9YfbUY
zRHNN90j0vwem+k7aTJMAnNkGimn/x6i/2/LTPm2IwPoU6e3FY+6BqJk6oHYjSt1nmbXSzMEB4i6
wct9RGabHfNU5fOi3JEvdxtDQ3agPpo5AnUTA6V1wSdJsy79FOIaVdKijH38LbgJyVNqHNCCn56k
/zT9MfdMUZkjuw9rcZ/gQW5FRdRkATeljkltSftYT2+H/CtF8Wm201RJby3U6+dwsfw5oxW7gnY0
ieoRdna98MGXBkyYEYlSFt3jTtN0k7jHKvoEDRg9FIflueFwbZELLM09OuHPnA539W+Pb+9FWxLI
CFeUc9VKzV9gmmW3yeHd8ISPEMdpoBJmVilsfGTAypI3BzSFxGZAeNWXSgCENdZ3jw485F0SBWAT
nXCKOG1R8f/Edaza9wz1R2Bxy1UDcmHAoiwui9IHinTnvVGn61kspOfSfqmTl+5sHjyXJXpfe/0T
/V2bqUlxsHsJBo6i+n1kq+YIHrOV1eJVopKqoWaylCHzWTKtJs2mTLijN9hTY4TG2hZ7NX8Ol/CS
SfMfbN6muhPbiYKud/WXRUTqp5ZgVm4qwOcDml0DYsmgS6LqB7uXhlygYy5HfX7p2MhiZHc2ATfZ
r/B+y7QixYZIiREXOR+5ZcRAXUWNvsXM9bWMqAliMxoQ2nGZLHi/YQ49HYKtgVTHajUWjYtWrO9T
ptvGj4JHzZYonu4RK9ZFuK0NIsCt4w3McOrRIWSWfthVq0wEnLBGtjWkTQyJOtNJRUfvwSciLGmK
bvq2W8mdyy1ovul9JZpIM8mjZ0y8yoc9QmBNtkaFzRQtsU1wI/TiWQlt2rZ2nr7U/g8ZKmdYyIU9
yufuf5fn53v931xD1m0xFrgqojEjOrh2XnjvjF4Xqesp1Crwa4oIjwcD9AIu12IKM3y2J9SdBGcy
rhPlWLExMZ+f7XC9Dg75ktGjxQnAKr9kv4KGXKroOckvhLLQUSKv+o/UJgVT6pF9oicV/3uCwjWV
Xvr8wXWwjmvZpdLSGhtwORIdEJzNLTITM0CjehZ4A69crA7h4Iga1Ldjm9rbBoGzELrA36J2EhGx
239CsJXznP/+/1jtoP9JT2L2n1kfpPd9S7oXkWA1sBThI29HqSMgdAdUGbRk9r08VJ3NUhYcw7OR
WcxXq3OXeTJuhjSdoAz2NeOBnqPKWxuGN0dN4wFUQGoODez39GnQm92c6lcrMgRI6s+sx0cCofI+
bCem4NLLN9B1zlqbn1Xc8RQ+euZdOuIWiIoPhLdtyP8BPr2qbANNLSYJDDU2BciMQAGFcPSUiIwS
MxxqTjqFm2HGJoLf0srm6c/hKEEBH4SQJqEkCyq42h+jn8cM76aLtDMlOLUEW91JVEF4t/OMktMm
JAZj+DpD7svlxL28uXkWBGbS77gDH1XV95McG+qMVtQ0VLEfnAKlnxzOfyU7iZczZzrMJW+cRKWY
uFOhsqzt3zdj8bs8tlyQouDMZTi92eQQhQ2jnD/1BIkleNEyYRCuL9Jcd8H+3V/Upfg3r27DLWLZ
JRZt43PKMv4MOWXIOPNC3L8vZcoYlD8PPdBqnBziE/+Q6Bg6QoRzGlaU/OSM6OWMKKiW06bq7gLT
lrUKjpuq3n19mGW8Vd4mgybR07KstHZ3h7EKSkXeHYlKu4Y8nnjrs7rnG/cCgKdizU7YNM/WjeQX
xaK6ZCOTJfgoEgnCrKngDe+odgQFQbOJl2rRXFCmey+0j9K9VkCb3cWLAOc73OW+3KPUXadsKiOp
8lmmsjDEEJahTlFuf1h2vnNu/GxilGnMCUI+RBwOie5zTcXzg03djWJ7BtG+Imv1mlEMnCEAOj+5
B8fH46rizOeOwCu/yFR4D/bYHnbnHsHaQ/b5MS66ssCh8oGmcHa8QD6CkezDco4RYB3hP+QNlPHi
/35qsUinWJkmlRgV7E6KKpOgikytH7F1q6TERekL1zAPL31R0W5sF/Hdv27//3flARSDRv4+0QfW
M/jIGqj1lHmcKhUaSyIu/gjiuETTzczgraCTMPf/ve4Rn+rrRx7L7U333a7UsSs9A3cvoRxUy8WK
m2wsUSuDDpm+avycUV9GraKBKjLVKYL/Ct2pEZpA7Ea2XijU4CGUZ1Kjn9spbLSsWCHhMirComnh
hTU+yuqslIOqf3YW1Qmu0QK+C1VJuri6pr+kVWUY9FoM439w5DrGsv7/phFVmIv7oR61LtEj2QO7
lRuAlaRVQ+3pG9z1qSFd/BMzZjp+X96TpTGOph9RVQ3S60eoVno8JOblGunb0ruf1wK3/pVRY8b1
igawpkCXgUgxDXRdDdIuPxT1RD2gra2kjUo/2lN5gsiCeXebUwa71g7SS062rVpCOI64Oy1Plj/w
3k0SXCkkxXUNcXXWoreSXd8AATiRhQ5sD3UlSoV6ITUBLX361V57xaFMxB5Pl88g8E7gr5BxaxMd
PykcVzeeVTdIkhqz7QySW1NrMdeBOTRQTyk3rE6HY95G22Ihjtsgy0nP5dLp+Mm00t6/dwWLT2MU
TjXGamxbFaxLuhACbdG+le6ktNcGMJ/kAUwGJL54GK6YHbrjBOSXyGUTZPSL4N6OsVJf3bUw7p/p
alt1VBXEGu970LgyvqsnqvHI2Ftd85eSq4rfScO7nykdz5EJ7FJvz2pob8GxuAJt7M7XZ8/NvUYG
7RYv73R/WwsKdCLHtuIi26NytViROTKrfq2fDxL9qtKQwpR61MOHDakE1kbJrLBrF/jzkveb9MM1
P0pWTxh2HYBkrYenmnOufje7uEF0sofCzwW/arv/riV6lSscp0QBaGMuiSUr87sIQp8w0Kc/SlpQ
EuDMM5O6IqeXePr9z/5xUTVzBMm+LImFve5I4MYL3X4heiINWwIVsh+5reacOSh8acElbEOumOyu
/3WDdN7/adzcPJl0LnRcPfMopajKpCJ6i1sauz7FtmMUCw9UVp3vomW/uq8CN8kno63nhRrbBbyG
LIWU8fz90gCjhp0Clud2jA0h/UaGuG6eIik20/xyr0MHJZQL2bR39rzuIR6IY1Fdtb+nH5n/4WW/
Ok8DZNmm5J5vyxAlpe+A8IHPDEruhdo56SXHrqb4J4lN8ERl2tz51ex/WHEeZAn/h6SdrdCXghd0
LvL3IXGk7Wd+x0JUhMjk+A9i9HVukQyd58tmpVU6QJcU022s0q2StfpoL/qTUUu1fwEuBQjTLokm
sitje0ky6D0w76hxHGcs/FEzTiC2qml+1bSDUT1eBS6MTwZ2QMmH90p6kUzg4Ys9x1vc5HvmSmMl
TXVnPaLYMeUjdNFYM/oOKFaljcFuWzVlrupW29yRziY3tWeKTqNDUF1Qd/V3QAmhZWN8kZAFje0y
noZBW6rZZmatT0tBmnLPD7ZjsSmkRKHxXX7QRJ1alN1BwCzvNsTNx2zwavm/HZwYAvfvHLiICCls
Leg7ghUpWcJtKws1BdVGenXknnKPWfIAHX0KhPhP6Idv7QK2dDGOUyJUxbj7Fy6RITiIrpdB9hHw
PaaRXjYkyrhlmyt3yuZHoreFqnsDMQfMsxbUPRxLS6uJWuWY00PHKaNR+SYJts8e+b/0XjKvLFnc
WyRCI5Zz2HgE0ix4oZrTil6kjD+gxqWKKrTyRt0R6LeEGByzqlE35jcBAwH7ZIsKGaENK/HxAdOY
GB4ogJEsN5au4bZwlB4j8HYW3wlu+LpCnsEw8sfH7PKe48Bshv/Ts+YzWQGITdlMV4uojIxxSw/F
YDQ3DwDzZxlNpACwUZjAN2nS0zUaayv7bIWYuOGbtM+CYdxL2tX46DSxHxhGdB8I/Nqq5i5ogrEv
AOvUO7WOZBrFTNQ32TUZuklM7g8Q7bSYetx7KkiP4xbTU+bvkckuGQr389ILTZN+77e6tDxe6Fjj
0U2U2jWgMc4uIcZC9K8wVpjf3KUd03msbIyuGUOejRajlu5odzBlGzszs5fhYHvoL/9W4VWg6RKa
S+TDpXu9F5JZNwP9/74OSZdDJDMiBlPZ/DEId05qKZHFx+T+EErxnfDHIqbfi6GnR/EaBMwlJRTK
VyBgVIoum1OfCU/Mjvas6s2vuMtvcPvV1nW/CFDrVf2Tjw10vT2EPXSwk/Cbs1e8cYRqTfA/jaFf
7ODMo7wvW7Jj82fBZ+dUN0zwu4Lqi9n4tlbJU3omulSg5Uwzd5rp4jLos9MNCrbRwDHFtgS8g1Yb
HUHAUBRFv13p4Je0Y/2pApOqI59ybfHnNWfvEsmrnjrKkmMvdcaP/cAAMUp7Y4Lbc4rSF5Nymaz5
7KchIqDa1OkGEPBo6Ilug5/4SbY2P9L+7mrkfN5Uj2BJmXgMqOPlpAxC24zSOqbqqP15C6ZqOYwF
21ExmfmT7ctEXgGDOP6NXLscfKXBVYJ3NsjhK1ngqjvdQH2wa0B7VlIpJD1xrOtYC6PGtxL4IusR
UBGmfY2WhY6r5IVjlIWZl80HpyqiHjFCxvvAb7gkMb+TA4ZpCQQP4gQ/NBLfoUn4aX1248jPx0/x
niypbNzsr4t6tPl0StPlj2jFNZzA84k2P+jlWkOtUEuCV8bun+43/kByKXvGMd0F2BFNn0QojzYH
W6DH/Cw8ZfFg7oIQzW3oiZ2n47NO+n4R+VcP+H89Eokdn4aacvG6I28CVhd2N2QXrbK+Hcl9y4C2
KOwtmWeQgc9pSOsCCxTs4B7Hvl+amcTUM8htBwLw+L3pu2z7aXwo6GtPgXOWY/vgbRzMyrDbAFRE
rsK9xcQtf6OIZaZWRmYlk1rtmq0QLcehGWB97MSq2+wNVPEBVuyauUCcWC6qAhn/iMlAW58jyGjt
Cd45d0xS8BlPo0dKH5wLUe6wIQqTjinP4V+GfwTWFZDSO8MMazD5vvHgLapMf1FPGGqMJ0Qni7VU
aAtUels8KSDb9iaFyyWanmSkeHMbLZe8Nem67D3XYrrxV65WVPV7fA+8Fwg9Pmf0M9RG136HxEsY
hP0SIopekzGWxxZ/WZ0zoIhgBSve1E7OcRni8LQyYEhEBB5Ya7qGXpw+iKiZjArwgk9Cg6fXVEqk
rDJlRa+Rzz3hyjYSFhcvbFkBr2fRqMI0s9w32Ca3dxv7/Z7IRNqFDHPL6C6QD2zPguSZNrDXPjWh
OVZWLgLea3JrvFGDntus3ZdHx7aKwV8xPh9wkcpSKqS9JIOTMp24Fccza8vNHwKzEVabs1hyTL8Z
uGospHaN0EMkoma5KomOZiy3pd9TOwZruxeAlveiODM0qWbWkHadO13zHt7BIU502hCoedKErpQr
jwppMFz6CnkeIhTwu/srZIdWDpBVOXSC1m5mXx13EKYwSp7/Y/c7mS6lGzqyzIg0mDWmWeRWzgWM
5i13R/I4S8adKWT840h3HtQeR7PJmXnxAntP+MkRAywZ5ai0IzcDBl50+xsTyrFCH+lCLUFkHPb5
toJmhBBQ+Zd36qUnUUQghtraHI7AT3e1mVkzYgsGj11/X5sPNglCNduFTRI02lNbSExn3xvmoZqW
3aeDXAGHiUsSc4Z7K6lxTFKMAhM8HzrkubZuGFXQ5c5OyRV79lRNNlQcaKaJqiXrEmbsUc8x3dOn
b03F1/J7bJB5sAH45+L40JnTKOroekqB0iZxaXUbxO5Ql+oedIlX3r+dZbJMoLoElHotUEXxcoUW
xrgUC6HGpOU1A9QliSOkrBF3xGPcKIoIWhC0dVmPhmhRCHfZ3TK+lUFwQZ1knpUYTMNdvHl1YRB8
FvQfRj+GUxqzjplyzV8zqQf+r2ceEwiTFoGUVXhCK7lKYA00F+7LDFD1Lft0QbAq42JMR6QLdrPR
3Hl7xObo0ofoUfKIL2Ec3mGSN6792jsy6gJapsnTOaY7ZoOWe02Fk6F5plx8KGs9fNhze9mv3+F8
GIwEZ7Wk1SX7uHQERy/HiDtrqy00TNAPH+LcXUeEEROANLr+sLRai6zXhwl3pHGetZx4QhAChc7K
xayl7HKsVVQ12vSco7IYqXkhFR7vWEmHfdokvWcDHggfIbWFKOG+n59Xpje9dq8PO+CXPPKtrQpG
3ZHUnF1NHgKMSl1BIKCV4RBinKwQAKpfoDuKSVgrx3ET7kXCY2ACBTprK0sISm3BoBzeJX+K0Jq+
dMcTGEBXIpriL2KyEgrUcAUYQXWgqtaZ4SQ0Nf5ad/uEWvvzw9/eZ+zjL+d2pldJMqmHjFQSp8Ji
SdGvrr85zcdrFV3yCmNEgHGBsFV/MRKL7GD+U45ulFj7ffr0v0htY9EF4qY8LKfLS49E3beQvRc6
ZhZkt1rkmq5HuF/4M0Xz0VWUnPr2UBCfQ43L16uritA2XeVhYt5L8qf4McYl68e5YPQr7sVoY8/s
G19EinoQ0+uJO1P2v4cqPkQtQ0g5VfGPXgDMrJYzii/iMtQZY1M8IIU1LLn+bNPFv/hLx/ePwZfr
THqYB0Sk3z8ixKh9WY7PK84oEXsOIQWVzy5qKoC1nvz/13LIaqlyZlkStL3PcVhJc3Ye8xvj+sI7
QHYA8E0QUKgtJ/RuxxiS41e+oML//TbghckFBUxdzJDIspytrn71c//rubY61wz7u9iUYE0zUXEh
NX0bPh6+rXDOjbKW3HQtkmyCbIQpYWaYjJM5BEXktVAgsSOctp4Q7l9exc4peKig4L6qqaVG2rPi
h/3Oc3uTK8MckuYag18nRGiu2pxsLSCgzOfD+iigO2L6fTXrS0NqNlPN6fNlTv0Rk72ZzhswlLLX
KGZIXL4rRd56NJ9m+EKfX8B4/zF3UkaBVfvuU2l4xZhkyjeFkT/Na5ET2c8l0I1oNkgLFtfvoSB+
nxvLIhkX9kHSlAX18a7sBE9Dx4p3CW7zTgdrXpsmlY7B8YqMuKaPzUjPZW5pWBAhfgDC7NSzTW/7
95q3trkz8oUcX+KkqWfRrVnPQd2ySiW0a+dUSTSB58fEJNTBFvDkNyVOyqUIBbgdltahC/Nqkynd
w7NfT8vsW6a0+cGZU9R487OjeScWO4QBKvVQGDJQP+VZ90qyglDRyA7ZlZc6h0D3AnAgwzKMesM2
AZP4PmGAlE7gY7seyeVWBU77zN0f5ueExdEADq0PxN5SbcoAsNcOlfy3n+ucfj7xKHAt1VezJ+ou
zwq87pnbjnQU8eNcIxAqZWWMqomS8sbXYTgymM6q2aJ3GWZ+AZIQ9jBmnfblfFLfnNB732SWTlKW
DEVGvu9AZKEew2RoP+I68xF8/ypSFKdAXCnLyrC5kLLh/gIHm4qsLVfgw/z9CvvIMlMRvIYzPMYR
zOYHTsJ/7Ix8LdUu/s49DUjXKILc4fhVLd2wsyTnD2eRVX5+sqv0v4bCUUMlVSA8CS45Zz4xSNOc
JOl02r7+V78HRQqQE9L37W0tcQl8J7f4p9QgBEbvC4WtstjR1qqPyNSy4BB/u79OZWAF7CkbvW2a
DVaOCzeje9ykxy/c7WDSxsl8UtLmOAAurBvs5u804kaILDMr8R8I0/cTQOQlnrWRqudlDFuyfyWg
unHq6CXPh0NHDnidQ63R0t60+mbnClTCHfbl/To7E2GG758LhGj3sjx7hknGvTSXJk2IqUq4B+6U
gR3I2t6k6xnEL+dAAqKXCl845HTdEcLfCrL+5uUHZ5v9dnA/jqKGFctMEhtCAFtzUSvgi+Z9Xk2n
5u6+/F+h/MhkHk1qvj1zigtHV+xvxSszKH53XXNjbWBG57HFp5fVTj3xS9UaiqJ5ErIBhflPpqb6
Czoj0WOzfzd6bjTpBWUWHw69KFbowkNlQThiSVqS3MOeE2RVfEqMvG8K21rfMYoDomHe0nQpA2QO
vuuZ7XKG6cUqukFuUcAL5hX/uNoBP/4lhBjvuqymT2wiexa9Ueu9fyQyEOf/1bRD85FNnj/rN0ed
YbzQNCTRq/7NiTpGmLpov4DHj6gPKIHcOppL1e+6QHRuGjHVxzxfkdAlgXTZx+l6EaODKCY6tzpk
7HH3TVngk3hAArPcYbqqTi95ZZADr9E6SAj5wqOO4vwX+05qa3oWNsa3MmjcBkBycQ/i7odNqYOv
ZE3yiUGjm/oO1YSoUHsVjGStSgD2cZXphxJoZrG/YGybKnJL/habKBQWG8mtZDWJBapP6A7WE44I
4SvXVIEHJXATEBezB20Q3NCNUH7YU88jjYBDEBVwy8y6FKQO/817tiddp43O3PqwbhumPPgQunAR
aBnaoQiJebePzEgTZZnP4TbTwjQ7a8OoV3kjP6iWfz7X4gNizguaFxP+sNIePtLsp36VD0LDzKIg
alIVMu/O4Y0D6nV4a0qqrg90t3gIKDDjdmknYZxKd4H0Iq0FgiHzrokfyXxotzn5VQ1vYsiCnmnV
XMWpvuiISVjn7gAYP/KtsJdooV9954HTOH11wRidRPQxgqWy2+msCg686eSlWFWlIjUusiB/ygkT
Wd0pjgNr5kwTMRt+kgezzFescKpQ8MFXOW+9ywMQVJA/I3I8swFiHnNZKyYo2COVy0YKce65M5iu
V59FAexCgtiKP5bGyBxnXHQSb+mIfNM2yRPbD0bMhEaZ77hwxH5DhfRbEw9bC5EGwzH3SBb8uzPC
9NEfnulj7qbNjuBxsEf4Q3N0imVvR78AVPvUTFv5xgIC5chzUoN8C4r+gIfh+hc22oJr2RB6juAB
UFY+/pmhzE9mHEI5GGJoFsF26UhJrWF4TIyngGSlUHoZKwJrPkPB3h+Ud6QmnRQldyasgmqUw1Uo
wT0fQP46VjJ9KWaTaO7JtxR5Fb7edLc2qlg4K80PW7V5jVSzJJfdvrA8jj5Wwds8OgBVzpgGLufl
WnNKWywDqmXIo9CULPa1rVYDzXUgPwzgs9z96+TyKbxi/mYY33PgQ/BOSyb7VwdaQWjQaSb/OWwS
o8/sZ4IWAkMpCioCNAwEoi3Oy1eiT4zyxwY+BJtEvAlkf9/tHBDnpnw+UdDZFyQJ4DCztz3rBej5
Izr5a8DOcxMO53TnmL1IuY5YxooBtVmeCyPXEBjl04G9Uuw3LZP+yFADWrXK23N42/Yjw5mUHXPn
a8+faPR/Y8uhxg9ZKWXvxnMIqiaA9/Rl5MvgUJrtZZi0jLk4S0nR08bjn0/OgmpAftUWr6yi0GX4
LkeAhhkcEO3B2qOjmVn+vakgiyRmZAhYRLSTvue/kL9w68BhSGw21wvvWM9UAqWe4c8l8829rJxO
05a4IJ+xHoI6SnLsuuQ1VOCr9cz40bIYSCkBM7fCfkxszMY2e8+VKv/7H6RYxzOShYxQuqKqnTV8
MNK/YxjtCGVlDCetx6a3ADIlMT6xwnHb91aNO7laiwmphokm0xm3qfxNglQDnhnCcRfmMaFC78IV
0nINGh4ZRFWb6VVjovxVN6okTTeeZxh0Kc6sJ4+gPJ++ALBRGogA6VeWM3aDTZ6x7gUPCCIYE5Lv
017VhMR3pal4lCknE0sXDnsqv8g3aBfoKEy6g3Bk3ygU0vR4Yn8phZT/NRn6C2xwLXkRE74cG8tC
ozTASuolGjtMJqHg4Ccum+f7C+ZANMn/dHvgDZ5UtGqviuEYFVwKHhKlbNofnOLf4+JO2nh4bRW9
2M6WeKna1IPAHQff8dEKvwUe/tE+WnuMa/RtISEB9kG28UAggQj60WjxGAPEkpwfi9dBz03Ll1wu
ozsIEUuT4cBG9zvUyuSt2ZE0Hnm112n4vIdvAM51ZuIy7Hva8Xmr/usKX5BVLvM8+EF+22+JMIJG
E23mHuGhGu1xq2YSAa3Vm7C/Y9h4mrOzIvALoNy81nM9JHiWmjmjt3qaVcYNXYUfCf3UqGqZayvo
A4v5baCJrx7l0M9bCUpgOQr//eNz2VWJAMB2dDkhjhF46IgpDMzc+3HSslI84H6Id3j5H4RW0DQn
KTM6Rh1NLLgNjXtgHpkr8LQO9BdYUA3DmL8JCDQa6tc4AO1UFCz+upCVb0Tulr+Z1yXfp71uw+LP
FxA1GL2QV0LhT22oScWlpgz/L6Bg+JRyuV54UtzDMs2PRYtvPNbeHRsV3yBQG6Y+FocFtolJ+iFg
Uo5C4uKpKy1yG3M4LD8knCktSboq7FQ154VBMBHVwxE1W4fvo9/SqO3na1Eq0eygbOjoBYDQMFic
g/Q3j9Cpx2ulluxNNjQ3HM1vjQQseqj6yfEHANfGPDfmdWCFK3nImVO/9wKTJiP/A0jbREySom1k
t/DQ1yMtuALW0TCYaPsGrDWSGBrA4V9rbRd2ybBdebYcTSY1GxiCT/PlXaZQsJISvsHceSgcNaoO
tDdHNCrpiaWklSg3bT55zCYroppz2GxGrwPjlBViu6+DsnaM20GNLG0Fsbmmgb89DDI8yhK2pCWn
s9LhA5HrHPV0fCXSEn9VDIycx600sG/7/CqODGCXxPr5VOQ4Xfn9ZdAFCy4YoYdbzvD+T8cR78+G
PLmU6HJDH1TtpI9/tQLc8YDXmnpgfF7TIB+SU8DpmJNZ+7vFgIPtb3AHr2Z9nFlwK4Na2MKC6ja4
jB9BBEKX0WZxWpJfzh89q2DFqH/mwhVOhoIC30v4pTRFEPXaPV8MzlysskKjjMn/dHo9zz+gVVbg
FlNIWPMR2fhLMFEVdqt65yBdrtLxC1chRSErermh4pq9JT/Yg/zRwFHEcmpOJ5btucBrZvnuAQ1C
2t7495ofmjCiUyQLF0PQA1AkzzxeN9mzBi/+lhlUCkLdeOsOVLXuYApbYwjsGXGIyzYvB7zh9t9D
MdSX0eDlLQ5La/g0hlLkrhxoRzvb3lY5zVjl1SOWWkvPCvQAZXq8WKrwXllv1ji4C5fNjRo6tYPd
H8AOH+/pSLokP3qEuW82e/sAI3C6C4WLawfvGGs8F9Efqh2MNBPZg2ckXjsacJto7gXD/gZsyua0
Yg9QAKT8TfDhzhJ4OCe/OuLuSEtr4Tt62myARU9eIbArcdZ9uOpSmjQyABP2hPUbcWqTV27t7bjy
625V0+Y5YMaKjOoqDbpjkMWC9V9OABxmUqvaaV1L96uTO0OLOOWGfsyTJuLeXxqbwi0z/QEWB/MO
nt05XuUC309iHXQ5dpRGf6XV1j+ggJvmorIdB1MFXVUrgQGDLAdVQBh0InzyuHfIAVjY2YaIUzB2
yDbxXfCSlKeujWbFQ1HmcYtcLyVq8dnPP6GZrZWWLkTf22Kvh3MP/n7zBnXWecmSSKUVKZ9LfBPZ
EOO1HVS0FIrj6xq1HrBKHN7FoNuMIcyx2xlPs0bB01NX/ea0MK09QqlPp4aHUWbT5N7oNBRfVkOa
ZmdWU3rj+tybWqnydXERdGDXAcgOAtoRXRoF80sRAhZZtBEl1akWj03zPbJnNjWRFH5yShr1+jOZ
WeKnsTtdSXLCQfgWVJfRWiZ1+zlqBcLwF0PGRC0aQQXLx+z8WdxOymnJ4dzjdihM3Y0HpKb4WiW9
WjS+eiGqQTUfUdT05laxP3hIRb4txTTNBeS6vc0QIMjdTZtHZCnE4szwfzKq0IcKF+ARyce/ETTv
3IwUOvv+FSFTWImJptbtw5NYWke7bZVpxBBiqzKDuR+Fsu7sa0r/QYxaYJYbC8hS0Wdp+6Z8hEtz
+UnHeghhGaqL5mPqtDOZtu7di2Tjj/bzJOviRwf+0n8m4Xt3BOPxahfze2cFVimBsvWjJFNb9tSK
44Fwo729rhihhyNy2IESuL+zQcaaBotTtboEEjJ5StllFwx2CdiU5e7AsHnNGWZrAMbnUW+89Xop
2mkoq02/O3cl90FZ9uG9DG3PaIj7QL601Ndm6vtaGPy+kqI6WEU6nww+DUhSd+MQPOadwvl9fzy9
FNFMtxqniIhp2U8X3n4ZMzbQTUuD/UyzFpd6oIbmrTzLFeFAu39rno4YExwoyeTCVDvIMhLHtzpo
jNfA6b8emptIGn4+My1uwwytUxTZ9USAU/aJkGJlQR7wSVnXfGVSMjC7Gd10+lmjA3oIv8f60b3L
C7oZQ/3N1tJcxa5eXnbQ8Y8IUdd94QU/ZO6ZLB+Fat02SBVAMBFi8mOSZIA/OTn6akaD57uqecDK
WcQGk2mzZH2Bu88JO33OBzYMG9Cd8zu/8WtYO80bEDPlcOB3UrocpSFDYYgMf1CD4yoZvP33ntqU
s5FXQsgL8vx/XycuIPmdaITyRHU+fDvyyU3Q77YYLrtirPPxpf1oaCAQN6ypm5+YzjExJJtsGXrX
jPipt0GURkXVkgB2NHND+ah0wsqCOdKW9VVhwhwpkVwVzFnZFVwzoDPhfQqhR6z2DXEm8PyS3Ss4
G+OcYRBKkl/7NA1zRN8C9IsCD6ijctJnxBIXz6e3qqUlLk0UzNO3byCq1EdxXwvCZyzYkb0msDnc
btYN443r/JHwQuv8jj5HqXUStyA2IrQDOFmKdL4UV8z4wPkvuE2cOzZwul/GlymJ3gqQfmU+UhW3
V7NbYZvtx46nfRPwBj/XuU+1eWHUUAWG82NizTH/Lrxow654qJKoUDadRmujYUBy439nMOfVGWee
mSvgRd0TpI7z/QsWAekQfoItD5MmQ9EKiDIl1yMYwOUBTVRFWvsMVZ+GMoyE7jXFv+FmL/kGP1z8
owuQNNQBDRx+Wh73krkS42KF6YTI+QEpLWVJ19FTcR/vwHWYREacqneMXTe3THV60zkaxcBP/Mh5
AVGmmvGWo68TBwREK3nz+zGRkV6PKocmt8PSsihnmc8QIpXqSBC5W/M1Dmy2KTId6WJg5Pwxx4dW
waYXZ0ibSAO69++l2HTFx0hitVo2l+xrvsvwxQvXhQN/dmTyNcOdwk+ClK0Sv33qGlPsQqtVUgt6
gjmQE8M8vikE5245aOfK6YNkwQjU/UeAWLoZ2eyouPtJqCJGKb/xwczzkJgRIhVqwMYRHvv3LYcw
0T3LYyb61bwRa7xNB8YCJ11km+XttviC5tBmsm0Dh9uwCk1WAR5y2Y/NAi7iN7tBYn/zkZAOs77K
QHEGZjHLlMtx28Z3OTb01/UFF9t6RNd8eqcv2E1nqJMbzHteIUcptyZrRxHbqtRLaUtiA6cvJ0Ak
B/XIajAKzcFsm5eQ8DlXI8Qt7M/KU7Qb2wVsUWTLF/ViMjIyGleXO2MXKeMzzLu0KJi42XV+o6Ku
zn56lx8pEPUzUmSsF/N55EOe3qaQ+MGrlce7hOoFIJaHyZbrJ8wQ4zP6LXf1K5sq+Wq5aCEB2ZbF
yHUoGwriXfl/TIS4FGWnrFImT2+Dc+gad7T4w+LSFIXK/9BKnQoWNDhmDl+K5oDmNuA77QqVPG/E
qgwW61jrq6zzhIrsk7hhHAetsUycbFz30fPUQlOussU4VvNiRTqkxKF6Hmw0P2DpfOIr7uG2NCTl
b0/znIAS2Sbo+uMA6wzd+D9P+ZvCUvH0q1nAr4pagaDPKD296iVW/2omJUjUFFCEpmpgDLdQsqR3
kzH8stzu9nBse2u6E8GnaXjvZYekVfDAqbdONx+ah3rKlBcQBXub2rnlWps//AIKA9Lyuk0g/l7Y
9e/h45MisUdUckGUTpxnlOVHyQ/wk0mDU6n1obsU+on6khuxVEWZs2wn5QYk+YZO8T5seKuX/pwD
LXMbE9X6Jj07dYF3E6V+hWCGoasf2mTxTxzRH4dmz6MvtEpSVh4ebj+aIGI3Xg/1RlAiD+Uw8j1M
iwtO8LA+ljvmMxq4n6v+kESHpxAU1HRHvawclzT40xqNYdY9BbuBHcEr+joqjHVLDx+Wk+nLMGK3
NTFiNg2anoXt9UVWeZsu9hGAT/Sgy9/zGkInVSh/Ek61KPbuf0N/DAxxZsDf39dHeXTBwYC43Saf
7lZxQOxMSjrhe1rjQWcCDS2MAFYTeybYVLqthMA15VhTaMRCAlFFAN6b3QbqUDaGr4tJGwgu8wDN
Q9xsNVHwAa2ix3tiNXSI+Lx2cqOfp5gDYYBiboDj6VlwPkc0O5NhqHqI56C3rv4aIBpXK5lP4IeG
zWkj5laIZszYG2RO63CMKc8ORhKtVGYyS0pnAZJOQNIUnP9FmDv7h8xds2h81rcg4BZ8VLH7b/Xh
QI2mMYHFJHUUFrytRY8w7HeXy26cOVZP3qy98kOygsN/oq08ChXhbJxU06XQW7A5gwzA+KJKkH7m
deX5UYGcRPjZ0JcobTtdk3opAkN7tOQt+ww4ykGuadIbZI6a1cAxwr9+9Cq2D8iBdrg2UsNluxlO
00B9cvF7jk6BA/qdDl+OMN1OizW/ZXHm1+ExTHtmZbJPjp+COoEKn/dn0GgnOPMti7tLT2fH5Quf
ANYt75qH01ufuaJ7KmJxkYclVmuKiNYZCeyBPHGnnSfXniCgvcSTTSDIlG0fJoPhTmHYqHbnQSRy
PG1Gp/ZNf/cpJE/jpfZz7UmSTPKRzHIyj6c+c4u64R5izO5MrygRNV5By70FUW2vPVWIHRXmCaY/
NKkwyeKp6iA+9ShM+nrjSbY5DOu/eb6DRxzWW9IfvBXiMc6obw9bYb7LtU4Iq81eDQtZNJLB0LLq
xqLrj4I30NRsp/0UYe0yc+SY+psyEnrPDZ+gB49w6UHznydibZncXMrP0CGMJCSdlzzm/nVq7TXZ
ssa5KAQXxf/EFPA5nzuElgOBAC0QlSzYAilOemOBzg/IUE1t2jsu8bPu79/FTOSvpnnfVxTE8+6w
zMdNumx22ucSam1Hg2Ab1uk/njdyyLsfByVZF2bGAqmbgR7ztO4oW12Od/rKWMJIO8z/pPbggDGJ
/E/6XYi2+7sNf/iD50nCdJ8tM2MFYzoVvrlEtRI9DLgwCuK5vdRXHZUuna1UOBxj5dr1xh2U7GeY
ULyQ6MqTEXndvOn8RvaQfqih5RzBND6zWoMQMw8w2c5fC9gcrLNJRkaZ85DEaeQQFmhsZ8cUqXXN
q7TL3ipNQ98Cup+Q46Qj2YWz33hGodztHA5fB5ViYLkW5pQ+20jGdSuRVCXK2WsWtE83PYYvJ3Nn
KtzNBJSnREspPBCQ+waxrYcJBuuzLyMa1oXhkRZmvPCjY/gPbn/5FmwtIyIWSXXLw8H5kIfzdAcf
zPzaksvoRszJzKFzRRIPt3ip3mwU+hsufq3nrjB+kKP/P8ZwsPvcbCpN0pyAqwxoQWCUjcFuYHiX
MWtJTGXL0F6jgmOE1FizT6ZLAWiNdGfKG+xx6PhaSw99Y4Yg7zZC9R7AD7TOJAkL1db6k4L9HBuD
1lpxs63GAYltpq/IrJSjknIgy05A9U2HVqmMKlDpfDYD64gdh2bXh4DSvmPs7vE6DMqxm7EdK9vh
FY8FuMdxwkFKmAaCfcyZ2Ve+48Hc2NHFPpvCl7SCz5DV0Nx8RLUQ2p5fRyLcyFLLYkBdK/ck6zrA
RXRJnK94WEoh7RaLUUj+hEZV39T7OCp9cMAsvF3RN5a0Aq8nFPoZW6rk6Nl6zB2z8dCIT0w425WY
/VorF13PvyWsKCEFprtzK3xztjXKr8Bn9//ipWGeDQxBVHMUldxTNoNxSRRl8UuuTPkJNSbx/Rcp
K29mRHoT0PrBYkiQHBBG4J0r3F+vK4xIEh90ki8+bBQSfJRBBsYLvuR57dwuHRO0ey8QvI31VOqm
crCTQcWhAipAxtyuHltZ0LTss0Vd1sfpaATLjohrOgxXwAIb1V4a1Ml6qGeCz5Zp9GEvDFmBWuqv
URO2sEH3xomd0AJOfsdVtMLTimItoVSQXNIUqBkLeX/0e4TgIcb7taw+8gpT0ARULIUevCNRKSVK
eacDhfSa+qSxjl9c4kDYL4mXmvkm076xZ3BiNEi4kG+9+F1NurpsWJePquVBXWOxGGEyREvp1a0L
mJPTR0iK+r7YpKYJpixXkhUm56HTp9dLLZCn4yLJzJQozDmifMBTEXylMMusnWw2sE6hC3qmKJK1
6RGbaI87Ef3qGOAahkg/vNkFhqNQSSCGUn3zozRSTdgzMJGvhFHJbxHR9SDRKcO3PLfYjOdItbPN
ruf7KG3JFr3gm1vK9z0M/bAwTPfTyLhpUWWEotqm7MXUdHoGjoZn8k421IattnFRNj3C1Gwc6VeN
UmFrawxNumolcxUkOGCbIs16dmlObLc6OE+6+leOv4G/gOwMvho1XVoB+FrL6XpG9RfhOEc4gLJV
8wOBzYzTeOPNCLFRwMJoyCmJ8Xo1QEs2EhyTSXYABTM3f+Lx5Q6GLV/vs/IOdJNlHRfJ6zgONJpH
HUFPUGIHvODCRQBMd+WhW22M7ZNl2xyGqZ5gDnWR8C8slJh617o0DOPxs1PxMWSxG+T2yZ2tg7wl
sEEFxf8qRYyCBZhJcg+S2waDQ+/mlsTS3YYWH3+OgByAiNyLISNkkzl2A6EMCrfgww9GgtQo9H7r
6WlKEd2lSuq96dxXHmcjQYgHFagm63vlTj/nNtCaQgVmD0oKaY5zGnmG04f9BHdwJxcVraxbl9jA
JTuhiXPXp7YPCqxhHfCcUk+FibyvGSRG7BKEL7l9C1G/JtxLUu0SIhQmWg6j1fXmX3X5fpkINFKI
8fAqDMNKaW8tzYdOLmnrH9uA27yg4xxwgmsbsHK2QnxwJiAioXAQDZlkwmHT40ByD+7LpVAe/Oo3
Wwb8fWFo2HbmF9BptWCeORFyz6OpgAUhcgnLjCMcDdhN9lZAJK0qZARL1DJHXtFLO6zAVsKWjam3
qC3aCm1a/iWTp3KwCOS2d57DD8EEPf0eBDeDxzzu2IboarNnWzxStrR34JiP47455gnV07nCRIkO
LgSE5GKpgzEncAWnX1e4NpPhO+znKU0mNiyHotvuphmJhNxFSAMjy4gPbAii1UXkREq8+7gMolEU
jso6h8MG4sjzvVfPvFlz7okLRf4ATYEi9WiNw8WL8AxC68dETR/KTwK6kSmnRAOheqcBAdGvXeKL
jNaiWND8uhNs8IBaC26wV2wQ5PgUjp5DOsRud7a3liy3Cjo175pDC99fUaqeHgOrx0KeRl32H/3N
+SNCMvK21l/Ungvwpu0XZUHN6pYG9oCRTenAy80E9kDXQTvzsnBwuN+fkY9wda/XaRsLP9+gNmy1
1MW1kA4Fl8P94kkVbSglpvIT02TEHc2T0k6CETM3UbA2zFPfwVXURjWXk8SxYfV9MLksBDReDfAe
32noXz4h3kWUBLEOkb3vJUTj+Cbc/Rf5dEfwtLxE/DWcFE2Z2PxcPs8iu1ilmi0fcas8AI5Nb4pP
y7ORpmJuECOlyW8UR9iY9a/d7D+2Qxfg36uSMsEff/uZlVIlpItJZNZs7Eq8N1Ovu4Z/CbJLZZJW
5OGgP2t6k3pnhe7SVddXIG9rncSFribAhafjabClkBmbDea4cGDDiPRujOFo33Gine8LcCgw0IQs
KA9Yp0v2rxVKia6YSRVfyBo+XjQxtarc68DyFj+NHssPW9gdNKD7c2rvOQSCea5AP0F2zuiXfNG8
EAzyMKoPlfhXxh9zaoRgcP+7CH+iBKZmP0hbctyxybm/Wk8LaYpTO8r1OiJ9xuskOXWkm9nMMYW6
flET2BPvo0Sd6YySC36TvEqQqzbt5Ysp+FSMFhkQ+MBZ8S1Sjm6vT+K8NA50VpxESx643KXCL+NL
8G6PiknNeFl+CBUsxNmHtXbBkCAplfhKtqiAP4rgt/END9oUqHd3New7QEftMw3NYKfM/NzVAovj
MIFkNIC08OuZlWiyU0O5sgNWEer4Wxu6752D9zDSxa2ZJtGJ3WTVD+xSVCEOptV0hL/uLt0Ti7uS
/Zb0n1g1oLuy2U2MBWH7Olf4gfXxBUNbgeCHG1GIZMeIKi8vlrum1wdPGuT8DLCX0fJhMqHZqHKU
RHgzThGjHSS+uhD6all21KA43AtBBrfm9bE7P1YIF5HUBPcbDuMTOfJBRV3yk8WldiZf1QrXkoWy
ceNeESpH0wE/IbXstJrJPumfOa5RL+8DsmHca4NxBnm4NhfXEakc9WzCr+ugX8zTr3q4nh9KpSk4
0X9hVeyIOfyK6NircePFlXSqAKHvX6gTDqkZonnQtF2RRvXiTeT2NQmT9xSTLnnsoooIFQtn15Ao
kIYeohEkcIV6NYcLtfTHdNfw36trkVqrXXtOxbnyFrlNrwiriLV0A8menHz5M5zBdDAF80bW7KQI
Xo26auTRu/VwDekSOMSbI54T6jVm8d8ZtK0p/pb0fB/OG5GBuz3XhKf+EguFKRCrSO4ZCq0LXaJQ
fcx18A0VK9hWk/FLCNqRGwHZ3Vsq2Kwqsn5gdaqRWAbOwfhsFOXHI6VofPRw7jrNLDr5JztXCaca
1rergvCSzvQsrXm04aVjkWhGPSvw5vidKgJ+NXNjNq4k7xGhmCFDSP/3maPRjiRkQB4weLvRc1Kp
Qb3ehz/HkzNh7kfatVR1mc2AVUMQGhgwRoDrT/Za+76aQs6LwQvQ8GpzVSV2rrprA2/nC+6oDnkT
TLDeFQ4E7iQMPNOCaU/xjv7gqBJHEnMPT9eEYQxFbfr2fgJtqlzc+udyNtNb+W8EdPgQFn8PWxR5
l7d4t4Hi/8r/HIaWPB2tCide9Oa/jPAyrhcL+MZYMCbd7TFlBLKD6oeD/bhWmg4Mm9TdiPoiNz05
XVdVM8DFK+8JzXq4yYdVMYkOr46PqymsrgAiNihztd7+of8+4rn2c8c6Ot0U+KdZpPwR05Q56ir8
SnhB0AE5GPKj/bhs3ektnLS7yXkqZMOvJk+gryB5id5tJwUDyglOnarHD0gxggnH7IOj4aNC4vVg
QO7NKr4xIWRzrBvtnRPSssEJ3wzayrf6o+oQGoHT2owDbUe8wzizjLZvGhTMr3qGrxcMOukbFRRS
ayu03XRGCW0cbX+s34BDHtMMKwwLzbYoF/7YcYfIckZfJjR1zc0/ZcArhiudvFMjCpAdt7ogFi6r
jPcoYf/syn/Dvv8y+7uc0j8e+98Z04SvwVn+wOOM2lD3nL+BYWule+2DFZ4g6jcXa1ouYbJ9GrJt
fKefUg5MfUVxR6x8cAs0ujtKUgYMFHcCT71LROoUb7XLTPEvstXzr8CN1tSbmr4T0TwEVK3kJNWD
JjMWf21Quv18dnsCFICPBmXX9Si8AD4zTIfN4C1adQzR584R5CAbH801OBgEa4HJII70N9+hh4NF
0UjzLczwB4phRcSRJ4oi4bOVEs8YxNLBStD+a5yB+QsSyXl6HKCsw1aYdTHD8vbIlJCtWsQznNTs
r7qQTCvzfO1pBoMrqR1G1NXuhMpsl9nu34XNoIxPwOrT3sdo/vdtBObn5bg+ASfhn2i8UGriogS/
sPe7fVTvbe7cS1JqsTYhIFU3DJ13GscvwdKmByAhGIrLGKl5QkNRgtiNdwzDcJiAyK16z+4IWil5
bc7aoK9g6jPI4qot3N3heZsaNN0I1tXKpArKeybqZooqRXLWv6P9BJU24WzL1GsP1QWPzHILnc9z
Su7HrpXCGv1RjmXfVKUiw2jC6MihSbPva2YH33SaKBhB16QK4zyRZQIdQKapch9X8n6syQu007yG
1Es+k1bMkbZfq3lPYrYvEsDF11/A7dblv0FtLCymbpQIJ/o57iAvObbKNeN3v4iwZTr8PUC5caRp
kyB4r1m0GoPPuCaF1i/UJP8qjIIrIkbtyjOpfTzzXIccfxdixBlH5kDXVKu+qjjPmVsiEAXAMyES
zJJiWdSR8KxJbQgyosPzOM5BuJ5V2Cvg7U+B+UvEwD7IJwYMJc8bIdleJNE9cX0ihgOUJrGvFsIv
QPwRPHGX08pg8DRYaoLyCjIF6OsEBiZ/HcWWiFFxwyBavswTtBFls+8jkv8N96jaOxvGbfr5ZipZ
gYk4f2Brn7Qmev1hLwo3mxfcKslw+VkVFwQJljUKSkFAQqrw+lLcWT4GA45CNB0qoJipJ6ASoG50
xEQioaCvit9pDBH42QBCE8wyKAHc3k1rxDWYBQ+FjsIbXNYCrc71gque1CRyk3u+0vSxp9xZEAVr
Z0sGJJiIYTIOR8uQe69Z+t3WOZ5uToxYuCl1sshwHVdUjp7ENvrWm3swZzXQxPES3TbXqThvay+i
UvltyM1TJvpHYRpoewNIkASuSHPZ0G6cmxnq6M9GWvMJLW7H2j8peQLMTnUZpqXk//c/aqFtb2pV
LohSUln1FotJiAdrAkPmofnfGZnSt6P/OKeW8yzdP8SA04hXJm5zGivkYaKkxJFBHPotWiWb/jA/
zELEX/S5FmA1Ix1Uhsp1/bxNCB2B7B3+IPY9cMzdf7c4rIHVi5yk1itf30W5a0dmop+4inclLp9w
BzsbmfN7bu6IqehmkTFQbB9PARGzNL67JFCqvJyvxV1vIKNYw+HvQ2NKLrqv0Bg3RMW+IdR6hrxJ
4Fu/nwFLLgntaRf9pI79s5nJgOtbnqGeOk+BK8BQlrwIFkG+CJxGPFMXqvXp0uUWJWWipGXAVJKP
PM6ztyZfmPsQoWwe3BM8/8brQU1zfmwevS3Kn5EAZPutYj38J5+W9y8ioLq1xokTtPqBkn6ObHFI
mdsiXtYs9raxJIa+n5wbL3MQOABOquLlnhQK6uYCEZiqMPV/mE+i+xlf563zXhjRN/5Xfvt9HQOs
7aHeLAG8tklE9oQ0U/yqTMAcIrmSQyI3umjAR63YeFTEs3QIxdPs39GvOtM5QPBMHUFd39qbrp/v
5rJ96pva6ZO5GWmt099YT8JGv1pfHTJFch/NJRZcgOxTUSw7RJhW5BSz35cS9uTi+sXCN1MEG30a
4I2uYl47vlSlHqogHuDn5yJu7XgbjRiATfrZ50Hpv6fGMEslXKPCyZnHmW2LWEZtC+tIcxCjmRk0
ELeUgTPnrCpPzTFg4wjdY0ll/NCjJiOG9lYPYGT2ULheyWLZPNmEkDslNI+xrmLPlKjcf2ahXGgN
nZXOqA8VzNoXrLQgogGB+52zUDscyUwN09KyPvdZESKBAshE0ND0hJ7mQMan3H1ZOd6i66KCv4HM
nZgERHNfSo5klI98r3o0BxNhUCad5C3Ri5ZcRAmxe0p7Lj+pXaFjkf4onsYcetOaz5iu8ai0is/r
S/bpPH4j0AnF83HAVODiSjzwh3q+Hn5beXRAnkDBmyXe/6V9lwsUhVuJW9ZZ7t08TaIF2rnvl46F
O4E613M2PeGsi9xT9ss7xiVis2sJgYs90VT//ZSFvlnKTy+EmJyJAL3R+8OvfwSDW1l6lI6E6v6g
rZhyfl8MD3h67oVkXghbhGXDBiTo+IjSx4WCycEihzlDtDlHRtUm9Jzilj7Mm0KtKnhuW9ZTXAaV
/JkZ9fgiqghhB5N7YX/lqvs/GasLj9QgUUp9B/PZ8vouehWVyS4zC14Po8dLPPlD8EYWHK7Xl8wD
ywbfrGspC5J1X2Rfk7V0E0GeXSvsRck5M2YXyZebvQb93HWNqH/bMxSIrZ2qiA3qWAxYztJbcYa4
5A+CIzUWYJUXGCMwIxBOjOIDSlxoiczOlmNjqiZ872saS6Jef8CQ9pyyH1K282HUmd1w1HgZ2zzd
pe/MbNwcKJ0J+Rm1GaYARbHYEgKCRA2hiQ8uU6Lo7OPYDU49EYmPZr6jSr5B5BVf9c/RMUG9XJQW
4Sy1HjZ1J0eglE47B7dZlDd/Oi2kEB8Vbcb0FQObPWX90JZ123PoHR6bM2Z05ZDtiScWb6JI0KPh
zCCDxCzA41s5oG+SEfv+xw3+wmqxZ0CYUTYinzaHUQnuEiBU15Ura5Jvq7UIqNmtqtKmNevrqpg4
eRW0z9h68issNn+3e8oySsgC8pFUXcSGfz5hhqBk7iTF27R3PGio1+lr6udGSuoMPmTHT+2ZnJe6
AY5BMuaLGsanMQBkIBEwN2omI9w4k3TwSLM574aBeY/flFBLGSc+ZOv0LMWaNyI8Vww28JNYMG4i
VrwXIcjX+tiL7cEqSbuLq6wS6t+Ag5FrPRNIgnGEKVXoCqUHBePRaMnfP9rPZN1xfYmRG+F+rRPH
YlnITjK76erir/XJVVly8kr7tq7auxhLD/9hWNaAPoF+QEuCODdnthD9jBHlKTmhsrQytRBb/A50
Cj+xeOv8rgjW7Wo1PouCKZ5w4XkorJIeJFzvEI0/GcJfpWjFHDqWKF8fL02EEgZqgHs6jG7MjG4m
lhUz5jXVFU+lxwBrQcIbMhSWMKdbF5/OGPEpP4DU4zVEYv/ValtvnpPkMp8d3WwG51KAHVEKD/BB
Pwib3r2PHeNotAnnEVYzANQkx15fAEWB0zmS+KsHQ58n5sTIGY1nWB8buByROe0s6yp8336FEAH9
XpP37LW3epNcU/xSnIoLbgGLIsqjooM5eem98ChTYHVjqV8oAzyy+hSU3DbcgROLcQWBHN2v1CR1
M/rnxEmo3cRFaHbcSPY3TXkP033Af949eV5gnmwZF+CZHob7ECtbrKzShQ2W73ga7UKVonbwBCCu
ElV8DTXAglCcE/2iGRlFyXlynwCzhSBdVvggnGv6MhV1KWpyAcfIkENnGZOwCNY9EivMVCJnttU8
ZginBGFtzVMc64ATSiDbFLewnbIXGuVTtfwFdxJfsFIbUqw8HCBVGdxaRs9xp6dE+uIrpK+p2TFe
5Xc5uS0mKlQfsl7OAskXPLhy4eXDjuxUGc3EaWsEPw3/xKjHC4a3ucJCVElB3zfGykdHvdXhA0Ip
AJv3NovmRmycPIRnh9asV5RHGnDhaDmSWj7Rku156Ok6SXDvlYqwiJW0JYBazxrOJFyteMOP8dCs
qW9qzhxUqft58zNZBxBwC84tjzaz3QtD/lvUrm02tuzHFAQ0Vp5tRb9aKiW89U+ij+BNpSAIYRMy
hlw8RYjCnTcyo1+6klZ2r7p6G3MA1Eonzg6zE+xtKszIWPg7LtTxi2p9PlBa9z7/+deQ9jQzTbMi
Z8I5tefT1ito2dw2aKXuJ31WcttFHQR7VOLqckzA+OTnWIdfCceGoDcX4SaupvzT2QygCO2WrRAT
cuf6lfJT8m60qiZRXAYFWQhYiJWfutcHhroyu+IF+Mg1eBRo+knnr0rOUN0w/LcEifEzm0v44Ihl
6E+5N1W94+nGrzzOQe7/pyAxfaWTto1ssJlbIJqZLPJx8Vsez93A2k2QqIrAjgn4TI3c9wcFkyGj
2+GP6+Cq+5hyKawY2vm5Oc/Gp6OVg+FPyFQPA+PcCLh+wP+2kqqYGmmjT4ZtmSiPuIIRMs0CTmYv
AZluy3R+AqkTLvoUkOzrC/NYqut96lelXV56EJxHxqelMxZYv5yZMtebpzVj5yva9/K3OP2Cs/Lv
vfv42MTICOa0hOq1/s469M/v7P93yiFWsQiFYOph6dceGrgz9drQBeSLSQhq2hjMkoskgGGKWr20
WQk8G+ZtecPKx38GEPCczaKZOZfmpK8LwvqkRcGKcxRNr/GYPxHZUBu6Ak9/BvsMSwQzSOBQVUZk
576uzWoddyhZXbvxELk6rA4b8e8gLtrMHcKOvSMOxhhZU+zep4E8M8wP3BJwAqXzuG7JHBKkarO8
RAhRwiL7dNGhkb8kAAtNPAZ/zGRk3vM8MCKGMF2Cb3I22WgEW9bNcNMtQ+AQ569g1qbN1yF0cFB2
eTZyjdYrw252a6peJE9cbXxtPUzDeO+ZNk+i7t9RwmjRNa9vp9erR9c6MDu5uyatFGuhWH+dogzd
UIQTplUFMaKDyCLBMX30cQ3tIrJPW+qCY4+n4yYlX57vdZH0AdWrtK9tkIWzuJvq1dMHA9/e2Lx4
4K0diMrvyU1p1tjkKs/l9vvFHuRxMuNdlhAoIqHwH04pvhGkbCEqO7r6Wt/dwcjwUXOzjOvmpZ6I
C2h0f9uaTYx5iCy3bOuR21OnTkIOMdl8V3H/8fTKsXFPxk3Q2UZqhBoJGQnlz+KAAr1TpJ8lib12
xIw5kn0OQO4fj2CKmf/Pa1EWLCGEtam8/aowDyuOUnezi/XIqkvCo+OAJv41lpfMH4gJgz3aY3jC
WAsJBPPeTzJGNRNNwr4RDp19qAbo1Jn2D7x/OGCuLiDILkMkt/+FE9YM09qU81+9CKzEyLCtRK9V
ZR+nZvYr65X6dqOrJb4l70f6XjtHU5MwEDA7FOcn5RQUL10Lp8wHKt8PXOO1h19byAnizCFqahh+
H0CndLKV0hS+gF8uXv7Cyqaxmm9Af6zDDBhIb61R9GhW1e9+ISZ1pzqa93BF6VPqFm80onhZXdTH
R8+s3XpjZrLNqE4y5lpVP93yzIW4OCzBZ4nONPKkskAFa0IxoZUGBf8oGceTRvVI3iAUEtxq3/fX
PoLf/HChBUxWtT7i0hlFVeXxonM/9X9iU/N/gU+hZzPfdW8dIzSjoCcwyzmsJLornBMJryiWR0WU
7MzRn2BUYsrh6WBJ5fDpucmMv4cfGTnbdXbgcXF8Sf1nD8LLCXdgEy+5fnPJckRdfoRKGLbuNG1u
HnMS/TUo+wRDX/ZcMuM5MzzC7E4zQQFckTz4Gbq++sE5lluc2irSUArZY11QZzZLxSHgLifoqRHv
QCN9uLr6wU9rFu2UXIisXUE47uBFSvO2Zag9I2ckyiGAwkdO8MW0+d2v6otbOPru3eYzayOdjD1g
sZLPF3J+z2z4WzJAAlFZlbD6AudfZ4kPzHgpqhgQ7fA+/d53zez7pXFjug/wVDPQr1dZeWkSgSwI
LmxwqPeOHXMbZRiF++tl1/jC6YmNi08ZSHSuuaxLYZb8W9aBgy239Rr87qogYumbTuPxaPyDoFcI
hIUHcu1twZb/SD4fCL5DgFu0gCG4o76s4vqCieIpGFScelAmnk9GQ1pSE61jPJjvT9tyt3D5TVXx
YR6JE+c1ouYpqB7AO56JikXdkBS2SOtc1hzeTRMH5N4FxI03XT3+95dW8EA6W8pAQXm2B/IbupK1
f9RamAdbAhPgRlA3yu8f8LZX1ttX71FQZXGMfjD7SGgHP2l9w/IEJauWy5MxvPJZ62f/ZseFRqVf
zER55i227Dvs+GJksv0gAC2i1hh91jjFm2e9G6vYU9GZ9LW+EXRgoRTfvBp6lcBJOxMYf8awv6eY
H9ePpvTvz0cXnqu6GjZGI2XaStfklNDips7KQo0xJbyVtm571qyFO4L71+ogIIVG9oZ8KQ9KJuq6
D/QJGrJwbS5FrOoFmfTydLGWEQgaWp7DHaSnm1W1DgZRPD6ba3YVTAJKOdyOl+YwDhpy8jWk/NTG
0/GFfE/Xgi2S0dW4Z8o8nEFW5s2WzaRvejQZrQ0lzMveJvY8En2bWxtpbUfDjxZLX00pPRiuGHYy
KHEfiAuHX3o0EwDoznwEzYtJW/64NF6Q3sskhUiM/6V8EwH8WP4hKDUu+QVE8kozSd6VG5MZW0Ff
Jliyq74kK91vqceRkyED4VKPiGFQd7GSH+J06U8NpDWstQOg/1aWfnTOQKtunegwNlNgOQLDlgn3
R8/A1OFY2MPX6FaQagA5zCP3UfiMjqe6ggmd1X/SucGjsxk3nIuv3o7fh02Sj04frpOf3Tp3ZldD
2FYf2NU1gaJ5hS68YTCrPw617bYVRX4sUrI021uScMpxdkJeForbqfkyW1kqJD0+Dti0lkUF9kMS
QU+7VFUCPA+eNCrVu2dp5zH/VA+nKaEme9x/1cxlX4MQVxEMMd0qBMkJ/Ug5txPA/A5AUO2mnTBa
3obgOPvoLIAE9AxhhqOK0bGeqyb616FMkcnDQbYSad1ajvcsNLpsWHpWQGe7mxwHzZCnXoOqPTSq
VFeWhjV4/aR/N4p/rbrB0MI0ok+/wh9RxUkNWICqEDxw6tO2keGnMDcL4GgpJrfXm5ylw5/BWokr
buAEvW2zMn7ez9+IRdCxNikxd/EQmpT9Bd2Yv5mXamhgdEkQQpwLanZ0VOrFvm4k+EFQhN4JVzye
Ry/YOnr0M4mDh8n6olmDU8lEcKXq/wTtXdGAgw/DMNJEHNh18Ll7LSbFNWfKXZs38i31zN6y+8UM
TgniH0BwyPd6taIqerrGMInPYqxsCTaIlJbMzvCgCCTvPd2O7yEUMcmWnJOr+FO7GrUyh8Ll9hsR
IWZ5kIiPur7VmKerS+rW11nuh95YE+HzbTi26DRIO4ynFM7LihYPeJD1mAIkNBq2LhQ2XSpubnGD
/YpifhLf3GaCAnH8GfEmLEoQB/X4PNI2W0aGrqWLoFHOEFCg0+t9wojJeHIa5yHYYpfxW4p5Z8hx
2kJ9CUFann22QzCUYd17pe7fQh9LXiStqNtezeOLogdArAPYdbH8fs+e7P4BZHTweQg5DkRN4n5B
DrY4mkpo0FGNfkeVdF+vhMHo1AKhtMEK3NJuGRJ3ItWx8jGdBTcxMgx9oL3yz/Foskw0NNDoqNbA
7drJGylm9PAB1aFmgv2rv51esS0+01ov+I1D1eAI+nWzBk3bw4fLI/9L4Hf9UsDDJbFgEfm2fFHB
Lp3FJPSr/E1lnxG1sKPg/POL/+ccmx0530voIF2i+7R/7zLf16WVRNpk90YAdp6CewKdyMaFrj3B
KA/Zid5LbbLVBvSCnVodqM1xRdROoGlTJ8AblmEH3gB5wcmbqbDrS6EsR8+9dmLcH8eoUlLTb9kD
R1BGH4BkoYbqpPSnt94RGSgip9bqdsR3srk+DCOMpX0bAXcipbV/R4d2tKNk4nGqRiarY046eC0R
x5l/KDChWR1FkeIKUzO6zHQOAa7F4/Tttsx8yH1PqCUHt653GIa6MQ9/jmnp13HvHdqeJXvpHCY9
rAOGanb5ZRT8qfW8l1MIWJ5jGXsSTosnQs3BbkLrXI/Y0MXVwFG/5h+o/5ebN0p0R7XMJA3wL/dj
br5agUzMwufNJFVijjDx9oDj85De05oZ4JnNwJ7x46sQad4LnHbwRAFr9REvVfOiOL1AkCXnwYVj
tnbbOOB0u6NNJF9HUsxmkR6T+/9YuDWNxgJcUsfOmxFT6b/OL3jfKssgI4BWDy7zoH6f0dNcYoLi
93R2g5Gwo3GEI512jC8uCqM0n9Zb4Dn8Ili5Rb6VQ6hMCOBh6o1iSTuaCmoQMdUk2ODYIYGpCkLl
EBB1BrTSkkSE+b4IX/GHifzzXsIq3XPrPZAt8XkTMzpEvbN8txZJA3eYzbFuMsascV00Rli7OU3A
9NIIPYBlrVutf+W/TgEObjEQuWvB96Aa+pZnAJfsaOYsGkSEQXLxHZhizsqIPfnJzGUq9HqYh/+h
1SEJFHLW3vT6ghTWciD4RpGQFeYR7/HR9Jw9IW/s9tAxFeMLZp5bv30bksDmyAkH4+dmGLG6J4d8
8tZ9ErL3GKOIYT6RhRMyPjevfZ6CZpuQKy4oJXbgpJ1JQklD5poEp32paIXzaeAdbaI3+thSXk5k
sDY/1/Oruj+d3Ts5Fu5NAHYSUK+UywqXxXPey167cmOzqLOBQCSpeUI814yyWqwHKouWvCSQotza
m2GLjEntJ4ptbCSTW6u38olaZPhwhKPmH+cL5WaToVc2OL03LQCoXiYNm3k8O6GAVGS4T4sJkXkO
cnN1w1ZwomnzDcoJk1k0DmiNVtof8mJUPpKsRj89mHut7ZUP2piSAQJykX2AMnnDCE+rsUqldaB6
s/9d8Xd/o2SrDW+G8/mKiAILUnOeaYsXuRB3I5rmkILPmUfR5MdOw/OoAfa84JBVG9umE5/RiWJa
CRBjhUm/sRDGSQyRa4NtMo780zfPq5jmchP9wOEReaE+vuP/YgpcLNNRChlH20XnRkPyuW2ZApxc
QJrL7NJTGdLaLZk8HNDtkqPUt346BrB/nMQxzutFV6lJYwa2qmTvcV6SFpDla63DdjhNzQ48aq3C
MmI8bGAsBg6GS2jlJfYK3XeUlY6S0wHFwfSDUzbIqj0sFLlHRZyxLzn4l2DFG55sh590YUkgJe3p
q8+fg2u6GBZ41AOS8OtrN5aZsBJb0guXYHpWBVPxKmuE7fkiMA8JamjHm3JsEAGwhVbpp18I2ds7
fcDkJmmqVIjHX3doutk3nA4SWC/ahWXUmzuqUIJBsX7IEQR/rUKrg2MD4MJlw7p/+6nKr5jjgDBi
CAZv0ttlJ0sko4lY84RsXjAfIC5rr/qRYRwxDxEkVNv03dp0khvqvXETUyOz/RQCmUx4OXQ7Mt19
XUtJZPLa5Cn/4gQNbsnp1iiPWLBRq+ebYfE/1TDVJghtJIRYm4pIF/4MbI35Pf6Qgah5z146KZKm
DxVhVw5sqp6Ig2CXIh/AVqwBvECvbOWBiAs4FmQE9WMLQLBjG9cGNYygD05siiRMoqvioeLV14El
moeR9nmEI8/XL6vYEz7gBAYkJwPiAlwdAvTVALBlUeZa6BQbxV41pxqSrtMGPQJQs/ZgIrUzMhMB
yqPavT7Z4+X2diIRL2FmAKn2dW5EE5vbj/lffH/eZPTWOfRC/rXHwy83f3DPzVCyepVubzvjzOVw
5J3euzSxv/MqTaO9nHdiTfXPL+sYLZpBdd1FfV68/UjAPzcvGa0HpBGXnlyNdnbi3XWw4N7hln1b
37aZHpPnf7hdahCXCZVNImPlNMcNTvU+a3+o0X2a9ej9ljHGYFg+55q+9ZxgX5LXh9Tj4maZBtLa
N3gMakTuPoLASUQa8DjRK4yetFi5jOesiFkUdu47zxO/LSpZiClLUyI5fhwcQpuDjuQMJ52lErG0
zhHJEuJJ82Rrj1uWg01Fa7S24sY6AFuXIo0uX9YqD6iRAZMkyT+ICBQdf5T0EM9H5fNlKu5xUPiz
KsnyYCYn3Qu937zVSBQY+d4HfAVkRzS1arid7PqHKYFz6BrvU3CmJzN+392HcnFxMFQ6BfwnuCOR
X+h2p8aBkuMuaT74VWS8NKLFk6AtKozrpflV1V4A7T3WbHnyQY6LxJDWVtHmszCscg1VRYiOFpyd
h6aPRwsrzBxh+Svvzm2Y9ci7c4sSERsuH2ow6mmOpdkoSpse7P/asymkfRosxjSOemde4mi3NULE
aQxF81fEkegxGw/qFgLpa7VZ8Qbl9lBKATo20GlH3lvPgV11ac+0uKOZ9F5dxlV45kcuB3+AA8Tg
ZfpNDJe01oUeO1P/4b1xRXZ8ErSKpAd5lPvNIW3tvyZkYDB73uh/b2pXAGtf2jxjzmveNQJA+JLA
TjEuuNHi8yOqsHIDS211TtERFpxrFQrzvG9RT2fF4gM4v0qfOppkFtEZIlaqcHF0sBrfLtAyOdXZ
5I0/hpncZCv/wPyVlw987X3J4W+lVCCnqeY+3m069xF6i+pb3jZ7OoVAo0JG7A+kzNl8+kpOJPnB
mk/3TcWgSMO6j0hXXDgJ+o2aGqqKoXnZc+ongmU4SxiqVQUM5DVjDyAgcmDf4+0E/SPIaJYJkgVi
dmdUWpcIzVqofUWPgKBWOHm1xXHSjSp+g3EP5Uu/Z04LmsumHtnJicLuGafkBz8uhRWN9rbZoM6C
zogpkAJk8fIPPfIYrAkRqoiHj5ERx9h99EpZ8Mj//eO1MAD0oeifAMA5+AXOQ6c1hyiFCNaFlHTn
RUYOsIKv24ag2xG+MMU+pJIjOhPI9nta4CkMFC96nLDQqZhDWPeXEuvweNBsbHEH4GYdA1MAWB6C
cs6nhe+0xSL1x+5D2VdJiToa/QuTRdT1ziPJBog5qs1xAkRFaaA5seplgA7JS7u1riSY1mFqnC45
RHIPwAQ/bcLuoT/BxRDvFmRDNPGmUy+RsDUrznBf843O3jelv/6HJmGfRzE6xLY6bVn0yaHeJz6q
4nEL4PMyIeicvTw8f1nsheSA2MWLvscDggHvql7p00KdqWqUimFnRqoBquZSK6YU5tQPEpMW6JCP
8IoQVwcs42GdjkK5g/CLbv60FZ0cCTQ/h13ZsLSlD88KM3hUBR0o5v7v4ieG+kIB2su09H3TLiAM
DC4OlHHz5VlOYnJ8szsu3C7zK6JPhnL87IwgmodZHZMSWerkSblCzO/bcsByw8fqtBh24v8bwe1S
mPp2bLUUf/M77XwJWeZ5y3ovqBvWT48b5OIgWi/QTqGJd7CVGUwZFp9MhABz3iGF9CEY8QGFuV+j
uywJHcCmGJALDFfC0blcifiAEkkRnNuvxMD0gwslxiEAEsKd90eZme/DXKPQPYqI6dPERtOmZkH3
8pbs86/H39p82rn5/TCiqXBUb1mk0FdwaHyveuKbwq+j3BBHYwd7PfJfozSBg/JwZQGuvzUJZo41
RpPLGEAvTCsRXbpeoU3LBszkAI8cVMuysRgKAgGdo8ftgiWkP9wCThherF6tktrUCfFe4CjD2/ys
HCZmSX2y2D1xQqixhseqDcPOJOahakFDQA2u2SSU/7IoOzYFW6zhmKy9O3iBBTykWF0kqdpyGXnn
BPI83cUaE6XhrHnBclQLLlwzCS7ZizgL2rla4SgdKDxd8MFLmQOZjpIsRL5jdLUynquGip3zhjyp
r70+gj4oiW4nIY24YRw54ms+UYYTovXIciSkFa6+1XRmTTz1N8FXuroeBsyb+2sQPPrqWnAjF1O4
iqXGQozGciHB17uLwt4DKEOiyXKnQFuViWvKEMUXySODFvmEVQHX4SPNkG5WZTbWZhAi2jrlAJ3h
yVN0KLYBxiSB2quYc77Iri+ilLDRSzuqSbYPj98Dy/bAADacL4K8JIim0pGG2BOYGncJ6NvSv5Yh
cZfKL/wEeVzlEnYDdRHwTx2DdHa7CdYU75TET52oDpTLachwtS8dcaZK/bQ3DmBj/hdj26F/dD8C
DXZaQt/esYPs6lQT5mVDfeL/W333aIf5xNLh33e11TpyP3QCdI0Sxie4XjTkg2iXERwdYmE5QFCa
AUhe8XY1NyeV23v1VWnKVEryby75kF6lbe2z1Fwy2VrO+prPRaJTY5flI6f2365tezin5N3K4V6H
QsXVxPr3fUBXnRVZc3EnuCO35zvycAiPHvupTIBYLkJmQUGGNJpBPhGEwHgqlcp4YhtfSUKl0cmL
TTOFTlXr2NYhiFt0tI87UXBtur9wusaQdZ4sQV3tyiM41ZGIe+ykmmr6x0JDYkGfD+nyUOmL7SMu
4j/+db9Ou+f0bBlp+2M5BbOWIbSJkIEM1WvKNpDNoA2aC97yK3969P0qHchfUMIsXsJlawCDrM5j
A116F+JWy7r6ZHy4J2xbzpUmTJpkIGi6jyQXNcTGNEyXq7ioUtjAV+T8rXPyKFAR/2tzt398F1Sb
AWwZk6M1RpqT5Yiktta0L3i5Id+ZQutgFAh1KQHpyLkNR7UjgSiupvtmHCiZH/BQmhNJ9JGue5C2
Xpapptcc0l9RcuXdSJGtbeIyw+G4RM+96ouPcJSGm/BMSSULVpQV1XGU2ruuaLMKc67a/xorat6U
IzsvnHwoxAE7PvRxLOD/N37Dhvy6jF9Eir8Q+4cuY1StH3Wc+rtFJfQqXQBqM9oUAPSV/iMyjvEQ
jt2vBd2LNCO8UaaD4sBuhDqYrg+WHqlqjuJWYPJ8j2UWF6MoBZEpyFrKFUBNrYm5IwTSgu0S22f8
p28jO5SEKVSpr7k2ZvLqRpa3YzDyFOSaVXapA9CYElUftXBMXm3a2XNwRlM1siM71bdjxR0SP2Oo
65jFSBpMD+dyWMrdDxJp2VKEz0r+r5gS+yl8VSIVOARSddwoAP4MeZq63s6hsX/u6urUvgSZPzQt
N06iXojDmRxrplziy4rJBClq5LpNm+ZdwyY9ihBgaXxdcOe0BJduHXn+xA3L+iOQlDCbr0cIP6DC
f2nmeRUFqwBKLKV0JtSk8zPW17U2W4pPsXOC0TYw/K+h0oK+CXXljNUUMOcB0laQ+ocoilgoKciQ
ySNvkZNV87Ju2OD9kDLPAkjbUdJ/HkwvSJRI9w6NL7jjUbKT/U4mzpP+sPcXir8J0O6zz7u9M8Cg
tT22fn4ZuEKdjH7jWeylOW4xnC6PdZKLm7Y/JqAblmdtv9/4JImup3ppwKFnT1ex/5LhQfQKxctM
91AG4tm8QDYPma9n1Ff5YzL8ZZ0ePvHk9oy+Y8RkTH1X5Hd/45MVaGgWx11SKn6OdokS6TsrH7co
ARhX5jmijuK/2AHsjGGTuT+g3qxeP7quYj2/pDhQ9TVBgDevdBEbmpmZgCpgch5hfScACUeVziMO
1I/emEW78nvVzTnWYAP3+PqwqilJ6aYqvR60zjnMVDABXfPEm8qZbP+vmqr3ZVtsiYZMzl97IFjl
y2vLW6IXcK0Op1tdvpK0ppa7ksptbMej2IGftUEeXzEUqh8qYZJWYCATkW50+/0KMG+aEwJFmuJt
DyDrbAd+9B3YUT/rRNIYyAAVjyx3atirQl3OjbOjz+0Z1TSJBImhARqUZkTR06SkD+kQHRvDA2IN
+S+fm9uwCJg0zCtyNyk75qTihFfe1k7XtAnxNzg9mydGQuK8/da2pI/fECO3Q6e4Mpchm1YJsxf6
Lghi7PQgCImfjBbgWAY2C10gofNwBm7YwQtPQUfRpjiiGiZXUouCVEwwyM0uCp4HA1ufP0xjaszA
oi9HszxVzDh57/j0yzi/QIKW9BvHpkx+Aq/jT8wtYYtFc/T4ybMu8NLKn0Z7xQ8lYNPty2+SP/hQ
2X0HmbO6zEEqGmMLHd4E32Eh74rdRKAznG3YXtnQILjsUkHZbhF1jXKv/4FLNISNH1h2APBswb79
bv8IJBK29scvHQ9SoY4rj4OlZMYOKnvDkMePL2ZIlkKmP8jMaXr/I+PAtMiWot4um6FWQHzEgC0v
XuE1Ed4QlfacA2tP3X4V8o0D00sTppCSlXOlEcS8ZhmiVZj559TvwIUe0g89LpcPnpK6Q3DmsYW3
hPHA/0CvshFcCdLcN0q3VI5viPLOZeZjF0R7L4SYJyjdrPdsxTNZeO61L/SVDnP5hrgBxPq/N5YX
7MGP6e2PWE0/ZamrcoR/a6ZzrkJkqEGLeiyJabZrNrg8+S6NZDoFF1izRBf4DlSl+yf+m1hM6jVG
N9/XH+hofJb8MgqtVvotC/KtO+2HaHiKW7IktWNAiSiKc07EnQleTuG8bPlDWcy5GLxhYBQUJ2gp
4zfitp8i1/bksZ7DpCQPR+hGMXyZ/8BkDewUKEx6IM3aSo02Z/gmHQKJM8MSm/3C0Tp/xF6hrrqi
yyFeWJ/zfWTer3EQoF7MabR9cESW7NIIG6lHaOQGnxWxtX9zg56R0WVxcPw6/LDj/I5MqIHWfGRo
d4OHlf7z5Md9EdfQgAQjtsLqZDgJ4oRjzPCQFaiHJ3UbmtMGuqUqisnNGNI8HUJteIOp14AWVJl5
DiBCw9zNgWByfkFjV3NcwQRVWQ3JBDQ6xu8qMhTeK47qN4gh3dJTf/1JCCG522XILgpiu57F2WH0
IXBJaQuYQCAyXO9eLrirx1pLyS3OI/oH1pmISq6nvKOF2KL5CcDITdfB7IGOHP3dOCQQvxpjxkcm
yx5e9XGrh2NxOyT23ZRQPEBOiDOzD2v7zEp/BPxAlHT8RZPIkQgMhdLRxUeJegWPCjBChdHFCZmW
sLUy9L/XX8qORxv3iuqwbUM/ze30qhWthh7ILZRH30MaJbYnjVTlgTbUr8/uNGa6chMvfcHFGiK7
9fnu+2qOLTdR0baZRbEeK78WSGwXnHZxE6rcVPaWQeWOWi7fuFSX4qvLzAAw2lMfu/vdZlY7VrFW
5JC4TQA2vT4Ksfbkr0qiUMiNFSMILnWl56CN2JmNB8sTp2AjUVmaa4Xf7c3tPb1cCyaShks096Ej
jNwY9k7Ij8uGEX0jUfa4fVvDOtZdXj+69UTtN4Gv8RbZyurhawiG8dSgJhAyMotGmX8kAR1vcZLF
5UDG4ZaHHN9r4S1iXUsyne/tRnG0zMKtt8Zl7HQoLBVA3R8njU7DmKDvHd/o85mQdoleoiePT5Nz
Xdk+Y3hrn8UhzuaZYQYZobMmHtsUKkTN8qmQ83ddX1PrMcYUoIpCb+R8xIqIYWptE4l/VJqVa0az
J+7rmsBKPulznVcjRnR/yAfBo2nDEwUWOm0cC0Ve6ayeUR4IWVmP9dTof19f2vkvVEtqBPfvf1vJ
BR2NtHyJXGyUHDYyNsn19qYuCfonmWs2rKR+aAba95ItUjIShCZlNTQOvOf9rgVlz6TWbP0YEfcG
NDUbB4PjLKL371IAY4rtKV+kE8hO4FzbTEn804xWEjgMQNrPGYEYwqiTZz10CeLQXb1YPuuoaw9D
7jIj7jrkqFP3XAKdfn0jUIO2dnCGhp4HgfrowEAsWK/N67KwNPxDwm3DIz/vA3DmJi4soPIQqnxM
D41mYSHChifIbkdVCiV1ShQPZ1wA2LBx5QGisEeVfycqmyfcw+t4jnAffRDMCR3DynoPeywkEn5v
uhTY3bv1cMJFsoCo12Ori0rDfTuehg98tIY6mwwPjbGBp/EDz2tRWOSWACg8KI2IeV9f5+XHROS2
ntkKfCFUTlB7os+dRoAGeKGttQg3rdx85Gb/C+LPgwfLo7X5K1XEi+HnSR8VdmxXa8cZiaNuGbKr
UWto3fGOCHqBY2YCtEV7ldn54zDDXygur3driSb2oxK30sGIUv2O5Tuhytv+y4yiohGxU0xeJE4P
I9QOABVXKFXHgkuHGPF3QX41Hf3soZGjDg4R6WclzYXRZj/S9g3Ny7Ja++cHyFJ2lrlxrgfhLVD5
rHDY8BkG7FPd5P3Ya6zKiONMk578x/5TMLXNurFVn9p6nG4owLn08aFZ7dHj0b4f7W0ECcayjCCi
0K47AcX1UW6JZjzXkEd48xGA0DxywklymrmlKBJ+gsZYUL6s2QfoRdg3l2i10R+38RpUlP7+HM7S
g/R9wAm8BNgchdDPIGMi67weJXkSVXH5zjudnJbb3rUWWnQMcQlCmGZkTfIqvA4lctvXrPOS6Rut
OzlUx43f7HWHqg394/z+D/JP6GIOKlqDpxaZmYhWFoVEjBtOnemcu0ZYTE/Pbx+oXFkkLj7l005T
f1lxpQ5jN2Fo/W/YjYnnZbMPiesr0SWg253GI3oCr3jCReQN0s2CrWptuoKF6xg5c+eyaTzJXeeT
cvBiFhshIPqBj4Y4YWI4QfjilGUazBVq+52bmp4nO1zaulEkWA9lhZHc4izDjejt004I21Rfh7SA
TAizOA9paHfLGQJ7wV40RGU69W+52LKkjcUEoqxROq4mgb6Rk2I6arDrx8a7467mqNIy7T66ZU+r
BJw3+bCBQvNX+sB7ITo6PZR1Zwm6jfVZgGoHQkGge9BGofRadMsQOFGPF7uEn/HohGtpEPpyVtfQ
9yXHFjp3VpO6DE62QrNfVJKxwtnw3EdDI9x1NTK59rbWFsVuYqhgKsSr2FdN7T1CFUZRrE+z2rPm
vqsZ2oupRtWwZkHUttYXJBJdT0USywIU0sTmlyyYlfbz8e8IDHYyjLfO8WRVMImpHHVdn/pXyRER
p4lxTC9PDvXGrWso7n1WX+iAOj9JP4Qx6Xi/YUDnXDvX0+6CxbTYg1QNsMGRjfUNypiTtZdUS9ZD
5q6Dro7CoFIUsrZOF+2LLC6AdDiYfNBGaCkJILNSXTEcjexRZQv74oPtQ1Lo7L4Llbb+x/NUcFha
D8IV4efOT8FZtLEyoAfqUKn2icusgloelNYGx5MdOiVGneKAzQBedO7hpz4haqou5Ax52eFu4GTs
YY2EX/BKseJQq+uisUgKsgq5Q2MDb7IDvgUicAV32kZfAkwlJCzrryATku+dZl+mJbadB8q1zaRH
OgvmbW/1LuIHYqjzH8VZhousb6olZ9bUxs/P7gBEXK4jLYbaeGUmMREjX943KmvhQmu5X7uqxLE5
1ILdeqRQyk8c4gEBMNo4KnVPYKsThpphWHS/dImfFyLiLqWZ+bg/qdVjb6cW6Gw9TNCLnC8zJmTl
TyIPeRGhbRSGFYqttm8cqz91Pd0odDQHi69mDk1C9E4QuBuKCyNrMTc/hVKswDxqU9SdIE9rgnW3
zGgwtU4HzWS+Mj/GwdilEPu00p+rICweTRZ49SGBXIXNHPRJEr2mdo4+mP7aswwvkHcNQk5zS3o0
1C6v+hVS/J4U/M6Qh+7gLrI8vkf2LHr3T1KPv8DsRkZnE8Xf0pQt4VdlyCpzBe5qdK6JM/NjY2qs
CSAVjNGJLjejeNxeaQdecPyyTpP90KFGj7hXt2aBvKIUc65fBkKg1/AE2v4b/hNNJKbeFCznxZlB
u6q2mkpB6U/i4clMF86L9HLAZuAwAlg39rqhDI73Pa4AqOVgaKkssOaHuR6/OBER8y+MQyi6ad8y
g+rJufI9glfApfE4TWWaXpGOdwUvkhET8TMFVipDljISwdDbH6K58SWvpfKQ2oYtZhDYdsGp0paU
KYnecWZtWkpX9XZTLBb4jgFu8FMFxYhXpT1fIaSf7GfKUAHoY8wnR9J4o79zER/71udIA8CZf5kZ
64yc7pJgSfUJQwdLme5P/wWlr7UtkV+H+5nLJeYxi/eC3P/6xNsn6/GzPPjZxJ26lDs61+V4dWS5
/uR4LtRSjnq5i3iY11FYugwNKUgETGX8mrNtzdp4y80DwEpANn16bdjKGt2tY9MjXyBl0OSXh8mB
6QnxsOL0QoqI0N9+oGPI9IYoYmddHxZX0OxXjxBjR7d+4rqS5QPmAZldEhIwlgE+mU+f8oKO3n6C
jYJRYrvf+/+GbvA5efYr3YN/ff7TbIWWN78/USG7tJZflANIjs+HHCLb+1cmTYmJhtWQis/fvDsf
qeWv/NKGieBAyD+LxLC41BDeq5ghUNo96YmHJpWkOAtnrXd4nzethEvzIx/iSNoyZhgWm1zD/ibJ
wXzVV2sjywFX0gVM3AMA/9PqbYw64Wr0qIFYHpl1NLbqkESEr9BSkJP+aO9u+2AinrKPUM6lx1m7
a9BRzCWZMHh2hbHNcqU1U22fNwaHU5PCtURiEsG2dcu+A0uosoVp4xJg8raBAo5nUxGnqGC/LGN5
t9vGDnvtQUcR/KVR4Pf2fnpkeHp/uokqCqhl3t2aIvBBNHc0mNnzjXPmxdaovCqTsiJsjVo9WAra
NOcKgABY2BEKPuEGZrUN6zDIpC08qt+HGurU2kj5MfmkCczvWV97p4uPQPrzva+W4vdNCMlTMqQm
isJ2owpWkefCj878wG5hysCkn5nFsno022yj/CX8y2f4O9iNaANCYd1zayZPOzMAp7KOpVdJGTVi
vthmwQrM2bkU5pbJBTV8CZeO/x5+AJgd7GG5bzD2FiQhrcUUev/eGIcmJgLfYHuLrbIX5YD4xBYW
OA38sXqkLjXLhWmngP4c0LfsGHs8uOGJybk5xf+bSJlcN4dEvnGgAsA0X+eHrBitkln+9wp+dEwl
RwC+yHp7svp9wVi39OVpjze86BSV/o0DXWDFeNZJekL2oKb8seco9/CQcZkX3G96C/PU+V1Z6rcZ
qBWPqMVlRewe7vY9Dw3yx/t1yQWiTOMJUlGHsjAy1BXQi7Hsc34Ua6ZflemWWUBCb78I+ZX0pv2N
nCmwegitTMY24zGtv/luu2MvZw1izm3Op7LKD0m7PSa3JrkjU2FBNBeTpSxEpbMLFBFpAapI/bVL
iBKaLIu9+p6+BY8DKduXDLR5PccG+LjzMhea9i6MQk9JIHeKZjZOQ8H9qL20srRDUGrHKP3YwvUc
xvNELvSm+3izHptJz8XSLOrm6KpBfdCNAk7cms6M9S1MSniLSJcA9w/R90bEwvO/ji29zbtLoXdh
l+XBXuM3eaLIT+AkOZY5NJSp6XH4IfLrKKeUpHRgsNlyOaQcs2osATiqvTfCa1gWnsfZ0Toy/qNU
+Urd4IKPLWviN07NbNxFHR7HcOa2Bj9qfYg1rbTvb95nyDl91ZSHj9FTJM++NbIO0/NdOcf+8Cah
nI7ZX+FFZKvVDCwnAB+hq9+0YPiCE+iQbm+N/Aq7jso65EQTA01ns03JOhvbcaVWBFRP1wATuIHn
swzm/XexSh4CW3AQIKDbTdKB3Dnk//bdLCxbCAAZwkBotBnp04FLg5CKpNg6PznZ4/ZaXjeIIe1Q
OzHT9JU6KitOOHrIq0iOzH4Pz7GbApAMO0ZY8EbRRm+lXZ2Bo6mUM5W3fEBUgoo7PPXwP8BWVC7e
odlZtuU7S45rCmNkgJyY1Yz5JVfv0Q5yEnRPVaARgkmNNcJXJ72nAN5JVWzBjQCICB9o9IbSfT8m
CVMnp+SII6+EsVO60s70NRckeH5i0RYpO1n8ooJjq4Pb/bPyp6LCZ+sEEK/wg+D2rByMGWeZS7s2
iwu6UGVgF8BjZj65bPZyfg5rq5FUn6MLsfZsXP+ykAuc0ETdXkDuXusv+4siAHw9TB9+RYZMAiY2
j00G1LbWNoboLB+kneB3f8Lb9cYRKYxJ4d5GmdfF60/b1GzFILTerPlDkkhOHsPTte4KCm8SijBB
Rty7lHdOAdjBf3CJ7Cvx8bAlL/87cvjKbi+ryrLg9UCpcjJDmeLZUjtOkMx8Uh2zIWBHgNnJwDH0
/YBHhXf9ZgEIqjZkgIoAHXnvn+prpQqgPUFuM9b3MGJvymEFdYxa+YGifaZyhw+jRRT6slkscLvi
ppXBImNS1bKEPXr0UwhzvHzPs4rOMTwp2kYD0zidl/MwE6Z4AvqrHKjCZJX9ggiHrrMaa08oDjdB
5C23UKQR0rO04LF4gIT16oGXGKt2lkiHwgpW4suRDjWA0QL3N6OgFgkqQqyKQLqA+Nv+rYqb9d1e
bzrNHEqbTr15uXPIMyrka5iqGkvaIIS/+zMn+J8g6RzU8tA8L7I2/xkxBgiZaG/mslfDjiUmT076
183sQbA8CPaJcEXwX2pblW43UCff/waMf5cHjCvyavkwXPxEqYR5+ar14OOCA/CRL6HD4z2+XiRr
3rRHj+3cuPj3MTxVL3FJTg8qYFMBZ8PSrU1rMcYpvbuqkaTUe8bLu6RUO4VivN1ycAwJujpooWWT
ztVTtV9ttt1uQquUHlAgQW867jFfdvillmzpq4cgpQ04PRFldDI/xatQsaoORrmfC/d5wpg6UPhf
RFnig16A+iYih2cCh45MNEy6hrKxzii9s4dgipgV64/imrWRWI58vMXF2Rq7ZmXUHX18eZHdoFG+
qFefeHk2eigJU5ga9CXP29NQtB/nem0OC7dMq7gG8IzKtod5DwalbaC6dHkHpewQiZAUdePc/oZA
+eQoIN6SE9sWSzCAFXPWWDt8i2Uzs7QSVEcvFq+ceJGQybGf4BFYgpAd7itIPQ9Cdvi8hPEymiBS
Ox/eaFHsao83CZ0Iu7L8pEE20X35O4EpLZOf2IU84uIFwG+IRZpuR9jOn3Ntb7CESsNShfex8p6i
UjiLMUMoi3IZkmpNsqsRZlp5oahiKkF8ll8z7rSi4u5WuZqzzPErMnPia7lofS2b/8vDGPp5VN5u
f1HelI+8YGHAJ1hLse+o3WStKrkrgKNosBrAhGQ6pYG3jy6123czu0LXcTuHcCMrYa4pjF2+sJRE
w7Eq4RNZLgjYIkT3RsD5dkGeHtLdZJsZADmZTXsRVhj6IzHj2eehnoZwQje13tfCTs5Jx2YtT/oB
ZMW82yPpEtaRnYUlODQ/PPQofMLHhi3JPHG4VPbmJJ8DSVmyllKEJO+tiE+OK6l3h6+Nh9bH6XH0
ZfttNLDM3B8+KzosZSNPS+2OWMIWRLX6qancJL3iamfyJpIMGcL161UmJkoNJrTPJvu3E+jzK7kh
Usv2DyQqp4d4nr3DVe0VrVp/j5WdMHi60Mai5xNMOEuZ/ZkzeMFg8EGGprQ38yH1L+2DK+z75yMF
+RMSRvCBsOS6Qa6Mxcrhh2juPcHDy5xWuDXjiWYPxgQOsW0Gqt2TktwPIih4rg8YKOE/L+kenlim
uJyzrmxI9Ld8oDwL05fN4kiNN7APbKsI74aDcI8elaOG5Zl2dQKqn4qOwGHXsgJrAoLIMylBZCaT
zbKJqXKgZusLUtDO19p7e0wWSpfUZewhcPpQH/d2RlnI+blep3QXYoo174Y4TeB3K2ysFCET0pLM
zhW5US8kcyWlO+/Qqwip7ITwS4r1s2QeDEK5nTBPipHC/nHPGHM42vQuCJqZ8XA6bgdcBf32E+sK
gtT9BobmzhM5MK+/Oyd0wMqXosHIHOEZGUZg667gpah31LdAy5vhXcyy+Wl8bQ3/vR5fOmq1l+O6
nN4tyRAV+k9b8KkXm5eZDUnI2fi1372WU19pac0s2GZy9cHB7rbO3sQpw6JXdMEJ4ouFdDwfzkX+
NcxJrKgRpN5IDVJclZBTXRBvOllRekIc2umj+xxEsBf26NKs9zZfgI72lRuE6J2b2GEyE6YJUCx0
bDEp8IuyH1/mMOd5IkuFaXF8Wht97SXWp2uoaklrzFubTgEGEyid9dosEjIWQAjJKaKR1XoZ46iW
LL/iLnHbwkhD0exlxTKpC1X0LrTL3Iqso8XL5Cg7u9hifCjcpLVm6iMcK71lit9kfBnwO3SAstP5
4JduAJ8cGfjgohzQSv+pfLFLCizNSHhavhUEiq/M9ydOPehR1BSt5iYq/zefytIvWJ6zJJLFc1na
D0tz2YxXyApM/pOr0Ztf5qpFChDO+tJLEbg9RuHuz4IGXPGCMF+UG6sO4/9Xw39u8kW89LLNVQWh
+xVl04z/l7RAKd9EkrL2y2ZuGdpHFMGbHNdtV4ZuMU/8nsidlv3iQJI99g1pK4lwsWTCsmyv9ZtC
sCF7Ov1smORuG6lgIJcLImDv+2NyOgsjGGT4Ks94PJ+vB0mtAekW1zw32v7BVYxyV6qIHfnCyy9n
LMOjeHf//vGJXyRgGuXo4g32+/pp2H1eWfR27NdL+UM9zapcEET4yvwxqk8hBGsOg/WkRm+yaLlU
/au24rQdjcvKE5PyzWwi3c10NHxRTdiwYfmaHf94ysGG9EVhnN00Ywl2tiyQzRf+b67/84yPp6xR
ZfdStpoQkECgXQzYRWdVmoDn1U2ECI1SKa3yPkCpitHx7ZPyLJq78amwNFT3spaQ3wsNdyHRqNZL
OjGY8NsJiyv87mfHD2HPIZTwPwRaUAUZ51pvgnD4b8xwo4bIE7h7mQN3reFo92yQnTVoe0RkCGDg
+WBmbUSrgpBly6txrgJmzT3ru1Irl40BhoLGxoHx45RVAEwsIBvX4qQoydQTjtQ4AxQVk0ibkIms
AIX/d8upGgva7SewtdqK6oNY8TzOm5FvwrmDJPMusf3lk89SjMiYA1WHlLShkO8XEMXt27Xv52r/
U90oQBkeMQFnRltACXEEBMfCcf5A7UdAlnIbbTjPw9GpllEY0BKJLsOaleZy43ffdCGF1KgV1uG3
nqUc5GSM5yRp7BK+1JjW7m5j5x8iRBqEs7s5UeQio+KB5s8rZiCHtNVpIFoDgXhz/uJ8LBOKNMyv
T0xd0evP9BXcfc0L/uOO1w2uFC959eZCa3hW3iY41quSkVSXV9yuJYyjBWnpIYJNXA2NI7V+ZZqx
qcuhGNTXHyHSpYNp2XIVMTSq6E7YAretAwAeu/nbUazGoqRUQRVQOLSiJPjgnTEw1wTJxw/Qd/zG
ZAHsQPDLr6efT4gsoTW9TkuAmnteUsGwNK9ZqOxWX37vfWTt2+MHM7gPyQXH/kl+fbp/L1Pnk1rV
+VacgsE19Z0aKARSCS8aKmjRcX8hJqeVSHbBpJzwtQ0eparq5UUyFJC/FE9+w/bT1KCDmI68QUOl
xYq9pn/n8xbjQKS+lgWIhHpNUpV5O4L59UbKV/Zyaf8y1kR6YZjRCEXKJYGveUt9aaJSgXP7ESW+
LzmSPpDfegK7PbQEeE9XOS4opli8SKwUCUL9BktkC08wijua+D8zNSIbV16UMZ+idguzEmaHQmUz
2jBl06i1ueQGrV4s7AGyK9n8Z/9MuY8a50BRhht/Zmec353WEDJRlsSAX16TVkqVlmIsiqTJDbga
0RTcImb/EfbMGIRwIIIXm6jt9OlXrdU54KW9XdRWj1EWWLKrEDkCxR/fAQ6yMdqu5woP8o3nH9FY
K2swiHJ+MJU7dti/WaDkQ0nz+zIuqWYdmWDUznTVcFiND5a7LnHGJjkEU64vM6hhisyto3RBORHk
i+/gWDtig6/gLtt6qW1TRlqEl8x+yRCsD8JPF7YJntfrdI79ygJcPCBAOfmyH/FcvNrhK6oG1ABX
CS3Hti7PMyr588SpbGSHR7mUXIipqcyeaT6AY3G/zbMLStozKoFbHoy4KB/UFNU27ezdGvhiU26U
jQw+LZ7FRVOUdila7Mbn2V8fXLJd8ETKSPOx3O4y2uuNDG2LhHSYaQCWRdkYHE2LX7PRJVFaDjjk
4cIQB9XhDFq8zGs2pZN0gsn3k/6fSYBLPWV0s8gfTQ5NVZwHWXQ1fYQdMko5/K33zkkVmVb9T8dQ
KfmRia9SXinAqJNny503T85VlbhJfEfddXjtlbWiWljaEXrhiSsBzZZyDUzmy4yq88x2YxerbTpe
+Za6yOcA+TEfA+LOkNFCoJ46aMLB25ri9HF759vXSIarE2iIKounF9sVCoQQ3698c6XiGdAG8GV4
H6Qqvzwlc2X6RJZfrgaAN8A+dXq7ETeIHnuTXdfnDXOm6WhRCcDWjFT4zkD0ADaDNXcgSJ2ePeC+
nGag/bwjSOzWN/YmeZpwRd+xmokOAO2xX7/ABq4AicTX9PoKiE1ER+PbLRK7TCN6sdLw+VHQFGeE
bqOexxW2ol4TnNikX7hR+tLhFPcdBNm6wYhlXcW1En2/zKbJQi8T8ycpa13fMVPIBABNyHel4WDt
v11aZqSpjqjUCS860dYqz2VSe9iWsXZFPprWgaCOGisBJGY3DbLGIZS9otwSmChYAbwfs6iVVOoG
s2AEmeSZpTLbGuCdBY9vNAkePguMc2xokyg10rpjNYqdIKNaAbDuZo4O1YiNzNuPb5nrsurKqbmY
T9hbrWEhQueHEPYNh6nZo18tA5Iu1NQgC4o1+f0cX8UPR+NjdXMwx9eraND5eAZrEL6aQSbYVpZC
q/rG2+xJOG6cWyNh29TFuG02qm9OqSYKmNlJiDZpD17xYwGChBzPwSiLu579alr1EdFEDl8905E5
ZiaYxHlb6ZFA8Bt55yQJ4pBGx+3Tek4SHv+fOsituF/6Clne2qo7EBYa2KkXbxBic0GOfk9V3F3E
w6txOkpCidhaAi37xtjAvUjjsIbg+g8B0KFJYRVY1c1QfUGOGkg3qEYXN1mDzrDg95gqw+BwrHQg
63r2U1C4rJEPRLCBBWGeOkzHA3AwYX2uLO2U85Ot+YAGt0LgdLJB/pljdQl+oFhccsGld4EVxjU1
InwCnHCXzVMv5ZdnFXg9ihL6YP76BwLqI3OEwsohJewJL34R85pIvh1W5RJM3PAdN9O7IViAm36j
a9CJZYISGoCzGMpRKzjHs/iyHq5ncBwukJpy38d7X7R72zchsuJK3nbouCylRMpM/Jc0Bv88cw3v
1aZkAah+u+NcsvRPtAGKfNcNBZztXG5KMobOjjZu+rSV2V98NmHFNq9kOqdsHK5cAcYZkmvm3mmj
0SvJtEhcRuaHQM6QvE+blnWeGxLwD7LLGHRw7b6AhPyd90xSzFLrQOHSfpuCZQqNk2lLi54CWj9w
C5LkMH5rhxSowLwiwB4Sy4T/hBlQERDHzW7mG7aQhq36zkA8xSjkvWPuAEEngwK6hXfjh6x4MHfX
4GX2Gnldd1UfxVpg3MXtxl8PoHlVFaV7/t4GkE4HK4h1rrjdTtyLguNDq+8ARV54H7Wckuiz1Hnp
agMQ7b026tLbHmvkedewVtpQuZPNCthE5lFjNwvafnA1/4xva9zNuAQ+NavvpkIBygEPVKL45ujW
V4k/4Isd6+PK1KmjoNmIdRNeGYgRDQCpY/l1+UlPAN7Mkglf9dddjIVGDhqvVCJ7Db10wBvgQ8GH
ki1khzIAw2eO4JB+Ghc7O3/Z9gMEvvT+ksjvvwF1xvfShEL/u3/LCH+9m+FeY8QhnJobXTSNXfmD
ZYao7o7HOxPQnvoK28yRZPAR9s4tyYG+oYQeVmA3GmRls+qfI/hpvMLrBXnPOu8AgG//yMjIfdO8
HqzOn9zktIPHPb2oqhKeow5rQMDlKnMZObWskSPzPBO23XEJCy0TUs0ETf47JIBZyXb3aAEjekwZ
t1fsjMxpeh86wRl0l43pcKq/SwEJ4zGqe8xfpboR7CjDcEO/8/9b3RejwzdKwrGXqMEfXe5vqJd+
rGnYz5gwD7YnrW/xLl2VjRmz2gAuKrtfWASUirzO0WJnUcJQptTY7aUx3+hyKPnryGrSa11TDxPS
tzrM/Q8GwqpJASa8078xpshBkXK2LYko9BCb7BXxEdtjZh7NxPiPTtiBknto6HPMsghKdN3BxKYk
kHH5rVHnrJgtwd9Mh1oocxSNcxJIVEylSmuZcx3q/qKGe7G9FvL+APGt48p1uRaeueM0nw1Gx+AM
yZuqPNm20REpXGDdy7CWNsBXb5aP0cHglBf9uryn5nS+acoUpxOi2CMXvj33OVOZHJ+DIkd58LqM
bI1U4vz6xZyV817ZB23v81WGt8SRztddnuPQ8aRGcCNZ4p5KFHA6MwxnY0yWangYNKFIE9a9z2hE
dZ2BZnGoA46iJXEJPVjm7jXjSY3pxUokOE+qLcBXJXCuC46cMhIiytTQ609WOePSy7HzefpJDv3Y
RWYA3l813OUGNYuhPhTYWs1apQ1+cZVGmXBkkeCgQic5ml9E26lOT48KKCZigGuAgst5DvR+7Dgn
t3rjcEIvmZO/GXUuLD+qu3niVApspOZOy6WPFOmBPQHL3NalRumvSHbmxbFcJLv4yMu4mL7PX48b
h/ded/l9W2UeHPPovvYzSOVennPpxk9UO/nLDYLO5ViAwKsP8sRVumCrcpJJnHQGV5ya0xD3/I2v
Q3ZfAMIA4elG3H7JobFtYKX7Bz5qWmfGjevf2joK43KmHToMCOMIVGZKQkalnfajKTDnhKZGlJGq
r5Nr2gL3A+Qq1boC8L6VsiPVShwaixO03VRAKwuTOtTHbTcX1VL2QfNrMspYCJWbwVGX8UMWHONs
IJULH9ouR8m3331m/1uU/uSZrIRf+lKzIC4GLeMTfcp9sG/qzX8g1VycHzw7jwFe2vGJ7Nkz/nmD
rIzEq9z0n6vfVVu6OZq1n0CSoaVCJuf/Fe2C+uB4GHjIas8t5GxNIz62M0mMXpwv8ezzHiVd363+
0nMU4VyLfoM4qD9q6wxb/Njmh1/222vwwufceUP5Lu4HxeSdGMraGTvuGS2UjHkQ95YFVRVJh2Oo
W0Z16LDqlcOswty6luAk1fyba93mvmvI3+UQsPHWTaL+MioIs0yGM8kdbNDWwSkyyzyLjabIq4+U
0O2B3gkVnz5aGMhdd6o27O9jo6U1XvzA5CHuxagg9b9Y+/jqLSxvNqLxmNSQ6uKNC9VFuzIFwNXb
aW9I+ZVcjGeu0n+++biev6t91A7v+VRvaoYQO99EG8Cw8b4rTEzXlbMGx2CBN5hButUlxteHZvka
2RLFwt0OPYv1a6shvfdOStvuVWy7qZuGifAdr4n+yXJV2Bu+Df2B5WIm7v8idXrFSyKWL+7fhn4w
LuSM2bJApxY8Du6q0Pridq7CBU+EHmp+u4aAL2dTz+rgqJmaIw0ZvXS5vgVocM8X+uCHAZXE41ck
uLw2LGiInFcAfGCCvQ3yTHSGAutZU2JRZ5K+BExfwrkzst09HFDRu3Ein9KM32sXRBM2H4owRA6Y
zzoGs1oVToJNjj+UnraneKq+YQcFO95JWdC87iKa3eeIJd3hHjGggD3+BDOrjiQ1e6MOMdzQqQDr
snTn+SiCmUqU/j3o1S7Wag+Qn9Y9I/C1t9a2mV3AenFGkqYpYsbZvx0lNXqE+Vq28EYHcCNVL+dt
vjI/wZEQOb4qdPKvpx61NHYA6u0iVS/kSmZA8HifRYfGIPTRqvo2W5geV9Ldi3c8GPCiMmlH2fTC
xU8x3hgDb08WyluwWL5c7Gm5ReVPOz27NrGnF6lz4tvKzd3nkIR7x5/JNlSRhmQ57PWqSuhS13tE
qghSYOprlgrlbDYpOI92ytgh5hmhxJiohrUz0m8QZ7Lns4qmDphvaY9VB+MJFeJVQ91pEWtoCnyn
yVcf8peO1mCeIr4DjMsrEPGb8f/HHjcZH/zotykuq5VvWhQtQPgI3mTp8Gva1Ko81MFpz0mnw3Sv
hC4gzHushAXruqRu8mgEkuG7qLqmVqiPeOKrMDR4aEdv599sezZFFGujjXenx71N4MYcxei26hdE
lL+aO4mncyMZLILJO72P06pMUqM9hJucshJ8l8/iGIcUDm7gutXYfrymliUURNzy7DTzdtJ0tQ8H
sPZwJzFhmVVPWOAMG/PkedYeovwSLcNQhEO6aqWqyhYP4jP+McWlrH2qPojV4EGymxN9AIpBuHNu
u1weuQ8ws73DvLZC455DzJSky7v4JEYLUVInTAm/HKWnW4gpEoKmEHWFo9m5vtW+nwZy52SorXBz
MWTruIbe/+xqciG45/HL8d4wBRTXztvk6Y01K46uD2K2PcrAmM+hGX/Kt0mxp+dfPg0yma1c3zjD
a8cpQ3EdpdowRH2wFkHdXxzign6D0gQBTgckS7Ng5ur6jVCfKYIzZwVm0Zzl0fV2GLPUjQBB2kcS
moKtZX0xoWLQJPhFIDXQ2LBfEzS/DcpYSLJytPyzHdAViCskb4GC2ENvGDSdqla6JA1z6tvA6K4O
opTl6DdZnnDFfqTjdBVBEnHwvPFXYYw+Gm4ehCgCmQ/LjMqzj0UmlCgohi8JSvpBWcOoH7yjhIW/
Ay/AddEQi3wgt4fU6OF1yieGtwn4BX6R+lhpHOhoR9L1uVV76A7bDfvuoegX+ObL4cMp8ZjGn0zU
72XpkTrfjrqw+t5uohTf+Sbw63dqlCAyxOspDai9ZXfkE1xsxxFyxX7oiviTcvU8AXAxJeJNxCSz
m7KYfg7SGB+qdjnle3WZ6XtE6vswDuuyRy4U35cqwZhX3zTzGixEEBSa9LGKydUFnk64A/psu1gM
CSJSKIMVzA6Lglw/0HQr2Ia5kGnPXlrMvEsLVz9gvPncHfizaWvk1Qbaj/5Yp1zQu59cBrXa5maS
XX3fT2V+lf/5f3mYYgkPKoIdBCbReafEAEDTaRDl1OH3X0c23MQeVhkcoKnAqx7cdXv68yO9rrGn
KFl95QUQY63nYFkvN1ELK87zB9D6HaRK3HEP3V6vkseAfYMCoy64GN1OyiPYBvd+GIMP/mIcPUQ0
k9JJn7Q1pcYDp2ioVIO6F9caNjnCGe5RuMuzjTx/FvAjYYeDr/V3gRSR4Uv8ijSVF3DOIZBr5R7F
O8R113zdGlumrJ5x9LBxRsqQ0bRpI9sOMdKg/E9FnxAXAYcCxbTKZbdxGeOLXV/8+iMjukJNzJ0Z
N7Yy5qxv9WNtEpaVsDqV4nUluf1It5C5+szNdLOUoP70odvYFF+w3UKrTfeNpo+CRGy8vP+jltKR
PTJadBTjOcShz0FQy9/XWh/eNBhnydhYCtum/I5k2kfquWd5D6G0o++FC3B31vZcDkpiB2SJYbCb
sbkphBZfAv6bFwBmzzY0/0LPTWf4HPoKrX9e1OM3pr7A1VJVj71rq0Ve9QjPqKljeg7rlVwq2+q8
mT2iGwW+/7VVf8FphQHf4gy/aZ2/4uhJPXkjM9ZzU/Q05PloLR6CjzP/BpcSI94VHVlGWQcNDY6u
H/m0+6d/NUY1+uTeFUyAXMj4rXedexakaygCyxRG6zF4a9FFSpTDSSoCTVXK32bNbcUGKe/9Ei3x
h/uQOIBA9QKC081ZpDKgUYq0pvEbRgyUUarS+CGWokCE11GtBowoFLYr6G6COWgugyshwdMzZ0Xx
qUaUSND71/xJnELBQHoL4NJ+UQ5bBlu/yVGQQqQOMM+qZqCYIOjWIsWt6GH5qvvtC6F8Z5Sh62kT
zPgJAD9ijXPyGVVAFauLOSI6wRwA4qF3Eti9aW6AxikRi3AOTZp5vMPDltT1UDNwrH+YKlipaqjz
UIeJvf8Kg3BbTAcYDMqbPfrGnsJ7LUaeA7pA+/08HkkanGRcu05q62q2ZkAwKAKiGTpHSQNdhb78
LOUlcMuoCCf0EfqPXKfWElAbO5WgThrdvOF+B+XC5mIy8fARj7+lUqQEX+MvEUZVI8hHaJsNTNWI
xsq7M5CFeI2iMNT0tNHeMbTQTAL3BemToLUWaC/JpQIDOKrL+x3urrMkcUgHf6q051WOi9bR/lGk
/7A0SCSuFw8f3umgejJiFx3q7MdLSMSZ7H4gK0YmciI4PdmD6WrdlKWA3Zv7RFb3pbiejge1WYMk
jZLUqBbPDeY9KP4kNq6PiZ3S4eLHQE44SHG1bk9CKTVaoKaS3C72kc+8f+RZ6x23Uuv0JWU82FcM
ixA3Z/OheEFM5IAvwVDAEa9ZiY9l8OmOhZexbawfkolFedrU2zasOI7VVE82ozzTEMxaoYGO9HEY
O3QzbJLrXXZ8oXAiqn8sx8OQKKJso1dIz5T++2KfMOEEt5j3Ew5bh2279dR772qB0LHtaN1YBn4E
IZcL7ApzsZThBkWknUfm/v/Ef9RtZH1JkDrRcERJPhoAnOglHKD+m5GfB6cFkNyhI0yBx1ZETg8x
1C0euW60E2FWzQoE/hAa8oegMzABGaGGpbgL3OL8rtyOBBLOrbdazQu2XUVdPpznsLGHUJHxlT/B
GvylBtNM+q/iIuwHGYHBgOSShcxv9TwnxwT/FUbePOrsLPbTkFnNwpPFjJUPVjaOupmg7Oy3SFqA
JBTybEPqtRcFW2lc7U8wWmMlqVbexVp4fKoi402FkjoCIFtDDSMpiUFZr7RPPUDDYv6wZOkAR9bB
lIA/Wyn7Y51eyWCvTV2dsmrrAtPRIciUA9T38UQiMey3RRoWqM3PApRR3Vj3HjzmeW/Yb2Oc4m9l
w97TGAdDoX4Xq+OVNgpppXLeZcNj22fINdSUwan0FxtBg9XSj2gEM34/j0HB6ScdvHjOq9iA0saW
8i48Wz0pNqbrEw4Ev0T09mUddEYzlj4nUd8hOaN30EMZucP1k+A44TZBLH0LpGTsxC16NnquvBxH
tPbfS47torCD8vxJ4vNWrB0YenC/W716b2eVPz2nO+3wJGkCKNiblRzMfj2ACG1e7pCbv8Z3far2
u0iVZyXwpz8rwpZToKPeRZaB7bNUmitUBgHCS7bWniilyFZQhQNBOZJiy6+fVW8qVi/G4JwGMSHs
33zQ+nEVIiM38lU9b1qvrtf0kUBe+tVxwgvFLnFsOMuZMPrTyUldIsATGkb60AS+VFlck8u1kWJf
u0w7CaNrCxroJv/zt1A0MZj+bD3I7zgIWfmyRT2QQlchjTWZk7Y8Ozau2VqgAiEJNmr6eLF10XaM
RBMu+5dPXZsJoIFYacSwjzPIrDe8kIETabxz48cgeDI6Pehc9e/Se8qrJh+RWCw2g9uYsRWhK17p
rVywV4+gtKXQvGLfWOAacYqYy7ZK72qMEkefQAyGvXBz1jaNExDEuJLyl8TCbGpToBS70L0g8E9t
9s7t+dHGTU534IQ4UVLy7VPxkz2hRO4GWV1x3qvPC04aAsBGOaWK6krVMpVVEZAHUQw51E89Jk3Y
ZME3S/MbKuMGK9r9RT9KvH7RUYslbBKaGKadXZfo/TXRik/P+B5ae1WUw50cC9U4UU7mZ2ysKZt4
MVe3c6FwID9JXF2ASfXhjV/ru7symcsAxTiU6ZMOh0oE/0AWRFqfJ1lhgDhGqQ4SbEyzsQom8Tfq
Lq8Iv5UGywD/bR1Psl5iWe3RZBKEavJ2uV3QRYU9DPPeHLPRQYJcFy0eLZOQ7CAobAXVClJdUEgo
iDfbAHhzwy8v0eoQoiv6HDzJqR9Hf8e4ykSIvExvEvrkvTBiQgE3WrGyKytiH0GsQW6z0jpKsn8S
UflL4dt9WABVIpG5ucdVplFg/DtYNFCc10yMsYsBrM2ByDJLu/JT2O8bMJ4NWK8bOLUONmkXQ5mL
WqbdRuCGceCEQLwRrmb9cRuu5GRIsacp+xK1y4Ejfu1ag2l4fa1lf0hfcy6g+8xiI/U/ssEsMV+p
9npidjh5BWSFrkLP7kBQcWbccMXgokeLXFvGbJcGadrWxo/vpwSHaaQaxG+kq0mGvi/T8Rj6xf41
iQyyhnX5/O8MoMALXZw2yir17/+NqfesIZBoqaF7Nv2Tuk52dOB9vVjUWxATBp7jfCqr+XkIEFAG
478uiL2lQ9h30XX3DEWlReXMDbc4Tl2PG7i/Cekgg1N43fpZjqISvRv5mY3AQigwjonykD1sinvl
AiL+CRN1rnccdzoS93FQkDeL6QvO+l5urZyvacipf6CbkDe4yP77W+DpCQMWyU1jEClfJuPxDJMa
CX9rhJJ1llGn+cNjUDcGBL/DDuTogNP/thMy8lYcJmaAUBf3ve0cviK1PU3jeNHE2xkLb7mrjuQR
yol4D1HfkO3QloqQszgPJq6PC9T1sb4w6amn2KQWyXaOPJHwl2Rsd2sZeTe68xMKr9NovnmlAGBs
hth4ZybPj2f2ThafoPQZv3GHjT1PYhP1WIdYuLM1byznF+/0v1X0mLRbxgLU8BfaFLDjpxZOebIX
i2hz0jFFt/QlRNOTI/rIfvVV3bB4haUe1+8L4a6rTzEdzOXj0IvFllVCGfUBNk1HeSVj6Sc4/mXM
zzFr3+teKewVtl1ZDYzwZvsnM6OUD1JTDEbBvr+IOtfA2UJeZxnSdRnukq4iQ58fvlIfigXRFwCb
1qjZgx3Nu68ZDGbK7GGHcwjAiVkhQ1Ow2q65+O83vtNWbGFpQ5s4QgnWVfrwh1Gzb/AKm10FmRt6
LbxhCMYY0/zz3+xsslhlXsKgwbpT6AJoKkrpmRn3ekCnvnmlZWsOx8Kw84S2oFEr530civWlJmTY
7twcxmprCWkB/47w5lHZfB0EqHwxVrFrZxJBtZOIpOM0xyUVWVt6xOg5NWX96b2kP8wNfLF69+64
dc7lD2cTD7A84CGpsVic5Gg/SxQrdsFzg1D2BcKNeV2xUoxrfvu14Cnnn0RLikcXptNMtZ6HpVoQ
BL4pAloREe9TZAhGPbhN7YWBonbHD87tJ7ScPNwK1wb3cZEoHXGTiULUOFK1JOU0AZ2/VTHqBbCc
x7i/GKpZv4ksnrRrJawhyBhUHe6IjG64Vtaiuaj/QXsugILUqaur83N7PC+YFwyUsLBokvQyrGll
dVR3QlSiCf249ckMFI4rN+gGpD3v2e6fgjDZ1qOUvkFu7qbw/oN3VQ+u5PZgu/AjFVN99rJU3u2F
mOxNfISZD8L/hdbEqDuwSwsELn+QS2B4zpenna5zr3xlTezvxhkeTeEDtb47iL9Kf9X8wFOHPMw8
Zq5oFFcwywu3EV+wIFmjWlzvB5hUH+3Yb0xpTLh7B5fxFqVEsn9x3ZnFG1ftrGxqLZ3zZQ9tWFvr
LSb0ciS8Syki7aYbLei9Cd1Z+u4DPAUz2kqz3/PssmJUqYRYkd2Sjk4btMx73FUNu2ThV7izwLnV
VkyqMA3Losjz1ju7MmrIl4I0nsMVniL0taM2uiEnwMhdd/3V9LHahI7P3IqF80ySiFEnLdigSHmV
CmwF8l5mWz5JF2CgumazohZcnjEM/DsS/jx1SdF7Dt1FP27nGyoLowmSHlUmSb3HvvjlM84augtN
Nb5QPPnz7msb2Z8i+IqKGJp9HXrS16ch725nlg8hxkPpnerXTrJr2rXGB+VOi2SBa7La9dNLlyHG
xnhJm7ljornQ+Fv/RxC1V4ph8JaxiZ2xJukccD4dRqhjjidGUn3Yns/nFvaYXVh225vJUViW5XKV
aoWDuxG37XSdrEmPKHb6MM2pYwYaEXC0TCb3oKwv95Xy2nc85Pa2Kg+kdVveTF0WzuxKIPC8Bbgo
Lggc2pFwO0W4yKBdLfvMe8Dl1zt3N1BrgIS6dfGePfGD/Z4GH+OHUV7wnPN2cHQsgUEx6MNMfxqS
Sl0sMawmER/sysY/CS7VL3L/LiyWqcsZtcTX/MlsrpHgvmfeTFUi1WXLC8nkYk28xtSYkhWHF8Qo
j90v1+NdoFiAikBbu8Ni6PkxbOtncLj70HAnos8GhztI5a5BmNokpT+J5ogP5x3i6tuwetRKya/U
XwcEKiNhMTta6MTdTEe6j1VTeO4JD87Yk+gBTTXYrCU8ZtzrEt/jDvk4Akz2bE9YnifhUCXen8WD
lZkMgmwG5luj3LQH8M/ynVPWH3WOZovvHXHTZL+tp7+ItoZMqzdzi5OrKebvftw0rvRV/g7hdFNg
1EcMZTuFbwfLUq3T4ZxNFOICOHVMSXsxdm2d53+EgExrYzkTHP8Z4u/h754N5ocFIqAyLzJEJSKn
RK+E2H8EeK7JNpNLkuXYUEs8qE5L83ih/2Vs/fq5qk79JkZ3xFKJFO+TYgNpx4WnIsw3Bh4fWjEz
Gty4B+0aGCzMZBPcNCbw/vSFR+uy793q9zUnDQ9bLl5o2mtFBAOloH3NrmPY9e7kyGTg0Tt6ZmGc
8GI6ivPTx+rbQNkKYyxV+fVFiW/MJptKvyNLF+Xis0FaYzQFGBl0EbpZgU9LriTrgdYgcA0eR5s5
8lPLhBS+jOKjPgaCpcqSiel3Sgqxgi9AbN9n+lbytawz9q8WAoNqUwRHQGd+HJM6lKLx3WxVWlcp
mw0BBJzC1BFAAHONw9TKVSCRsnC5s/Ztr8xTWOKtyV6HMQjIterLPbapjOfoDJmNnwIdP4G4Sxf7
1toyBo9LO/HA6XYXKYHrP+RWRUJ0YUYxLizyGsR0G4NWdpOLCAaONFbw8HuOFqkSJovaSeHS+aXj
/GByIXVZT0eyknbRD07jj/AJG7OiuuQ7wSmGujQBRhAmF/O5EtN/Ajvq5+8w4ccBzdMTGLwZSrCC
yZeOH0EH0M9pIJg9Pmgps3FtJz3CmfDNQ6TTgtSQJ5HpFzeruR7oMQhqZFIo3ip2j6uVA5KuWRGW
WzWEgN9X7VHElsarfXJwVf0QTEHB6iud9uioTLVPLFT722NJeCw4+U8VpO6XjFmNyEEXth37CEWG
yN8I0Wp8v3sVmFsfa0xGyFmh2Jub+dxkADOpZ2wg5JV8xIE1wxYXntO0QRXyry39gJNGG1kC2CPf
tSs3O8YOrxKDSdFZJhmaikbH6tJ96JVG3gLr95MUkICnM6QIxUAEf0G6xpjg7ygcK2qQC4j/3a5J
qf0U88Z6HXYbTHkvRc7NeqhalK2gRsUxabELXcA5rZb3wx3xZOm8rMx70G6Vs0J+zix3APfI+G68
zx0NvzAhXtXt/z8gfPLEi4W7g9DAo6xoEjb6dCYnDQ30CCMBM43aSeJJapLKYU7hFiLwu/nEyfJJ
b5MClQNqAUIMKT82grLISuhcCNvwQjiC0J+nW+AdFag4zzSOOGnAJ5JfIVRzIqm2Ir+rcG8up8LO
adm9Ezw6X/V5TI3evIqq/QZAQfm6rHJrtjp6St9B/JTZUvdAB7WfMmJLGXKl5THCwIjUNUSp1A1m
dQcWcCJdCWceGKT2AjHgXxUW6GzrbasHj42340kNvwuqxuijQKHYSisauTeklGKFNlQxHVfKcSF3
kvzj+4E8OWxnwkoT61OLZco2rJ28/got9UexCZKlBP1p8JOeeSNl1jGLrnO52sRrKGs2toRsLkko
+VHRkYtboiy49nZA7ly5kWHr0MBS8ebPWTj1mBQDETYDnV0hGQfOeCc2BL46Vu7PmtMZn5+h26Fu
HUg+U4RuHLy3kTk08tgqaVyzwQSFQE745mBjwnx+VeMDotH9jZ6JmVmHjNQ0rORX8RQiHfrR+1bz
4YjXoBC0Co+5eTx0TwVvl9+cMA7Tvnc3KhEYoKzYG+djJzuku/4gPM545QfDdjYR7ZyGf6NIbzhu
fVTshFaF/oq8PVbB+R29m+fc7vCo8qe1LppmdM0rR4EJ9PrqHBnnFT3amgdXPSS/wuyJkE6JZ3y+
KEXALEXTOXhDnYdELW95+Ey8WbRG/dg3NbqMOUDWgRlFBMDb/q0V+fC2d667xnjtfkGK0+Dlg58Y
DodC8q+uBZf7ISrnjXunch8XBe2o5+ET0dGDjUxF+/oaVZpT/wTdpEVU+16APvrCCa4LNBOn+F5O
cuN1C2A0h8dqO91rhDJ2ue0aCSNNThSLXncmJ2+wNE3HG14I7wHgef7/mqZ+9FVIUwS0dwf6iBtC
s8KgKXSUyOpyKti0kndlV07GggZCI6PjrZjVstXD6NjAu7GsedLsDB+O+36/e2yZKMcQTqjIanV5
CIEJ5Y0rHG677F9eCEmSoBnOdicQLX0pFbd5/phENs1SFtzuEiDxrqy0mx659ObGbmgG3gLfySBC
fFy6FGcTrJmCrwk4vxTY//0hDW8o7QmxJmHKTqeFlQDm3C7gKbPp0ABvFPQlbAbS5zWwxvomUmGT
lkFyTMDLI3IINe+rNYpuq/UojoiW6ByAauurkHGN3PPcqUwhd41GV9yStCOw7rKAEj/LLgwlqeKq
ozvts79Sra72+3YGCxWmZzUBm5JYi7g7mQJ1BpGBxG1/ArfNcZLxP8ckydRwHqj0o2RpaQUFseYZ
a0/C/yOsrbCiCm37r4Fy1BMpKhKn3F3qKM8O75H6UhCbt9Ep41/6nPpNsz0Q9NK2y4/O3CfAcfPu
UHsUIRVEf//eXTqvgY56wryJ4lXMtnwui/LRAjf9twS6IzBuorXYHZfcSmcfKnM/NEgVJ1kYG0k/
tk+f2wBqe3SSxVwVHMHHqnZNobSiQI4G8zu1zCCkp8d9rj4fq8fe7AMG64bipIxR8QUwnXXt3tXw
ndL9orMY8KBvyqZPRi3e/d5s+M0bKgWDoS+nI3V1aoQzDqO9whflR30JIkujMFRgn1TAQvbiHyk0
DHJ4Zju7bptKfzjdnUb662rBmLhWLQhcbehXKqIMtYOinYTs+sBoH0W5vy+i+QDT0yUVYmfdBYkC
xT3ZGWe4mXlgtJEvNG9JXyogYL0z7TLPZBJNB62VcbH9c7BVJVKdlbRFaVIybid9ULqKmtv5muLs
pDfj9BuWHTxx8ZgdBmqKbI5chzsivwkH0/dcz1wvpqFln61g1vlH5CkC2JTm8CZZ5fk7mbuIozHH
HRMQDnusWoHfWe7tHQv46m3hy0bnKwlKYgUUXUrbPcMD8c8nafCvLNmK3z9i5hjAeKkH2ymewYsM
x3R2BZhNDXCcr9+AROGntPPUqMNnXTCyXrXosPbD42U+PkvoNTxp65zWs7Cq4f5Nbfm8N0Fk+Aso
XPfNelnnH5ytcPXxX/hMjZ5GFyBFaD7vmNIQZ/TrFAHqy4NEZnuPPWd/GWdZ6FIMwNQYEwwM/TLU
I6mCnYPPVNIIXfYVTx4vt7awGdAgxfxSwX3jKHoounrQgoixraDD76sdSF/OhqHNuOnIeqxkNwFh
lp4+8J+uta8Yt9UQBFoFjxWHjafAXdO77BGgIdUQ9agYCNoLWhbgSnQ+rRqekgQ1XnbAeyrrrmag
tK7zAzoMFBTZod5dbo4B6fNk/YwT7bdQvGJ0f0VHYHWMB/+spxxhscRG/DXqi5CosQ3C4QZxq1ag
olZr1tSGqLaI0UjztlNRnyBVxYHmG4n5v0z1k/dnxFSp6r/zLUvKlxylYihjhZWQhdCqtftap+eE
W/WCeUQRjZJWVZgpxgYxlyUkPKlOztq7ZvsNNgAgT2USpeb1PuDqaCBQEUvfGjLhxhzBPP1591rP
dYgzW9c8NRwSWPZnNCorJjbujrqhv8W12l8BrKav/EASNIq0zvDffAOyFyAlUTfom1N5DzyW2EsC
tOhdvhHfeTDs8ozfhJqMoubi5q7H7wtsc0UO35Xr0eBJ9lFq5KA1E47bmw6Gn5Fh6zBQ6QfsC6fc
LsIJZ+lnnAEUXuFW/7GFsl+yJMbNG4NC/6ExD4Onv2bLVeVV5+G0n8nTXkywOtGFBFzNSzJGAOVL
dd/RXsgGaA67gzKVbOfVcUSHR4q7sc60CSS8ypiMbJx7HzNsUsrfZNczD2uVFD6wW11oiaINi/Vo
Up6tGTzXysZUsGHorOis9++nxByR0Arftv9nzuDGJK9/Y4YSJrTzDETHz2SdJvruPGH8SfC9zUa3
eZC5KCUJgDlRBl6gJ2WYa6FcVHtaWAT95Tn95G5l0P8OJC7UXSBAs+bn0pnTa5izbOEAUSvrL0oj
1Py8OOXBsJYQQHTwsuliI762RGxgzVLfr3MDKlP5sIsx6AxwOeHfnvhiqRNSPYEdhKft51zqC23G
mvYIxMgSQljEJAmfOO55E57ZJhvWdcvQ2m/4tj+rnmWubWhjx54F7yS0VOw/uSrUkSXNCz26OHMm
yvxRoFFNavNoCZJDcDbQk94O/c0kZXtxDFdXCW5CrE9+MfnZpMdwx2X2PT/pcbIBXH1bkewx3AKQ
4qZpfLOO6G50dv1d+6lElz+3QjYilygFzjch0nQlZgL0SiN2ujR/bLJ5Ogsl3y3w6tPhFVvyV3OQ
WzgOfe6tUfbYF8v0PCYgjt9BDGpiTkcDeIny0gpTg2tCD7QfepZzVF6y67BabI7PKQMmkVO/HUnm
f9levLpS21YICOR7fA/jVih1Aa63QcxuU3jjg7IoRP4As2GIvj5O25zhgYfjiSD2It6SkEDM10Oh
CyYOrPUNMiSFLCqGj6Dx0cJbsAsPlQAF3PhQk3+2+E5uX6jxOC9jZ7cMBJL30bIVBWV6qGSC1Gwa
LcoPpoYGkUKPT9S2nEYwI/RivgVfbFwyVkmiHRdegEcNHpE0bGYcHAmJ8DbeQUdwARtz5ymoxOFY
jEuiRF+DPUtqoT6RXdy6h3GVIUK7PhcYhobubDWcc2Zj7drFLOqaWeaEPhCUGLjt3kiZyZFqbjrB
hHhZVop8RkRAC0SHZSk7QOGsrPLF03jWYDWBMJleWqKKC2H05Xbsoh3cycyZvdl6a/SJQUF3sl/A
S6CKAclFhXMohbyrfRMfVDjOJGRUYnI+jHytXPFb12mwH0Xd2ZwEtbw18OYItuwZLS/A+xnZf6E2
nv75IYvUKJvVy8t4jDLGLvN0/tOrtoMr3ne1vFGZtba9QcbSA6xSBzV86aWHd3ZD0PZi5JQgeE3j
M/fDEbwTiy2+1XD2/bRR9LNTxSXtHsVloLO2IJRibElM5s5/76VVZBcF7xjR1AJNfN6Fst1IfGji
qmH8rdF6zmeAmfYZHLxqvdLf9/ZZPvH7kcX7tK0Cn5EW7JZQNq4zeR1jxPyAN3FVaRl+eni335N2
HTUU9BQ3qKTAacOKbAtLE8Q5FYHrBao8CZtKvSyADuYXYYXCZd0db5MtuMeGB/Ivh4eN8N5cpyF3
faYkOKWigRhJOYg319wq0mJeocqJ1enYlPBA6kJfgqUnx2nKFfFWbaj5w07HN+BV/s6Zvvc0SeZm
3NyPiDiIjqy89VI4yl9I6nUDeNIAsx28bLspxbfWVIszx4OvZLGC8DCK+FRXOOwPBVCK6pEwnB22
Zmi09iHz2F2KROsGHPlg4F3a5wjVlQz2QZeadQbli1EBRqGjUPUlhl4bC3PkxyGo+zJTLezb03uT
l5jwdqR4KgUD8aizJ6QF0EJbmfIhtKdrEiXcInGGKTzhLGJkOng2r6RCiEcoPFtuytVcUq9dTGd8
vDR2QpSx2poj3oT4GNiCjYk5IlEtj8lozuOZjUUP3kSI8bH8zVJG7CC3XLniBnUykB7Vl68PgMqL
ar5C3PqGfqjigbn6844IRZxNUjynzKKZ0mpsb+TihbW+XEsMvdXCRQw3LpMt8naVfF0OIaG29pcn
cST9vJzzpMZ/Hozb6LVpywOLRtINVnhO5DbmaiIwF5la0LFC40Y4M6RvFfVyNfRegDgL96ov2K2P
K6durNHZbDffXykmzBm2mFedNDgRPOcTi9/eF0Zhy12ngNz3mPuVudOJ5LJfWNgkptPvQmMsAxql
3/8UTYrqU15pKzL1tqEXL7pQLZXRZbDaqErVMM4zQlS8fqaJQHokF+Sq5yuMY6SsYgh1cPhyD66s
lVRZejhJJxixrfy8yAHXogH+nEKho+eHXdqDiz5Dpx/kBlHVQlgu+tDxkMKDPax9CWrg42qvAfST
9wqb34lkDOnqoZ14pPekzR+7ObdMh3I5Rzp/Z0hoqrTbvv5tPNQS5P4IAeT7v6v89XYjQNuM2YR8
t7+lIjAfYJd7MACn/5T2ovqUbRQFZQzSKzY+PyFIdHp9enmwjOrZfR9w1pYQ9Xn1+br7iVMux/w9
FqLclxzfYIkDH05FHvXQuzEpNt2FMmtaT9bWgDne7Izm8BFZ2h8BLxAbDuk4pugpu/DAlVt9oKK9
t4K2MKtLlTvDjxpFx8LG6DGujpNC8F0OIYV0Rn/kkYqA2Fbi4t2qJZSk8Jx3tPKuy3QbCf+WOeVk
CIY1I/2vdJFBbxXoSlFb6afpqWBJejJYPRnbnSzNYJOLp166eZ1g7gEleuf13ZNf5jVj8bb9IFCu
HZVw/SsSsDtNchrbatpIhxcHAERn3MVCmLSsDA+44vJN8wGMxM5EBwDiUOVqejhBJAWG47giutt8
LPIdaJey/2HA1nEt3Z2KGZMUrx1xdWH2uYd5I1p7bfPtxyHQpkrKrPSzZTKgJkGk8pPhN3kuKhlG
xfEKZKI299eox9JYKzK7WyGhednfB8GnQD50d8Ufu5O/gfHNkb1qdOzlbMLShUIpCEZPmnNvMcaW
qDK5tnkVBcutraEHBV53lqQClQ1rJTRxg6D9niyswpwRlgQxC2eb7Ih4aryc3Etdioe2jPiFHMut
yK5RcGZaeBdJYxyaRmIkImDtbbqFQLTItjUGqMC3CBImgj0POuXt+z+xQ/WAp44ulK3YEYPM13zw
Ll74R36++Go/N5vR9wbzSFvoAw9imLingtKgqaX7t8H2sXBJwdvq5/2vKCA3hQRB3D3hPIzAFdaD
9NQlSX6AqoLMmvjwINjcUpaUVSnfpNEtySlXyXiUSJUqSl6UI5eBaxYG1l9O8Y7rIUD5ocGkGlmt
emVCo0/p34hrmkLX6bcJregYT7L/qgeSq6ew4+Yq6slO+YDj6s+xja/eKnyxD6dbKNWqJqyaRsMk
fAjLhLsjL0HRBwD9Bn60SLb6NV4qwZ02lhcVi/WL/boUm/EsYRbzqhZ2CMfghq/inc0hv7N1OmgI
+1iZNFBVe/j7NB4OzWGXZaEOEQszYSFexyNlQSYW3MWjM/DXw1YduJjE87/DEY2qe+/3UcxzNxFL
wVf7znxuEwuwfRjZsFdxMgg0cqFkxxUjAqgWtT9YdmUC2ozI7zzD6qwAWoMi1VUM8RMB9P1uEq/o
2l6lN/lWINKFV3ax1TKPThrscroYZuKbQvlnVfuGD5SKAcYgUOhG61JzO1Vl9CXFsfjtZL/Vf0Wm
IafgLRpUpLHuaNDPfR21fJcKGV7tOrW74i1RpkrMBoCJdCKrccv9MAY8jyuL2YIy6se7xRNjhZnO
nVI3N8n/nQfCtjv/AbEfU/xokT/Gk++iRGmiR0PGNF/o8RKddjl+wGEYMh86ZafP+QgPpe3GjtS5
F/UNPcYKqJIAg7qXArUrMBMpRDb4f4V/DL3mBdn22wwjsvLguBALy/+UMAcjrqHCaTWx8RZQqST2
JiJWHGaoTztI7ist4K/uhYkDg3f5E4auGE5+NeU3jW3QpOWv5xX3gh6sy8fgSDHxqiBPIlNT7E6a
Xe0MG6hhIXga1AoALlATouiKvGhPof6nSQCJXJ85PkkEDZjZJXcfASDmGiFOeiVjwSxFokwM1OjN
cpstFTUHzMjmHvxehDw0sZ0BOG1b57aznqwUsFHz2bhPfkWK3sAOWTsl8KMa8HXdTPnNqIInDCEi
hAFwtb+XCR8aqsLFxhVd6sxblhQ7x2jmlK5x8xLi4XBQc19nYui7DW5NmChyt//WMbiGVF/Qr7A1
r6QCudUeef2sWI5eL58cso/0CZoEZLt6f5qH4b8DPtorN6ESxTy+LLvFEPaDHI9M7oSFReSF70q9
5QDjYuZTChdXDDNUA2t6UuvWo8pnK/vQTcbuLgpuxJ487jUu2puwuh8GqaaR7HuvmlltXM5x7yaJ
B77arFRMnbIAhzaV5R4EAPIVf+xPgbW7KG4hfslKTvu7tT/z7RLx/54o/VR5HEDbA0IC/irnQ5Mq
uS76L35sSaEovZYUer/J4cHYBSm7Ej1/5PSmhM25Rb4+TFJpA7fVeR/OpqFZ7Ulqai+GQWxfKXqy
076KWYiUx3qKmhiMn4tO8S/P43w7Y2NqAI9kgnSSQOMibTgmFTN/XUzvnpk3ya8jg7CWk4WWZ8EB
vPmzPzChv+Te8eE8XCT4/PZvz4X9HM/PCYjTTW0I5b3JuqSzj8UY738jyW5SKZmFrpURl8Qm5Bn9
T2viyOV0Gn7fLmEFh5OelqlBGhUDNSNkLmJZuhhXy7UuyjXH0mr1tivmBSFpKktTdOptK5ZHDxHL
9LEFkhn68NXttMmi6KX2J58qds0Pixe+9DgnacPSSk91b8sdzo4jJBeBph3Jx/GHeyrZ6TvenF1D
tFvbquRsgMw3Ce73sKxLonPJTxGSMKLXxOqxrc81WtOIfeKX942b+d8DPHKQqg3KwGZVFs67h5fS
0hsI1+lVx0v9ZWOhio5agj8RpeUNdYsKJFJIoFHvMmhpb9GK0S0WvbtZNDFN9W66Hud7cex6EdCt
6akBS5aVpzHWYmfuUWcR4AQqKkhHSYOGLCRT1CQZGmom4LtmgrvVg5M9MNnB4gbaxF3ciraWrpxf
yOch1duFL3zy8fjAq4vpO/DCKtQ++4JY5EehJ1Sm2gyfbzFcvuM54eBxDiB8C/3thfqUb47fKoZF
exF/7aGdasKRxq5njahjQB33O5tRMAyZmQ9xMkwEIdkUt5Za5liZI1SYhK06s1q+ONTPcF9aHafa
czUyw9eo5bSvruj6RsqpwDMgiuT6xB215yQNsSQCuYcdURi+nk/nZRqQbR0IDj1cOU7WAvm/eciY
VTQPympxYzzOsqzMj7S7JVOZBpXk85ihm4KgpxLFvSvGoZJUdaRQmvq0lgk+AoY2uvYMF0IXRXba
X9tvHHdIYe5fwBhyxmpJutPUndD3Wm5U86bJtL8IPNQyaE0GKfCuRb4r5QTRPjZSZiJY9Y7sWbjg
JPF24QPj/5EUPwrIZFg2ECJQb68LVtS+zeXsHygdXu8y2YkLMWi5j0Yw8xRtxElFv5QdYhQ2tHev
45ywLn3KJ6601OaOA+XdIg9tsR9UQABAp7g5VW4Bwd3wuOTv+V/UFLKqeb+MYzX8qAgU3zsmnXxd
fNCideZa0d6AJDL67bTqfsxmgrekt6Zchbp7ehcFlF1fACZU3YuWtKtzEDm2FK/Yq3XngqWn/es7
qFIOr/z8vVkk6JRZoVi31zf2FuvrUrTkCYK+0c6r/OWqjqFi8MIMZ/gBVwRm38ZEE6L5qWAGPuzV
oPIzVYqTsyaG6Mqp2CsUxeXYDLbbeq2uXz1JELwyl8X77ZT8vA+HFfvvGyBL96bkL9UDQfEknGD2
jqebgCpJ/9tcaPnKM8DxIE2TEJ56Jk8SNSB0RB4VrywwCMhknoaglGruZU9SbFHTxyYFdiuWZoeS
4lCY3NmdbdriUi0PN+uavCFD/z/EV5DKk7XE44mgINMY9xMW6tza1d9HSHgleEli9xcZfdlvhLST
eFYMr9kFRMlN+4kXRfiN/RsDtnMpzYkdQeqJe2IEMCTCOOfSvRKzC0VuSPwzu+R9kR7ALs/jbbaO
Evxw94YJWg/a+cAHQ8UpaRabes34Kn+On52tRHk3p7HGiQltWsyTIacgcBgF/UqR62tbJ747ea/j
1fC1Odgsos/VWN6iPGdFSaBEhrVzRlkTjW6EHS9yzDokw58jHpiDoi035DIRaW8j2GFQqVx0Sr6x
xfRvgiUcH3gW/4RUqBNSCEeV5W5hL76FdgmGCS89Ddua0rQVGBmgc2FTX239NC1KGuYRKwLEDYAn
OAAQNB982sllTtz6mcLIgSM9ydp43WgSKrNIjSK0Rkeq592DsT8P+6WXyLq0VNAUz93GAGR/z/+P
y63EHzLfF0s2SKYc8jElRcJyF9es5+qjHSrHfTdMbFpsTMbIMZLQuzSojMLp41Gw0lH59QA+am5U
8XWMqS77UY3SEMWHn2IDWd5SIiQ6f+RxXzUP38a28uoEBHVDaAzE4BXwxKIQQfDFcE7ywlHug6bl
4/Iri6+FWZCHp9tTdJBcqRfAW4yYbIzEkPdTca80Re1kC1vTAmSglDn0fMwRBidSSZ7X4BKUJYWw
teIBJ403Gd7g1lMnp7VKUIFgBp0FA4NKsdGIte9lXd20R8yC89Mc4UIi3I33+W6Cwf5IB+YxfRbl
QKHGPE6yDoRBPDHYJL+yA9iM+uXM91rxQGVm5cjD+JRZflibvJAq0AAjtIqYQgrJa6caxIHH/GT3
9QuyBrq0cb1Klo8DztWOxNjDBYWsEenO7YzMtjWN3kQ1GbMUoM1O752c0Rv3/O1rlk/IC4cjwORh
RmnTepserS7TpWoZzhZFpcTgaMwZhWAO0zecst7jK6yw6r0Vl35QF/aFNYjDukIZwSI5YFDf/IYm
URlsedxBxmlqV7jiv+rC3GRj/Vwou8YrkiW8k/OapZp7Fq/3o4RjTqAjNFY6BoEMsd1fPmGWA8s2
GSLhIaKTGJLxtgUP2pNIzyPV8GkkapMGFH2m+CCL8/AWfY1JABSKMc2n3N78QeoREy5aJRji8a36
vBXrNYBmHkfw2Va5GH+s9LBZETMzUpsgCw7+Ho9qvtb8sAdRhkX01MRrh3QMf/hDFz7T2cxGQGV2
y85en0r1r5P5QlXUv8TLKsyd75/SI3x/hJyeHV3EQJlRAo55uBYv5gpBRD8qmoc3gnftHYHx0zsZ
T9foGXlM0o8Gh6/gYZwtvdNxxa85lN7tH3xLk4KIJbkHlkd7gs/pL15fEfn5H72lJ1zBmJDcMZzv
3vl2W7cbdomsS31ajjdVzKTzjdZrlaYFYIDbMVFANgb+naudrEWQoOmVzXIA070JCI+6lOK9NKJg
z3MnGkSFqRO3++BM+7Ykyj5fI5jdNy8RA9h9bZvjf5bLxxy3hgqYrHFUxrIhXXMqYwfh+bLG71rA
zBHgw3w1bttG//tq14n6lbByAy2ZKNgzwZPPhbiiO/Yw+vfrW8HlUzhA12nYM+WhkuoNqT2rZWAD
Oflo34gcaL/YC5VRdg1iogcdMadIZYibZr+EpuRBemvnYAmMNTz9LNnQ/OctYipWiT3VOG0VQYTM
fvzYdezS/VdbR3zPFbz5HZqgYZ0WISCqdr+2pk3NcIviFyrZtreGOHHHm7LR/LfGASbqOAdNwSbV
Kf9GiNL1xbetR3XuFP19NPw2ibL2WlfMabnz4Y8s/sJSWD1Cf8ZT/p5MKQSccYzCGXWtQVOxUTG1
O678Z21KofecA4RvcnTg1o8865ZikfsszlskfPi2hQ9b0eR9Xh7MTupF5OC8S/L4ppfiwuZ5Vcgx
sBdbXJsQgwPMUzm9dkHokowGggufqHl5+YGHtHPd6ta6KO/zu/2B54IhVnb4jO2GWgd2XgMFYaCi
F80Fakp4vHUfIFhhT3mIC86z8B1fxLl12MCbVzNP2HR8cEfzHfB1M9aHrQMf03Nq+WSfS7fxOspJ
Fr7SuqPc/6W26W7I9GnqSjwx8kpS+0YNocOxh3ye/S1PtBzGX01vanRwY30IRBTN4adAcAxZSUVO
VDvvREukfrKT6oKrLLeT0P9e9/7H90a5kICusELnCoumFDS7io/ACVPg1ozMDAOabm91H4GOQZep
OQt9E+S3R8aOcHsu5vvHRCnn9LSpkLXMJXUgHXdyAbV5UhNewQWCTKfG9Dxq1+8OwMzN8UoDWE9w
pc5uVqVYxlzAi1Btdoq1GWbbE6yHDyjgMHtAuSVwzQG1wG/RfGxEn+Vu4Dmhr6QqQP05z2ziXPRW
sAmW1nyiBWjmMW5hNqO+0UpZUlBqubBeVEtCNzrULdpZaeMd+ZcQK2XWjEF9ad90XQTsWZQAHLaP
oDUv2ACOySQ5neN1BosI0OxMmJvy25ov7DWoDiBwR4sD/MZ1ilhHhsnMPrzV9on7lSyTMQvrgG3k
gBna6wcZinUEC6+aZ1DR9BTtvkdZWNvcQaWpq6NfO5xn1O1R1DcrQ3ivbcuc/K6aSeQF6fte908T
qhDYEJPGjkG+2LOTnaUOlMGYov+I9g1S3hftl15FQwpdbaHQJtVq69Wk8OC/PfHYaeR+Lhp4B3u9
HN2bh2UkfZHx0okoqviKFH3pWN5Kd2HZAFEIdtdLHDsZ7qVk9E4T4FzOtYwlbuiF3TKOmtVaAMd0
Hvgp5dKvZ1TRq1z0uwYI26ZL0x32rkrQHiYvYwdT0Je+O2IQUM4tLLdez4+Tgmz4bqzdQuYkUMIM
DHNmz3ZKGfEnlPVMkxAWI4mFqwTN2o1kbD/lEJdQvDEyagdtynXcUyhDluQeX35qQXtrZlcDX3LT
Um/uDZpU64z1ii1QONQt/yR7CIHMHfsLdBhOQK1tAoGeCjb8kf7mXhv7WXPhKkbq3D2cyeibZeem
ZnSWLBId+m2a20BgvfBzn31s66cx8XNVU8LNJCytrMR3Hnq/vbPlMzOgjYgW8PcWfIb1mMtU/IMu
Yg9pKDICGcybaEXZM0Xliw55v7H9JQ606k1M/r+mIr87KiSw+8TUbH2ukI/iP7tPNhrJGblVSk+w
iunScStz85ZNC20qoZoz3KpA/9n26YjkzYc8w6tO7wn4h/zddPj4MF6WuLfwaR4RxlPulujmCmUX
uujjHiH4mDcjuWq6LTnm2kP0YEQvd5CVxnwxSh74W2AV0/vjl+k40YWJ9+Ii3H3XA1QHdgsHiv6N
ewkcFh5wmgSAr/a4vmVK74sN1+9cnjQFScPkJDduyGmSUAwH6LvpfZY9PgcHVlVUTp7KSHJXeyK/
vyuXrbeW1eerAQT6elwv5RLzMnu6cCGP1OXPvdUiYB88jzwAUtUMCjlwSSClVOJuBH0zndPeq54h
gmAE6jPK6gWalbnFk/vKMdKWMTIkPjCg6FSPUKHlRA7ge/fpDrcNLiPia9VW/lRIREWpk0oqjVaB
24inTzkgLgJTEwHO6iP6e8UQE2g0VGL7T+GUjqSMCNT87GFkGhiiOmvavZaM4ev5cD4zNW7tACmF
g1T3PDm5lfQtKPTzonHrUFdgJkOZ5z5YlRNY58PeypmokIsJC9w7e+Glsc/Id3GAV7VRq9Ab0ZGV
qctys2pGs9vwX+GpoNYdoLCSKTPf3yyhtpx3Ml6KEq0x9570rgBv5nh/ILWXHsb8sF4j8wVDR8ZC
wyS6mrLZ/o2l+hlmJrH+rKpFRzX8pb9jtRZE7c0oi6vbGHCmf3hYD0cc9JWrc95aNS9NU8H4LVOS
pVAPqrp5pDSrq1nhfUH0rOE3ALx4ZGJtPHgp2FM3ooocPd6NCXsCKuOg2zDMmsLYOinVuTyUPHBT
vyFfX7O8c6DeSU8QnF/xDhYS7bA4k7j6pR21xRo2vqiwljMiMyDjDCbBzGwcHw3mRK20CjZOAhV/
MdzmvxRXUqjFdlATJOcUq3XqmF7gqsvjo0OodlOACToJEJqSqCmVvcwcSpqBeSQqWLzsk7snFqze
vOEXXLpv0Zscd6xz94+Gt0iqPo02VL8KEnu+WFQA2pvt+UowuC3GEtbf5veDSaJc3RWRq86zoWB2
QfRBcHIABJUEJEpMD9GQwlfKiiBvtOwuKDUy7ypRHh6EkMVoVI+O6VWTCiUXV/vJrrY+F7xDkOI5
/W4xNM33pKF/6QokCs+/q6yARaTqYX1P85lBmgoizizE4gg0sayCbvKKgdQOwptFNqF6uQf+75XB
hl5/q3dzFrhPp40oC/MOrxUXxnvPwunZYNpf1STUsnJK+Zr1/7dYln1gf3esKmaP/9w1fMRwrSPL
AwWXutWqSe3PRTmuAQEqCTyas11AvUHRAjNP3jtmrRLFT4RcLFzz0RJ7HE1WmMqffXxtFgGmDK7u
tF8zNpkekhS8lu0E7tcZp6FO4zej8AANlWjGcEFBSD6R+lDwLI/TjkCiUwWLgODCO6tp85CxzM00
JZbHrUmetKnqPGCCrSu7YH0ZXHwd1D1EaOviEUIpySjqpsnsoKP38CvxRLGKiF/LiXrMtlKQ5tBZ
Sz31vY5qVasJOc4CJqKn45rmArH2jDNEZ0oOgEzKPx1qWtMcvO82/ktXhi+uyghA6L5xH64ArHlp
HjX1h0YgE/lrkGy0IuBUm6n3zgIrr+Uk3P1O6qSlw863yovRlW9GTqKdRK0J98MjM5KhlhrZ+Y7c
MqYna7WEPVMBrJoxFS3gilYXYL2VUWuqKYqHZpi9tbcNvmKgHo04oFG+eU4cKyqqUxrJ2etLiWTj
MQ7c1s2Dtq8UlzPBWb7GR5y4Jztg0SZnUlqfOVFV0j6z+IK7mDeQ+M80CRd2ZQmASF9x8UyKvVxE
+u2kcsmFvq3dz4YQvq7RTC4PfT7IlisvPqOD9gmSwnWqQ4I86C/Xe21Rg1UpXyU74kC48XM8L7R+
aHP7HmZWURtq9218XskArkPlxedwEhYl55/5sWACz/00w7DniTFxWwDdgVSGJyHtvqSN9Zso2z5d
/G3oqVkVHAxKwXv2EyyCy0IwQn66+t1X6Zi26K2zNwRN3yERJyN5o58qceTpeZe1QbmgoarpFouU
d9sCWfPzE8iubRJJy+aEX8YsG2QrM22f3qZTC3wpt9KqRd+zdfI7XaFXKqoaZDaT2Fw+fusZHDdf
a8mAFLfNLvxUlk9i39UiASfXlsyQsEsKDE5W17OYZ2/0t6fXZcdDuY+97bg4+ex5NMJf9Dgf+bhD
7maW8j6b+HQ/Us0aMhKT2Sj5gHiyKbOs0ish0DCCdyoG5yKxmFrqwl3YOMICzgT97LGLb2ZILxWf
gX1DinsqKb4MS8ZckGVUeYttI6/Grav+9DflJZ/sRd9hSsYB1XvEFF5AuVlYgs1aC4MYYlpVTuWi
0an9jFXAnZPBu34ZV22fZZVW2P5507Lil2n/vBFr8cwI5rcXcgPs6gH2OtswpZvf+J5UJtOxgB/7
LdAsxXXEO4ydp/P43Cbp3TXMw/m8hy3BEwJZo/85nXAl0KiuiJiWEh8dVt3cuKWrqDTYAM4XfuoH
UTbB9GqGg4y0sfKinRpGrH3KpiSFShW09jCrOpS9U0XIkYV9/P7zoFf+WFfOaJuOCqvF5Iop7Vf7
grCGarKBLw89C6HysTEMSHSyZ4f36AaXkeM3fwmKh5MBem1RVStNjjC24EoMjXW6PS/PQXURGAti
K4qEm1cVYxPARS4bOW1kob06KGpGltm7d2oFOPwHHV2zDD6+x++9smc8jJYOjhjybwoNdmn7sMds
W5cR4nRFSG9U+njlG4cWbyKnJaGkKh1MsDYsAFjGAFWfZnI3Kh7s8XvJwm9FIK1G7l8rXt2icYCk
vIRMWT1ZwZTmDIyAgaZ61a4UErcHnvE2VNYv2mRkXFnm/j9t7GNFylu/EYk2IwzxkukzfLpfn7vy
GE/P3LLwxlC5qQTxabxDWmfLOPbzM9h9DDR/IP1Nn7FznRuBY8IxEwj4wjqopUjzCUyAwdPesh1o
MVbRmce0lPtAkweHhkV2jzIAGi7/p469MHvQLkx015tPc/kxKuE1IktPSNmjf5uFJT4+kFd5svEJ
JnK+olu6hy8XcZgqpUzKH/ORuESQA1MWy46vWvRzxBjo+4pVMgKPn3+PKAIbWu8R4m8zXFuYjBqF
o5SUR4N/v8juRSTMHpQdZwQw8O1PzzSDXfQ9JCUejM89SY/vcDXOOXUSKHz82UGnCM45sDDxV7+9
2v31rsYYHNiSierBA9x4VNbiH65U4z7+JnSFAdSgnL/ZczbYsvyerGDBGLJewn997EgJ89A/FW0r
G321mfMA+MLMvrfoD3RLjRvlx9O5PbenMxbCK5g3SLvW0+Yzcfo0ut5mOuRZuKNEGj6U3N0dfA8P
Y/kNHhfldQ4biHNuK3uD2rGgZeOL2OVRjHXNE3xUk3OLetZlESUygeiE4y9t0uIHcdATBD5hp0ot
hQkPMzgbUndHm3f4IwjIHHzqLXsM4/b4VFKlidcQ3BA0//vUSJd0rtQgnN2UggbHRc7zp42u0yAp
VTpbq9qiOQLeVHd0rw5wL7NTglCf/hMkIP8V4Jco2GaXOsAM3VyHLBeEeGH6Z7kC0E82pQyl70lw
m0mahlM9Gr9WPOjZ9ZhtwdSQ3yPATu4hMU+fhQCTcTCWgHAC0RmZ06gfUEKh/pZISOjAbAG1KdzM
qlUSLxBAwXh9W5e4HHJV9QANtHfEw+WR/e/V3HaKIcBBa7HwDoIM/zKKZmRgCwvwL/LeeZRNgE+b
OupbOepfcSlXJpIVw/Mj2bd9BpC4BQeCX4ExsOA11u7pD0sWQjaoMpTd+kp27+g+q8GE7Ep3d3eK
XaH4ShXBIK8dsEyZpXis7yFkN8MyJUsl4nHWOQ0aMsWr75jb86/bPMbPY/qkjPCB3Hpqwp3I8mY7
ENz6bpHFH5RSpPkrKBWaBOxlLRFE9hQ5MZvRUMOyTR+eyiADdpI7/7k8BTYRkhEpacavHnPUNk62
wygJoi9dj5CH7Pzd0OxkqsAkwLwB65Uvt9hue5gmZM78fpCbraf7oOnznu9+8AgmQW3zZNg5XJHd
FdB6xo4jcuX9FaTO7dR2QqWEy88uq8z6cYyIWcF82r5Dt9Q/ylfBYl/FNGIyFZc8ppb9M7Lvi/6k
6JDCEIwYCtV7fKo+YpRcUNdUrR8q1at3bu0ftTH2e07Bm6V6/hxd0pMIGsrb9vUfigoTDa9GwJg/
d8dMEFQHkPd2Uw0HxD30ErZarxybtfG9reAJxq5auisRhdHq1Zi3AcHbyEacVgi1EdgFw3iX7qTz
T86czcYKqEclgsm/k1CAJUGK8sOUbYgeO1ysQJgVyRM4Tm4k9bLu4tO7FARN9hZ1FyxykeqOw4lt
IIqarKK/ww/+dcAOZYpCwNX82bG9tAAqOZpRhHmbQF07RWC9ztSQrXovEUqLDYYhSpDzZStzCklC
/WCM9pBj20qx057yJEzmwbCmP5zCLe8EpJaIESHX/Jz8B2hwa/e4mP7sAIpYKBE5WiRcZIlg40Vk
Apq0Mnx4x2HYNI39Bq/me8MBqYtAteJxhkFuBslRr+VJuOcRE4C8oT1asEmCyYgB21XdS5Wxcrxj
KIkCemeaipfJPkvNTJN21333vvaLJA3Dudx8ZT2ee7L8dUaqsgn9E2HcG3Vx1vvlfvX8iHvDhnDU
VH77G2Egrx427wdEbS6buvYhwy1vPxmaDcpHMRIpi6mA9levf8Gtzp+1VVnnBtfLZ91yqG8ugyAN
80vUO7ntHnLrXxIUi4npEIiH+Zvh8DL0xgUsoTQ4zAzkdX6YnTPTFsb5n5Pv4uQBVYiu+VPLY7Yo
g2uxmvZwq+gdBmlh/wWCnqs6iX6hYWt07tP1+v226iH+DSjAfBTlWwdosQkwAu+VhjDhEtpIJwmG
BGFAuKcdMTunekvs23G0FhL228HfUk/bPW35/a7V/4RYJiUrfY0I8F+UKLnJzevzDqifQnvS6fRM
0RdI6CPKdAseQaEThW3OMqRcmof6m5ml2HehYJv/9wONgkIuZrGRKB0jR3dMPWOMjzixNXa/Oyjc
8kzXnw+wyuyBL3nKvf3dSA7HD34WWqBjH8irVaw5GYa7qvS4EkgRb4ny+xemRqaO32kywn4rRhmN
vVkjM3O+FZZpJBxsgqUvVahtGHHjDXcExH0EsJzOKlwgxxguK5GU1Eq8OcYlDZCetRqZt9ta7NgK
ilcSbW6i2BJTTVazWauMvGXsm2ygSeINar2OW0Wv8ORgH7sXewlgw+6TPhRGPNGPDBnOAtfPfwJA
DnOahB4aNfcPenMNwes1wjn7+gEifhrvhK8QUDcf3TD6GSbioGp+AcOqiEyfve9cAGNQZW+C/noq
vljw2Xu7AnQGlPzOs5QUdS+3J+iEo7avjk+AiNvtWnQQHaSFcp2mAc8HuJdhX7mX8pIH7QW6NsNX
B5gsDUdswRpyf03y0R4GNUhW5YJ/Yipz+h3R3DOuiApG/jy83WgwNJE+U79Tl8bkL0sve53isqqg
cJiGDpZztdsR6t9870H60T/kwv+2yUTej+35yB/Ec6wQPutDwH6JOV7l6IQPZR/UsbLKaP25cMQL
Y1xCjeOrlrzDiXMYLzMrYloDtea0iUf1ZicvHhY+zAMzynFj7GEjdSBugOqnWtnaazkLi79fFWc8
V8YbzK0mnCGPAYZrXc0SQD52AIgjPThyoiLPFOVlWre0ZieZ/cwHWnh+Kx5OR5b5RPSkHzU2GYqa
5Ov10rWRWfWVH1V2lkI1RZ5r85a9wTW364BvXy932vmb8H5j0ZGpAL/NQIEov/9MEyW6nj2rVSDV
Nejm2bvsaErro4ZiWJ2IWuxbsLP5LHSSyKAwJGsToIzFSdB4rmRXDyIEI/UO68lmOkhABvhtXXNa
G/WVDKL5vM5HONP9qezFs8nF/JX+En53NmpxFKwu4FXoYGz9WSuADPigWSPSkhDyoXLKxNr9QyXc
+W6JCie57GWrDhNzZpojD5CblWdWA8zcWyu3vKAmPXLZJgXbaFfXE24/9wUG8YwzbXh/DXDUW6xt
hElUBuawpimul49Vx/gZnKdwhbHg9SSUVTFk/MMPCKTlX3feXTiswB3UYGfg2kV1M3aDGz74XbNI
OqnmInNdmiAwNxI/AjbHbVLZQhr11LcAswjo8iQBMG5l3lNrn4jKuSSW3t+ALXct5lH53WKg3JdQ
7LXq3+E9rqf/IKBcZhmDJfYufE8vpq0uY76opZ1IuAvG5pSJ5/v0l+wy3CWTdhSvhM/QhVTy6DZM
soptrumGqN+6yaRFuB0BJwncQc7XvEtHX/jg0Okd0ksD8EDwyUGT8WZ2awXOaAllUlzG2yu0qjBF
q+vqjb7T379UMWNL2HAkv2H+QRVYtQe4PkEzepbROs9zA4+Om7LRY+bLiBU8gQZ/tbHIRgcyUqd4
kSHTEuBE7P8wamI2h7U5qOo9nmg0Bq8gOjMRRw6Md7YFj5wS82eqaYM2y5kMdpxSYgorphESh3W0
Yp5d/QRa19/iwkNjQaouzgXYElktR7Md1plB4JbJGCgZpgz6pU0ZwtasQ6tnRPq3lGU42+00tA1I
Vfsc2aw8lLBer1vWxir+12IMwS7RZmYRltJwpo8vTdFu5Pl75mPdjGEa16nzlqqY92OM/7HaDZQ9
tfqnyq9Epd6PzwVaFWGOJkZ+e7fzsnC/qUubNc7z+AtErbuU1iMHjkDauses7vZH8IyqIIeLQ6dI
sJ5AGjUbHUjSFDkZG7Ch7XnhnGRZLXJaDp/0ZUkr4saZ+KDcmxaWYG67V7qjwDqEML7LGDqZy9Nt
QoxLFyUstwDHRZNXv6m8KfnpderdE9nFq5K9yq15uvQKnltCL3IJ/pjYP5H7H7v8kKkeQdhIhRSS
ZeDi7fzC9A2DmasKh3wtnTgE2EnY/hR+BOgkCWDJaF1dEdjpCwelVAocWUnookhwguXO2/rrC4DK
Qtgv3Jo3WBLCZkKQBOmyUsY3ZUl2mxI4ys44qhvQTorjj/k7bi657lQkaM8JsgxK5R+6Y9z/LfpE
od6axcGl2Sya/oxvlHixFkgKVVPiL4H9HKeF1oUhRNpFsOfUfTRBM5cRnqVM63qJKwfdRlLPpIYs
zjgaj+dNGeSt5FTdZtFNm99hPE33E7K3O4uxK18LTi6EWBLGutP66xlBoibczOaz1/0tljx2d+A/
uQyXjYQIiyeX8RTOJoEg97QYzIuwt/gjbq8jdNEvqcKFX619MVch02q640fd5FLKKFkOxd8NJ9jF
amVgJrQRvAyUjOwSXhT4X5W8v9s08xd11RroD1DeTDQbj8Yx6kXB6LKborZ0uwUOt14HG6wE0U1C
mA3ctqcceDqjQhY/icAw3SUh3g52d7WAC3417yNq1bIhAo0wcHCcl2fefae4lJSqona0TYuRquLv
VfDuPeTuYfgDQ1t/7fmqSeKqXcwklW4al9P4ruv5eNwp6u2X9ds8ab1yJM5DFwEWHYpDpB/M51mc
+qznoJBKiBlVnwzIUMEe/PQPTFCEt5XM/CmbX46BFs1cXu7m2xtKe9khog1d0J0R2TVQrvTb9zR3
xgb+hPlg351pF0Iv1i/jwPlRx59ejE8eB/nbNRtol7ESi/prDPjR78ddAQp46I4yMHR9tNGo67EH
ovQo5xEmJo0QkU8wxLFxGmuvnF8NZS2EVbrW1NYgXXLIjffyiRTd41yCOulu/c6bJWsqNUwQqS5o
LZTPyn+YNx1fLKS1Dmxy55K8Quc1lJxUkQ3tB+KMrgrRLKyfthViQpv3rkRJ+Yaaj9cStsiKsrZN
i8fjMuFdDAy2a9JJKEiZQzpiGdAZpmsSMEfQNxqsC7l5Hi6sqsJPsLOdKWYWcVNd5hs2Vcl5gCGb
Ln7OPpYepvR+RHPHzi13iUUuhA0tFpSo6UtAazzQIzrJDxpxIXzzc4LVLunT7Ptz9+ErcjJg3l9a
YCbxdcJ+xNkdWoWHnFGUq0/gFJPR7jNCbYuE6dJwx5zRwcRKkwhVPEkMepb8Wgj94i5Uy2P6IEbW
ReEhqS9yItypxJYaTVXx+h8hF2hy1fbDSZGOJSyEfPMsyCajBw9L6b9iSjd+rGnqsigx/DTmrHqB
MoPboxVOVWdcYNRw9aTudlCZVlpvSaVO1V1/yTkUEGJEl0FuQE3pIunominYGC7wCjgT4KqH3E4t
Sp6/5XB80td53AZTygIwNnrbTPgEpGCk17yL32kpEBgBzN4ExvaQtKSZr6nRy7sGUXBfjm3F0jjR
i4US/2EIZE+BqouQWrZcjUDevuQf+BvNeUZb9Rrj45JY5evDckyg+PmX5pV+4O++kL8c5Gz6pDR3
9EnXS4kXXa/59G80waH3WUDzrzWFbxh5lBCuZsdo6nnu2Ip3lLHAHnBcgbq+HGRtxhXZSPH84MhS
+sJUZxci9BsXt4r6WXyMhO2kc+xyj0yGCDpbwgCoSQqT66jD2/lUDU+WKU5vl1l1+dH666svGuvu
/cyyaqMx45e6hDpOtrQ4h+B2eeoHj0pPL2leFkd5fWW79cqC9SIl+0UBesT2hEOrYqenUQUXps39
G0uVtv0LV7HkEl9Px/0s7ixblN8vzGb4VAeaJCNAxUryvIzajxg0UqkGflm53SX1XY9voN5t9KUl
SfAcR3PNufopg9R06slirQ0wj4a5SBrqmH+mX5xy0NJ1CCySvLAiOH2INhkQfCgWaD+lsypp8efl
AsgmLPmC3byG/q1AfYkF2lrNqbo6lsRSxG5qq8hJlDoDFOP15pXkcwipYF208R8gGGUH35juBO5+
Sbjdh6N+H074gnvpwHhwwM1uhi5R1jahsk+7KAKX05q0s3uJHRSQehuthkMKxFGk771qxmGy3Ji3
AMeW+1FbLXTrNoXywmoFDMR2xp2wSnwpqy2BsVKDaIfcZIo6bZhYvC3q2Y4lOXRDGw7K5n5dVXNC
Nd/Rc+4sJENytxENgbYQzbUXgtJit7QyKEWbT5xLRsEquHllNwfqWHwWs+AR6CCuDZ7rF/IOrHf6
EvHdPZT1FXESd+6XOM3MEL4/VlrE+oKl2/sNbNyTR/75TXvPGVTjavJGvpoB6VI+5O2U1nGLTpyb
BksC6rcdX69X6KdIdBWzxswloosboxZyAkUlBG+VGmUCybNA+ciTlnKbHoUErMkSD2th2D/lQhXH
agutm2n6GKSD/AmFbBX+A7mQVJj24Z5c5dd8kZQfc/Fz3Jz3YuytgYBs1sxjAkA3aDB18wvfDubS
pQ/yj9wA9042XkwoZjYghu4v3EnjIWzHzcfJHzdhU8N1H4CiS7nv/wR1zNxYn60K+CBIFxYP6hsk
KkvnqBjz3+uAinTYbEpPj+AMHV9BVrc2WJvdOAwW1Z05z1miaTDfEIrcp+I7vPQFOoXgAvBLLIBW
7PIGuj+yQmMfVZOouSt/bmFIiv630UT01pkxXFtTIww2cWVEIWGknOIhxNLdZyrys58Obu8sv9Uf
MReLVJSkJAeqhcs4eVaTvHzB1eReB1yz/g8uzWyNAsRv760zIddYwBHdxRyt/ozg/qh0UMR9hBpS
ug4iXwjIaPlaoqbhREJSxl5wOSSx9KLic4Ytp5KutlO/EmXpoYJkg5NndIrl/HgxlCIVfrpmLR/K
p2UGv0giNU9Lomire3HV34r+3BaN71ueUrsjmbilRoEuWy/tSZWYXKfmxj5H8mh2Zrx2tla/xtm8
yVaO/sNYx1IT2OxU8DukQnHV9SZZ6jatAlbmJfBnBJvlHFCZYJ7x0s2lCEntAf9/cqOWbq+q68Vw
yVWBjksQl6zKX8H2gslA2E5adlFuQCqNi3O5/HJpkk9F00uRUhkrDgqUAv/Hvf/13WGyDXYQcMxG
IIHbsOFTsdxR+NeMzIZMvrt2QHrBHxNaglz8UXIsnP0mlffCtjpl8RMqXuXmNcn2ChHyYr7kwf4Q
dEOXccysrfz3b0eZi6MWkdkaLpNQ7MJ7rGSfD2MVWX7WbCeZs1xH30Q+PR3/mpOz6jt7LK36ng/J
XTlOt/C1jDvgpe869YlCJeqZAS8XBqB89Sl32O3OnHX2QaJeJgHEdScwgoYo7ZmPF8O+9lGr+Yrj
/HMN7pQzHVcDFXlRCWMP0R3HVy2F/4Rb6SudQ2LGxfNVtW5nGJZdufmGj5ukPdjL+Hnp5yscbkHA
Dwxnf8ydDVh3ktBSKivAZqBflEoz5jFHnfsI45PIHGWA8eX77jvGm1xLY9AFYaiPppAUpbxDVdAz
KoC/o/n8k6/R5pcY2xOsv8AsJp29z8Oig5FQBFNQ07ienyV5wsq2+Qc+lbuQ8Zqer36H5c4ZtBr4
CxqGRxDLsvD8Lbj6v6DgvKNvEObkPd6uIvoJ11z4UGd9oRb8J9abhKL5DZYxte43tN3ZBpeWo7vL
xX3L7VVE/4UIZNwx/hVfTRoeuGKVR22sa+EwA5ZVnsE7sAG2otxdPM2vFS8I4SvWY+PFOoFN1B9+
YW/AOUG4ZmC4cNqbVO3e2Iw5KBJhCwiaFB+p3T4koZdwgDZQYdUKkcyKlENrY2GXQaTuqzN7Qqx6
OPH7KvF+DIxHWwToFCZRdKQHWWqGJeQWjEus06TRPRoepDItXp8B/fIXGBde2UgTVdUW5BdOmATe
s8hxRL52QJL1BkbLt5c/ErafaC5BjhyhR9FsRLOwgREIujKkB8BMRzAN3AYrQVZSWhkEU9JCAF9B
kzuizZU4fEVhWU5X1UuwqmL75f8f0vMlGRbfL1u03ICJzYSAv1ahsdIgXyQ5tQv+4Sx8R+xCVEgq
bRfiTVXsNRRQ2ZEu6SRGBxq0jFiyMkVjvisoPHqQ2vhj5J0yifAhgBenSlXP5ALJ0ryyF7HWXxSx
n5AkpShIf572Z08xRObNMxWamRWhBHC1Bov6EQ5W2gkF8Nx7hGrtAqTOLmZfByJAaYKWOgRrBDBa
6J57E6zMO21jXkZAoWaqvysEQ0mYFliWNmDB5/s0Qy/0MABpW0CiCEXLWSojqtOD4mXIY2kiVNWj
DFzAVxeXCc50WE1uU6UWd6OZ6JeVjaMmQYC0mHRHSfDB5j+R5oB6dj822NQoWQXGBatxD96K2JRi
xoRrq7HUWmsnHxf0Yw+PnZ8gAwkWXesq9kyKv+yiW8HbGx5kWUj4AY7qt0w4hs22zc2OgaJuE33J
zcCN0PvnfKKQLr4cQp0KCAq3PNslzURZErlz8vWerFQmkPTAWHj0zTt2a0qftGwcAkL85+Z/zBGc
a9TXZKuvk3t9wBCbUFR4hoGh2oBASpAJfE1gKt7DFHuKx24GXyFkvgzdRUCp4iPyumrlFZ2NKz4G
1G3wxURg6Bc+HkPE0dfyv7breWy/+8GDmScA8pSLmsYwjF8z6VWvprrWN4qUD4cCabRTw8AjCAdQ
gXRl9/coaVA20rsngJflBxFJzTRzIbcVMbjWOhufkAeY6ZxLgTf2NSarbeyz9mizQ3wkyZOtI1KV
qfKIEADrjqxyj61Hx0S89XT+sthKor7ZXb/90uBKMO3tcjnQPx/Qt5HefehfpuM2cFghchWQ7QHM
0jfHLP3kmL0uVKWl4Y7N5Vt8gUEg0lwlLnP+JDVwGNG7nqxW1BbsoP8i/fSwlPIUrj8IBOXhOI6m
dUDaksnjRP9K5VqeGz2xIfrjAVRWWKXDHgWSvh/ALIFgfSTvWpOFNMSnbUGhraKb8vnDvyibCw7u
kfLGtXXC15fD3ksPILVdangyRokqGpMoYmbcM9GzVpI9F7CZgzpJieN82Z47xBaAzSZMamiyUEuR
1XoMuUPX5Nq3/iFPYZPs46C6weAywdjYi/RpFSk7CT1IcdW8ib2oZYuydnnZ4iJ288s7C2K3e+WK
cTyKyU6syTVelCCVBdJkSkBBzpq3+LqhyXNtSX/IbAvSAaV+t0ibExvyhga+ddW5ZtdgUVRQ477p
a383seFMDfro37eixH5yF0d21p7poRieBD9jCSsiZF0BaER/2Q3PsOcc4/dh+tub2VEdm9Mp/38o
MuePmMl5uOvKAv1SQeAOHv8ycG3POKLuf3ryusEhaDpXpleHrrAlgtq8rRbrLzImCbGR4+YZdsag
nSbHZPDLi9pY3rCFPt5480MX9PWAvNAADHYHYdG7omPukwKK7KKYWsFw7k8YoXvOxB7ZSdCVuCBB
OasIlAs/3vR69HywMDfIaMFw5JCrbeuqYVHRS6x3IPsHwGUzEtOx32OwAnmNPHy9NFfHcJDIbFhj
4bodhr/mYK/EjUle0FNrjtPmROXRrUgKFwDV1hUl0TK7+gJ5gLADRKUmdQeHF6zmboqQQN1rn3D3
qJ+ZK0Ugtdj7QtYizd8cXjWZGt+2y1RXvnsFNm6iCrktE5a7r0fcHGfTNNWKcVLX43e/kItCRxlP
AWK812aklxGv4l7wo5D1TEFXnXdJvQG/Y1nGX5bOxtLdmT36HftTcINX/kXVTJVmU3X92eNCU9PI
/2cqKifQ/Dn8a9f3COwuCK3TGYDKw5uh28R0LURSb/rNRboGoNYqS902EhPNBewkcWhGrACe0QPJ
EX6isXV/RLIlbcPL6SareLfLzpTGscMyrMqui6j/go8kvuZfM8jhNJW5yAKWlAzTCOrLxLwvO0je
4E1ecS/IRrqlv+mg7UOKZxHSCQwEmxCujY6veJhQZcoHjoNLfe3fEMRcD5iCvvR6bXMQedQ7ZuJF
v0U0JEH87I25PxW3x2DvgOHIuBHl5B9UVCggcj0DOblEZjOKOXY+mUDQy69grSNL2a5OE5tZ2dsx
43SFA79icY1ti6qa/gr8L0JAakkgbaW425k/M7DefiXAm8ow1+SSFLWpeA5Ytr9zMlfuG0yAx57b
GTmYnYzIPW939hxAyLmnoNwx+4SN/GxQ2BdOEYc7PydvhGr7BP0rfnPYWTqwc59G91c023ot2wCv
R+hXkufS9MfwI/54PRO7ancmRIRpnrq04pdho45uLKEmB0Wg4vsfDQAcYSMsus02EMdsZiRQE7wQ
VR+w3q8Y1IVd6zFRMzFHi32trEA9A22FM1pT2jcD8o6wHEYSmeKcIEdHl5LEI5DoYwQiMwXcKW4p
1k85M1BxO7YrG+vxXOUk/SInGrmNLHrWJSdql/T6+35a3P5uGzq11LKzaVfig0EQssCu//CyNfXW
cEU4BamnnSXzM34ceg9oxXu1oROa3+07r6rN4tRxcATuT70/30UuFYw8bSJSmNHzpFuPVBCAMcOD
JVe3p2HgyBSNz5PjhsxtXEMUR/BviM4bsV00J6q27toY2r/Xczf6xetN6eBnVJong/ltAVFb1E3E
OcIcrChn62ZTHUYtcyabh/ptdW7mjku/ZU6K6vg+cwnmb8BOdoh5viI2PFa2jpQmqg71gQI64H9t
dBYGTBmPm0HGl2U1h3tDvvKfloKTOEybEh4dgAS21iev4Db8GJtmgaUVIE3Sha7Ni7bAm3z1zp+1
gr30PjO6EPllMkQC9ra32iaFffj0E6ZrbMpbDqDp/JkRLau7TR/mClBkQDVCW5aB9rSLN9KQ5b26
5HO4YFzfv2bvTGo+ebs983RjD75zBaELvLzh5TFrNoMFSU3ASLVWXXC30tRBnmm0ZhNJzeI36rUc
xVZ7gTrTXsEwxYX22V84+VkjsHj6I7VIWHFBU2eFmGOUSiYpqw/WTFwmnQArR+D3sivc8zio596H
+lNMy6xtgzeMlBwIgBwIJP4e7LExhq6MgYeQcv1CKoBI6mUmONhgrAqdTL9p1gu58Y3QgxM1B8kp
NQWuhnCOiCBo9PJHy1MN+tl/DJ4NT91pb8u9WUlk51Pi38t0OakOITu5LkpyjSnF1wwdX5PQ6Ugw
wYqycwkfIlqvxQpCKf5WfpmJrI2yYJtNSRGGZW00g2v6J4fc/kHPG5tE/ir4ljE50XvKHFpyDAAE
HJSwlwt4T6LKL88SKxjplW/rcHU/r3l8RpAB0ycXvO2dUXdxTqJoZYnpIVdBL330J8oppj/GMSAx
uGZ8QjvnHtFdaDFrTFItQV5vwxixXs5qJmFYPYorrfPcaTeSLDVBuFEriABP27oyaHGPAjbL0XG3
svvwo3IR2Vta3uU/5eBtxhduVwWyy3nIP7pID0jAHrnKFMcuYxbxO1NtZHR3LQbBx9L/aTl9F0L1
X8vLenub4uSMxMkb46J9D2HNbqyZXHHBZ8WOc/Am3NhrO/+0/in6JNLVhQtUl0+l4dyVG5lvS4yn
ygK/qb3fONSlwtsSXxaAhHE7RHJDBSDAaI9JLobJeFEKS9qlg3DdobteDsRy99RCUlKVm2MQfGLZ
qTrKaHOFq5Vy/BNPeGyM7qvN1iq/urU0V/3nwszX4NVeU8GeVEcwb5aB0ZrgJnM8AEXoAmhyDYAn
FZY3y6L+s/A0p2SpmFsssV+IuVuQ79np36tn0tipoRkZg2lPzfrfpry6unU0ewImZaGnzvxUADH9
LhnwBSS46q7i9gClhSZIrhMHypkiiEQraVT2q3DDXsH12u71yN9Ch940RxVZaWEpAWTJgJxt+oeM
RauY2cg/3Ott996YjsC4VRLvuqR7R1WtqnYJunXcDNOoTegMSjTQ8N7tTZgEobllytxGr6fBXDXc
umPOKsLQv4QCVsK/g61L2UH9jMCXneCDMjkbLMaNfD2mw+MiI/vMSgRpHAf2AUWs08ME88rECTz4
qE/U638IFUKW54kSiWsncg4NJmQT9jRWW+7oXntUg1v+LunqQ8+OEBahylE0/Ay/GlGTI6J+ZW59
1UlDLgK9gXOctdDYjIZAZf7t5CCr9dOkfGQtzPnP3tLto8+uKol70tKfEbYS4xWRuQ+/nirCy1kH
hoSCzmJozkQ52H0O6KFSBrCSpQKLxwltAK+f04f0tG7EwDeGjGy0UIK0SJPT7sq5XjSw/EEp9B2z
6XqCZJ8hy+hNMpX1U73K6ABDYeG/rdiCcPtFe+3ndruIJ3xKCCHeVrhoDHxHyB4UmFGZhkfgBUqQ
8ngB8YECoAjX4EUHU8ud4COUGhD/APm7VlEZSbRqQB6zVDk/UM4Nij2w3mKE2E/kO82EtWvAQq2m
H8MGyurEoURHmsVTpPfINEZSiOdV66GuP1EJnyzXEP4kIqxdwgkdC0rGkwc6faedOcgIljFqV8rx
OncshIwf1SEhKj1NXG1WTQSg0/pVq2steFKYCDv2KBKmfhpibd/ueVELlmzekpT0wr7Kaiv46J4g
z/eC66rwVbQptTX+B/+2nSZZ9i04C50KXTC1X8kDQkNhy6VlgU8EuC5733pGIVXa/hXR8REjfg1K
KywoNlVrF+yBLQVYQvLPxsmoOe5rw7Kew2nqqkqUHgWXHx81We0wk26T7OC1h0TcXH091y+pYc+7
nBF8xkYYegoGofwlSSsKv95IgmHDj2NZ44s4/9M0qpvEvqywVkSqccD7R0KOhSili7nI91vFMCB8
lQOLomKScHBN8JlA8gm4M1t/rzvUunP6E2wynTyucRC2+D+LAdRJ3RvS05neZ0UpTwdOrS4NxXB5
HHC30IyFU/YIS0vBEQ7tcJ3RGgdHbJWseasWpODGMjnFuwUQmuxD9MdhpFtL+Y5Ym75oSHzqEgIf
IJhKkV3uWyvaAms2mggXSekl1YWfLYhzFnQCJv0vzowcQv9JMbWjWFJjDer4gSsPL6RPzRpLd1Dx
QnZJtlXV3F2TsqhINUXS3iwXs03Sgx36LDahX/A/K3hMKw1FL+vKDlINi/R39hsOsPKSIbsE/Ti3
yczaYNeG7xgT/Y5Ds6SuUEz5rVoW1cK7s/8xtgKep0hh+8jdk7fvCuvrMBuuENmbXYWDhbhT53rC
hAiUNZsmgMyjxQsM+W2q/UmRfnprIqMWUjoGoMokXbyfWGkwotse3LxU9e2c0tuUKRo28tJHG+Ov
UrgcSfRtaqpwqD5zIgh6IJeUuVr5DACCSQ0ZOvnZou5u+MDuCGjp1GdA86aBx+3Z4jdMnjwCwdkr
dMLBCl9oX+NXoueSvtnTa9XYNyZko+74BE19E00YKWe2GpfT4XYD9RcaEMPUi4KVpUHOLH8YZBhl
tiWrJG4fv+51iFzbVT3tGaPedF9el73FQF5YKFmD0LWzkN08t+tLZBX7T/VCMqO2SHJWgBSwZRiF
KG0Vww2t1UdANQCBQP9SITtTE1MxFelAdctCUuvIpBQi9vvh6HCzdIbOqBgi+oGcwOmWOGEYnqbH
/2yVw5n809pAzzpujKxA6M+V73OgDgF9/++PhwXPp39eT2bVi7cPVdOc9FnFwnJHLVO+UvBP89b3
i7JBZmmkFc9Ial5g4uzq1AisQByAIHWthz9nwDHSvnp8Ioq5+T3jCoA3Dlvqm3qRGWgkUWqungJl
BEa6zWCLixPLZZ9UgNOZVwG/cr20/e4jTS3PhBWobaogfL+mlo2hdwCkdrW6pHhwoWedf7pl+BIC
NJVdF64kGnB1CUJ842SunM4iexBf7xEtqgAw98VSRIAm2l1I9QQif7yDrRgRsefEOQ9qZTuylJoG
sZCxghgMWDMy0uQc3yAqx0Pzyd+UDLJBgUgbd5TIA7NN6BVuAnAJxqzXUjyzgPxmifwHiCSRh58p
G+DtyNs+nw2O7t+nLNNfC1bjucWO7AT0X20ZG/ePhKWnOamAasatxUv2nKOMZvFsxqoN12WrvdUR
3evuMpBuP2qVLSg+5lQbMXTPmfK2EixanDDvca6ZhW2Gzvo2lpJEJUCUXM6z2xmyDnsrGm4uYjiL
K+5LwJYI2Fl0b25U9nO+0m0FghGNGeUyJ6Lk1tbAWG1Ow6OSIk1lfKShhakcCspCga9L2qB6RDmI
a/CoCbZvL2uAoiBxbPaJE/6aQV1fIHzlzoCUnNHRks0N9K4lpadB9/Xz2G9l9j11pfx13okiMpx+
yBh2U5bj6b+C/4K55vYQI3iqWl8Bknj2Bc4hy0hnPdSLCif9hJ4QsQCCKbSJJOBzwJrlr4nmuzZl
4CCXfYcpmtNrybo5TOCaTE45pxRm3+vmmlC1LQ2NN2ta3PJrqgrZf8je8d9QbhLNFd0L7nwf/YoB
dmJldwFf2SSo86deP/INwYnqnd7fO/PB7tastnlnXdh0iTs/fR6itLNShCXBAB5qBrC49f8kM2Xn
gAu0J/3q9VBiiWC+MowwCzLBymDAf/x3l/aae37V33l3uu3JAkkN6fD+wu46sRNQD96NHwADlVqP
qA2l17U/db8SZl3q9SMWtzplLueCSNSOa/sauTlKRMK+jKY45tCHPvGSTZ9gmFoh6nxXuUr5jM8T
gJQ7hM912jTEBwI0MZQErTM7io1ms7hqvjFBosASwemNNGDYTtQ/Iy1u25h1WTsnlxCwogI1Ou/s
s+lA+6IMC5Pvm/62j5+Y8asmbwmdxYBKW1NRnJ9TKu/C3m7qIhsQUP87EDq5PzqQZZObMXo+jdZO
JDj2GP0gIvggOlpL2BCX+1Fp0AdkBAafhG78X1+0e+sROlG2XmRROixcOiTwCFdREJn7DoljJLxC
Vo39dyoooMo2ubsQkT08Y4l+nVMcNi67za0VPcG7DqF+9Dlh/uhkQ9lwPzj8hPXJ7qW8J3HJiFuk
MIWkxwwYi/eyqgyh6g0v3s4/WZWw5yWx9jXveQOHqrU8BguYXouRg1NfVmkLaiOZggYmJz2HUcOR
kElGR0t3IDLWLT0iws2To654gqykzWRnJ2ijEe7Fc+RkdeilIbrkP4eZYv3i/fSk1Mw9NJhPjJCT
YI5KtPeYFogpVkuE1hd9YVqkuqXp7b+c0V30fpL9jZjbAjU2ZF9EHui4hrzRv87TZ0YU7CKlBdsk
FFtma3k0R1ksAyEizcWla7eYP4nSXoB8RaL/vHNKYs2asO5ikLJPI57udWxYpzV5e/BAgD5xKhOm
OOGqSSLtXA0LV/DrOmCRftUarH4P3dOKrNKhrUUVxyhleua0YufmLabxbe3a+/s/WL38ITzZnWf5
uI4jT7hUI0K5xzZOWb9Ib3fADN8rJQZMm+S41EkphI7bdrH2x8tLUl+PQS8eaegSXhBrjTn5G70a
brGDux/29XSglRkDKhevLoXoQ/1u0Y50lBfjZnflEThNo2XPQMKzA2/GD4le2f7Hs2x7hc9nZIbn
HX7xn2en+OSuCySE/yo0mi54asGuayvueyYyhKpXXPJCjp24ZcKXPygCF82emXDV8MxC7H5gtmVw
JQ170JBaai1nYmYLRbHHx7dfc0OE4H9F9YEqtolhlcsOIyGbtL2jVgmwB5FHy28E2za8RxpFwT0a
7unsvmrRDtyIAv0fnTJnIjfFUhbhsX+TQjZHsrnM79jkj1t4/r4FaZV5UkeX04NZngQ13NwahJGm
f7hRZbJZ3iVSnnHUIk+lcQ/obDH1BUom1awVwke1FROYrT6SgEgpFybUO5AB1x24ZxRbV+L1PktA
gqpRn3HOFqfjLWIiUDvtZLKge96Lqe1CcUzj/MBO+OMOXgxmLd0KC6b/eoPEKKrm4KE0fICxo8qd
jRWelUmIRZPNCx/Mr6RObOTUTmvZ4mSn2D/6Gk/hL7ajBc193gV2YCzxpSVnFnHP6FWxEjiV53Qm
ZM9gAb9gvZX/JeCHXNwBjIZeU5XZ1cQxb+bIcmdbZjz5Gskk96ueSwTWtAN2lTgsN1DaELyWpAdh
pNiuyCefUpoWllm+GXs/SPZ7AAECSt8SWd2f/d53lvIsHiqRzUX6eWrLMWZLy06NWaUJKW3zfopS
SkY4M2FfckeJ92QBMrI5SrlSmt01eLRlYhdN2oVhDnIwqO5QwZBPA4Ti5FVlx101iWRkYRFcSM4Q
JrZY+A5ESuBkLk6eIIHvdPvk5Cr3rEsPSgwy8vRsjtwszeLAeO7xYiEQiudCtDiw7lxxWD5DfuQx
6UkJXH9smlsD3re7FtV8rPB/7SjVtqZXT6APdpcXT0Pj3l8vMq4lJOJYIuXjj9xFgwkKfgsBx9Bk
3qs8h5gC3Eg0kDeMEwfImRjNzud+EeqLJ5z6P5Gr8AULCOC0RPH/GIhtvdJe+OSjRZ/bcAEsYMrM
pRl1JZbvGp6AtBMYR51sv4oN7+2BcF/koRdj3j+XH/De9OpGAHMxyXRa0KHQM1V8IbdVI74vrM3/
Q4dXQP9KH4VmVx0m2v6ji2Py6Dvn38AJPpP8/NlkaJpJI9cWsq8nCpR4yU04c8mGdTzbyn8q3r8C
p338IPmIbVLnfA8x4t57lR+q5nItArMev8Z4dgs+70BhVZ0afmzLCz9jAcAiqWsWeEQTZqy+zvaR
olnQl8lPUFK/1nIcr5/jm248dW+1U7I/LZUYjmUkwzTWDPUYS4jQLKDQuHniOngDY6W/DH/cV75C
kKkAx8f7yFb2ysy06OgG2AlvKLj3/A05Yv6aPmbGm2kygqRWvGZ5nZV33COfua3zVcEprYub7FWI
Y7CqDrDbVI7Pw5NWOdGgxDHLI+ThKjEcZ0V5La8MZKLgkymUVy5/qFztMv1inNNPLgOO+G70Fpxe
EDshk6NPmzWKyVhsIJ6k92+moRC3HvQbgNQlF7M+3cG8qa19MM1z5uz6VuCR4YgSkMXHsfvWcvuq
UHrdyjBNkFAm8Mgtd1CetfY+a2Oskxhj47nmpPNmcE1zJPtAgT98qLmBO42tHeH/9KSpyIUKUht2
jya1d5J++gx79kntLTNd9T4dKY4bscUwGESP1zOMgLF0aYOCzIVYXbLU/QkHMgH7LFkBwC2epzb1
/70dyKxTy8qg3C0KiulUyErrFt8NHYaHGnlHun9v2omp4dTA6hvY93zGLF2S4Jkm/SWJ72PYHM1o
F+70eE42fpNeMOxnQ38hc+Z5TuvlY5AaOU9mCdy6BDdKud6fxOinrTYzyD2dEPnqFN0umrGt3HXD
h7UbhLwSBB4XdMUr3qy2wmPa1zTOaxKru1vvRaK5nBqhWxh/9erIOvBn+k7IwUYAm3rM2feu5qHt
4SwC0PhAFt4xzaF72pTT2bdas2UGF1l48AjrQPD6YotOEDRtD8Ja+YaAcz4daW67eU8G1idQOJfC
CsEOfkfDY4TTPpVPBKUtYdqkdKsZWIL3eqe03MtdGBL+T6YxZdEnmiD5Jovr+hjW05DHkHXmdMDY
SaYC+9ju9DM6Oc7dU8XYR3S77nYog8UmtqcsTLuC+8k++6FNViwr9ZAs/p0D/65C8zqxNoEzgjVF
kSTVH4EAisB53GBVo76NXpsvNBpivCSv6ir9kpMdlNOsTHEaVj0SrpcSY90Eb3pfBbI10lemHfaz
r/dIp5oEZ40jsV/0Gdn391ylMjlAt+hYoiU7oESHLmb0L1hM6q/HLBUZUCyiTcX/oAogOIzuR9kB
5kDsoLesjooo5oTRzWSa/xaHCkkFHyj+ieWNNhC6/htBXz0pJ6bB33p3CQzyjexCZzJ0aAg/cwq6
uYxUSomG37L1Psbqw5kfzcOt4Yten+W0gZ+nj66MW2EDeNbeVigASwbysvHSOqr1wL4RppGLNEPU
HDyQiNw6CgcyHBizuAVb60mxdM1CfMJbPY93Eek9z2YxDteWvctvJ8+zFOr9JfaYUp0r7uDMaGSS
YWcWWqUJGbPK6O6IdSKeJoKCuwqjTP8Yz2DPJCLPienKf502iaFlj+EA4fFDEz1z+54p1t5ZaQDR
v+A95w9dLssjMzPvWgMcu9wCfog+YQE0KAzXbnTmwfLuWJgK4RnBPHRDUgJ1aHVUbDJf2+LsKDKZ
hddkYzO3HGEm9KG/JMV+i5WqItfwGvJQoJhmrHD0db1aPeWwwGsNMy53c7bSF09NVXG6HzSUDtKn
daNiE6HVkehYioffPNMbJmFXMOMRjIZXBtykmCRx7xbxqjVH3M9uPrSWpgVUG4J0W5rXbLCZDSyH
Ph2CPOt71KW6YfoxlGeVPLIhg4n5yQ5zkG8SnDtA3rknZ99p0tCkQ9Fd+CI9hAITVWNdXHel9HXa
8QTTLNXXWo/Y5eyoExPPmN19UI2/cvFc89b82VLXuZALkUGC2cQYeDCLwTPwhKWbQB5GnBxMvaFe
TZ8bO+GAeLsOH6WWGQ3xzw+0G3lVW9gF70e7DQWDuc4hs3D9CZa1yVo0JDj46oX1j3iOhEvRixBU
+rOoGHQv6z0nrsTrJGhe4kFqg1JeZaG1R8WhbjA8t7ISyD5luFWESyQ+pYoB+Pnxil8Qqi7VZxsD
56/dFWCN2D0AVT5qcYKVKghIIo2uEEbkXO9lpQG61UU0+hn0ruE6MftoOKI8Xis7HidUy5yO6sEX
HNToknG5x3GErw2NcFQRY2Iz2WzT46zIPGRo+V/zxqgBv668SgJsngV5hZNJa4+gvKK/oqKDhoZN
IopVs3o3Wnnxl6vg4lVLICqlZGXetLXBrSJBx+KWcUWJaWQt8Q7szoykaY+R+VxCStUZsu9uwwyz
EiLp9MOuR5mldlUscm1YZIodA09Vqa365VTDetVycboAwcE/KdNQlR1iqO9WeBauMeOk4VYImCXL
Rh1fen40JbQkkAEeAzK1q90aUEKqDfVLakcydNDHYqvnZM2jBscy+vPlxikXlFNmm0x57tlCrZIr
UvziTvpcT7Z/+SyRvuwJxmZ+Sj0abbRroqDL4OCCtF0QETgEdRIo6DYhLNn2o/fN60qVyMgrThbb
N4eKwf9rqMMxl39yqpqJ9iUou+QruDjCZDzKS7lGEdu4RI/+Ht8FTo5/UztrteFT/mSCPi4jvfMr
rzrcAPtbSTHtgAzYjW/gyg2rvSM/O7Elu5oNjbMtrevPOqvehucgVwcLmUaS/C1pQWVzi2Z9dFNR
dUcNQrrPlKbLxGzBlKQCaoqSdmJq9v3CzSAh3hDqDiFFl+NvgmxbzewqCtm3dSUAY0x/w4mSmdKp
iSxTZOei1REVgToHSvdfi0Ld/5ejn5eaaD37JzgOvRJQgX6f+T43JI0MFUSvhxavw3R7hJHk4AHL
D8k7/M+pflwYTxxd0PO70x9eNUSK4Zvaj9fbXb47LViqrfwprOXGL+73ZuxHAubLqnljvs0TkAPR
u7uXtXaoIV9ZbmfUZHAsilTsm7OrHEINhsoKQjZ4gxPBUMiufJhavthtzGB/ROm2P/NbPneaaLCc
LqYzBXjQp+xtuK08vJUEQvyanTRRX6SMOj96HaTRmtgm3o/vb+I0cm00TeyqsrIppcxt92sUdR7q
HvqTo/jPEVVlZLqz0S7MdwZB+JI5jthHN3TMXmD3032yz/G7GdH+NAyZQSzSop6I6Ar+eEqqGu6d
tZ8MCd8My3EsGerVKJH0aoKZA11EJxZDnj3R/O/zr/IwkBZqqP4tnK1NPZbsS6tqvZwt1aprdEjf
dBXsbPKm/8JxRDR8gEBXqwJIW12lJrbYkHbQHPT4gTJwKhhvYa036zqXf24FO2tLd82qdVOsspiL
nMw8Dc1qJKuy/DnF5wyt6Fe1SaLK7tygEZqwqoIaKUmoGgu8tD4eiH1Z+p3oMLxG9jbU5oFEHWxb
E9Z6WyWzfSwT6rZpfyEa5jKzFKxHly1wcgAilDSmYLCiFm+g+s4cThbDOJmyKFELL11iTfbsFP+m
KB0EnMWjAHK956ebk/l2euQDRBZygodKsHWgbugi+Kb2cQfEVIi09OqTRduzfT8yIb5Vaym9FoyI
oiXWXS7HSvXK0aYQt+/y5ER41wUOtiRv5FJSGEE8bnwisfqmVav3/S3fwWu1oYyY2Ku7ekwDwkHa
uoVhzxu5Ekz830X3Yf6Rcvs/1O1ptXq0ap/VN5f3LNNy3CKAb0PkgN9iIC/KdsntzwhsfFxYyRsX
USCN2zRwMPx0gBoabnTQkK2BoUqdP8Qvc91iJnJPNUjF7qTfxxiLjUV39/IWxtEutVekSCHqDbc2
NURi1+X4cf5DWJgiUY7zBFIdHR7uDOqzNJFlmREkhCI39yGA4G5OGoOgife1841nSdBrsQX37KfJ
f2pOEH8R6UgqqwQlA8b5Je0F33hMNMsgBtf2GHMDl/zFjS0xUawCnfdvyh2reKbN7yXxwwnPrPr5
4EJPFh1I1cA60waS+Pf7KHWwpJy/HH77u30sxOwxXPYuJZckK0dRryw0cNdtbACAsPnwM5tuNiIn
7IKXdK1Qt37AmkF4FSnGdPq0JQ4NU9X48JBczpoADAOz2kNJo74JTdIMUSPEWh6fE4Bhk1WMYNJW
wIuozZyyr+xX3IHVr1vZXam4UxGnf3j/KsMDiW7RcTkEV1o9nfU4XwwLSfjec7Lz1cwzCJvcLjYY
WGVOiZ2KT2PXfuBrYrKN//WOkB7VF9Aha1eY7/bhNXffmlNjjWidFviam8FlmQN9Fo0jTbZHQDjW
yMPEZQz6q10SnFSBoFGV49DcShDxc0SekuJBZPzdVqZ/U4kgT+zVDB3uUNkGBKpaJekGhaoWTJ9B
nkCZDR/HZrM7YTcrxLWTmttqQW/2GxWEs1yl66nRisiULdmmNXmXAIlFlj9UUz+se431KK3cdVyA
vL9WaCMQCrCwWO0SZMFepiMD3JRqlQxKuy/XSPudKrE+1zrv+Ewe7e+SZOgcTJeRSYApY8vY5iaX
VHB2hhyp8z35Wmuvbvdyd84FN3T9qwTsKf9sBl93s6rEEe6Vqa40faadQhaMPEjjr/KBlBLJYNxQ
azdsNCkT2ckDVPcwUnndKHC/N25DYF/rmfw1kHMicLym640rA1wVnGm1nFAkNoMirRmZOVtoJ/gU
SvMkO5tGQcYGuT6XJNILiQ7V20vB7F/2ffFm0tPisX4f8hVcO50UCvkFGUSzEtuH07UmzDYLOQ/o
vXvQZyi+geu9TrgFSconX4xs1R962iyYU+20/f3De/qBiFAV2HKn8HwlleIT/EhCRcyXRUQcJ5gQ
nUpieHi94bKJsFd2ztQbCr8XccIYbnmSZ97IM45kML7bo5a2jAOMgLKwRyY6b5voV0V+IZYEerWV
3KQ6F9R2+UjMZs9hijqpkoWtluEumy4oDg6QuaCEc7X8dUspwFKFwRDiOWzVPMWaiRU4r+aa4DUd
XJ1uCwbPRpUBtiHMnQ7DlDiLbGiocNqURQzKe0EjQmdIewqyeHGYNr5FMvQ/ISBYMkl9d5udZsVq
VwmwdhAuLVMDoZ69epeFfUeRXYtgNSdK0FrmGKuJdQuWtXF69yWyRBs3F2yscK6juYvF1YSSJFIt
dsH0iSG77pU4cl7YFCR4lSg9pZIMQUOyMdsxbyBgcesMHddGPtNlG+tMdQK4ag0ZM9MTDOElnt0q
YJW07fXzhHuJvt/eWtGLe7ZzC2Lfxht1vOziDEYi+t7RNKGRMAWSq7hB5IodjFjTTEldDS9+/HOu
emrp4kGCDx6CIF3b2Ulu9j+LmFBo5GDwdRC8GB9o2iuSTFj6QN76bngSFuDFdAMJo9Jro4ZTXrT+
XNvWOlOu8rISUwRYu2lhpWzU8hs8oNYdlq8wrUQc9TCtWc36ETLEyo6GHpvV9JCBi88I0shDhF/L
Y0+FD95LpddXj0iffeXhWPAASYYb/Ka32tcYE/CBclUf2RVRl9t7UbzKlUjHGoV9mzweVZiyQQ9X
IUVuKtDOeXzwYyENtRXKGN+A0XhHkrZiNxtca9GqJtGCI7nJLIW0lIZYUz+3V3xL3LPy+n7awpoS
73+ZipcE4Ucqv5jrgKT4h43rJCcp94cbeC1YDxq+BajOebsomfOoT6tiKyG0Zs8xCHXjD4Q/leyk
RQ5a1bl/C2+TdSpASBP3N7j1r5LT0lT1n3PWsGOfQyvz9olJFi4a/Snrk4wyuMcmj+MzI50GRDxl
5LTw6El4B7euSZICuE7Q5lrESD0jJykKEuAWvKWiRNk/yCfTjaVi4TANszzKw3FLLk7HUUK9mCpA
ptIEiaFu35UXKn6hEMciqPsydqahzjm5oigc1XfSCcYa1cq4s2l5OX08xwXat4xyFw35HOwpAJgN
UDYa80pCt7oBWJ3V4VU3LhZZvcWehS8aG3ANIHBXcn+oFzQIlIaEN34WJbgJqN/aekYDmbK4WzYY
E7N8RDaw3xfJIJVbM8/i7sTgm66adadPLkejjJEpB+N8VDtDuhSgPSe3c30A7oTMV87tf62JwfCE
6b0KU0yMKKw6T50KvIQpTTie3HAVFhebwQK3v2mhd/o3V8RX38sNHffzurocl9bVQgt/aKQIIxye
nW4Etr0OKG1MQ3IpOsOI85+f49jxBea1Hf+m4ePiRIYEd0sa49NYMxxoGKNeVUYfFH+BRKpTDppv
AVQ/4ZfSS1pSOkQHYRLMqxNYs88DfpvJz+ICI1lTfW0RYPovx0B3TXh55KD70Op95VQcD+XU4NKC
zaRjSi9QN1sZT0D3RsQ1wH6tTzfAQAxkdQLuyv4MLd4V4xKILlSkXXuZmI9T3HSzu7UEfWxJljhV
ITMy4tWdDwUNHEVvnM6zxOvKHiQS+og9Ot6n4ZjnYO/W8aHyD5vHVDtSoMTLhcCwAC4Kp7NR/l9y
UiFSVVad0Xr5U3IYVeWHoMw5r0PuSRniPpgnZF3GX9uksbXjUF6iavish9Q7LMHy31h8ZKLHErWF
Bs6CpXTC9/aOLTMKkBcFK0Q8TEUhoXLoughZDPTUhrbHvVqVT7bHKdf67WbVpxu148XNojRGwW7/
PDIT+wWufZnOHeaa2tsEe7lbW6s4/awdALDrBm5uxzMBXeM+BImicoGx2pqh5bWOldlk/U8Mmg+9
wu73DSc/gAUAzEqv6bnYCJOJOVIkfwWh738UpA+pPKgWVvKen3pF/0pPjmOwvCH1ut/bf5Iat6u+
Y4ekLDyYG8DkJQr1WMyU17SHzMrSjrsq5xTZOaSP/GlUgvUvC2J1oTD9QCFOh7eH7dAKkl1ySAfv
IrmDNqjGaLHxZORb0EjP80L1M9r2WEPJUBqjlAtHRFnaUDLAo5aTUqJzx5YId6ZV9r8cTuqztdWK
WcwZLZ6iS26djRk+Up8aJXO/CxCtH8bCQxT49Ro1Iv9ZsxXGP7kNL58TKqhbrkIglpyvvKdostCL
Pt3nsCBb+ON/KmvuR5/Ju/O0Mm2kScRixANkOzY9ivN3/rRZS1+mZ7G2e+rDjmYeKSIYf4O14oL9
aBlWZjSApFT7QTWuPBYjBJ0KCbvKdAdUxdnz5Qzas7NHuUv8J1PJjKhPXspijMfQUl92xRHAWBpO
R0nOVlRI5KYjSPC69MKXog3X49NpjrFTQZu2tHhD+d4wKnex6d0MzCWAe/uViJfgNwW9soc1XtzE
aIhX9DZ2am4Xbgn0nKDWoRMwLJcwRRrJqMqUC0O+YL0tqfF20wxzBvviuEZn/4Fv4OBanHw/5tnK
dyNe9dWGVSs3YJXi2NE/cdG7fg/ISmkZncTJDu+kfCRUJn+BvdCEtprEibIdy9teLkk45tc6UQde
j4zCX7ZFmqpSD7NipC4egAP2KCxPUUhCFI6fPJ09WKVMB0M3OYMtSKfH5Su80gBDf5H3zMxy6q4v
Iup1G8m2SNYiOopb0eeZVDYyvnfs9q209VuPJuZht/SAAxO/5TaSXNLaO1KcGo+4YIHfy6ji5N3v
aDurw2OpULehoYnrGEfUlRj3ZASpXHrX5AvaQP9vprzLeKem2oTrpPe1VAHQDVvufPiIGSx+hdVM
Q2ENhA2p8qX4f5J0aaY6raYeV6G4gg2fMDfLymta1nikGKwv6y+ir7/I1TVOpkxC7ulVinpMmykS
xtgERUj1P+a1qvH/C+0Qhjey8zLyX7sFyldXAOhRpZhmnl8Ob16rSO0Er2Rl+jvhSTts0rNfn7FP
WN9XqN+H+Oi+yS8TDfPB+EJg6oZTSa279/BEkSjj75MsuHcFY8i8/lqd/vzTl9N9VQ7e+DtVf/3x
Uc0CPWsa62rea0lvdd4ZxsXC1j7j3M59c0S62LN9s6sFcAdn//57mvWsrzsaqoFN6yUb/uVSAAwh
WwDiKUFh03I7oGh8jKJRrq6F3LqmCYs1uVfoV3mcFc5WqvoTPzfsKjHw+brv2HR5Tw4dC2zQs/Z4
qJFsh73XhCnavjeAwq4GnkR7ZRVdxqIhDAfnftjWWdE/R1kHDEQkImJYI6o2d7T/EwovODMIjKl6
7ZWgjLslovXGRixp0RJq5ErAmzbuG2D/AovOhVW6Z/DXoBrcHd4fiw/gYPGBqMvz310f9WERbLgo
ar/N6y3xz35nIFEyOJpwFoVPobtZ2X86qt+YB7MsG8OAA7srCvqVC28wOTg1qkyPFcs/nhJRREya
Vp69e4RS9z5vjxhS/6Wu14Z6x9v07yGIYyobFvg7I8nC842Fsl7hjgQ9Bmx/BGje00PyyDbT+4g8
do7TR6kb+m6cXyoR0F81mWWomR5jg2oPEjv23+CdQ2FRFNok23cDMkhSV/1RTYyBxlaEdl3FaY00
O+oCyPqSYOkk76iMEEPEvleh8eiUIP3LSv8zHaGCN5cyPcaXI1Sz1k6ppFaHhzsL3Ld5AhfUS3yO
nbqr7s4QlXDZu8WqCkytZfr3HMJvCVmRiVeF8SmNfuPF2f94Ms6M5YW3t/qhHsjMQ3GJP8zz92SI
dXiFZNtLZOVPSq0gh3m1r93ARRsV0nhNQWz//1o52398r/N5GjwwTSwGRGGzzSUawdrxJHpoYIUj
Aih7ZgIJz8jXAeAWCdFU6lQAS4QqO1eu7NFOB6ayyaQ1FEuc2TdPXBSqwKd18gMXe/m6TgE5EhY9
qLV75L9bFrnddnDgKn5cpuEUuqY8Y/7iTPWH9wd23szAFOpCxe8Tu16l2+dLLPF4gfKegsXhNYr1
94fVAw5/JkxrtudaKuK5Ap1owCKJootbnljR7pmD5k74VZV83+vfCxhXD12bCF1NQ/oaQRuttB6Z
o06jys8rPK8k6s5ashyHyg4Gb4MURrFwpvc5+vvXaRQmkeKO/lXsoCOFka36xdn8wgiqW2rOz0xl
Md2CwvLp5RbE/ZED1x1O1gsc8inkOu7Y3E2FzlciUmUB4u/11u0d85PXkz2yZaNSWt+nwqWiCOV1
vnZ6FPdshABjmScpqKbgrEjZXbimKlQr64I8TM3rrhP6XBF/t74MXWDPgrumRDzEX2jJG/HAs5Y1
0sg9t3qM28r2aBzRL//w/OBKFuL6K5nEofwx/qeH3S4KYxIvg+g3QpGfyQqShN4vvjoD0X6Htsd7
j7RFbsCJM+nUY+8kpbcHGi/RbYQKwPFqPD+93R/98CjTDcrGOHfIN5w8FEfwB2TDOGXQ0wsnbMBv
iTX1FSFYT5wk0h2bz4sXQJrVPV6NQkyqEMvz0cBCfZVFyvFssuj+eSt7BBBPOw0KOL1sY5K89SrD
FMESqV8EZt9KhO3EtotXs/DP2ZbApxd2rh9q2NlXBIKG4slJ8Ywck+9+yrZuz7a1D7kbdaPrc23v
rg2Ogg5xfgxcBEK8NC1fjtrk5I1yAbjZ6pBgJXo4TzQd7QhHbggyhovElZdLhBGtRECHqFKaqXpX
3iQSZV0nu1c65jB9j0Ph18JA9virS2JVFA4VGYyA7r6iVWhHEDtAlbUl6nb5QQ2G1sTlsyx6Oic6
YVJm0rV25k1KvnKWtf6JeepT9bxRDTCH0MD+bf1pVSHDC5htAiVV6mREBhINn4pci5llaVwcV3m4
ZbKydIbToG65kecQUKGRDvKUqvFHomjKBB8bwDJFaHk3+ghvd5FgbHtxehTUkSozjefYOXRmEHa/
tGM2l2lDh3NlzAt1avUo4/wyEX6mokW3U23w+OjpexxIiAgWY04L43kQiKnPTE4742huSv41J50c
zQeJ+XP7fJcRxdU3Q10igTyAgcH+X9g047CFuFjFio/N9tvc6SkCgX/LDOPKDpYsYGUQ8CkbMVom
g6mEmEb9qrnlBOAohtPqTfoH4PiVS0W1IzppFHGKYWB+kQbmBDW+nwOqiC2liQXB1YXYHvJIRApI
9VnLpqrneFbBMTM1clR0JYRF7tGP27cwYHC7nfSCukEnjPu+P9mt5WCWJv3fAry8sEVbhItiJzzx
4dWZBmQUs8d7rBnTeBLY6j28vabQXmCYf17vEm3GQv+ldNJoQ2IizRGYIEghjsgDzelnlDmt/AUM
ePJuI3zMlGjsg36EZzJbFKaXMst1uAc4azmJBboiWZDUenN3BS7bBAUHIOQg8bfBI06AG+mkxhLt
g9s9YHpge2Dhzr53IokTNu1Mnsl5pGFzvUNGTlnmSY2N6qExJa0qUMzyaxKWkyNQDN/CbQrUUibj
kWY4qt/IpJWrznpcmmuo5DyVbEL+xtE+3jZRcMQ1NnIUsqiV1uwvdYCAAplYyo5c2keeqfvV3GBW
FU4RYOzCcVK3/eyOtceIpaLY092nJGqEb7/Sh3GynOgKRXIA/2u4ztjbQ/oi7yRoEDjT00ayiM/O
aVx6wIDDVPOF7vTI/g0GEMBWq43hAawZX/Q+B14Q3Usw1NFi6TpEwmMCJKVg4CiolhKMOg6AsZXk
+Xnu/pY5EPTGCSbwJfhC4G9Lij2yqQBB1MEbosgGaqPd2IgvsiukGyyFBPtF1tvFs5UUtctXEzg2
dzM1UpZ3+OI81RcKGSO30jnjsaDuOvo3yYf4IRP85AhZKrA8yiBjPeydDS7jza/Su+ul0lDHenRY
BGDeEwpOZMGBHxhbGv2v/bwcYuSH/f0KxuznCmVswrav9bnvOdCiGGCiTfdF2AcVA0Xl8wPFMAx7
4BgJLPEPW6Y4LfQoNuuT9zIElRzN8N12craWMXZdY+I46g+CpQWzkDIiw0LFJFTGW6+OhZ8YvjX/
QOPUin4FrwGU28NthlGhv2vZ/DCnFV9gbyIvdnnBAPlCrVHMv2Al7Fl8AobMIrqsfuBUk+QGVla6
PcoZW433NKpwloxCGTbO1xDB7GSRgvUEtdwD3U9ldv4vPHF0syqd/PTTUeAtsDE2L7mhpB5jQt+Q
PEyuvewH6frTRLmtG4kAnOcBwZX2fTq89HR+0/el7AcziqYI7gKNogtuvPywrwfAoop7crknvG7J
5/tVLn+fk8VMlqSYSoSHimKD9D7TEzGKRG0p2XV9RzhrW3486qZzs4PDUEdk41/5AUlDhDQv+s7A
P9dhbdkqT9NvnT7050dGUxQ0tKHWsA2bclOLsaVja25PZmGisVID3tV5/0vu34MqPTSN16CpEYEA
JWt4eemT+4+LQon8OPSQzetPWrT3ujVE7EQExHCPvg+5evJ8VzE+EERIdWagm34Nn0sYZd/r0NKu
AcBaZQjO64KDim8AI8iL3lntZvHeN/dyCke/DF1yP4c2ed8g2bEMIl9yb7mGz/iGfH9j4mplTJxV
bd0qh+Nr0wKvE4orV/GhK6JZ1/DBB6pXEQo4DpeJkfQ6CVoEULL84lkOtNhTaQtXCKKeHiX/I2NH
3PFfhZCaFzHIr/0o2pN1cWzCPdJFb6F3glSzXQqHBlPgAGtHw7ugMO+ExT4pSCe8MHFWvRDmu5zV
8YG8tk4QMzlk029Z8Fh4YdAaD0ghaMe8UpS1i03EdDHhGVOMobz5+T6Vz9dxE/d0UYC7mMKTHxBc
B1hNwdkz2skeLdKRoFRroC3stYqfPeHOM0elgAEhxlG0k63TDE2gO916WHdC3baTkiZ3EmpsEMyt
q32yPY/tPUWGh37NpSUfT0d2Ut3AwbRdLGRRjk4H4vV+XkuHHSxFoYk5GPJrgIuWAjfE8vw3LlgL
SLABPEcnhxW82RFI0BG8gt5sJof2vG6Z5TA8sSP01XcWzkqrC0MgF/jP2ruSBuG8zJ5+Y1nRc1vJ
b9t+AabdNuXE7tDuS+U5Z3qtxBDlD6rRRxYniNAkpl2KlrHqqpeTVwFhaQzVd7ukruHDvGyuTvB4
x+fOHcNAX4fuNjSVZ0hGOj+fBKl8CbgT1wyq+2qqySrdcN6wz4Vq8nop8mzLOIcHRkCj4nxlmr0I
g/I/JlrKRxDaLXwBHaV12uAHr7hHhhJTlV5K/zH/xjE+EWgSyg99D71RM2F4lBQ+UxibbpiVgMM/
01B/9OfkpiheSY+ZpC8YXSemjR+U0uBejg3obx+YX/fVyo/MzBdLjX0OM0WbLLzALV87wkd6xkE+
Gcmy9aoi6EHw7Yf0tiSrhtYD4nXKqzM5YZMJBnSTMuQAI6r426GrNEMhplJRMObCAEJfSmhgLCx6
AmyFdw+Y+a5V5tq0P0xYyZ+3K8WgsxEDz4Krd4JMB+amR45EkRP07TGBQxkSKJRsgcpMoN+Rietj
DcXMQJe4UyTbUu6Ut3/zyMDxoTr9CSwvlKleZ3hYJl75PQGwQFymW+JKibA97WEy8285gV6C35XB
HK8ACD9IVeVBVLemCH34u1YsYUbXrCYjzubLv8bjeqOc29340dXneiEif+BR8vcPPXbD8VyRBDwc
tqAUqxmhIl+dXJGVrZrFRBw3HpYUOy8uZMIm7sMVKktUtOgtNysEJX1eqHBSat5B5Xg9J3rOsI5U
mkLNRsHqMfYkq/YndTAQEGK8YY5SezYQ5XowOOqgbGAjZ+J1hERgC6D+YVpdeE/S1rdADF8tAitO
/RS09hP49c8m/0u2CQreq5+mLVrOoZgwmKYjEIt/zAbtg4BcUgmgekE8eDkWIr7KZoDVkzQGOnN1
u70AijtXTqVax/UitqO5yH+5cfIPZUBETENSFHUNZ4EC17rSWIFR7+orSoGRFSvw/+yMV50DRhIF
pm65LDnc3SGSjFembEL8qjgiDNFxzwQn2WiVj6DF4r2HRXRXTaOJRCzoN73q0yU81adyXybvj6Ea
rYS1wVF6dtX+MgYnuYXV8aPdsI1ChzRgfQVzsQ75Z3OW7bBtfXeOk02i6/Er/yJ8oaYnFJtP8e1A
1F39ZNcR5SLra2wBqaMo14mSojEbgefEeMIY+SV0/kGNlnupcNuFquyYbb7wHzQAjvDmsuSR+zS0
XFuq+lhj0cr08mc5W16JbR8vr6F31DoBULX5sI20F1BHFip2/EHxiqQ5pIRm2B28sgZFbZIVljyV
42bI/FgBIvf6eEead3N0gB1phmz9QabPQm5BUHmeXd8qFsjqLMpyiDJ8DQcJeZME1JbXmLeE5qBR
qJn50ty75EHksiF3KzIc80Q7Uj1uzQ+NYXEJb64Kx7oai00dIS7z5Pg5qbc82qNrA1K9t6A2UoMV
tWMeJ5kx+ZH8IRC5+33UFpVDoPatuW97kJcZ1om+XkrE8LsYTfsFtIi62t0RFjEyddBpWh8wFqe4
4OE4vH0ETehCKy+zAy/uRQpdwHy8GcUyyeP/BvaqCwav/bHHN+klWUWxnc1s/bEV2L7BjnCycawd
jKY1Ngq9CN7uUjiisHmtmz6TP7pk+/cdBKdhIHkazPyKML/4RmMb84xiIW+z/hxZAZU87rB7woML
iUttoENNcjMMJPM7ANTPpXfV7N/LrpHV2ZrLadJy65bFaSTjCpINkPDld5+9zMVcMQdzL0gqZ67d
3x0ocwPNIcMCBpJiLVDXMvEgRQLLA7EiqRfXROyC+bY0/cp2qdYxlAzCZmuCmEU13iYxH6CThRUJ
Cx+JIW4M51RIM3ynlT9pf91dZRjxoJOlVR1jUjXm03B/iTzlzaF8gmXFoQrdfJYNxulmcyjxqzum
oUdK7mbiE0oTtgMYSEia96N95pCZEZ0gcuMUlpuPU+XU6VPLGZqnYc9YGO/Fubg6aFoOsURnes8n
KybEeAiENeV0eDPGvrGKin7CoyGRoI32WluMmhhtK0k6ynOVKv+a4iRHtDAa/0o4jawL9GcO8rax
UcrS30VeD2VuuPDgiDPzU30SE+2vRVIpDm6I9W8F4v4F1xrPRrAw800pC9DmPWLfnUmDI0uDz7Gl
ZbY6CxyVtFsh/u0m7ZGycG2rzyLWYR8GA1kcpRGEgskhU9bRDqmOJvdlTCmUqMZkZyw/rHStWj7K
br6GvfHNAR2n9ajXrto2xpt57efybGyyNOw9estPiJdpDtVWP5FzErx2JCV+VHq8fIcZU3eK7Gwr
F8zP+4RTwhfFDEkZ7swvhcRAoDAKr0V519Zb6g2hSNudkDRQG/Uk+qfLTmQg39neVtinTiHv0bic
lrsq6srDZeXoVBmG/yRmuusba97YEW2eUbfOf1969ZBEGs0j0z3TT1/yB0YA/A7OYtrpmQld+Luf
iZH5Ul1rsQNQAmyrkNUBO9eCVzTZ6P9BuSgdbdngOKR4L7fVwnTjHSmT05aCfy7t7C9pYVIbFBxp
5waVk4Ff0kbFz2wpZRNt4B3sZekx5rBWzpvHPnRM679BaR0bqQdlYULnClgz1LiNI3/veip62DvY
cB6JzNtrWxeVMrGz970dUa1Fiv545iJaWu+yQ5OKrQoGzyvY5DLA8LoWP5r5wSlH2IndW7atZndr
R0u8E8LaZ8j3smLiVK031gpG5JiNz8OfPfMeNdtCrKeT6S8fxfUNXKJnNMcPqHJgqsfI2z0F0ICK
1I0/xjCq6P2UsZ2f3gYIGoCsd+Ma6AEZIbqamLoXNP/YV+yRubQidgwH2FcKa9R1EU1tSsz6E5a8
F9lapw6jdNKKMf3iTaaLe/5MkyyLyGwVadu1W88+un5E8iXbFxrmanXfpzoXrX4aAekWZBSIawAb
5gGMLXJSIMFVBmOJeuETsrBmCShU0BuvKsJ/u6oExeIO9WIgacgO5onBmJDrzYphQy+hKxL/lGlh
sV5hIJ176ZDy9XOgh6nrgMufH/mhDM/ISlY12z8wB1sw3e/Y6Yxg8K6E+4wQjArLVimivI0NvaAX
tBrr6EpKJ3JIo/XNygE+0m79P8VVunA8JFmFR/NP2f0k6mu5KEpDewDq0c8cX+8KmMMZ0NIVqGV+
lAU56pxwQZ/QxdkIYWOY1cZFNLXJHpR75tZvRcRLNFLhggr49qqAYjRhXmBIRA39uECQv5QUr1wy
5jUYXDgItjUwIu8CsDjOSixXYVMc0hZVvZ7n7GWFwPakz9bfwh2jhhHCPUcVbpMuwCn6+4Y1gxiM
4sPstZ2sPNAfMbI+iIkG3yJWeZaAqwB+rYi/5BI0nWwi/YJGpCGFGycLy96cmfPkVafdMxM81BKt
UwsC+OIjBGISIK20ye3XGOZfDV+Wy6ZvJKZsKMUImeEGcwnd9UIgC3cNfZxtnWbiMgQ3lYxF/jsZ
a2/Pw9FO7FstqvVQKLtaXX7t0Wbnjf0Xnn41TnJVV1RYPq2/yoabSwlnZPPumZL7yt0U4xdiK3d5
6D77l8hzUH67BBqOqyYCpc5v+HsDmzWy48sw1VNXHhgE+0UwZ4jm2kWa/Scq7n5BJvKyfz+RLK3E
DueAB1PJxMVNayIOEONsJ9wJcOxOQ+c0/UAlHYYCkwrxPtIDXWeSXhamogxD4d+MLYIzrFj+KGXr
V4AjsmtlD1OK4kOKGly0LuiYt39BCEPqA9MZaxoQJ7I+E9MLfDNz0TSl0qQHlLc234wgAV/TdFk0
8bhG/EPRg5lnSaeQ2N+xGhfABDuscJMZJiVM1PXtIjpQedc+aZ6sx8BpRK3Ciw6Ng0TguovlBp/z
NTSoaGSzHvaq6axn9QDJLIsbEeHk4DBiNoVwGSODRvqcszYGvlisSQAq2Nu1CMAciIGSARf20P4b
/syCi4CbGlnvgkSQVTtYChY8FN8Q8htc1FPIDGjnJHe1WNVUgWp6huU2j99XWEK3szx7eRvElZfA
MPiMgj+vDv66baLa85EX69oMP0hrEdy9Yo/BQQ8I8/ROWgvIirBvl/cT1ej9sSlT5zb/wtn9SycA
QZ6iTQBzcmensKLp+nvoOYuOnLNF5uWVi8YA57tEYcbhqC9GADUQp36agctEaQGGRgEa0tTGJVmV
/0ojqZwZWgl5qZM+0dKawVTt3mhEmdZexgmIceNkEAZAUSN4yHS2WU1DVX7cyuhLn0lP4TtGzyhV
A756az1lS/3z0TMG5FWs0Q+IylpDctbKIEiRYzHECjp/PdQ4qbXO7nZoOy/c7jHCL5lHICJ9WY6J
rKZuP9tkqC50v1rlycJbxCc1nm+w3NKJcXISBpQ1sjQZY74TKivOYbOWmB6c7Ci8O/LkbkRPJlSZ
SW4h/I85CfQIJ3MypaWR2ijK33wawwPbEJm3euCKtKXrtfQcx7C4PMe//b3JKOt9sZFAOiPmZgY/
j0SCrJmPT6fIwQjxmsjc7HriU5iueHRxuBIuavQ8JUpP3m/7pANoSiENCiGPTfw7iljOCWrceTXY
s8t0NegniuOp+H6GhnG2EAnIeIlcZVHtBkIv/1YT31RcUROA6YuA0uUpv6H3EikYfgp0CQxD8Fnr
Qi1zEX6HbyLcwgi7ZN6fNr0d0mHNuXyMUZ9QFoGaq0SgKZeKyT8FK7Ekfz6Vh6ZHAjaHVwDM4Q7V
wD4FEpDjaJDDSqBG+vWQTB/SLl7I/NpxRvSU7RlCaZYNUoxk81cxEhP9p9KX3BLz5qLFlGJR2iUb
Pagt+tyPfEDbdbsSdZ95fdMxWc2ME5L5EE5iqDPbuyeNQr8H8eQgKB3EEHHDmTu/lA6S0twx7Gsb
yutYJH1fnaV/Jzmv9RS/m2ulOoB9vtMAg2Sg0zw7Pl3/0wW/h0PkCQBcVGkzq4KzfRviBrKhcbOs
Bc9rJWQ++40ZmRSoATtw1du+0W4cU+TzTKKOJ8nrkLBrQhZiuzVL8t3pL6uX4qunHonaS1Cxk+tJ
GLHVvQqXYmE5kjPV7dVj8gH5BN7uPj3BZrp95WhD3eOFxv2zicguIs5YF3nYENolO3aUBlChUVhb
fXp3Uynr4pm7fPPk8J+cHPG8u0Y8Ic9M7Md91DIIKZSHn7fCiAbHtQIxae+KPpoV3ryvgwnFXY9V
Kly3S79UiFGg5GUUPk1CRCQfEuHFVOIcROH6na+aD5reMv6cByoaRllf3d+HRBEU4jRuWxp3WRGN
1Dpi00iMThWUCdegr+y6T/xtUq/n9h1NP0W1myVAiyZ465bjJQclmG8waarF6WiR0zUzST6FS/NN
DQFnmAYTT/YiIP7QlTXTc5UhCqQy4wYMhJAB7l5J2X5dONn0Sd9Uc0XsKqVmf7wuFt1ZZOztp9zp
OTaHp97YVzPIiLAn2kxVGL3TmGTJ+qFkHHjW+4i0vC/9fTY1B8Oj8DuAu94LanR6NMTN1S53rJis
W9ttRhZCZSdF7kqW24GAoJc4zb3l3EiPZKFJOF2+ocoKFRm2msqK4dl5cmBUilHZftPAAjLMCd1o
PSdqnfqe5KU3EgHhP4pYsOogH8a12Is0BEQVIhPw3rDTFZM8Ec40sopP6RXJWu0qa/3bgOWXlu1M
fu1CSGXI41u2dLnHT9gkLXcx2nU/kIn+iiYQKZXUi/ao0dOihqywP870/34e3eIRyszkTEpoFwNU
asQx6cd9MmYhVejAxVFTu03jwRtOBji6b9MJQIx4q5JqYK6fKMiQUVAnjxh7WUm31B+1/nM1GABP
NtG9WUNfnxWDlORfZ0OytrjsX20IJ4DvJoXY3Wx50qwPRW+83veh/4wgiwOe2Wlr+5/T7UMc24bM
4drKHCkSk6jlC/u1NKIfm/5djgovw7mjJpvBaDJiuXnPsw/PjQ7SC/QV9jfLaIMEXCJUU/GBKHmD
UTwHlMIAIIYZstJ++Avfc+uU3xii20TDX85MDtnwAas8Vej3bF0uWFad4xvNl+ytX6374rVjtedj
1C5mhHnk7x4cORsGV20jZhfe/8RGWEgcW4Bsv4ivXVrdBKjg7E7mOWquHuY00dwv0SvBH0oev/kr
z/zt9s01c/UfVO7n4kWijMoZYQlYNE/AyALxuoR+hrKrmraUR6qu4LUB1u40NP2/UbVpWFxu/Brr
0lF0MASHmPDq0mOOYaeq4bVqPeOvZXPofBreHx0SBNWQ/rSCfqvUJ+fssd8/kOazO+BIBF7H0Aus
6ga3qt2WBe7zdICiG9wfYORWwTJUqwRHpSVHqGsQIjQrvYaaUVQoNgn70BzdwRg1VXTVLqm51X2D
W62+SG6yC0pCM7WN3FIMYnDbVP2Q9cW9S/RI0I3qduiK2N/7s2mo0SSkBVfRGaIUoUiavpm6GfYb
R1gIF1U/PRseOvXvUq901O4J8XFYQb4VraUnmKdZJjNb7K55QXp2ZuhWkjPksvVKVCdqQuIiqP1z
/LJwLERq2BXRBUnLEvOzWVK4OjZaMP8ah1LN725QVf1xRPNyWRbTDbCOQ1mVL5xd7e4snqwViq81
43+XR7SMVSWpWTMqoGDb2mXOPrIyqnrQ1BHv++NjDYlavh4c4yC/Wxp4Yi4ng1aW4pHeNtlc1ksM
U1cc17HJ4EUSV05ZCWZD4SaT5b2SXdSSeIbePZGcaSNZLTKBDhI0+qAuVje5kz6IhuTpQPgKRFHK
KoBOc1mE2dkQqbCgjgPn5Yb4jITFLQNhmseq/a1UQCafTYaW9K7Ddk9shpEF0FZFwlHQMm8YC8Bl
BTfMCS8h1whZ1hwZEfo/b07X1d+nwqPPaHwLKaTI0q7HkeCSp9Y0dHUHMFmd/zwktAf9LajFKzKO
E84bgP7ueqcr+0B+1IfoS0gLftCrsEo4J47QLfpH6WYQ5YE92lHLxPTk0lfxemky1IVH5NRz4k8x
TCpDNI4l4tJODjG2N8nR/Vq16/FJQTi4IJl4InCxKZj8x4aoWosv7EOKXdx/TZgYbhOgwwRWVxJL
Dne/VBofB+L8SoAFGYW3Tmfj6n/RU8M1RjthsAkb3DJRaw1vudc+hsCU5X+UscqX/AwIl6AJ9ird
ztyMXY2FGreFKr475Ed8iRRdxxa9Iq6MIzrDeA/S/M9X2LUqaAEazLdjmV6Nl0uXuw/xKQGZVNEq
Z11XerEg7Iv0rCno4D4tKTTsXFN/pIaqAWncaVRW6zTB7nlll7kF6tsth4JWsglvqKvfoZKGkQjQ
2ZflxiP9qKQZlrQmxlE/nK90cUVrWVYXj/OO2vVkZSWm+XSvAbVDiXvAJ3L5zcxgro/Df73lWk6l
RNICttujgoAFfGK62bFOH2vI+zrZJVeVwDI4w3gxrtz8pciVofUhssOlFQQRBOm5CGMuKyYECELJ
O6nE0+qecXFaq8ochDpUIvHZJJoIM7IcDZ53P6unP1/U3e0RLJUw1cv5pBNUT247NhIrSrKCmnqJ
0pQLA0MgSxFRMmmGyt1uABdy3pe4J8ELsqV71VqDFUB7yXrbmcbTjPuBMgQSWECSEXJ88t/pRtmT
ECgQpUXJP1Bwc3NwtyzC1P0fXYNjQaJd5eQsIUdjlKuvq+TMP7dmK2cZ+scSXQgRj0Jq6+DWfkIB
vzog/yd6X1XNrVzVGmawdI2YxLZm+vUfCBu8uecDTBroqJWKxs63Hytej8H2fK0mQRGJOHLVT6g4
D7LM+3gmkkkVnmyLmamZCK4FRSrecub2JFfvyxdzYcWhmd23fcjxAmQ8kwNWDZrDbDxQxB4IvBjK
VuahOOkeoTBclIpWf61sOoAchNiWOUduQ2XonVSpw6EbdW0m4+QDjQlpu2LxTDpSbqaa0WpYCjHV
K+FOr6UX/XV1MgxQpuIc3Hc7SLX2Y7bQU8ncDsEuXYCgpS6NcImSbfpzHwaPv9Po/snARDvSRp+b
SZjqZ0AvE+GEwUi40GziQh/N5sUM5nosIs8iLsRHWRoVhBDy/YP9DI1xHW6QKzgLZxMJQdV5Jzyc
D4HVf/IYE+0NaORcKsFtPF+Hc8OIq4ECcrr+T1ydX6j7X6JN8kTh5evWmf8fI1l4ysmZ4F1NXAWG
WodKKyNPVb9HYMHLDy+eOsbZjs3S8u/24TpPDEvYhKsZhJZXxYFa2iLfIb1nkT1hE6yEH2mhX1wD
cLqQxpVNq+JXv95wu6Ly2yi7lF5yvj8FPeqfEZgsg8e6NtiqWKUzkkzt0xt4cbWV7wMAnVj6dGnQ
p2FHE4vmSX/041ZVmAKuWCYQwKfDyWDGbBjhegnfK2oMerlIINHqC3oCQj1gDxMoNs+EPUrDJc2K
JALXh++FlVVsVI6MIvYibKtS4Nos6OuieE3BKWAxIpo0FUq6sHG3lbFlW0SPRq9Ww6mbxvLYzAwV
DHCzJS3OZ3cu3nbp1H3Sx/uTEpL6Wsyz3DyxhbQdWMlkyIuBYIlRY1BxCt6MP5sn9BktZjy48U4s
zZ23IXfsjpgJf6/NHW+3gb+qxnKoHc1xcBu4tg7ray9YAMDmlVmOsQstCebzh613QuIa1lnqp2eQ
upkwdo97k2gKL92KMEubtxtOw0jVnWZ/iOWV2Nth3PXf+Wvk87sEvDEtcCr9iv23Hb1qVwpkp5Hz
ZBpY4VxKuts5yUwhoJweT1jW5taoWH4dn5iIviKHbb2RV1MYQT8KZ14fNzhQj+f5S68q+qcssD4t
dVQABWPXqdZ7bsOMoaynpfY31/ZdTGSamboqz9dhlUOQHsYgR4UjxRfwK7rGoQ7uiNakcHqGsCrJ
KAAn85V5OK7yLRxXM/uZKosi2lh/gpi2LentTSTWV00PXm8dDYC8Qg98barOegWdI6pXMwd1yV41
MNln0eyuik0RB7ooA2sL2yRbt8Q4YZxNC7hQb18gTVX3o6+NWFKWK0wQjk4+6jXNwCIqzfyPihYs
EA6getayUpMBOFiNkGOOenCOpECqg4VQxD7A4L+5zwhf4tJJK1GWuYy4pcgxcAKo5R/qkaB+PdiJ
FJl11sabPjPMkkZrvnUFwRFTpboTbX1xTB6BcBPtD+oM4RyTZGa0rVZvLQqPGInrlanp94fEJM9J
vI69J0yoP9Bp4nnFb2mP8a7fcP2YOlXezTf3+PJKXVOB3XWnNF5lXIn8ki6J727EayDXXENVyi2o
ppRiHyFYpVK9GJ77O9R+JLqxspTgZaJnBGgFiza/UkJyexbIeedQKd8HXcNFqjNjp+AO+PmVYB9W
NbckLvYO7UFkXZQnRjcjKgWsOHBRKF8g1BUvCK6Fzhe6VQddOlEq5UYruE77bF8HqNr9y5OvQmam
/FnByOMVYdiMp4V2Ac4/AjrgCxXq8CdONREPuA8NeaOve9i6lCZZz0mtlIkUJ66tJOHSBTtY3Srl
sNuqTh/fxM4TVFjvUR5vkkoMzDYtujGg9kLYIhkN/jUJpAaf3eWPSYuVaOfla86JK87s3mOXvBr7
4k8r0FRPB93GHfwAuxFEdTUTbtkT+IUth1iNYRSvuKc/6YXHT1J8PYcG161G4JD8O4EZYF2EP4B8
xfmKZpyXS5g7jjPIRMneJO16TifXrXs8sGs5sgPS6skVUOSi3cHE0LDxooKtKkRLJu9pFkSxuZ4h
G0qSFmyux6zUILjlx7WiPwb36zrZnquVJzvAMMWW868a61J+/ZO549uJiMrvpb6Hd1TrxvYwy11l
wLLP9Q1Z26EVHC0YDAk4xFOCmcVcGyUF+U5W0jGbMSQg6suWisfohL+P9UAj6b25zSwSO8lGvb83
siGjwH0eHzfnil502YYSWN9W0j0iNq9Ev32CyN7QTCFbmoza2F7EP1KNFAbUnrZX5h2hsUfgaTNL
SmUt1Nwof3s++KbLiYuKBgNO8+Tmkt4kbIs2w/5jE23JQecUfPUY1O4vhvDPqxvWGvkr1+mrqjum
qPLxndE/ZG/Tt+tvkPl85WqW8kROv2jUZSO9gsEZ6RZzR0U1xX6w/fsZK9I19vNk1NKcjussqorS
47k3asULUKN2pkNm1M0WzFDUxSHDoAeuajxZoK+Vhr4qVLLGQ3HYW2mXI7wSjM2/useJA+QiQ4bE
4W+sCT0meLkP9f5ijKhpnCEKvdas7WREVbj3tPek4xU70T4fXPoEBaKYtJQQRbMBeSXgNbzbdRgw
KxE4v0Py4HfyZha9RVkRgXvX8WKrYCuYnoAwyBH9YIRUJ8J6WWvCwfvskDQgvscKisjLycqSLgyt
mwmbHXxAsBDinTPoRffrtCwxnfzc8uNqpU7XFxcoX15uoTSZZaAUfvax77y/SJ1KRvJ9efzVUbzb
+X5h8W1FiWYZTM5ixHVTg3QyQhaK3kkdptEWWi/gSW01scAW8DXg5wHYCbOX6Cv232rE0oMBSR4q
uKX7buG3xRr9r0vLS6S3qDXxKvVVFaU1LxVJmBN6htWJxn5bvzjwY7MGQ1P9MS0ub7buj6ADIW0z
/LdpT1eDiIgeX00oDHCtaOxU4tQi+z/P4qrHFUHMpBStzOfU6PxA3twnlC+CecQyUu72BM09SSky
ifkyIVOuqivOQJnuy8vVdL1uEx8wwq81wK22g7libNHhcJztbzekR3n65pTOycj7WlSuW1tmD3lN
2TyfmKMfsF72o1ebtrk3DncL1J2PRZoNpeTXfJpu39v6HKDOJjoJYKnaUyD5lgb9eXBQTqd5PGV1
XBudFTZESOD89Qt2K3WJI9HNAUYnE/pjeM4ZkxeK7nKpOBi9PN+xUB2YVZul/Wc7WNqqEjM/q9tB
KFoOBaWGq9gbE+ZCqSZ3pqywCdSs8YLVOJjdFiQ3M9416ARG/7xbRAAGkNHfSFQ60O47vIlm/lRJ
qzWvdy0h4S0aCHPlqvpdhnybmrNmVAxBwpCY6Y+6rn/slxSEyc8CHmB7XuDvQbT/TxewuurRK69R
mVkm6MFXpiyb8omphkIzk4rZV7tQMAFLrO4zINV8HZ98rQo0kkVoS/bvLs3nTBlGGyuMtz9KFLEd
1CAQYbos2loQExgMnxbJllJG7hQgoJqthUcdddqdZE1q18hODvKlqGaLg6Z3IN1g9kx0T5tN2QYW
3o12NjMbFFnBxLo2PIBjT810b1DTUG1HvG1+2GGUiXTZbe8eua9PAx5N2rCb8sm5KmGHPpGpa9gQ
sSiTfOR7uI9Ie4HbVudxjhWj7HCaS9qh0zF210g0TXP9hMf23JZO4l4uGmBz7JI7YLD3afcKb7MF
xRMeA9hcOebAwvF951QUEycv3T2fsPIno2rR4snmYHSsYbhyHVCLJdAGIhJl2Xbox2oIX6qKsBnM
7ex+VKxN6B05s1lbwdV+Sk0rmqTf8mpaU8J5p3hifr5ZlrQd/ThskltV7traXE598ntBv0aO5j5Q
zl57hx4HRfqQmm59FCwrHlV91Fk1ci+7PeA3zB9q4WZ8GFzcXtrxvEpbnr/dxiYhYu8xSK63QIyf
D90Pn4lSO7NSEI6twudzGX54ZBiEJc2oc+Ol+tNlKDnrB9QylqUgzS46RIpkLPb98+n2DcFEPXVy
/z1/wBSloCwJEeCnLC1br0sTNfBcI/KdkCqM+SYpxqDDqpPm7NFrls+EGgZvcJN46dSeQA92Q8Gm
kP2ZXHGT74pJqZIOpVmwCge9DgRrUom+qeyabSc6ok7C2zK0ud28Bt3MREFWw9qMpLtCXC8cSBVy
sMvXZUcz9NrMs/VBcNx94IanWOfpjGJj11AiJ8bmRLky2w/Q8bhHwT9VpVK4BdbOUgMu2pYIXWHK
Swo3q81vWUrkZCln5/cv++OwCdhg+rkf+OLSSyWbIoO8CAAWemfa3ca77h+uFjtntOhhcX7eY+aW
evbzsQcIh9LwyIj25lhRfaeLk1Gfijm2CF4IppdeHW6cfz7Q2OmzMAYhe8pFl4s8RZWD+W+OuLUH
Ea59APpcSLhdzVUpYzz3bw8uy6U2Y2J00oNbR4tyiV/g5ZPY/VCKwjDiJEzRDN/xEUneW3Trghfz
WBzafq9TXzA7n1cVxuq3pctyNFtHAxcGxxTbH/jibRtntFyuXCUWZDKzG54Bna2y0NHc5iXJ26gA
3g5cX73ecl5xPrSNzfEmrbx4HOaiqV68DrfkhLRr4YIZcuBc7llZK6+tGB3XMPOojF3oSylfQqGu
SlR4SVjp3XAAhUebeLQkAYBLFknBuqt/G+0U3BRwJ8FS0GF4DBZsVM/CdEjgRQcwBRcFiBqfw+DN
2ycuRRuQPdXcuExvsq56WYdkWR/gwKFn8m5+E5rbUNdFGenFs8SlIw/T7L7i/7ijOjRJNJ7Ehwdj
s3iL70A6sT93POVtiLqkFUWSm/UpGCyree9YsEctSSaBVgfyLVYX4AysVrNIWzO3iN6UNx3EOmXO
M5njNmvBCBh0bAUHV2Svtyr+xxv/Hnxvbwp5d4vbtEkP/bSicpNyafoevDOBxYnBu4xHLk7LSJZW
PMOgcnGE023a/yKO5xEKdTifLqd18xkM5c0JI8SV5zS2rH2qucO5btyh/BiXMZMCiH8fFTVRtdOw
kK8d73/F8SBijCT/Or6GnrjKDstbaEaD3DsBylvibInX0IN6mXrgFCddhi+jMkHYKNREPTyjgLSj
1nkin1kRfdHPqtJNG8a1D/3qC9VpaCPhsoh1iqdv2M4du7jRRtdkRglT5/rHoANIHw10mHjwa6tk
FvF2NtnGP+W45dImXFXfhRCWxk8JnQAjeDZTShFvDxYXRB4AD90VNaOGih5G3CB2LiH8iTF7+CSF
iUWWT1X3eRFfNjIx62siAK6QfrmmKz25JUyQy/KG52Nj5u9L+yThOvwEUO0Ss/35TLXSuWF/KkHF
wuU86EcbMyHh2q+YN0/7FnYhfsQ9+E1pMWQ3i6bY1ru7xm89PmtZfyOAwBpFp/AKZLBxDL/ajNXe
pzcy54h47MKMjFXlkgfdWrt9A5jN8OTHPMacM6ZxId/28WRU+FwpcbviaSd+mPdOvCfmIr3pmgnS
Capt2Yt/U5qdInHdA35WF9a4QY+nHQXIT5rN0QGDkl4XOHK1f5dzInGmF3cyaJ9JcfWOcmukNgrG
lYgDZQyNas1ChOmq3uU1JHsb9WuE518XDwesKMVKP/YqQArgurrpYlXO0+q+UQnwFKP/DofBPoDO
EwO1Za7RCVkY4Tvu8+9aUTp3O0tFKnleczqLe3G0ElGPOMje+hoXUPKu/P/X/V7jyDVdh5I8hbS2
GpJ934IfFwWz7zADjqYrubmGWiVeB/rCB6mNROG0kh0yO6Rpi/TzQoWEbKf56TfChw++iSOS9IxP
Cr7iIZhcjhVppCS9+xvAlXZO9d1lM9fqGbf3Gc8jWOi+6q0fJOS2ou3K0qeImw/t4rJsmXTLo1q0
JhyyvFwIHsoyP6tSMlo2vSShpJoDlTjaZ8wIfM4H/waUv6SzvMV8soLkckXvVZDQmNb9GoRy/Bpu
mpTFLs/SbpQhwj8Upd2980LVuEcGP8YVU/hNqsmg/SN4si6VuynYHB/GBrGpc/p13IkSK8Jk4TLu
fopuGWFhvzuYr7FkH4/TIegiP/M1wZVcV2y7VyRTLu1AooT+y3wPCNl3m2Y5Ww+Oopuv/GzmR/dB
SbDslTx+biB//2Osjioql8sDP6YEDOdhXrnVnmBj1DdWbiWkrvyEKfjaHSPsheUlsIMWFVX2yw9s
T5AWwvuJvR6LXmrGu4x2Dka/qRKWl7QflJMXKSO5tmKHpPEmIePTB3T3Ea8kbIeERIH9hcgwF3Rb
kRB+1NcUvEvfGav7sfBmh2gbRLcei5ap0VLBtcaI0jI1uaKe1vdJg9qbZZi/tg5MrbVp960sdrI3
/cDKdcS/pZZrEXojQx6AoZ7tpN6tlW5V5IbZz1aj1ovotnU8TPMrPWW2aAItGi3u/rOyfvRn4JID
qbm2pj1UPGC03v1/mxdFstD/7OBxSnD4vDn29yzhHgQupcoDCbgqzNe2qFUQzcbfOfjFSJVhWJgP
o5VMlzr3TzKzPgT3ZQwrEOmCuFguaoUIVFfx+/j2pMN/yC7SX8OHlSpbXriuua3DLSLf79mCjawp
Q8snIKXPZYAt9lpzh9znST92/SUd+JEl9XZiRHanf2URm/UhOdOjhxVgxKSyiDqmGnnWiOGqNdZQ
cDmwXlYX+ZaucsVXqJV5C5cMGmt+FtGD7vr6jr/RVrbLc42l2XN7PCIzjC3BwB8UAIGDknRoJ1aD
jHi6mImMO9YBBblUOA2OfOsw9FRKvzMz3DLP/ugNGh4lc0KihXW3/CfU4LfeinmJWa/hFpquBYLW
jSmR3s63E3b7M1/1nhauGXeamyLRJ1zGHoHj/3bJhlwKFF4OgUO75wSGdlInvqSd9INwT3EQgT8P
ztRiTHm1GV4Z5Zu6GntdZMcb7uzNlWPCb1ARnHcT0Biwutf2Q3WbDHgvLO463zH2vuillYyg+Rwm
P0rmqOhjSFav+RmZEWgq3raNIRvq6Y6E99Kjm2gBSes/JKVqrZF16LU//9f4b2hDsMsOd3dW0Wdh
6U+GvX+BZdUnt59Dsvf3LgOCKI7z709WWx6TJ72Dc7dVcBBqe0o0rcureISGsAgYRkOpPULj71i1
IaOE0+HuK1oK/9CHc5aBmEn/g+MZ+ngjOuNNI684q+BsyoCoG4g12NQRgJHHKlfMxUgIcLSQZcoe
pQLlXnnI4rgEEo2vPjXq44tZKEt8Mra64ShYI2kPdLHiJyPztHx/hLEZfFY1WvWlDxwJWA8tudVT
s5uoYTAM3KLeMdUoLwX6DdMxqRbEihTB5J6cMyXSQCpmioC3REgctoiNWlDmpRfiV/mcnayCRgfQ
NIHPhfNy3jwmGK7NmJTfoAANL7wLDOkrGWxiG1IyeHOPBL9AIffhEiFs77kavTGVgb9N70kq9q66
Bdej/x2kpAMcxZ0fC6xDjUjIuuehl+oqcvBwtOjFE6uBmPxxs7Pj6RPO1TstbUKPwAkbEoYNqlQa
EihARE4A6XQ/5XIVRn2If8qULpqEpDzspxIUnCF7T2X5ipayuy19DngxhAvI1nsGvy38BlwHWgKZ
vV24DdSNbVOrIlU0znVmBFFNWZfLGAAcJG4Pebd7Eu3DyUnjQa0W0yXPjjk9lJcGyUJs9mtmzlpL
+fGcrW9qj9tjIobrKysNE9z7DbpCriDhgg6KEnFeqlWzyAWbAAkmX4956fFLqFP0komVqAtJ4ao4
VdkvDi3wLd+lEUWh7CCZgBwggdiMtk35vSLylmbu/ncOFiym83hv4H9Hs3ToYNrkw2O2rbg9B0ri
Anz8z194qsgKsWRGcN3Skju0I7b5IbNL8eM/ybCdO0YmyZ/LCj/yOYELKusRbBpf9gyNyLHGoDMt
+u/SrLnDcpdSuFrgVUAc/rqyZ++Fg35Fb8oWPruO/Qo4hWJhls7KXfW0Dm9FY1xuVW/FnIY5bm7a
IEOnPK9Ob9tFAbOIAKB8y4DpOFTDedHHQiFRnUDKBIyVQdeFS+cslxS6vKk8xESGzTeV3zoK+uno
YQMYyTqJLDb52lJAUX38qKWG115H+vyNSPBlG4SKbk3cq/LTXBSBDRup8yhVZdMIiXK7wRg+3dvR
FzszTvzgKv5hogp4HyvYvkq4f/cI5dGO7hUhpRQua4TKyimbx86KElnv0xz3U6ot+iw0fiNaS/Mh
827YTw8qTfYyr+JcpE8tfETPb0NlhxBcb09AyuSLVfRE0hRkwdxmsho2pOrm95SxZX1bAx4ZHhhU
QctamySMJZFx4CFBkcidjcQ2eMb2sZIDEGzcGF9/l+Or2N1YHq10/8qR12Lekb92SQ8dl5fmQ9az
NICLnxqw0Yel1xNi49Ck7gXuJBKfOhAhvr4vO9UvBxo/BFf+KNv/8qFquKdrz0S8QB7prom/tTPK
Lg6PNlfNiiO9D1D8P2HnElJ39hvP1a6sNmKJoUjkwMN5WXk1TPaua6CW7qOrLbISu+BJSEB2XTBL
n4Gs/Rq7PQHCWALl8UYYZBC2nG/L5bxCtrDoMuU7Ry1zPwSjDfblb4n336WU2YaH2LsuS2MreWb4
4PgRGgru5hpDZgiNCo8Y7dwFNdDSGbrsqyfvsQVj0G7coWzGNsDf1SIwqaW8jGh4oTYNUhtdTc3o
+qEj6f8pjC0NOCFRAlczZJuvUkUoTXfhSIsQe++BzyNAJTx31ycdFOkZdtAtoRwA72Np6DJDIIId
Z7vkAfj6Y99sDfiOlx+R9FdGCXbO8axptV3k0WZ55TwsJUrHEkLYF09SVU5FBSe9EazC5M6Bd3G/
Es3Me0zlarQ6Jryp2qTQDTff3s32E1wgH0PpmwbEVUWJrKxFZiphROKbANeULnGt1fuqXWYEz8yV
rVn/08W+/1n+d1/ToJJc+TW78Ozc7BU3OmMrAvWkz1wCcys/EZm5tiH4pNgIGxRpmQt4VtH37r6E
mo1HR4CjX1ozmmvseCSbmu8FLCmJt9Xph7cxjiXYFB35knibzwqEAzEBDvhfN4MoI7trpvtyPthw
AvPwhkQALVSTByc72ICtWLdxvYjKVHtT4dNpTZpYNc7DrQid50Lkd+Upasw5Z3ZgFVdot+rSzRzp
+J9jOH7sxfDoamvb1sbwZzR61wJT1NopLJRcBcuxc8ragiKD2psf8ZUszTCiJuE9dRBm+9zaHM5m
RnA9+19C80W3938A/u3YKVbWfwpOMyprz/HdsMuINBT4jxFjpCSsCHZjI5b6oOdaooz/b4TwRUE3
vQ9iJaWdVRdTSVofU8JrjGJk9dAWz9K26nH6nb0g9it7Dv3+0MUhesxZL/l3aIeC2w62SwNZR9rn
vXdryeQWtnZSZm0eeWTgcf/f763XGqeNMExYukLIfSIkF/YkyyLhlq+4qkDHM7/awplQSjQ0zIDY
yD+vMegBtKF7iCHB7ZA/iNKuzXOTb3jlduE5dyCQJDshdwyI1DxDDNU8foRaIklMfwn65iSV1yjQ
F4pNBC205DZsYbJ+j+V619uIHWwaazWhhseZgMxUpf735FI9zDNvM78Beszo8a6BD+UEoYjRqZaW
oVctZVWUIbNVSmC0HMauVO28ytrudaTSj6I3WQnoDTNs64Sd7Vs9UrHOJ86evwikypv1ViZSG8Yl
ZW1eEMGPy2QOxXBlA+dqWQU+bHfhdok2wHGZv+WWkxVodAm3Bc+cAt81KAQ3c3O9T4ZHW7iRq7mY
BAPnZTmKwsyEVxo3CBw7+rZ0o86nKrcp22EroLqBb5s8LnFsSjCQ27/zB3in2lMzDZYNFBkZUU7x
SZB5lXC4V45kZ685zgoZr81psQhAHHVfrb162rrJ1vEqbGZV7dCMvV7I56GEgWbkpsAnmhF2YTuk
kH40RVCJZ/pZJYO4nvsr1n4qILQj9NemNqJ+Mu6bdHDWXLO0DTimE/AdnsuCOpSAdvz4mMMsry3U
JYRDSl117IzHPO1GuUGh59rLDaiCPmzEDC7BqKZF5+PkgfqsHOkoMmnn7v4bfRM0V3nLvFtaxw5f
q+Zi2MJRtVeQc2zofJbDPZlDRhdL6wpw/GC2iDxVbpWZLg67D5USOUbo4E4F6KUoz4MFWsUAmHw3
JVPPM7lOSqF07h1DflBMkRh3QSApE7S7T55oQPKVrCFA0e3VaLf62OtsxdQsOGu/8mzeFmZJfhHt
dUVY8mu03as48lpRAoginkccEBdEcK2XFMi1b3fZukf745g7Ho6y/dpRIKWJ6QXfauckifDolhO9
F97BVSVMhfEJltm+RGPiSnBSrWPcDS0F4EZOsgPYDT5CFp5tBMvPPXDEBcHX71TnaHOGcN33fpLu
pV8dK9B+b5z7GHOTxUmMZ2f4l+uiclr3AdwBUtlLAQ6M67g0rF+4kvn53ZGgMkFJhcaGkkhkTWAS
73OD1gvU1ljlRs9S7yrUmvfvxeg8KIOg/MUVOQtpFmIEiMK4kBJE8Bul/VR6rUOD7KyKn5QM/2ZI
ZoOl/V3E0SQI16JKLM5rMutxopcnbnt2S7cpup+CrIwiHQDbzJRdzzXNsa0YMelGBoJp+gVksnNo
BoqbZtj+V098VLsOXBiB6ZgA4I/BVjJA6QLxtvbtyqqSZF0z4f6Vsc7ARcNwLHcYskqRHPmfMZ4h
Xne8DRM4HITq94XhGSsMTCeQWq/4cy1on4Ut/Y6uch2YSgn2ZIBywT2uS5r6Qj38wa/5vuwQaqZL
ypDpDKewSB8aXrHG9OdAtaEyROi3URvrse5yqpeWoPBO6orWKjD2GOwT0wiansToNNxEv8B56vua
iyYwxqwpnhKJeqgDrbXe3aQ2yoKW6kcJzqNpQInl8tToO1Z6k3hoFlmMGoa9KruNkab0PPVER+1y
h9yqFuHKOpa6/O6nLjdEkxK0oOTlRJnySj8REqfo8tmg38HSbOwAHM7ExI18c3PPPZBj289GjZ+l
mYzRfG5f0tU/qnYb3SdnDitRDiBI0QMZks1TWqwpxk8RbUIZmqHexmcbA27sJR1kGOFMXJG678OS
o8oRWz0nt3HUM0FnGWaxbPB8BOs5OlKWKSZV10vx784kWVcgLEj1Ogb1LzMSo2xsQPh8i+D5d7HI
5eiCfSgq2B5/nfV70+1/esnAMegwrVMFZuFXh85HGljxCIw8Tqm0+wcQ4/gi2GT8T4mp9hoI7FZn
bpad6LhlSz6kkAGNp0+TgAmAOVWqM6yAlprzAxLntSopVBu/Uk7BfJKzDUbVQHSImOkMAx3nnId8
zHePmrL5UcKUQa7UvFWOcFZNZHMJ1bqMapBLiHxuoT4E4K9Kz7iePwXKmtATtIA6Av8RANdDojZF
qtD1Wx9KGOsj0CFo9X8zqe+hivT56WVwt+gDrJgp1cAu/NGEFHzdXNyiYmQGxvjXlUoUXO7HM0oZ
wQmstg1Q96nHLnSk2TWnTQKLezC7H6OW+d1wnk32SyPasIpi8DDaA/DW2J4M2UvqTFczcIZuCEA1
BgdHnuxXgLtvzdlxalnqKsf1pUwkbb3D4Txc1Sd4t4CJ0lE9dGiu+aFTnkPqRI/7WCa0zvz+j1H5
IsXxYmdv7JNqD/ap0K7SzqRfFaSVzBt0ZCFrkFHz1xEpKTl2lZm0Q+Z73P9y5Ora2S2nsOu50DQo
GHN6rahOhvRO1sogRLB8EakCNKHx/2wnvuePDRV48/TuPgDSPkkpO3sObV6A2RwFLnRbr4W9rXOM
2NsvEn9U2jS1QBBvG4DoSRMMyfF+2uW4Aw95oI6b893ttwuWgMB9UdLHP4xEygc5iWXtdj4vQ+d/
uBQCwaopvPj3RUG6lhz7zdOjl7pohtHxKU4btUdzAGClNH96hqUyyxWWk98HOpAb/wJv73yeiZEI
6x/j373nNd8ZBjzcZrI3pAB+R4lay5/F/dAONzgjMzF7bWcEq98wXl6AVIfMb/JYlQsXEn6XmCgy
0lBJdmOsgjnsQxinS8luTQwLSyfYK5XH+dkIHi6j7JOVeLgYY9KR1v2qxz3tIBy53LU4u1bmVifL
KulQbdg3w99wwY/rW1mrp1UZgtlQfgfwyGmJobAn2YUO98CvqvHH7Jyla7PNZD1K4KNN+y8h09XG
qAe9lhz4/QVoRr05N+PaKr/PYqfUNnxYxYDSMLUe98tZxdtrud7a4bUORJNtMNS8VFqWoxoM4GI+
dyk31tWfCFC6ceqvnqFvv5Tz9QOrLu9o0ic6SudFxrXc9iFdiumA+QDdfB7508bVk+K3CInXX2r8
3A9dl9kOgAvKw0Rl/L4AzKjkb2/v/HzMBtbWR/FXOyAQuseme9t6D0CQ+5Fj5U7qsB7pXES3tMkL
fNQjH3MhIlDFedbj7P4/y+0GrJDTFKLoQX5I6fgCT9cMiYNURgOXl6SSBvxkh8e3CXNV7LbOVF/F
/6Xuyn2tBCnc+c549ZL/L0WsXe0OkLYLCnL+61QWbLSTXzkcYTuN6r5tQzRodJawN1yfhNYhKpVo
FkEbF1w3QoPdjjDxEGk/GSSChxeJpHkkrGMLSzFgvQdKjZdbCTjImbvoKrfn769haocgvKJFlWLK
5hR8ci5w1bgBiwzca5gcQiBkMjWqdtUqnD9HrEkL61bAb6fmuwP2fJVeOKnaTV5GSNekFGFCNz1T
eDPsZbir/Z2VuPvOjuTQpn4+87O0RMbTbWqPQqrm8d5FmfxjN1v+WVXzbOiW2TAPN2RKKFQVrUQT
p2DbDbyJ/wNF1SjDvOvRboYypL0cNmWzHq3meD2V5BNPSWiw/bJSPhR5heRW37P7QGY1PYOx1x6f
px4b9YzyJvS5WqES3EA2ERt2et3ElvH3t1oTGPTqoeWBrHT3Nqy9ajjt4TTL2eTcw1BHfnFX6FH1
yaUsjkyEkccc6pmwwU6OtlRRVZDEEBfn1SYrxgaCR7iUyEa+lOjVJ1VFU0gQN7SjCezV7M4pYJ+g
DqGFGSxfr1hJPLEnMWwxA7BWMcE3t1mC+5IeAqB5xkLaAhMGQikfok95+QfxmPPvQ1G1aA0uhja2
tBQcEtccIwkz9yRh80R5gb9AHnujiTLUTFqfe5R+qH00h1KXr/0D7Fo2AgcAgt/+VYYIsNUZm9kX
J/8p7v+bZCuNBzakpLD/JJdSsAUPuNcZj1z/qv+corbEigtEt0Tx3zpMYdQED8gZ6M+pkMZrGXni
I7tkdCqPrKjMLDvNNaMcCePe3NRnCtfPtEF1VLFE4qjqiSNzeDfJRpzKrfTd2eCrggon2VlP33jW
5vIv/yEVFMNvqbTY3AZfLT2wjbaIiH6TdxbqLfAG9mfo+IrjqBCPUrcJJIdsDPrKvqEbuhKyeu/o
ghvGjIXIvSmPU+beTKQz9MIKxdnLic/FTe+iokedGNy3C7qfrIrrWb+m0kgdHH3ZMYzI1ClrJ66C
frtcON1W8+GSv202RmNw1gXq4+UN2uWxKYxm3IP5cJNaIkXbvx2yM1FROFiA/Nu46dFV3spt+BPc
3YUfB3iMfTNDT0sKwZe0OudQ5dfr/w7JgPev+fZZeYCctxZWqnqDzG62Wqs65tGMV4DaS6b0ykhw
8hZQmaX/e5pPAbh0+LEt1nfXHIlSauvw7QHyv+DzFMcYOY2sn3rrkNXv7h1QyqNLBA12pya0kxEt
Qv688+XMKQ2bAKFyBBxx3S1JCRnrEiz+0es9g3iFmaF7nqbkZzE0tK4o/WEa7uF5fwOxdku8p9sz
k4JhXJQiuvXjQYptPoFbdfOredMLY0TGjnqGpBrA5aw+KcJJXqrA2dIlx4fZGpfzwOb1wgVnCx0W
GeepAv0LE72hsuNzmf5LkX7Z9SmfQ6r8LGzTm3XFZDtc/StFaCqRYj74+36etDPtjVnFI60SdSch
cIiUHjP6NkCBYEm5OHw+tjymTvk7jyzMXfSxpJt8wgmqf9rCldxoUalX/HiOeQfx9YLwF2yccSTo
I+NALY+pzK8ulcHH565mYB32XnQ+qDEjfn/H9r33m4eMevSQ3nTNQhA9iskGcY57GVFsll8EIceX
yC7CSKLlz6EXv9ysIxUrCBvEA1FPfhNAaJ3cyrlskJKei+ORCFBpAFN7JBOlT49tZdyIn5lbkdNU
W2ldFWMazL225E2PlxV1HE32xH/5Wm5R75pcW2dc34P75IyTpJqGTXNFOj4GdKXJe/Kt5Z891snE
t8QCTK6nligNGCPj/jFznx3xJR9isH28BHExJ1h4AS1dZA4j3WIb+1DbqjF6K6OkBx8Mv1hdnZ8M
1xy9AtQ8VeqfwijiZIOHIxUgztTHMo7/FW4hpFfojESKSYBIXiWS5a+LjRV40tjTg/0n1mGMghwR
STVEGZcKRiaX4c3j8P+pMfk6Y8gOEVUe3zOMyAGQ+UPIOTehFZ8nnVeozcySEU4h0AMGaThnZunI
e4lK9AhZjhdhKBBQDW44tgdV9zAii3aDjtd9I9bfbhTh1JQOyW9nxy7bZBFSzKmLsYEeD5R+4BDd
QmQI2nzprXFNcbeKsyvHWKuwCTOAVf0hIOQWEHcr82ncqmWnXoAOYhRTBi1nfYEIdOasHKnDhjvZ
mXUsLXu22XDzqpQ/CaztNwE6IFWiJijQFWxIApKUnsFlL15cF5s3xsLI0Yogvh8WV7CDdjiE8MPC
n0mHC+U9Ryy0qAC44ebCjE6bZ4DfhTacnEb7uhGPtBx+3kzdANLx8JeRu/F1ZlMuwUfPv8b2r+rw
PGAXUVxbCTLNlkXObFKv7r/U2OWBTtgNVoTLp1SeC3bl85bhLApa/DS6AMjmhTKfKCFnMFqiEo3O
vcrFegU1THxVzu67TxvPG++64MRFK1NU4eOIyuk+0PNjOijfwLbOEpq+dMCjlFvx50dnlMUPrx8g
/eQiq05aoeF4/QVgys3sPwkbSyO2fXcIb02qcDV2megCZj4Fa2uVxzh7bYgC5uIWNX1IjwxXVfHF
I7991p8ZvUOZtqwGq2W/AM85TPLWmvzTij+2ngNwDbNLA52iITn5o1Lc1DRATs/2Wl40YPYRykFb
1yvjVZSdWgnyoJOe59+11Rr8MJfvhgGRL3xAoaZgAvxSjnv7KFqjFTtIdbPENXaBM1MEUXP14p9t
vpgf3oncS/mZ7mGxk2jhtNCgDxzl1V5bLSDOkQQO430zfFOJNVtePDIcjtBvssihHy504V7PfcrB
90otMhC/Atij9zp6R/Vyc9DRGVrjSCcLBAeDLlxKVqf40Pc0Kke89HPbIVWCV2cIHq9WfGRb4HX6
PUSYiuxZT7FNo7VIlBa0QCaooH5U5aMIpxzId+eRmzgxlV/0Dh2Pr7jEPZOBfSu2DIqEz8ChHrm0
xrXtAMv3/a5rTbA7YUGGR4UhxAQRG9t/qjaTQ93Dw1ARNI+Uzsg+iYhn8QiO8va4Q+mzH5261kqJ
Mfru1NrTBa/9Mb+zRzKsE5mI4jYfZ0HFWDu6DzZdD/ZEjyw/0+/Ov/QZZHV6duITZxUyr8AT0mje
RFCfQpXOeaSyXZ/FtQvnp+OVlPv2ZG430UwlH2GCbwGourmNiJy1bpQ12P68lU65SJosXhpii1Yk
GyJUvSqk++KqsM9bcL2/q5pwMDJo1HeGogKGYJq5/eLipgGt2Kp7N1d9YxHDiJNIfE3W/19bBFp6
OPWH1XZ//aFB8E1msjvezPTq2PPawRNzQdNm7GvcsoQFOEEMoAXss9vi1WLTxGswP26WpyWDc+yi
Mh9RiYOiy9LJH9zIVwDVwpGMqgLJ6X77ZQJt4WAq3fwowxV61TzCu6VJdCAD6UT+ZkGJB4cfqPkL
JsApRQIEt/hT2WYQScZ35krlwQynJmOw/uiRfRxxUFZ0aPRLui+digdUqi6Oj+PIwshwzry/Ae0R
Jp8rPFDblk9/a+ZZgpTgYbSrjGxniEsHwIyj5/stXrTIrJL+MavargfgpthkVHjxAlOwB9usnh5/
QeXPoDpp1PlXckIRE9CRz4xD8IXITdwOGwRb6m7oqwXTm7UY0Q/9iT7ejWB9Lv+XI+b/SiihmWot
dnOJXUAt3XdptoW6qm+0vk3WjbqCVfoNAbPgqNquMsMSatcqBiwL4Tq90H5fOX3M0zGx27ozds3g
g2r+gKUL7F8vewjO9FZGOOBMx9kJ57Jioiwagor92KZd0Di2xKj2Lesx5qbxAY7EEpAuZjyea0s7
4ZYso4nXqfzrfeJKg0X8sq9JUVb0+2RQP1OERUIkqMNnkRxqBD/SJK80UxFSVGDAkT/lA/erRAgo
xuUaHJJIvEeEO7Z4CMe/F/3UovlFa1qO1on0c2h8J0COoxlUWzAWjg5u4HpKVt+t7qREe+XLV8Pu
55qsWjWaow+InjawilSb9IY6l2PBqmm3AL11X6B7fLJJxJawDfYJbEE757Zhh1wJeT0z5UkYXBNp
beW6iAqqWVBPsdTEfmUl5Trt8cDSFn+TiA6S0BkPgLEtuapx/K2UVRthNs6IJU/jAnRwds9aTDw3
Y3DB9dAlZAdk3BuJyFkQxwkW3g918wsHb8Cqjj2FxAkeMt05FfEBM9orOgl4xaHjoyPUThetjM48
AkkO06LmONdDPzCP4L6v+HsiAzRgWe1U0kxqUXAbK08Hz5ztnKk5KeDoIe8klagfYNaGBHSw7R0I
HYw7+cOE9j0Oishcl6Ks+/fAdkg59cirkwXhcUVg+RSTTXPuo3G/V9C5eX9e7MatR8ET3r/xHNZT
3FbsyNdZTTjnaZ/ry3+3xbYTmfGwqGb71H1nyJ8WxXV+qKyMI3gWoOd47d0bRyb+RRAwo0tJlpOx
cmX7cWK9efqhdGUGGk1RUZAu7d27jsH/Q9N1C0keK59f3fS/x2BnEHNneZv6g8W77InV9wZMLwka
jlG5BJl8wjyYdlQJuW6UTmbtTXlGj/YejYQjCWaPfApaJz0w1LOnvO/kzEqzL9/pbuJkYOB7lNWU
g9W9mxTqtp8Jh+6aE/23XNwINjMmSlSoBX8gDDR/cOsNEWhZ/VVZm/rhBHufhW3uti/jQleoJIpM
80YA/f95Dc8B5k47iGAHy0WSGL6t8/v7mYncY8TTYRyjaJNTV9XouPji5bO0BEQGKCs+tZpAp5RB
8zRM4Izu9WNObOavwMDz7oe/LPSgxxnoNoxOW5SOH1tF3e/ENQ2trmGMhpGSUhJBZtrZ6IY1JbRZ
3KiJgoY32LqjlFnHDLRjVCXAeuFvm2DbE7IYuI6yxqvP9Q8soEofZybjqcycB3ta1emnChGci/Dw
GnKIwnERfak7bdxHyMtjzIxE31509tbbFAC8asR3uDDDDkHT114cM2KSUqQzVD/sZ2EQFU1jOyNF
F0KpNvOuXPpgDDb5BnGDVwAXTZB0UZkIuyK7CsQzSEknjUatB3M4rSU+n/vzRfOJpWzK8WK46baL
oUqd6qMrae7H5AVS+gfCxEcVqWD559ETEjdorC4wdcrbS+lbiB+/ToadDdepILpaa/VjlOOylKZe
/BDc+CwD/ph1Xk866W2g9ZrhoT4I/SyyIP+6BTrluwxf/gidAwF6WSM2TRLiUk1QWbGl9APM6zMj
d99ML7Hu/cL0yA1nu8e5CI5Xa9VqVR/mHqWNaphPt3I5F/GTnLfHbm0A0I0SBK1lU2Wc8QVQfpI3
kgZ3W1VDlGjBdtyNmaCdvL4xj5rvnybNmXPte8Azka7LW1twXITBQvQ/OTkp2rtOB+TCJKOrZxOI
djYAwh/jHtNXYTOrYUgf0KMKeZIickHQBSg/XgFv7ncBsrHFx3AGjizYAw/fX8XHhnkztpT0gHGi
UsrEy4SmzrmCJx22a4jFxR7oxcTvtCRYY0FC+Rv50CTRcVNPiBP11jP8ILsx31fQ4mCe7uyGvQff
8TXCuTl0wVw6DVMZJjzGuV9laUb7D0bHNqUaJcDjkF7pWoXawDYxzlGPQSlZXwLGO+AUySMzCEBi
xxaHayAbpBsOOTKf1Vj3R1OzwK4PSBi+FfqODe5PnyKNNJMSZj+wMcf955tfJxz7AE/dtogwqvhf
73/muWiRVZlk7v5GpwsvReNd6A0Fntc+tCj5DFFhbwKCjw7NFZHvvlLAYNqrDXBQGxKSW4USiE54
PeGXKksrzg0LLAykHU5tLY6UCBXt0sX99tGWpslNmgAQjLKl7IZIT7PPnSf8a3ssKgklOcIoUsvO
k3g8GGQNhDY1GHyW2jRaQx5yphvZ8s6JYpQ/5JTn0juDwvfSUYb/FDn1kjdhDn2qdcXqMl0hSLMy
UVj0FXfytyG4o7Yqo2VPMR5EwyD0lJUQtp3+6rUMjPzxtXG+cb7rupTWWC0+9TbzqUECV0S3QCYc
W+TULCd8Ibp58bUBmIgiDnB1/8k2kYRyxFbWITO0HHKeL4oLGbP1jP+HXdsgFYUzOs4iax7VJXQc
xp4kkFTetGJn6rdTR8Lrtz41PEkwOmTbDaciQ2nfVQQydmczsrJ1Ed5wxn6qrWE6G32IqR9IEg+b
KBOd2Jx0NTiSXwTqOGHStCsGRiYxhoqayoFpnxBiaOEqprgpzNtArw4FAsCo1uHwvicMmzsRhcf5
ghr+acCkZb6oURVZzBuyXSwBA2fHFChVxMfp2KvYxW3S4Jfm2hFO1/cWGlvwz1TB2FY4lraReYsk
8DLmFBYly6jM6gOKfau9NUEh9Pz5JYjeZgHpd/gdGQvuaXC2XDhpTSlcFDFwZVNB7l4s3rpw7HgA
FjOZnF4o5Z4QM0ZZmRiO7gsY+cl13vuuvC2kza1JZOXJBhj9bzUHKvLonVEU0vRTYFAQcS1NVpl7
hEwr6TPcUXCU79aogAJFXOGaBoGY/wSzl5u/XPKZCWLWkPCOywRwPVvj6Ms6txboeC4c7ESmsxXt
ZV6EXv2eIJVA26nH0+h7ZNila/B8jz95mYoLC69BvhyBbq/BUB0+IiVDKd691PylNUFNrMRCelK2
0YVnMsmJLoAXqM4qqxgtXOv9/JDFnZcAEQu6wUyh4gchMdur1lezdc8mmaEH9LUDsvJSah1x995R
6G1wunMRJVOcR9s06ZjYPNNGOc+2R1QpbYZchRqhnt+/CKKY1hR500ZoJ7zD/ZvXlOLcSUW92PzB
Rz9MsDvoLYe71rZkF/KhPGaYq6iXOs6qQihbKaGsO3sf0v6HvjJAMrWdrP3NJrZaI7IXcXuBvhez
vs86O9QxaiihmYcfecywEypxQzEk0ynuBU6d7vSyqxzw8I5FsPELZtMMFSfR+aK+QJhiWE5fviiF
mzpQBMxoUx/39QZmy5DNUZ/qBxl7rCWKvWjxKmcC27MFNiJMHAGIATmi1ZVvPm6oSAFgoYCLtAY+
SoSVjd8BNKoWbXlcghR1x/TKT/FLDKohxlJRYEyUsrx8aCet2D2Nr24o6YKg179glLT0f48T63WT
3wRIGbyfJ6cvJyL0QkXgv4NbB6F6PpN0aCXDBEWToghXpi+HmyTZ4a10t4LAbb8THwyil91liCrh
rbYEP9WpFrH5C4K1s7Ra0eRJ7XW0qMj5WSEa5XCNyd4OkaoiLG4H8oCdNYXXQX9/eyPC2WUKxWQy
o5o4VB+jR27yaDrGMXCKWzCMKxAXSIV+oDQrYW3ndBKpfRHZaZKgTJrBklViyE5zL1HnUdrXqd1B
a05cxSdmbVYBKZt8RqKLD+2/0mmnPS/p6fH4MnJdWIz7HlyuOtEth9Gnb7B6cDlBQKa0w3faiErB
Gvofy6FLj5QB9KPTtsvuOL8zNs078QBUvCMi7KVQ77QrgSHTZAYiOxT9OF/EjLY00UFMpWxDWfkK
yb7aTQ+pmRLUPuxBM9gc4mcWzbv/IOlg+tTMCbr/VAlEaFEOGY38qYcfW6OOcxHWOr5Y1bQHQzJb
6yWPy7q27N3JTKFIDdLjA5oNL+SG7UHtDcl/RMZf2dFq2Zs8cSedInFOqXrTVRm0WeiEOuaNHwAh
TbI1oO5AmIGG6/ZUXDzpBY95Tr/GnPz9QoXGbnd4uBOJBnZEvJCOl4kvmjU530q7hGVyUnJQGcgR
gGrH4UtNHAvJiSnuCP1/hFkVW3fCx/p0eOFgvQvtWzIjrhAHAiHjAk7Oy8/ElQmTtkfl5No8U4eK
nAfo6jYBthmML+71ngP4tKads/q6CGMsbrSOFQpLSooWWh/ggO/DlzUrzmBJmeTdpqWdso9I/LJf
756yHCHiBnBz5xwhNbHjzZWg3c4NCzJcLBYjnHtgox2zM+C0bmGHkWddaeI2mn57VtzC6pPxCVkU
MYgwdZdfI4uYSNhVCYSDMhzuWiwvHBRek+klu5Nkw2tNPOVMg36G1gaGmpYNLm4yd/Ll/BeIkidZ
Su4bP73ZuXnfIOLIZ9Iq9sZLJVhgy5teN6mc4bv2c9EN61qIYipg5emnvZQBeZ5okX4JWb5ihGoD
R8nPebpDDflv2YU+BKX9HuQst5y//CnmCqrx8j+DxDXmI+XT31XjjAio2fkvunT3m4Zq1HNFAQu3
n7TmSDMKm5843qsVyTVSIWUJFkyIKXLdtqLl3WDG6O+NfPWg0Wlr3m5iT7Zno8cpxpGH0asixPGl
w550BdsZqI4f5ovR/pzn4G7zZ9Fiyaj40m2r2Ua97ursVCxn7CVZHHzkPesHSXn9Jnr3LzpFuUEQ
UWXv9rnTVfTy8lrF9dqdISvseolhiyB3d6hTHG6B1ReL4bDmxQse+RSJGrRB60xe/WzZZhSs4rVR
KWxhj9DoCGazbiBlWb0M18T2uE86yYFOzQ5wc+6sQHDuVIsmwpvr3T+Zl2eio5FBhIgqfuwq1OTx
7Gdy8eyQn+bS47Mo2h7bdfv1bZAnhWAnsvieBUlJKUqEzTMJqE7Z5ysd2pq2y90TosOxSifyyB8K
54DmvehpqUaom++D0A4e67MaxP4gvBlAZvKwzNl8PGz+eGjtzMaArTXWic3A0/7SmRQ3pMGIwdbZ
0HzsQWU1GrpBWuRcmQ9QZ0MxaLwbmeCJXZsewifP+7jIWwPudhjCAtWfjotfUjkHFgTYSKci6t0k
E55O59Woaw9u7Qeg2IlTjKupzSJ1k/JYF+p8doiMCdKqd94jz9krsihrKEQjtjPuCWL/7JqvBH5r
EC6h6A4niOInhr9VK+vzcLTCiXXG0WWYH/Q7Xb7q8RinPGJ5rN0jsOkvfkUaZ3rCJmQ7iPIFQNAI
3uYfC3BuDWjwjZJxaGJ6zF7nPLDFl7XyywZv9sQTBbBzMy4ksmbD/oIuElyiQHRvArmHdhhRw8dV
Up2PZV0VDNG1mAyMGYFOhTYIWcHYAodGWZfg/GMaHgfhUdh6mezKnP7k4azIE/ReDN4cVcp97wIj
7AfdJBW7ssLuRVccucTE2wLkeF0SeGtrgx+hn4ePuVxurcmKMOASaJUuFFZivNooQTxfa52LT4Y8
7snyTXchz3IiUwsbJy5X6LYp3+kBKFEAEDIN0XtiZSpU7wjrjHpdjF8/pcBjYWQxADEL99uQ0Izf
kXxKXSfJfNA19YaFYQISpq7e+q1AehC+HXVqPOIWxzFdEIBWJva1qh5+iZfJzqCO3cfKiutpFaGW
EC4HFJn+O9KkA6Ckyu9Ey0VQCvgX8Y7uIyv0bjZrRI4YM1Qo/xaLBN6yB/NymADLqOzsvGs+7HcU
5qKAs/XPaCW3AUxBRAQBfX3CN/gQECNbvvjz0GDiEnKe1u4OOP4UQenzn34RUA2/9201cxTQx2hD
uZZWKOlsE+vtSTxFkB+FUuARYXAvr+JNSQ1SAthhIdWkvlD6kACau2h2gn1QZytWbrBCmgdhE2qS
/TKP9GtzDPbjoSzwbvzd/StY/P+kLFjVps0gwO30tbhtggxzvdnrJC0jwL9v6Dd08OcQgcfbBaXN
SJN+KuMZvJr250irhUuQqpGnhjRb2CseJdcylMwLodrCOe2VNDzZFo2jfAaWYqnAgcc1u/0NvQnx
plHqS97pqtREQfnZDRa2InFET0tUhOqf/XWbN+0WIUgdQibIqTlxqRXmFQGoNLmUF8DAJ2nFRhBF
YtyFZlmlklWuqokqUzh6gBawRJFYcM7IQKQfBBmyISpLcCtOljUyK8ta/C+8pdEVcLAOay758SOa
UY8wsrXi4wRMvpfmGNor67W0IZmnuxt2DFF4uI5gdazptppYUL85Rym4Dg+Z92YKy4klu3iYtKIf
Vj3ujMXAOpVDpEsyiT2Jsbe3Py8N1xGCmNLdism2uxjDw1Bj9MMEjcSupa5MqB+CvwmWZPoawN2G
/EgNr0kIT/lUmrW3t/XosF+GpobDxSyklL2Oyc+AXmdyelqWx3hOojHi0JwzhbUtgpw38mSoXbDi
nOwumqk0JPzZqvkecPHN+Y3nDyOr0KQy7bW6biOni1pk4Di958rl+0AG3ijAEucDmpFC6jsX81nD
jqfgJWJgHmoxAq7rRGXOORizpoi4GCO06kwjQynxFPpMBxUSkkf2w0QQIkz6RfsIEZJTAIOUmYiK
6llr01J03lYKDTXGRsJUG4jtQxYQGOprXaRZwMjFYJ0Bvs0sRk/a8C4Qrp2cBy4e4LCdMlwdpY6m
RWCrgfRKbvhxpZCNnyhWk5SjMFjiA0j+pUf5uG/QEwOPGC/gWihsnnSCxxZPQnPhdeNC4GnjZfqR
IeXFvpdaSPZ1IyjVfSG4Ah8gFjdofHcsPkMZYJn7SLNNXbG+vTei6Cf9klenQVA/euDCuaWFUjES
IrdEA8JXMnCTH1cB1m1xHFg8fDk0ZBpUbpNQVuqSfVfXCdBnNJVqLpH+fV6IBOcBBvQjqgU4/jRP
I2SJ73kp/GIGlgbtnkpEq4w8qUZBRg//dCCE9hv6u7Jnohqz4CtbmBG54L9CybrgQFRLf5O0Y4mb
HD8uJyeeAlmBgiKTNn5cPfRJKZIUJJVVyNDg13890VdXzEkwyp3u+5uKJKGve/5QSTOD8nysBeoW
/pX48ym2fkl59wImk72j4dodZAL6WA/xFBApwGIOw0ohbtjJxmjXxVpCvPCh8/e5Wphi8eEUOyYQ
mEsbpLBz3T9ueWWh0mvL1dpMJ2jKvFVHOf8FLvPpHKZFYmKTF1Kr1CLuZ6U2irXKXFedaNxCZ4/O
yxcqUNXb8jeEtH3p4mUahf4wETwCbETMVdEi6jUU1bT3otAhriOOmtA1y43MRksnEdyR0iRNsZi6
++wdOOcdRInVpbUoslXVrSzFnN3OYC4VigmQ8kMe3XZYAq8uJ/xOMsw0ww4vr9/xO+t8q6ZAXaU4
tbILMNejbTkN4k4V5+gsqQqpCF29qUV21nBfyzPJtZliBQw4iHVnRPweKDQJLILX/byq9OVe8Mkr
6ZjUXMomuZPpgeGWmt7ViEYKVXZdyd4yaEcEwjSD3+RuJFbQjja8Z8RxKtLWyd+Z6Jyg9HhRQqGi
y+a4ZyWA6VXuDRRpQIlr5JPtYNeKXMBhnX4sz6cNVl+SyvK3ebPiwcw5JojmRc14TihOaJQXyE/H
65tvEHrePqdmklKolKkXGg9nDrCFst6iEYD1riaNH99PsHoVYgMI5LBbyST3B71yGPcpHX/YUqxg
yh+THRGwqqyWqAkLPOfpnPmxThKonCuytK4/M682s7nE3hUU8eaUrTfCQIxxUfcJjULjznjwpjvc
OZmmFFreLdvUocKFPvRsQ9TttLda8zDq8LAvuyZT+RDljhovINtHP6HDBlyElLqd8jgXaNSPbP0G
Ll9p9ebKClkYXPGzDFS7Edr81EG9F0eo9lM1I6d9+XSCRx8acw13L4EwEtFpmwXv2cHZ5/JyhVPe
i9zUO7MD1ks0nctJC2eZjmj+RG8jBeYqDnjzRQMq2M+5HoxPehiCr+NI6IjuLC9Tny0o4LiFxxNH
W1t+ltLMtdNqt8Z0tIMDtuG9pFqenVMNSLq6Buyv2Tu0KqhaXRcQ0scRPXF03GNnIVgQjvKvUezx
8RfAz7y6+IpKj1EI6aNT0x4hTlY3/qEzSL2m/5xZRz0vxLn0Muw8CH/g12+GY76oGULvcbM5swSB
PzgOES+VWUM01GrvalrmWZbJRthzc4nWLfAnv57nJlKBTlTVRERnxhV5nqv1odeNBZrVbKC8uSUf
YHkUCZI3rd1B/KR0MSz23ezp7jY5xhtlgnyKuyZAPuMpF1xP67XyPfkNPzTunYb1yjbHWuvXDrmW
2RN2FUAHv4AoX5o1aSNSBaxhnjqFpp/UWT2QwYs2Q+R4OvYfYdV+q+A+kcGzASnAIJIPOVAhB4fU
AcRKc9ZnWR7T6ri57xzw8TRNSf+DFcSXre1v1OxkeacLgo3EMsxhPkS3dAUgbdLPaPDXdW6Oid8x
Un1NJ+gsmRjnr1bfv5nCckuBfnLcCHRIGfB8Cfudn5GlGSd26iMdt/T75OnDMNpAkXBrOf+2m1qc
erC3+CGR+EzfMTkoSiG7/1HsFdbILJzbEkP8ARlQvmW8XSp3YTLZSNjkVJ1Vj7o5i3AdhO3nkuMA
tNdVmtjSzWA6LYs8f6v490DYdjbT1uB8OorCo4Pj7PZ2IHS0AH09L7b9xgJT2sezgOYaYohHWKpE
9ba1JW/9OP59X3ogkm1/WuvN50EPf5UAX6Tqe7CFeB0yDHqzh4xqG6KS7HD9iGqeJhbBN+O3yOaF
3zkzNBCWAn7UjR6GhNoajpqBZga6AWLJxpn7BnSUF1EGc3Rn2GEDvhNbYk7DQ0CWu4fDaWytI3JD
q2CnT+GdyASp/P2HiPsBu6kZFi3VKr+GHdtSmJFxH+FGzN8WEY0QboshtZKNHNTq6SMYdJqcaYDC
2DsQ+BCLBNnH+82CDwBZsSj11Vw1/rH7XYyCsNsCSWt9DHE6KtxKOsxUXN2eYwkWp2hOduV9usL3
rdv+UPlR2fp57IiP7t92FGhWjQNikLLdVtptw4ZiH+7dFkaRXGZeeKBVYD4Hed+w5z6xOzov319R
+VlFX0KlBLiTjua6zvoaGZdhtpOXBkpFTWRokHn/50sPHo3XkC5yy1FISpztLkBnMbh4gpwUZKWs
Tjx6k3nd3L+f379IoI98u94G5eH6kHyDzAelC1MSrmk6x5n5xm5O0krbn5MV/zNBQL5VzUDNo50B
liDhxx0UZ59q3O3eLNFoeIGOPGuZeAACUUWXRYFaSNFe78S9rjDAMTHP+Cd0jDDI+I3JEduvZyoM
sgH7S6kMGml54RXgOk/KldM/Nz3xjaLHr+C5eLkHo1avuACtMyzHLyHimWv+HvHfPYdQnIz5lCOp
Nrh0dZBF69dnE6L7jZDhCajMISJCpdU/3yK0l8bATP+LldaJhoyCbxuc+33IwaJ9o6liu7eXf5Lu
4AfqQCdhMF3gHqytqCbfjcOY+V5ElfSzjS1lJe0Ed7EsZuMKGNpsWNhlJPy7CRiLbY+IW8rcSZJp
4eVktPcrqzuxsr0+2NOY7YPVJNvGzgZ92Z6hWbN6mXxewUqqbOKHdhvYXlLRordgekT57N2ElzMV
r/dmEP2WyRyLtuqoSI/YTUmcTtk6oWTvDObFkwDUtVI8+chL8OfCG78JYvkt39HM9KKWijL+KHgD
gUB6bJM4cVUP+pfSDrWglvi2t8YRLgznPQqdejY6Pw9tlflfMqjJ7iSFnmqQxQduUJh7zXIe5BWg
Zu9iC/DKW7Jz2oJ6rOQTCbfUSvm8QeIY65h1MjBtHKQWnP2pKUurCdjttfav2hLkwVAGARaIJauv
epUVNVBjCJtPCFYnX5OH4WqxZLBemRowln+TyVUBG14mKsL0joAzQDOz8sBHRqWNmgXxr4Q2x5Uk
Abx0O1CtrlaE/321y0V+ORCdUKz3BbCWUP5Yd5Q7E9nFIWXyQF2/HVRkB/MzyV6pUoq7nTHI2C3E
0BSwzREeBxzRvmHqE5fFtCP5AhH3NwrPa17h7tZCouPcbkwmVJDTN8pcivpUYhAGUjAbszc01Pbx
XZDEQ4BjoTbjuHQBUfMd49XMGZBjQTMWCUOxPQrc/RYBto19ASBe3JfelCZ+szijpIZwVGxHkzs4
RsicOJtUVjMnFV74c9wD6z79sOoW+2rMGWUyBZSephKgTosPd7rKS3cEXYH1Q/XiD7ohbzNzhlbl
jJHk5S84mdGtaXzXwBZLeFbQKt2Y8TOqDYhZ9VsGgytoNIqvCwv9mj+McKAzoCue2/1MU+ftvxTB
3aRS1CWQa8LZAJKA5Bbj9tRNHhtnpOn0uQvNNgVUvCEdpTU+KS8aUOmne/vC4ZGor2y1Q15FkGwY
+88pkHzXnO62OlMszaDk+VymZ2HwV//uJIORNn0hQVSjmHf0I/J0/bkfVEuo5zlBqqgJPl+No0Lh
qppLaxqJxVBSptm3II3sQjseZ/K3JxDXcNw3EiuErizlum6KzGfxRJH7HRnU1W14hzbySUaE8TSp
YqTYmt2OEQSFxNq5xnBqTAmCkP7BEpoePi1Na9M3ult/+hT4DRAPrtq1TgZKu7LlNe+FVseZDB4Q
DHqCsw3ZO4leFdUE6wCfv0m4iCxtLYUTZW+Gz+sV4gvMEkvU9q5UbkATA0YYG47mil9oHBSB7sxO
DBaoNAmYsghn+6CSoRKewR0XwstAs8prZklGO0ucfP9p/5g9EOPxmqsq+70waP7Izx5GoSZqStuj
MM3g9Ntw86YXYHiBLkJ+fbWZYfSSzvXnkgeCbTeLZ+VuvesGnSdNlvbngZ1auu/T5wEmiAwh58Yd
eQx0QenuDJtMY6xfVsCd88TDDtuL02Eft8mw9Gwc7UI98b2C7+2WnlA94+N6dmkya4vkDF+cqI52
Xmw9Y5/rp+SjI5ST8BxMZ+lLtzNv4lSyi6WrbXWPQZpAidQBFAEqrLwWCYW0Y7hbiWgCJujV9X5A
US/MyZpCVqcpXqo5tKReIs4Fo3iPpPUVLJqA+4OXXURfRXn9n/Lm7rmDpaTyw+Jjt0zi44O17um1
s0C7yygbXaZdY7xYdguvN/NEm+jKa9UNFyw/IDuLzhz7uHu8cBW3DdEtBVkiDDS8Ja4uSh+zPxZy
0BRajvvXeQobmcO6bdT4vymcnF/OlwtUygsddVXosc893ag0uZyN7BNR14631oXlRYzvJwsIMw+F
FhYg92dkhtR2nWcplYdD6T3vC1btW5T3QfqHO3q7Wyiylugp6owZ2vsi3kx1l7IrpML/l/tuEf47
Rd05t17Ldwkcb80PzUjucPekav90BCM1VmWjJ+upEbFGw/AiO2sSYdnWOpBfFqDWWvRSw60gVALT
5Om+jy8W3dRr+WdkA3nsxYx5r7j4yo/4R6FKZHbOv6VZAjmE7pw0sFzgzdFK+L6BKHrmAx0L7ZXB
n5OiL7dE+GMYwp46bv6VSlSt47m9uEixdd3ebyi+GNCXP34TzKTeTTKKAAHdkkOqWzXv6fIrfMnZ
/b/GaLIu5rFvYM4KyNO44RDOAKAmTpFnxnlYHJDCo80hMRAyhJ4y+FrCfFuruP58XTGH2oxbRb+Y
HybhJoTTeYpLsyQ69d32RW2KjUeffUziMNBkymu9Svqxgqlw62CCtIs7F7zLoqZEcPiwLEqC3zzA
8OuVF9Sravzi0YlW+6+ySPVMzoH9zwMHu8bTE2NPAnP6mBu1dC2VhrcW//M/cwIg3hTOvvnH18RC
zs80eUW1XSJor7wd5oyIgiGQWMKdUOnackAZq8/kSYJZ3UD9FtuGlPmEnC+gG0jgJRg38XKjNEdu
1XE1BzeI5A4L0quJTOd86gqHsCJKPlKA8AEft/MpnJ8tLyUnRyR0g/UfCLKuNhjIwjhpag9atB4f
lIGMwqX/5f3Jl3S1Xesvcj2wSpl6SNW1+kf8ZR9zMs0oqa8J3CLlVk7x80uOOPnLhFGPZQAYxajx
M3dRGF+X4SGzbjiaTOC3dQy/fhRbJhNfutjdefFHEodM5R7UuCj0EFpwBieDy4UOMndPJNDELCJq
2KFxrqYUX9AndGvGZ2i0bWEoF+jKi0X9pWj1Mi6d/mFwHzW7zWpWjXjm3P/pgsDiDmKvbnQe/8Fc
juKwHsM0XnR0aWBvtRlH2/o1tg9kYcJETVjcNLiBgBPILMTejGkP5w8DK0IhX3fEb1R3Qdq4yON4
r6BI7uqB4fAYFsqx05EiCHgoOK3je6HRBxlLzX/Y2IsRyNscBJVE+uQfL0qSM66i7iWq0rcz1MWC
okZUHSqnr+RdTrgoQY3gld4pkWuivRgHcWDSBnu6YwB4Y4VzEhGsGFDP7c1/A887lrit59Jg/CNm
UMzy1LcRUy7u6v+uG12D6JMBxi/2bryQ1S+e6nE71W24zVePB7jiFXys9UYuJF6IXHkPteSfZbO2
64gTDQWNbfCOGHQAqoxswkRxtugDARqn8WcOPZ3WdQ+LajYiktvGLbYEfX+a83feRc/0WNzf4zRc
35PV8/Kgabl8CLIkIek3WMpbbE8go9/lWtwsTHEYonaThZFzvr9UqGXqd2N2zsRrZyOZ7RQph4du
0q362gJ48ll1KQ/QUUXtI+40HvWaCo1ny23KW1JoNiYpk+RtCN8UwmJVzWk0mUlOGJwkEv3ehWzS
jzriw//EwVZYk28ZrXG6If7f1m4BdxbSF5WUSD60qx/YwQsVR7HSqD5WS1gkV6WcnMk/HbS3FN4N
R+C2eGZ/k4QLmVJEk9InWi86mxNWqx2VYLIlA64T7SEZgcH2ucsIcBeBl7Qy1RxiBx9G0h/40xX1
/+1YYVUwFNyfj2Woucu2fX+IdtuPU2E9cBqEG1RrMrZEFx81A8qS7cVRliPqniOJfFucfe4f/Tqy
Rucf4L4OC/VtYmsGtSB2MRQrz9YRm00aITiePgeg0j9gb7LU0zhpDaKVay532FAKsq3x+BRyA+YJ
bjR4DSvh9EPCfWWDUc+t/wSHUcJTgMMZR0G8novf7pHAijh2sSyTGklDKrJ07OIMzOP1OHa1j6Nh
NIITZJO/UzlJ3eWbnd/2WQ/h8qPi7/1x3QkepM5+oiI2Q0rGvSfRblYSPHTKXXbPso0pqTg8a2Wg
CAT6GLmD74DhGvUTgAQtnXUVD/UI9XgSNKL9aNjp+dDwtSQcSb0rqx3EUJGP0nuBVPB4x/IDNmuf
TJqDu9M589XfDcSaIXNCd9BUe3R8sxS3tSanP/FhFyYC/c92XaoIZhHH8qO+2BGMEIbUYtyx11oz
JZdzzP1MEMhprv+tg0XqFj6VuV4IJLOQt4ZtT1b6FuEwpRdaqBUvWvgiiKxBQv5zxfyvjbbos3Si
Buv+liUiIG//K5uEMmWJPsQVSF+2U+pMyA6+BBHG4MSv+QEjRm2bDZ2M4yEkYaS3thaLzpwd5bys
GLfDpJfaV4kEWbwSYqtjdBBXGMfXuYTSiD0JnhlexIZk/2vzHB9qrZLfDgXqN88NHGoI5uJJi7Gs
zW30Ss2RzHBJGIasHjACjdpc3dqxKiVXHC3ugTGOdMf2icDhMZju+Zb8klWO0AXLdkaN6s+ghA3D
+6h3aGkDzEj3kY4fIztvZMgYkGmoymcOIeByeoLSUudKmEP4WdnBJB9MeMVuzXqKoeFSgE8R7fwP
mq3r6fC9V1CszNP8CqpO/tAlRqB30H4amrfu1q/7XppebvKANrTF5Z2SFs/Rb2Iv1yK9z4XYQRwE
oShFdNgKQ0dOYu2p2cQcOQ6ResKzbhnNanX+SIWufm49IPqGvcNdV35X2JiLfKzaCI5gRBhjI10J
q9azpJ51V9rKmrxjYl1Ikh6rOKI2yjxTkcuPY4xN9hi3peVzXkp0dLpadSbXIFGbhRgymbWnHrHz
tfEC05sRekbKJMLwjaMVTP829u1qcIraCtlo6RUBZD248W4+hT/irI0R2ZxbdBdV8CvzUchqkKFd
MSpB4y3mEfOdRRfvKg01V4PrDTNNBPykOKLN+G7eeeio04UltzPTXyOqnDiFA8YvcTskK5M0jpgm
hze0uJY5UXT2JXbVD1BdZxFR8RpIDgyOvIBgM3k0zA3F5qZ8i0q+VVpIe9T+zXgwCpCER81Dzfoa
GtsHS+ZybLtK5ELeyEFawL2P6bPMtnoPXdjT4J6jLgemNFCkBm6OhLWa/xtB9cbW0Zvji8SwsuGX
x/j5PSEHaAMNfGs63kh3Z41C9aucY6SHarCgi4OQWomly7nUK5XCkoIaH76ozH8LcJLCAMhsv4p0
dek93iQicV9IgfjS+Ejn9TPlnw9BmhqQMseR6myBH4eyLGWpMYD0IiLozBxFGvE42z+fFPf++UDe
bHcLBipaGyy2tdrfmpWgeYxbo+noQ63RmocTALZ3X2O6nW5KGi/bahxyaul4pf2bDifnGoJ3OID4
XqC+hz+P6zIznk7WLEsKcIZcad6owxEKM6SdwASaggWmeHyV/wcVp7dnUmMlanCsA5yzqSwCdq1P
BpyRh/Rsnq7NGO4Jj5vTtQVdjk8BySxsiWlkLGiT0Kx4C67ljTO3DJq2ssHkrjDqiWjvH34Y8Ql+
pcrJxO9WeuvTHZni1uA548d6aYgG1phYaxWq3WDAwCBzSM6aN2V2keHl7wk4mevpTXgmBymt3T5f
kqxTXp5MPZfN9xdaJkgHZs11waUd8zJOakrSpI99PlSlKE+HC77jCeayHTZNcq7ZWY2XQZaGr2RT
o/KfGudx18AZ3GvGOHl/M6EuC0hXw2GIirJAnI4fdGvidz41C8bML1Ah+dxSNYkytqHDvh2/46DZ
tytrCIxJraiPG94GLErH6pDBdPUqobnJQWOWjYbXx+YdPS3RK2TTeXNqJJlKR29i81IoaeZ1JxZ0
YuczD+c060xQgvEVFKMe4utNx/7mlc9bGILe3F0PjimilId4JcEsOiBjaKlOK1r6zDIYITOXNxPj
brlASlbDCwUZ21yqJ7cePicLbeOPPo6s4YHNUlO3WHBeJP6SD5b1AoNerbYDfHEMQZyGQgoN5uTW
NcMuEsK4En60RMz2qmVJeyhkUfh5uZFzagQlYhafU/CsObgXyvFAwfw3/K6NFSyq4X+bWjpbjkO+
wrZ2sa2FC3VxuX9XQ4dbi0d7cP+6JNcTYlkRODZ3r1iVg/Y8tN0l68aJb0JKWDcRKHcCPlN/NGab
pzBk0niCIpwLCzvL+/+Uakrl2dPhFHlpsq40RtRn9Ws6haZ5emtTq0rOC2SUu6Irw1EvnGTY1iK0
9/AZO3i9mdMH2SttfEeotpxtvpy5xlCZfrAKsAtpnLA5yA/Yvkw7g+AjJqe73xerFwfu6WZjP7RA
ZW1GN6SMaVI7YxnI0zbYoLdMeyagKL5Hc4CiS+YGVqM+L+NeNRtp8WSIZiQz9Kbt5ZqYUOsfIERW
ThnvfZxbKSkJICLJVwLw24BIm2exdb6FE5B3XRTPAcJFLmuy5FQ2NXnU4kuGmCEsROmu3NoQX3wX
VgFHQ9NEwbUxdAIiLHExXMLsymm4PM75gE/ivX3NA6fVgRElnw269Ju6m3EGK1a67F5+xLw/O0u5
ss8Ond0ccmQeyA4ghFK6uXU9GvTqEqTmoMLiVT6PAOXxSQFeKL+ppwM3tFKTI7K87PtZC2uUddhC
JXK6RpSJkf39jMqxeah6+WAm78k/K3nj7g7CQSLYecuZyS9Ek+psOfHgjC6ou/tfoqTPrvmOvtxy
f99IzoaMSVvX1YTM7TWwu3o7q7fs/jZhAL8Kn0PqbZGfnPCA1Grq+0vDcoqeGUZxefmkyxY6FlVh
Ls34D9EW9/yUe45DiRJVvw67YeFekXDSK2uh245h4lWcO7kYy9FVhBZfQuUEKBVIDftfrtxwYIDH
ZeEYlp7QqI6brjForUCh68KRrCnz9cLV8LIADigkNgRtan2eKkF513Yq7fWCDCvwMvhKUe9ja0wE
LAOtkwf6Jksi6dqmk8LOONrwHeAxhIKkEM6v84QYXBEhgq1p/mDUnJJoDoUi49v1x2qLvMXUsicB
i4F05RbqlAd7tH7/v3ivcnU9zFexjGQUhxyf62vlal8ngrQm1JYthNtQ3YCgOx3bLh6+iiyUdSfm
nkTXNJU6jrlMk7C7Hjz+li4A99DfbLpqlXH9XdPJBMayecsvWW2A0CuffR8eM/RPKlC+HEnGStOb
HKTrk20cSwGTJ3V02t20T0PKNrgabU7h4TQF0LyJQ3MQAbHcafEJdBTqSlcBqPmb4GOU2W5YArW4
C9xbByfKqFt/ku3Ps20fReXUdepuwDx6m4dRsGiRnMYgtmShmYfdzOBg4JV6GkAye1coiYr1hp+r
HV7YGzvRRkq8JJVvAsbjcrjEjp0eiusZEfqxBVUS5lhy9IKWruqOG9X3PW4gZzFEdtmeXb3QxtxF
G1qx/B3QMMWl4cVLIeOcGw74rmWYnyasnjkOzJHa+DgFQ9awWf8FsxyWdzNQViE3cq8FJAc/TJju
9rAbIT2WBW6JB/LDP2pVgpb/0cliJ9SUszoJRQGFVdUjvAqmVg+URYxLb6PCm78jT0l0xgUJupwY
4T8O1J3LMdDH6v6cHxyRMi/I1CCYtlHvpfRaRls71omUQ0cdyb0RDenYXm9SUFR6iHE6bxYaFk3F
cTqS+bKwibfWvIv3JZgoYrKKTVM3SB+QRvAH85yDbQDqK+4qN+H7nq+v67ZlXaBe6tm4vZYy7RaL
xS1NODtePXQUc9loRuLgvyQfKgZR2oMdJhTalCjefuI9l2xZSE8m93cL2edf0mIgqzyB2EltJavg
dnvV/i0jbyWqxmB3/PjSnSbh9vrEo823Mc5ieu9A635VDLHLPGWZiOjJ6qjI6XKozb3/wiAM9s3C
QKeMl5dwkCMjdWMFntBc2TXF6wSRBA4qT1DQTM/ekZQG/UIu+qVBGa4DQ9jhMRZHKs71wtXNT8fT
SHhH1A9iWO1VZehRalJJsjfwvy0mtZtuuGPwIyp+EN6HTa0pztXIbxjnz85hoaHzoLPD7BouVVCh
tv9c4ZVWQvr1ncyCOgRUaFWu2gECCPFuX6b39TBat9HiFpbQR4Q1qH2lr0RPJ9D8GeeJI7HI28ZH
gla5FWgJOB24MqeUEEZvwxj2fnxx168DXhZrjCNv4g4txZzOPQa0jU79T1/SHrZ1fcw3x3msy7Ho
2alR/XsDklbAG+sVGvKGrIierv+zn0QGV7YbgPCJ17+gleVkzp3XnFlf+P+bUmpxi+nEJUskEFH5
8q8Lhz9Iwf/BOqVIFZJ+7V1hpiiKeVBM7a4xDncZ5oz54a/GIlOG/nGqpDPg/cLH/VIXe/JrtNKk
6IbdJQqA0EmDlT6wI7sVrGPbz9elB9fzhs6qAfbVgtYvvJHGFZfn8G0YzUrMQY5cmol8tL/gxicQ
CeCbjEEYvLugmn53SItpz9wrcouRJqhQS9+yITyoBTKINFIX6yUM2jSqWm9DLbQ18VkYjS/86Ofb
pcKB334vcsCEukfVv6OAi2VFgry5U7e1wRkOACZra+vulczb4ATHpGJb93tsTKW1yYlg3gBuBqcR
khyDcu0HBC0f3H3P/JaT6G2kmyEcDTn9rjQi9L3E3qoPRFs+JOK98PSazFQg0MGsZ7n6nn3dcf9z
7MORy4/RMD0Sud8nDU1zrM9P3hIfqekNnwq5O7yKyDlGWaKzU72V9o5MxQnHY0RdbsAwjqdBjRk2
nX8IL4I/oMzksTuGj5uhIPoY95Wksdw5UKNM2M/w1zCvWtlma+hu9MgcJpAucUZlLX+0WiLuvI6Z
3T1rXRCehi8X0UzLersNPFgauaXFsDYU57SOGHaFWZdLOQw5/F6u99JLe7odKqz3wltKq250ZbPi
lJRIvJGiNxsYLCKHq372gcssm2tysHwub/LhqGPS57YbFfxK9tQFhKvxLZikS4fEioapmFCnizt0
lpGgtb4IF1ypeyqHK9HW1qyoINKI3785doi/VdDyIMx4NxQU+1KADhGgBOFrjK0DdGOsHCFAhKbW
ipW5EktL6sycr1n8BfGAc6KVVACuqN/E+7JaMN5JCaa3pdnoH/8wefFsVF+fw8PIzaHqXCYo41eV
H+S+OyqCGzK8XDvUwZ3wDyBGQuRXQYcuAn7S0k5MSnGZqXi8pmCwPI26XV2Irtc5fidl1YYsO4sg
gZoGL0L3bXoXb7frIrgqRpl2avDzu4Hv7mkLsne8qyMx0EYsLz37PKuX4dPNdTmswfe3mROX5P0V
tVvyYF7XsqPDBRmk0pIxRAlfYDskT6BisfsSiTK1r6z/FH37LavYgJw65VGKVTuXEW6euy1xZdZ4
2m1PoPoMN33W5zYChSaT9hR7hORo4DPInklYuPCH09fm5XAr5/xFbqZ2EcF5gbF9iEJ32mgxxsWX
RyGdDuor3wKFKesbjsG8U9rfOppgH1z5lKgaS6oTSdD5tF2X0uVApOe4bErbf9ob+Rg7tLzUwXUt
RUi0j/H0K/wKpykWsPbQUhHZh71sHxuxr5MllKKvTc7Ylhv1tpGUmnBAF8ACuJqOuFScXlO1Se6R
mht4/yRi4KMP2E+B06obC6gDpAdL3pqLxWESsY5QBfHiEgtSNKBeZxnMm7yWTYYBlt4ZYlQG8D3L
DoeWfD9MsU9I7bI2pKrni/zKkJjVnGMvMb4k6I9N8htkCloVWTWu4qSp3rxxVux7k5Th9LOnEbHJ
UzQ4mMMREezo2Nc6ngnNDyrcuBOEBaodkf9G043Qmy9GYIxrdSvVFO/F/xuaxX4uuax23fgOALdp
DjSrqmNEIf6NP3XxBBLaDzwP79ChI2WVYSQIzt1G7+CxApRayEdXYEw/g59AiT5iP1ww7oYxaJbe
VBSSYx4qN5cNKNHy/vgrioxFiTkId+jyhoSq7sg/QdSzuVU6k//x03Rk3TH2wEBker23grWgzPf0
sFuLkP87Orv2ynUvgdTErd/jGO0+dPAvPGWXF0Q/s67Dqq+Ec+0OlCJaJnYMkbXzTDgfWycaqnCP
YdAO35JPJnnnPKwWAWcE9h+LfwcKiuMBw8eXPCwR19kUU0kBv3NaZMORc2Se+MbUTgLPCZBOaqKv
+WGqx4Fav74dM5q/zoJHzUTeGzzoFCxiAD63WvN4abd8Yx0AAuKPjvUIXHbFsb9NZjhevWRKwaeu
bHejEe+5G8hZRhRJAGM9fk8A/GLBuLwYcn/IFUqXVQeEZloX9XXiT2LY+86SBgOIc4/rxUE22ubb
CBfFRBOfOQ8FkPdwuOLlQRMJRGRrXuW+mfjtoWIoxJ7VMmSTgUapQllFJ6SR4b0GhEjcJOtJg8OU
vv96xgDeP0fmeium4iVXv8Q7Sl3def9XwyPoMet+AzKKKW/HuQpLoOWDlJwYwTKqYdd9yxI1dOQT
LTjceUw4Sel1veTbstuLAuSpkIb53VGShcjITzkOYTKQ+eeA8pK0GAgBC8+ypTgqbAJ7OFGkb+OF
8wAMM62uS0wQejwZOBVu0oza4JHXC9Ih0jsPubUQJfq4YEUgLocA2Hrd7QnCr2t5rypevqZDLRGb
fk5JXVrXU938ZGo174LeAee4mbUwU6Yii58mEv6gxdTRi+GjOg+bUehejRvYtHP1g/5oDzq6FBG0
WtiNrESJ71qwuhGbwkNAwAHlMhhF67gv8GnE4Y9mgzzHuvqSbGuLSAM2mQpwEeLYCb6bguNS5MHI
3m5TE7GIDFFwWTlp5oSAx0SKbU7DgTTfJ8LZ56sgxKIdObQLLOHMBbkYEjqLI4Kpg8sUh7FXNaiY
zcSnjqli+4lKGph8kCfJ/NGRpLkrEpp/MwruE8+eQhE5qc6NwsqUZZop/ogSCE6TM5o3+za4BrHg
q1fx2zL53QnXVAkBPTdb+raFQ8UZoYY7uzK7Pr1HU2W44VZ4qNb8f+iJvk8HUeKzFcxcRC71ud/S
BUBI+GAH6f5Iy5+aAiUUj24YAzgZzjiKpcSuP/b7hYU4P0bdt64W0tGdJSdbLsBYIaL07s7nGwmN
kFmxEdQCX6nIfo4wxa3LNu++7a7G/vC/MXtO+Svzl7gb/RmNAv2z3Vamk7wTJgXzC/Q9s6jGSPyU
4HVnNXzXPSWBnBaGJIB9/hVq6RecomzMBzywPqDV4fjIaAaruH01NBka3JGC1ipO+qoygk8v/MyD
jFjCMzIeO+xQOOWN7pkU2b1secV1flOGBkV8W67AkwEEX9gJKhVaF/xAbxnvRO8pTwFS7nyeHsGs
zQIBmxjPnTGHkaFiqgzfciMSS2Hhv5ccuKIiijMFi1thZDdjioeaYMcJmM7PjjjpPar2qZ4am/2Y
TUu3BnA+G0cwJslw/EfbHBYsEUXYrYaBNg04NKU3DDNLcOSpuhaoPGsqqgNw1H1f1DxrUpSe1mvy
1NZ2VGDNCrPI65v7woHS1fmMt9j5E5QPlh1EJwM4BBf8EijSt3vNJ7PeS+3mHEli5ZYaC9dxV8OE
m5mgNFOe6x0X6aA52XY/DLM3bMcouSqnok8DSc5//7pNsRdHGh7EzJMR/w1hkp/9wMnF983CvgUC
uPCuf9w5KxpTjH8/HEXk9sKUwEBHXcGoA74vVEaw3+CbvQTzpxXzUbbRkTlpCv5CdKVACOBDEOR/
tXT+gCK/62qoxlybaY1+tAhzTU2vmB8AplqsxaK81/jNpOB/nobM/wF5ggj8kTeICp/9l9AliN/w
eTQierVpuPs9kqNxPv75KgwOZ/Do32ILRN23dH+1xUKywVonbM7diVwTkFCT8rFhOPrF1kdWTmGr
uzvzRy8f2sxgUZ5vp1/BbyVH+PfjBt/34zrEFP75b/IUvcF/dFnHBQXQL4u/ZQGq734bEoemsEVd
trPedEPyY1LtaP14cU3SSdvGwb7bKvkdwknl4CRLwqB/kPs5x382quyimbpGEnb7eF5fEpYnIvne
7mXyqbKWGq0w8UE2KfUosEtwWAFUsNbH6iAL4hLv1QbGo8MgVqJM44RX/sTS7b/W0RFL+YEKtwat
TSX7+8cR4gkofG756jsXIXAn75qWs6TFXzU+eCirGOrmjCzRBS8Pmbjlgy4KJi4DTiXxVxBSGbAk
sgWP/a70WGeNBKBsfO+FGNvttMlCOrNuHptYNb+b8Iu6NeseLISqRollKA39EdUCsBh9Tqce9uj0
UHoLfwvCqQsaQiH8ze17fWY0+n2jLzXRXNA8dJ1cNBHWD56ywJGtNRi6KwFpiHmqrmZPmWGw+e6K
e0BjPEUp3AxlmVmhgygXehpesDkzx0pN0UavEyKtbjFL1DFrsw2Bqrsi7Y3oCQecCKJtXM/uXcJk
W900xcGyKZr8U42HVlupQ4YEIOBBDfIsKVWEsmDmjnqlecdXOnSDqN0O1imRFnKhBzrWx3Ox+O59
WuvOtCythEamgFehL1FIMxz7pe1/APQRHH+4Nuttp6S3ZkK3Dyxp8+tz9nWS8Zk5j2s3uP6+Vy2w
0kD/HtLp5io/R+hADevn8gHNJC873hiltY70rcrtkd/Dq+Udbpn/gnejFLaJEAJjdBlxKOQaRCR7
n5GF6qomPELo6lvl+iOxZSjhAteCURHkMBXNRxJ/KKA00vv8uzBiNDTrF42U/NhPozU2HMGSYYgx
uNT+wK1InidnUdCV6k15zFQbaivqhJrg3G5CeI9Rqa3u4MigWbAvPDiOMbM7LJBVwNckACXyJeQO
BLcuCPRyEHCxaq/tkAdMODOt+Aw1VGe+r7UVbcLvqiS3qR4vkMsaNPMf3YSELW1IudstIZ9cEIow
1hWJZiZyMdUccezrc+Z0M6kHKIooxiZXvMAqILbQt+CKZ5wHtOJCkMUmrStcK0RX0g8+rUsXxFK1
9vezRrZ9zAYinaYaXqdqNxCkXgrEWJMp543JVsPC0UGVirZF/kL+6+W1YcRgs894lN9sE057B+NK
xIpd+YmOeCUaSiQRvU7Rmp2IrCFaz+ZBl0hI1QCwFdVNhW3SxdaTU/CV2lrKmrlhwxMUdAwhXdfD
xLdHwsp1QyN00GqDrnYBeqkchoWR+VDj6KhgTS80ECOYLe7KjKjdsPTOcoagUH+8iXamqrQmVT7R
OYzEraG5QKHSftb2XBbWGsHwoRortejYDOI6xgbgG9+vCLx7iAH2sjSFA47b8CD4zLWPmGkrtVUD
nCme2Bf8/xYMecz5D0mUurWJXiBbAVAsRBmvY2DBsx8n08AoOfN0NS4Eqry4LpnCLShAar52mc/+
SJo2T6DZwlUA4TS50R3YPuTH4rEtt3l1Odwem0sIxDUjF6jW45/BPzH1Jf18Azg4dSz5AgVeXSkW
yPA/MRxjgS+wxOg0wb6ay9o2OwtCQQ18x91NK2ghkX+rWvYk0c5Jb/+NreU7Jtix0IY4CyJ0zmTE
z3W5ULh+UBU3oze5t278DoKZI+nQ7oz4S9JDFbbZJug/WjcKP2Uqp7O7OANkouo6vpe+2231fwk/
3koiaL+c0DUUyV8DrXjbuvdez5NFGG6IDuMR7IQfVfounlVJPvWPtVn+AYR3u03x/8JOfhr6Dlqq
7zyKEFlenHceP1RHItvIAehCn8nRzbwd9rB66ur4StZLzz1ftmxtK+kI88qHWggdDNhg6s5TfsUn
FEsNRSkZ9J10UyaVU4lyaXvsx9BG2ZzFtpLReY/7o/SIDwXF8B06xXal5yH+pRdlqnItyLWHjfqF
KB0dgzUo1QxI8dvLUZZi/XvAsgJOYroEGkVfLnnmXGFTJAZsu9bWb/NLGMWc2pnjA4aljt6s7V/x
Qlt/N7b0hK/4J6xT4u+ZvwpSZTttVX2LnvwlO/5l0QvMemuh7pnBMaoK+LJBrda9o9nSYkjqBlkF
QFj7JbEqLXo6s210cjFyfDaiUMUAJX2vrvmxwPKZ1eCOFCU2lu0cDSWpfojjFI+9APdbfCV3jkgc
7a+EfY27vZxjd2t6YE4wuEkoJtMebZuEtpPjxokgSgFHQ6AhaI4uS19YwlPtOJM/H0ap3oue68Yn
kJod05GrNdUND1YZ2Bdx1do8PAp1kQxWsGIF+EVrtAudS7bOUEhMYEMUofo/9Ey3J/U9291Y3QyM
3pQbDiz4ZAzQi0f7VP8fibOkGsz4t2j5w9zIuU6FLPLerjmGZZ15xEaDYN+zE17I4TvWRmNyosoj
rEpu8ZRt8zREo2qWqntaqbSNWlxgF+A3c3NE1r88s6nmzKB5K2ruxyYO4Wf15kKbhzzaHXcK7Nkr
EJlZ0eRR+SldHbv6nOkQWndijYw5LIZrfI+PuFWcZXZ5Kw5laEiUsOLH3xZB7qARPkRFdW1OqT1S
yq/2f+A8ynqmsz/FLmfBuROwrY/o4X23sTfJifewcSaiBqgDn3R4XCMU7kw9t2ScMYCinyXScoKS
1n9BMg6UuWcc4WNgkiy/SRUmlQgg/mL2lYlAaHjy0hE17LL31Yh1lYhzCtof/9wsQ2C/PIF/ZsK6
XfvodwGCR3Bm22wYL79epvHWKAtTsPJS5TNX+z1jZI4UWhMwDr5EMLITvX4KE+XSIdpaRJ4wi6zd
QYWTvqQHJlQdfPch8lMmUXWwbrkRTR/Oz3XDFTktL3KcJnw831Nhg4Bs2NCbwdnI9sZxUfpJjCEC
iHcB65v1YC0ji5ZvA3BjIoOtP7sGKaN47eUKUT7YeIEwj6z4tWmlc2eX9e5OG+ddEehWFaqWfgoi
C1gpQN0IG8egDG64ADpCnnG9Rz+PQ0Wz1WCXEUp5T3Lp0QHtac/eA6OI0fMPqLqEB3hBEx4g9tSO
Nh66brcKsJUb6ow4+7/WpjT7q2hMSmdMVreCCoVnewo9b8e3hNTbayUhXlqS2z8jYPMxUm/pj2Jp
8TY5ixToxI4u2Qq8Z2oawXt2lkYSwkkLgec+ARtJrHWyDfRl4vskqHUAQCKP3hgKT12Zi+6kubP8
1o8RnzDoQ0I2RA3RLkmrTD/eH5OY9bws0X3Ly8qPfly/A+Th/NdaiISKFnKhIFoLN3DFMyyqEcIs
M09hZm3dcJLjJkQ8Wi8NkLoFD16AOSPq/j6hPxkLBW2iz7lAhAI4qJLIXrhtDclS5HDZvhNL7rzh
9o1Z6yIboH3TyrBReby66som6sftTVybK41QjwVq2kjvZrOsMn1rGLKnpbEJMkOLKSmpTygZyjyf
AazpH+65vj/JP6NDH0dkYP2kvVVFMn/KNK9O35Aj07pbC+scCxdCPERP+0SOFt/MyyqjmqYAhULx
Bgv3ob1IIuiaZzYZcQyyYeDhj5jFBgGpeyWgyW7+bwmDk10oXsYn9q0x2HpLlO012agjZAEUerja
0r3weylT+PYTk+dzvuNBkfMxDgMZf2ohGxG7BwQOdF2gK6Qwzf1B5uEnlo0HyL8Uutz3DWdwrHl1
F7f/o4wHclTUxAvgaBjo3wNVpPP5ZPfM/Vp8bJVv9kZMHw9I1tjAomvBtOBtiU8jM3MMt74JdOgw
UkAknOmldlWaU8hvVYWwsBdjmmykIr4rYQO0RNTnPjf9uM0PQqmL45ih635faExOnzMan2ybxxwa
ONGXJmRbPrXhwJBIUpKembiL0Peb3ZYCklVew52ShwxCEXkJwxkbuYLipNZKNhKSspbv9ucliCmV
FrxwFzrupW6Ip9QtXPBBtqWPB2/KK1SJ/n4UqsVZA1hfka1MpaYcNQCsr71RUYkv5Uz1gxyPY/mT
9j8yL9SAaBDK1AUcq/ifjAk3ZnFA9Al0CHYsmGHb48H9Zr88P5cRiq7oZlV65/41ji/8NBEwBz5E
OYWoFM1CB1PZs9oeUmVprKIhb0wQnNflt6EqduoEzvVdNBBu8V5R5+z9wv7E59GkgS9Xv966oLzT
WSDLoKlGwhS8PRYGcdLEUSZJnAQRwwG2OQvpBQCzrlisfr5n5DH5RypI6pR2Y/2oxvSsVasytwGo
r2/B+jrwNn3+jGxlHFh4tuWY6secFNuY2OTuMsewKXHNWhB+GNDTSbyVRmhlPVo9ssTe4OCCQJuA
WjgBVPIsaj2AqPMv2f4qPwkRb/EuwKl6kpe6H0xjzMLbuVCwNQ2+EWidNjhz+9H6ZlFcR45Nzxq6
Sb/m0ZM9RAT91LQVfUXoOrnQNEc9NFAS1hy4fGWj3Lug0BomW7q2OkH/o575Q+54vFO4WdDx+7Ww
7CWqvTWOFfWrdUZ9c0VeIyqJZ4bsUYg6v51dkztF9Zot9ce5oAbgXLhB+aEt4IaueQx4mEk50ycl
9YD8bThp/8XrYakR22ARLkvHL1UgAVV9GTIACgbE7YJ9gZ1t/XkxmCwaPOOTzA6hJmRhyYUnB19g
MmDQyeu2ViGiEmcGhdUr7R2k19lU44MsNlORlhrSfT7u6Iw1LLlUAD+8IRRG84q7ufOCK2HlRSd4
dOj3TiUdGIkw4H/Z4KIOXe+xtIC2h/GrSr7l0NBWJXwJuNmXD5ev0jBRzEBWMZR5oeMr0k1VY/tW
DLpOx5YxQhgpC09px74h3snpsX8hxR5+HQRnOFCFGBBOZYyoULxGzJ+2oc67ZfAaiqlznqtxBnGR
UZ9WkI1EaAqbLMzfIh6X8Dz8bMwmncAesVxv6YCy00hQmBdFd8GgWc0alXilpsuJsJBwrKbjpaX0
4oJz6hsWJy9XIs3BL52lIbVmhKV9+H40cAE5cuQ8n+I68+ihQV/DNj85SkRhNIcFYWTMiH6aThlY
PcHZay6rhZYvNEaYlkUyaoItVjgx4z7GiZv+SPydbs6Rg2cMIHbYk3Ai/kUMQo1FDkHCbZPlb0yu
DlERRn8BSZgNicmnNF1lb3Hv6OWeNR0h1p/YzwSMSNEkgkYh51JAISa53lSD7Jk97d8jRKMe22RG
85M5m1O1kOE1wS0bRZjbQ4t2p3dGR5Ps46N/oGhvVNIRA6OI/3B0DzTD1KtaqQS+ozqIN7GD8Hak
J0TV2Oj9t+FmB7tNJ4JY0+1x2kFz7N56gr4VJBTNiccZa6khj+PV4+Ouu9EwbGN35T08eN/wiLKH
o96lAahlaDDJY4wniM7t7ZN+Vk+E+rfjFUfS8wFWXiFCBHU4dBEAZs6GtEFJKVhGTA86yiDIWjUL
3EAEY6KLSnBzJKw+3CLX0AwADCiHVO0FpGOYgAzBIpLBUJqrZJ+EXZ0JSrsN46RZhxkwO8qXTEnN
nB6MsJean8/ho6oWUeR7MumHuV7xfUWJxi+rfvcFYE8CCTGJ1wG6E691SOitsUOjyGyba/26DSpm
3N5r4C/Hfi7oswxjH7pkuxIUStfSw3bjCAA6uJH4a0L/cwjNVIWzfFuTCv+4CvxpX+CVkAW8U4Wx
ks64yNIIas91kiE5wvjjnWOenGENGvQOYfioZXu+GvQLABN+NYixKYrStk4tOg1heUBsSOOh7JTm
wvTXH9ftWW6en7CffVlLFf6/+DrxlylXNs4pwftymTsGaQJm5XzyUymwl1l3q3ZdM+A0tkF5bdbE
hmax/6wSePy5vY/QplT3VCbggUMTTP3PMedw3xCJAHgzTh4WQtTbrs7xvzItC6ghuJXWvcaa845c
EWOInuOebdx0WGdBJEj5ObLiEpU4sv613Kz08rCXdOlTzHv/KQKibUkf95FnvSO7iysXOh+yh52t
2IVqk/BO7pKKwGvMmYVHmhCFq/yzk+g3ZFQjtatiZqviJYU3PzxZaEJQh+GBHRc5JhRXTijanuWZ
Dr+25FT56hZEEH7aQdzXf4D5zGY2XqP00w4RbtRr/AQlwYDcm4So63uFcqSKfpgGsP4bJ7byvs0E
xUCTDquFQNJ3hMULa/sMgZvkmq679lDGdBVkr7GuR8vWtlURIqYKuiODc6j1Kq7RghaOu9pnj2AL
xOgvQmAh2Ls2T/a2IzKpLwyL+cu4S2pWW9CdyDsrIB16rO3Vac3iM9QGaTYkxoP0itkMYPipZ1vH
usQZ502fhm7ep930sIy/E/k9M7Qg1Lt0uZW5y9DJG6pyIA4ZQGG7DMUGJNvytAxj7jhL8/DYijeV
YUHLZw6v/znNLu6f3YLSQGdEnqWHrsazkTtwA8od0fj+cPq7ezQxTQ26X9HbnYzmNSBme9w+CKUk
yUwAA6ATPskYSmqqjWh2aHJPcW2DS3P364vLXQWWxrRbwnBXTDW891akY665AzXhFwxj92fLpk16
2A5wfiDnbNDSzqqMg0ep5cUufpjCdPeRsFmi+98lqrw8SZbs+6toad+SqidNld2oLButfNfUND4Z
IWBmGjK0/4GFll0jQehfM1MddFhsKnaahy1RK6MxC2snvXaUbnJtL4uPA7u63NAlxIF92qfqXsM3
ipY8vMXJOGM9Piqx2i/sA6geMiC06DDtiiTmD5S2X1VcasU00bmctNCr8Ybf2M9m4k89JjmyRSzZ
TPIVoAxBMI6BTXaftcuWDYHjV8n8iznfYbxiWnqGj25b6phEh8W1WudaVHs91VdcXuVTuHG28W3M
SgMbttHWeeveyvtQsKw5WpwrAxx4h76zF7UsatlOjbG9G+sfMx5UqvcPHg2a68tfaqf0wPWfMOZj
FJDOwD05FHEijc5AqOl+BQDRmcIb7RKI1ep4i5zrC4I1ezYcqlsSfkpJ1hGrcZo1kI9SlzgJ5Xjf
vycVKGC7tqzmYRaHhTuFwGTV6ju8+GX1r1BSjL8YtLw+V/ju5nNZeBSuWjFFC4iFEb0dEU8OW7D6
nRzvAGtnI/dggeT3RQVK614QoqS8GH+KzlRAW0H8/OywkEhvozY+FTaUHAGseCFVEGF4nxi7xucS
w5nGCaiktHm0n+5cOc5sYw5hZL2FDk/mVPaD4TVf7i/NuN14UzyusY5eICcezphshymrsGZ8ymWY
T59lYCEZ5B/7zEr1AZJ0lXWnB+vNZ2b4mdsYsxYWDzUvgBCKAm3S/lwo56JcBKCIm6o8jDpo4fjl
YioCCccyLHlD3q0PoC+AnEG8eGJmUT1s4Lnyx29v8OepB2lfw1NvgABf1j6P0yEIWNb0YNlUo/Oh
hC7pt20/Sr8bKDl08Wn538MJk0zRju9lcnh7zXPfh14TBCIoaQfCgled1zmkw/iMcBWUgJQSglKB
w3xyLk80afKdLTp94s9a7TqAC/3Nha+uqJZrDimauKOdp18/KAmn8j74Hb/wdg7eCWY/ex1buLzv
q3FhB6IesyEM0fYjekfDmpCAhLYSFcMcavOZKi0UbtluXgIAWznpQsSTrDBNp6oeopVo8BDGK+c6
RrJvRYSlVOQ3WvFsc21W6DqkhWcV9rPy4AVJ2Gip5k87su629I9PJjwr5k0pkRGTzgNodhJnQnga
vomgvifOU/kZeDgd6Chm4dl+u+bbrGsXySwW/zmGOid8XEvDtx3HOV3NWGO2W2PpTzOPi3U6hJck
atSUdaKX6EBzJpLMiEN6ybf2jCuHf4yJ6CilZSTmj1DKGIGzdomLs8ZZHVJlYr4JeV2/uIVbEG9d
5BsyEZ4g6FeoedXDeN395noVMPf8rHB6487H/n3oTDEensCK7tlBVTAK0A+6I73HDWQuCF36mohD
Q4JEt34aCj+OvgYQ9jiBbnxlQJXccNZNEuozC35EmZHWNNcsCD9S5sudr2szUC+pfnEwFEJVsTSD
B4Pgc5lIwyFU4P7j1B+FAaUorN3VM+Fr2D36Wo0Wgts5BVNjcx7/wuIS+0ebK9Hkt6Xka2Ezi5EX
7Yqs1A1wu3Er+gVzz7y81lweFFWLUEOOrLvsEODXTjrGOwXbav7UFztoT7ekCzh8lWUDiWY+epeH
2UFRhXOyGIJ3JPur6HiIL3ga2sgyFri5ZSBRMmuVDrlCk1oc/9bP3N6xxBQCiDTheYjOad7j0UyE
PBAKsi6ehYSy4r4z9Qw6KyjaZxHLI3hTb5KXSZjaiC2lZehoyZnzNlpqMpFib7p9oHee8g1RMjxp
Qt9WGjb2pipkIPSXYLE815GRZyk2Gq4/HjU4wbp7N25QpGNp3cMZypcmIlcMam+gKfDywmB3e0wX
aZ2iuwAVjWTtiz4v63ohXgMWmkD8MhtojJV4JOPl3JTpAuWNxVqp0Ret/9ryqWG/l2HpGiNDCzxh
JrBZHnFwskJTnjFnQOHET2lD747fFtx9FU4QK+n55TuItaHBRZhdDQYF7l6q8V8OCNikNM875qlr
ESBYi+dRfqeEc5b1ABBYe3aaqHzLlyJxhrBHaS+5ke8oqKvgaIOOA9xzsNoHfXsnqI+o4gh42ggZ
sXw34eYogSORIac1Osnk93S8dVJZBewBvo+HBEZdWMCSKC6BN+4qW+IHnFJNn3y5bU9OM0gdhxzg
xdcQxPmFPBT5cD4j06EC4rb5jK1oOqsi4+Bkbv42H5arFpjrdYfZoYCxXD4iEL1wefhRQWPNR7Cd
T+zTqgIPHtn1/jw9s9zaOS9Ojgiu9n4v7gNCG9wzpuLJ4IMP3Lx5iW52ic9qi+dy9gv/h6Ij00m7
tq4SZnHri7G9zW5Y3s5r5PLiDQkLFop5jY/hIkjxNmN1cRQC1t1luKX6jwnp8OlS+chHt8G9E4Jm
DQjxW9ZZDbB1OM7xBL18yM/AnB6SNdWSwDx5+kxSRqrYy5zsCc2+Rn72eJ+LvTLs0LZVmXKtlOYe
wWk4qATB/oI/6sMlSj6qNtsdHzaCiYv7/AROu85JAASyY9eaMB9CAMrf1QebCQuvSv+/dkxkbtpd
FYplWvT8iZB/lk6exA7Jwq8t2etObPqpoLZEsyVWQmtN9croguZPWBRME826EpFo9aE/Bh6/RFUo
TkosceKkSpc9SGTUiRoPqZ9s1i+jn8dC1CZ4XKYwnPEnnUSvXeM+kRIa+NRr2OL3zpVgvphRQwXw
C/iWZrCz1/4VD5hteZZyWngs5XQ0jIp3IIsNUDoEqg4zVQSqPCyOduXWilb74+T9wC5O5aL8MiZW
5vNwMbWKT60wM3ygM1p/agyidhUrjqEwHfSmMhjGQ90Zkp7RQHDg8AWKrCRLw2Wx1zMrYFUwUn5P
eEFLkrCugSGuJ/63ED6Nk2YBdXgabYzBzDTvwLG0MXOKWv2EZiaj+EcYuPm11mHRrNI4XUiesSFa
aPL8K5z+2/VUP0/wkfJYQwtJdUaHcthXaTlYRcTKdTmFse5tgRt1Eu8mtwWyIMAL1V79v7VteeCv
zJvxJnMwKDeh4Nhg/tmPpcacgPqT0Hhqc2vDhrMizodBApAOl93xLQO3zpbIOKYRJ615rcEce15s
LZrLkM2E+GwDlWKLMq8cCgIBOcl5XXMb5xF6+/mOD6P8yurJdkpRz11VQ2sXuK43+bjfV7TyS1Qs
5QwelTO5hx4NSezK76FfjKbIC+/YL1Rj/C0Wk2gSiRHqxsxWmvnreF1EMNHo74Qu0MY8GGzvqVxE
wM1RgakefxLe5azmfq5ozsX/XA8g3bSrb19oswbaqUpetNCx8yqsFKxIiA4nuO9kpcPdlHSTRceO
z+7q++yYqnbYNgiFEN+k0KcHDuTYS2ZiNIBsgdmkHB4rR+jyzC6T/RHAD0jF3i4rojb0OZ4aOqow
qoZZtaGOdi8K+DHeF0CZMcMyx3Zjdq4FqKiYHaUcm4vq7Tfo8EXW3FRHrBUca2eU7qE6CO6eA5+A
kVOGMLJOKU/eFv8E2y69Mci3UclfemJxmd7DVZBzAzvcExEPcaxSoOhp64HamssWfeLax1hKkO9r
8cfe1P32U+ezdXpXCYJhlOs6GbbZL+FDuq11/zs9buyCL26OJVTOK6zsC583NoAQypg1WgO1OC/w
n39G9g1s/tmZrX6vQqjRABGaKPnuz0yExLDxLaRwCcISzvrIsRnQ6R3+zWibFAGMN1QpGTcv97ZV
GT3ACPdfAWF+3hactBu0/oB72tTzeBmpHNSOqpDvGvANh+hCpiTP+30L3QE0Qpxug7DTUC751MRy
xT4nRG9AWTyiEEjHVvkc7BxNmTxUKSl/5xNxN7m/zJTUNREcDLO3kKZpkJCo0TXIIRfDpe8XxaS0
RQm8DsMrCG0yPXpoKGibte197n3iAUkI4qAeaqk/0SKmaeWRh1rFsQkzxHPMcc8kCwg0WGL0x0D/
G3xcHvlrqCQx7KADGTUnVvGXBLJ69zgvnPPLqcMSy/r6trNjp8so3o9qSFiBHg/UeJ46V6wTfiQ0
iJULbcus8yGllIOMQPxZsA6XDtmUhWpbBp6NasCEeTP8Ju2FGgIRgHcMeCBn2XFUkUf4YebkVnZd
PtQMgdh7hF/9ZcnxuEhVJsCunMXD2VVIGbALQIm+v+R1Sge7osJi/ESRPF4OYdVBtCmlcY7LcMun
8gNytWoroRq8F1wZCXSWRdr5l8n5kYf3YsDxTEgcweLlq75273TNrPAeY4Jrf8cksxB3HMFyJMPT
UzNFdaDrSDVZuZ3+qYrLG1MAQV/MEdSwRC2CnJIM8M0iOfm4XOnUzU5ECzhuvAhlmkLm28RonXcR
nLYjkLEBoxKztbnMj/FMFcugeDJQkoAE8cQLMdY9E7n2b9PFKiCHHEE9m5OBfmaaDEdsUQqo1/5d
Cg3xLCyx85LiUQIuUVt/+mhwv1i2eJIUUYy71ZzJUsxt2GwKogRn4tmiMEl4AYm9+bo6ZS4WCPEf
gGdz7sQthj9Z1M/920QofNDt1oMonvNNi244BLJrCUEGt8dyM5c97GFwhAGHJI0Aud/+X97NfzkB
tV76tIZnlFHsL6ieHHf9TOYsisUMTOtjsqlO9iQwIJ8gQVRpwxVxTheV+qkXD4OzriS760j55clA
f8puugnHIpb5WIbCjjRkc3G5weI/UPQiPKH4ldAHkKTYKrnKuyh3MYLLZl3NPkZOnD5t9leNFoRA
YxqxbHqkVMr3129meB2R/kgGmilm/R02B6kVzG8kRjBD3TDUlrF6/8+EDJvYy2zQHfwqw8Jxy0c7
TA2iH5L7ExawWGkYqgTjH1bMHTR2HqZpvLl0qXbH+QBUzFB2TxEvSMSErt1KZ7YBmDxicsnFHgog
49BgzDGPYX6ceeu/AGGds71o59uaNYctXCUIs3+iVyWkFquZJUrJ5Yu1maG/PQclMX/cWvWOpc6D
2nDM+fOC+lScwaCOawPAr1B6WfdBzpfnTm828KuPArJCIhUY1l/7P6SM62GG6J0jNrXB+a33GhxS
xWIIZORdlqfVYMi7bkUf4SoxnTSgceLICImNYsSt/HpRlEKKstuYpp/9djX4ijgpictu1kyKJ2bh
DiHK6pexYs8vFHdv2Ulxre/Wp+V/xFe5ZEVICTEuhNifMZffIVlingRqrgL6hXt/O3J0+LUBHuz/
Jstb1h1fJNK0akElOhO0jZPt+h8PS462q0S0Xrkr+FBXY2LvfM3Ki7jYfCq5ss8sMjAbJgqd+2r4
omeMBrb7zGYRA1QCXPnTxKNVjZDJ0Xclj3VgLz8fc20ZyOM081uzTdjhfDN6+seuoqS5LrJo+We9
jOE85rR0YEEuXGlx/dKQl8Vit4WE1fqM+b/wZtwKYe8b7KHIt3E0VemEQsuc79K6YNytOKT0Rl0e
cJHIy4lNNjxkyOqPxLeif/blSc67WAVs8+YWmvvTOsgAEjNp8fEnIVEjGpSQTAzkRQef1W6uvEkW
BakVGqGfHd12QNnGfYHf2IeD86XNMi8cjkr7pVkCnbvknj8LJFoYWEKRToud2AFrDnRReaWjJype
Oi5HxlGNcRJEblWyhMPPhrh814pc3g5qODhE36WjWfQirVedQrQeX9O9QMA85KFJxrYfdLqkUczp
pcnhrc31kNSVs8QhNRVP0C1UYqlmDEd5XWOVCNm6J3FM3vq4OPIAoP/PnaJ9wWxCiALwc7nWMO4I
iu7oAHGwUQ8X+QlbHBDpbgYIm62XmS7CDCCCmmtmPVnDc5i7O3KWqO37AypX5veFHfFp+hqx5n/+
TY0kBOm6POd5OlpSXIg2jQv8OwlaJ/iOcOI1PRvKwacq3M0DFj4Rl67dOF6b7Q9jbhfgDVBQbgwV
dymtIeXtdsMmp5XM80JhMnuw9ph25iqPA7oK59yhLvyuX+i+Rf48YZs8DbU1tIjrhd453MK2KZ83
zxXRuYWXG+KsQjXUQnYy8DzMIlExKsxxcqidWPqs226qU+D+zYL++Nxj3anseAzSgLlB6p9g1xDU
J01fy3Zhfh00teRFIgPWtTMNuwo42Tl3O46MBShxzA3Em/doTdyoXQA6Q8VHXX2asl2jf8MyYb9R
rBONJ21+0Fl9+jJby/jLdsftsxnyFaZM1BPGYBsUl76rDtDjcio/5KKfPPpk9n5Pu6LzX4me8Kvq
yClhl2WPs6k9vcqFoy+I85WPc5e4kCqXy5zy83WvTPsm+YxRiW9qzj2po26OaVRHfwUORi+Fjpvm
szWU4CV9JPOzfn8fFua2vgiBjIUlSlRqw8DgkcI+b5VQyHdyoEN2WzgiT9jhTEyUJCb6eCXlWCsg
LnBEWk6JYA9SgLwE7L7FPwG3ymdGKGflT4ptbredWlR99GCde2H1HohdYTNvQWmJVKSgD8AvHPRG
PdA9Dn18oJ8tuCXPBRsZqJ2fMRy9RVMPmdQeGdF5IPO3z7GJWmtewoZr4Rph4bnhR8quzgjpcR/K
xO97S/yae38Mz5hKnhd6upSvy5TYa8jfksWTuR4TIZLDrcmWyjgTHdgOEiITKKFI7k/CNHAxEdSB
ZEG6pC1UbKFisDr/563w/NBPaVdF14F2yO0KUqFMRNj8h+S/Kf8KaowYE3ba//rd3c/+3RjzDb1E
wlK4OwltWeVMZJzD91GWyil9eQ8dveHdo9FMAsNpKrY6Lj/LLM5MHHiL2+eKDbBCj+yJxLXWdvlT
rWa2afaKuZjmfAyE/Fm+ShVVTz+V684DBSXvQxx4LzwnJOlKMH2j2y1GHHaewlFtjxnetPZrs+R5
48zU+iCT9bpg3ph4e+nDu6On3DP5cpjpev+teU1s2FuizC//GZmlnJR5JMFB7E3acIdZuGImmwDo
HzTuybTulXdqiVR2Ftokk+1/NKMqaCpvWZOcfh8U8mpqNmLTxfSKNsk80722G0+i9lyKT1bJ/e9k
hKBSn8BaaD8T4auEiYNpP7bV1Hnn70do7yH5eQHNan0jliYeErp/k4orQXoMvWoLwMGTPCmnv/KP
8+OO6n4JEpIEdQIrNQ8z18OOCTt2C2MEV0hGxVge74fvGl3iQsokLnVtbaGq8yT45JmyilmDQisD
3xN7FMke0EYwsf5bI5tqk1WL2YM8uMmRN+9sVTXpE4vg4DIJvJLjG0WPDpeffAOPpMPv38Frj4mh
AtSQmVrwmOUuGA12qbuBDP9B+jo5U0B/BQWijo8z+ULOrujym6cE8JCz+brqythR7TlqU8H9EnVU
r9T9G4Bw2h3mO5vVtUJL9bfsccPOacjvsGEUNyapwz4lKgge0tz8srFDMSvXgPhVsXunC89BPUJ7
XsXNopGyNh4XHB4rMKH2Ax3eXND5s8D9NFWf9kp3TT9KfBsU2STrOG7eHvwZt3sBZr1J/1bvhnld
mLYbSJTvpXKJKkeGGHtfVPsC2/pfIa1wdJriX621t397zZjVd+Ofm6h1uU/7D8upF/nYZ4wdRlZZ
PDS2ISUez0kR3zju2l3kA1T+0ZTRFoggceYLoNvMHIXX3XGv+LJfqpko4hm9ImEg4OTfZGas6DRK
2GyQdavY0nq0A262ZcMna/Qrt6vP+IWU3qR2m5bXdreLUUKaCeJcyVaKS1aPgEzg8XG8IAw+tLd7
Oi7u+gAOQ38sVzJ1Cg2SeYSAejuGX3QiMCN9cFcMzpYdVoR/3qoQidEvgxEfLZdo9AsWMjv5ghDC
rvZXHRaAYtHknp28x8a7gxb3FRem+GVqbHJe932YQgAPSK0ZQm4IDFjWruHyI2FYws7p15rFwVcE
CrIJvuYRk7YvAzK1uf9jrjqq6fhXZC9eww1LnHpWDBGW5Gvm+jUv02sW7zlB+ZxbFUHYodiooP6j
3bFgOpvOwogXg9ELk0pqcywNrjgimp9IKH1qKFzw2XYdqHh7K4qetC+jzkAEErQhlPXifOM1kMdT
e0uMEDmAJOBp0moMDFdriLpcdYC6yF+aLRowyqYPIlQlrllKzIKMMV6vnDqk0JC8PpaEnfEeoI2u
MxCz6JLmrymAAOGyyMp3e4CSzPe3cWbNYq10uUF4HKAHXYkQ/gIpSLKqJEladpTUUG+LpGVWAsiC
AYWl2kxQJ5kFPcfNreurr4urB01RYQIZNH/u71gIn5HvlD8h0m3+EGaWorF5fcLYgKxEMb/jK9HC
m+eG7+MQktr36R0pK2DDZT/h45cjSpYY2vHJQ8ExYFd9oT8A1/aL50Z7EJeq4zaw90DQ8eUznhgF
PchJLqIKLLHInWuf4LzlYBfjq8nwE5nmTRPkgjk3c0EW+h9ZSiKAIQXGYigFkcUJaoXclLwYZ5oK
N4myUHsy2vRnRfwvh5AtHz8kZrxSKehiuCKWe7gSWh+DfdpX3Q0kOSN0vqVzyG1ddtohBluG/m6Q
DWSdf/0/6TgWg7XArWWrfRjeINyjZO8kDWdmMV8fq+G9I2LA5tOlUJ34VwQ13nLMrL3FzY+1k4Bq
of4JC4HbUqMp/XcOuF9NU2Sxs8+ZWMdce9Hf1+bkwaPsyqtKTUj9wehYChTiFDSdO7mJhQ1dLWjJ
kGV0oegin0xk8K1OwsnXcBVXmbKthve/q1aeukngDEECeXua6BdC4MQl3Ndpfx14x+Yhwobop+uP
fEKW//BEnm/0AKQrOSwWnmvhvab4oStZJfmKf7jdf2RAtww6Rc29rDcJ8gdT2QuIn4nrxuSgK+Oi
eYNqv69fov9QeL8kDevceNKh9yfVZP9BEhZygNpN5XnyXXHDg5pc7B3YoWQd8HRDhHm4n//9hEDa
1RZN9rrwyqgOgIVPduAhIZodH6HvZ6A7T6WurvL9JGp0v+ksVxJ3wKKR9HN11qLboUdGpE0BGJRa
XT9HLIuuKV97Du/f1WrXEM51cNSOxEgn3DnptJ1pdLPhT3IkR3aVA2tld/tq2Yakph+Ijjlnv2TH
yNPxymnsQLPFfyAFvX351fRLdP+MWUuh3pIAIcKMxz4u5i7+8BlAnAAHoUSF+HplxrFT0E8TDaaO
Gg2SinKFieW51L94a7JqhzK1Srd7rEAw5i1HJDIa1hTZ194z7fZmPIlXYw9E/By7uhcMgFzuSORB
Xy2Zk9mu3UmAnZOY9nsVtoyGkzMCiq7Y3naHuNaStPzUIaJWouYgXqw8mFxYoffMGMfXTXJ8+4W8
/fY6/ohs2kiq7YcelROtgqj5pWKoTyDpGHBUkpky8SmWZIqr5T7cusEXv97qTPRm0Gt39KcdEegC
TsDzpoJbL3XWhQCXyFtvtggjjdz2HjzR07V06cHn3q7fm7VF1hzyTL91Zy8BVTORNxFpENMZnYNl
icGZgjpaHLOXYoSlUtn18D++X/DFV7TUnCiWNrfV6AiEfbAp1JpvXBorTQ75zgiD/mZfDtG88IPG
pT8w+wYwwS/xm19UK0UKhC0SkJwAHGbtrNDcTO5GnEK2fCoUju0Iq5O0mGEcbgm4Zju80tAHXgiN
ChXoY+lVO54CuZvei8Kfx7cBbTz8DC8D4/tyaixFPVqmGN48aWLMXwVBSYjqxFjxlj++FIf+WJ9I
jXet4uMVh21iIbj/X04DD1d+H+dCErE6DFYDxkEMPTHC1fSVv0m7Y5LBW9cqyosnyLAhD1XvjeAE
sk8gKxG64DmfpJHUsejOz7ksG1c+MvOqBOBdSLRRAEF9KZu8VdjXGw8XOlmjBvZ3uTlK767/T+Lr
nYUBYQVxfSBc1Dy5nA5WxFOKZFHkjSCrR7FJIYk62VeyOQ9vvammZzirgAaf2mCHn6NQ1VwdwmvH
Q4xoW/Gj2wpT4fX2mXDJQYJc8vL9iqf3Pa8bREXOUa1iiUN3WFNc3N8V1UU7iBMaOBgjy8IpHDqL
EuyNKaA+a5SkpFjq1W0Tl3PM20bADwcHv87Ji9FNyLVLNKmBx5sKO35hSABb/LRjtXymZB53czYj
/+pVFA/LPJwvR+6AVmMMtKxLLDIs7pxZ9+pf2RI5QB6l/c/MCd4SafxdEUNhgG2k8/YTezHA7uFg
dQob77hDWaHiTp6Vl/s3xr+Wj3jgFev3rJry1s6g8R3P7GhPVj5OG49AB37VFObPJsmiUziqJZfH
chc9o606FEoQrFnvN6lLHljA15iegpqJjIu0XFAOchz7HL26Z+cB3jNxS1WI5KuUJC62Tc5EHdrM
ydbkm2B4cDR5E62ljzo9p+uaf6NOUqDCweFBQmqlln+oGdSmgLCvLDE1U6b4X0ihmzCM24LQF/K+
+lAN7+svmVVFaoZM35i+xoZD7fJl/t+2A8MZh3HpvkWppz29fDYpVJzZkFppOwS5Mgk4zD7ImEG1
66w+bt+H3hKNzGDI0ZrkVohK8mjd4mvGj2xozyxSE19XVM/221YRj/onUneb3mgeCIxcE9vqS2u3
guogNnw3WLHM6RHyznf/kZMvdppv1nfu4m4m2rcSbqI4mKdf/5j1pUF5bqhUaEoBz8AxFAcSORZs
WwV6ee8LbezJZQStfM6aBfiO8uQFi8Iu3XXAm07B7+6bLYiLMSBiNaGIamB9z55tRONEZp29ya2Y
o5eeKjzMEWtMcNxKuZA027LVHP7Qp1WaeV3nxqK12JeY+DKcbQFPOo74a44uf+tmaJZvp/70bNfU
8+TsCaf7hNPCwTNydajTUV6BM4KkinlFsSjyZiFdHspLIY2R9fqHsY4dnlUwUXw/FGt9uvK1R/vS
BaQigzY0i8FfSIkEDxOWoPm2etewixIzkA/9co1COzEUUi7Y0iG8CkI0AGgTVYehKDnUs26EHXBN
7fd+sNzgU+a6N5vxLks7f9cceIuz58B/W64IgNAGO0ZBuk+X4oVcKcmZA7rFwWSoiK4dedAyDxi2
GAYaDG7i48a9uAK+UY8Is+WzFF0MaC9omO6TWMz9e0H+b0BQABhDUw0CCynrMaNhgOl9Whk7JG79
f9CTWMqVMEt9fXB1CuWl39jNQuWSQYcTMDW8jJvXyHkOfX1gxMDU+KvbdOvKC0ccttLnIcLAeREC
w3BQ7kpIV+ncZIAhYlqO1Wc9l3udeCAyW8+cHjFnYm0lIRfowYoaTekoqpGcIQ+k89wldCMWN68T
kcjmlqEIU13w73TslofGyVTJNFFWfMQjpl2iR5FesGf38JVrO8GfmfGQaJauUTD9fMHiExzy9yut
2AzxXVy3lfnXwXQ04OUDM6gqwujF+7A2z6O69JRrQw6zojsHeaZWKG6Zo0X402km2RzHRYtKQFZ/
dWgPfeZX92kkMARC5vuNDQKe5+UL1/TEdt6tpWqRlOHMR5pCCsJ3cvHIKCUuMDL0oa9msUBBzE7y
6hUKKW9BIjOz92xBoeuwcqQfzgMRWoHol99HFEvA010AA/qIxvv4gjkHJEr4gdWP7xeqIZy7i7fc
L70Mkt28KXqzrjnPTbk7KoqUPVkzv0vvc+l+3ArtL7tNYPdnU/mSX9LIM6I32LmyNZUHl/edf5Tw
JyOSdRlOYdN9y2NlXBsuGTujf2o9J9B0DuPmAeiZU/1hSSZqbITM1CaP+BS4nZGt5CRSRkokW0mF
1YqvMA//EtvHjSdx1UAuNZTc5WIX5SijyiG5vn4yMs7ugOmKmjIBIg+730QojrVioj/qgVQNAFEv
ZkPHqFnpeSUXAf7kINlI57ktEaiFG1UIPEit4FNUQvY64KZMKMHr0JiFsMsOv+s/HnPlimr38lQB
pyo7VGR4tlHHoB+tZWkv7eRlw0RnWHO/vvyH5j3Rwl+j1W9CQ511JyEmQtVJDhuRz7tLKtT3ZX0r
8JwLpRRoBnuYkeiv6T1LUAmgrrC9n/EGIwOfrshwv524+KddoSivBXmARxFIGu3sxOV9a/P2mfyM
l59VwVyj1ENkHsYxHt5i5FPcvHItiwAQp8DwLXgrfG9JR1pnVV3B+Pr7LFloU0gxy6qW8iXQieo3
ztdxUGiPCaBUgU4nz7ZmjAyX8b/A5QGEuOmfCTq5u2cgUwhs08pDbxmCUjDkgNTItWN7U/MhizRR
NBhttcVwQHE/RwXxZxgyY3EXaoZlPWmQCNCUOBDPH4NYXFxJSyB7hUf4AHut9kjZC5N1SsBTsRf8
hFyb/YDklKgDm/ddSxunAgw1A5+4y/O4Mff2ZWLQD7OMTTmzGVzljk2aqw5sxSAFbCbKhkNzADoa
H5yT88sBXsdYOj6JaTZ00rCvVu2X0Agz2HGQolY/CelKuMNkav91R69J/K+T/vxwBOKULVl2U0MN
NILCLc1MMF6YZpkAfmd/h3GBIRDxxYNJkW4aXdBN9HGSuLYuknDek0tgJGcgYi2/bqOz39cEUfN2
6UGTF1tJAoiMWk3E3sQk1ylcntPDfJeDQPjlclyCZVviYFwoU/Of058cCGFe6xuY8LNhdBSZDKEX
C54u1VKZ6xW6L08orvmOV9otzcvhFN/+jSCJrkoldKOrcgAKrdAUKSNmd/ohJ8xNYf/9xYyy4zgM
j1b2WYihRDgAY2lDwGpcXudXBs856m6NnuNwch5Os2iElGpKthbNNm71R7PkttLgYxoGfkcVC4DK
3i/BtCs8HJHDLCfgiXb9Um0T0kiIC4gX7eG3Get2Y0oXQpVx8HkQlx3YCSUMXz/9kJwVZkT11n7k
CJA2wYaCyNOSJ9bKDRTT/eghGZSAoCw3bUvxdr4cRQ68efKu0CKVoEVvaei7NWaHp6Zd28kYpDqw
FvZsVYcXZFUyMkcoSBZnsbk27mTn8hlwflPxb5vR7/Fd7a0zd/45I9kMpvDm7e2MkeOvlApB00K5
XMW6lEnmvP5nNmjvzZ4++gJc2w5GuoCcmlVFeFkQK3OistqcuDRdwPHNOYa3o8pF1w8Rugyk/kJN
4B74Nd08TN9feu2gEM7DDKaxEiujL7DK/DFGoDBsYInPWp/pLZ+tcG1RtY6BlGtvzs0glVWmEtwJ
AE540pESEhoJYqHX9YlsJ3PTupHOp2PX5W2yBYCPE2IE6E2zEmrhJa50JF4xfI4v8mWwFSYpNmEe
xymWr7Ou7jOGU9fVeNLkgyxxBkq3G1eY3patCIDB+bcizRT1uBvqGGm1SYGGT6Que4TxOC8ZvhA+
hOqn8W+T6a8PtY7wiKrQjt7duCbUCT2TLhkTAOIpm5ApDAfuqUQ0hq6wSaSGsXY9OAxnjxc70L8J
HIGvZajsRLzTfHZwDry3o4a/xPOaQQTNoYPeJCfmC60HGsbzOn8puLcvBuaVNWhvlKjTU6HrEJms
A1e+w5cFVtgx1Q7hDObg7/cyX85oJ0DobZcfOLJotggbwUhXOwjlBpqSSG0/4KVCcQmPZmwDoUAy
W+7/fURJxNm1DrV8duXD06vQ2ZDRs3jzG1PsAeaAHekd1AIDOlMvaqsK22xCxNqGAeweJ/8XgRoO
1LMHzYEUFXXNpwVb0KlXuBuCzT+6ExNqPQSatn8mBldML4hlk4Tmb72lI39vzRndZQ7PYDF4PFnn
KZyBaCSaD/sbDcVtbZTEhwDe4w6eguuObKunEUSRS+3muvK8GVNjevd0lqij9fRtmXhhVbTo6bLH
+T19CCbuWHjgqjmvPCFu/6jg0MWTLS+31XbPmtITlxLqufNmByp9q3uSUHRiq2sB2h+u52rlJE7q
MacDQpxD12ZYQiAnHCFKxM/8Qo0kwfhdC8vZc3wLdA87+7rPWt0BYR7D04GZd60bckCIBe+au/k8
SZNkj2KPNlvThld4IppXTg4v5nN/Pe6y1XeLP5YuZ6/uNcSO101Ew44gtu+HsLM8EudAvSebHI3H
ZSB46PgLB5+z0UCIrzRRkLft7AXZ8t//tlmKG8KAQYNXtlIDJCFpZIOay3g3hSN0u8Y0q7CuaQMu
kCyLELY/JH2Be03piTYlj3CXy//bBSqDfciWvo061wygC9kChtXpO/Q6ubMJ5HXImkeoDReF379U
sICRgkO8qmJhkbXrAaqZdUTuk/aUwxB1Ox2fvFdYOHzo00myQdaa+cOLit4n1ftciuTPWrx0cbJk
CsBQqpKhkqTrbfbCLjKjKYfReaBsJpv6yJ5eFFV3f/YjhRdOcH2FMpOeq9VF23x+qd/HqU11CYTn
0eVFbdV9tXPA7FaV0xkFYkzDmbRFOyCnmJTyzGQ+Q4+RPVD21hecQVIPWgXPdeOdXpsmNjzxwSvm
XF8KfTS95FITmPHmeyEE5piea9jeS0m4dPWu+ZzesWsrlh/qvadUAXAZYQCyGoCo0Eou/Ua0iVCB
rY7By3zhsHUVnesSfJboigkXU2mYj+nC8Dbdkp0FxieZoyhhbbmiXhicElWvvxaW/U4hEU3ZdD5J
3lgO30NRhrJe5Wp6pUiU56V3Jado6leEXWk499LhuIQ15vJ0xfx8dqwsTR9BWIJmUeD9Zr7t1LH1
AqM6SRqUADvthRyVPfwJrlRck9AnMdmhnzljZfYlUa7qY4/Mf65hO54vl028zX9UY+/7DOoWVwEp
JEfgztpUk55mK1E1bRwoHYr7haMYnmXMoqqVr6CybRlXvvqW2/5oAyMnYrOaGOgmOSsqcKCJ4bXh
4tRPRy1wFgRqN3qYD0x38kfcgLQaahPgaidIMv3ZQfB+9XYHYivndFvFf94JiIfUXM3XQPQ3tHWT
G/arN7rfFjYMHCgWW52ZV1k4/NbF7r2imZvEGH8D/5pZVp8DHwTd//Wv/OcDQSi06n7EU0oqg2bR
+FHLEE056SvTejTejL7fpthJZA2mJvVLMuB2h5Qti3C9kNuB73vPcEFbKV4oxQt0J0WM8MQmXOkA
r15XRpqCU3DdDofPax7LDLyBFG/GGabQJuvHDgcPFzuyNMvbgSYoFEK+OKIxS7nGdn2701rMC4b1
CySIfX8WSthdidH5ij9JcwRO7Dote3p4/1vVyIJEedu5Qs6VWqv5uXf7W4YX3MmyV9DncZCPzfYK
buU33o/rVipGS4RzwxNbvWlUHm7sdaMxcm3hCftEudlNXR0JbnAy6XIY6TZXVd3HeQXP4SkRULbo
BfzGAhPwIID11xiyO+KcEPGxuFMYEF9g9HHkcyA0mRBhxE/LIXeRwFjyCcsLdbIL9NPFcVDwVvUk
p7Qvr7JXTdbK927fpW5J6+OFe0BUM/n7rVfGRhbsCQa7OFhfAqPSd7Th9hmdBbUK/aV7XykT297G
ILNBoGyf2n1QfLEWI8g3H+ip21yfz2YExXojyg0nWsrPKg0l36luptevbZvIWkxA9tPRaaAnkLan
ysJuWkDxTNiUftLV1OsL/SHT0yATgabGvZx5udDWAGn2VuCe5XYc7pqcZ6TLCr0RGm/2ffcdS194
sj6Xx9pRO9PAxiE1R9fkEvMNFDpVqOD6ciZVlkEbfC9rva+2iMbRgf+/2pa8KCQur7bE+F0gL66J
A+Rgx9UbC6U30i9Hmut25vLmnt/8eRz0awN/DeUICcT8MB2aOiN06A1ai428Am/DoYKArUAMt6Sg
B0XmDmHOMqds3j8zJzIPIrehKnR1gLizik38BPFHtzHaitMRa7XmSW1V+Wow5AoLq4iO4XegHcGL
0Kmp4UXJcpJPMCkf8eBLhM4KoHrmmwTUR3vloNOHq4PO3KWa+ACdjItnwjzB5sjpfGYsloGiIVNw
Uln98vmWfZUMx/vEoW6QXI7VgAyW7rNYWPmPFHFEOSM+6qmz3W43ENYcqDs9hsmQPX472gwDaJap
d19+M8P31r1VEixeASpxbX4uNoYAXNJpAFEJdqyq4qFme1zKZ/O00f7GUMAeqxVVhxECh71PFu9q
BIC7hagBnubGnL9FQySj6u2mOqYaNcSP0ltiCEMSRRLxZXR/WvfRXdEvoNMKew+Z+3PCdUAKEBTz
Oa+686LWUfUPub76MQhpQoTJEa7Sb1KfMBMgKMtvoiDaNt7I7wjhu/uVlrfEqw1ye5sVPbhM8qCZ
cgEN5SbiHYuKhebJ2Ax95robWjuUL9mVyCnBhan+sibWyqeNkIBN8KZk8r2UUUWsuwx3yBt99vLI
/dm/A2oYeddK1MOowAxWmSSlTT7TxDWvSMgoxzy0oG1rrTaT/ESuw+wNyp0aijCCgyxZWMnsFr1x
qo05RHNolHVjdPjIHsdXu0qJ+exoUP/B/Jha8HQXhc8vq+naXez4cuKtgeVYpey8pKsepJvCLz/H
EEUo2nxO9n+N6yC8LrhkZS0iW8RkSxHIhGLfUFqv11qZ1u4cwS3y21C8sM4ktOCYQW47k1YDVsFJ
iAsRC/d5iQyxj2hd+eOyzO86N0ygBxFPzhHHAwicKg8hyouwsqluNDGKVzz9jwNYZjP2M/ZxEsv+
mY/256EaZllIyaF72p4FBSsMdIe3qu043qKa0ipRXHhF6zeV3xWVapHZB9+awtlYx3ESLgEY4Zrs
cq8IYDYBrOBow8iNQ7AviwQMFefKbeXczIoD+Jqu2Fh7PEKVU28bDSrtGigPBDeIstqHKyk+BCxT
Csjka74du+8Q1TluP07HwqDcJcfgq+vG8NcVunfemIFAd5FiIp7qWBwhgXWfGqwrqr8Po6AIGUPg
aZ52cz1NWnr+7tfuH7u02IcBvBsnXJhtXwN54fHVlnAHO4F0BsWu6aPM5DWLVUwT4Fz9F46VSLuc
H3QMbmtlQgEf9kIg56AAMbe/m8M9uFYpW6DWRJmlsnI0kE+kHTfIk9UvKU4WH3xmoVrugiwgG/wD
AW1jFisZSQ2qNOqRkXtLC0ezB1bBqIuYE88HVoEOABB1wyexQvW1NH+NWp3xJvAGUo2yIJhOG7Gz
Nx+pRX4liI7mevpFr6d+nehr2+2Smmu9z0PwKntCjAibwlriQQ9EpRytHvj1e2PQgsIDzqQfcv7z
j4KHztL/zcBNR8c/5/CeKdMganbIoFgmxCeWIKa9IzOcOApjqIj5+AqIY4lRPL4I4lRc2QkJ1OWY
ffN443m+olF6YAiBa2FhAreSl1JxUtQMWYv8PBHVCTsrD2pv5fb++sTm/X30dzr71uSmqTufXgvk
W55dk65wxyRZ1QOWpwHY6iqFwqZPidRJDHqYcxRMNdDpweZeY1PaC8iKedNu4Lbh53wEE9YODWRG
UMjUHqFDa6eiJPwiHyPXwUdXCGJHLu9I30LuIbVh52OdMJDhpd8x4mZb852sherp48kCBF014wj7
bI8NAHrwoYZMA85jWSjUg60IvTa8Z32NcJudKdaiKReUHjTML/NCDDE52zykchRRQ3Cqsm0lVpmO
60XT+q29OK1OAMVRQESJpm+FtHPNDHPiGUH42wlCaT8V/h8ue1UVpe5CQj5nqHgmB91y2maS4l1+
JTlFpdgFK+Slje1xlnPBu5nT+7E4WJmberKRUAUxRt4WwZ7lJNE97CVuLs5BWTHdJCuGAto0rCSt
YHoZQ+WrvZK9YogpE+OhIePt5cPXZjBe6odU6Hv8Qczh8TjA1N7OqVqCHxJNiF5/s31o9HKsYptK
xNGJfJEnSvuh7xuo7oPkqlSaGOuWAMBb0lFY8S17pw9tmtZ4RKw+kuztG/GUilJZDlxX0ZL3lSj1
s2tbhyqhcbe4xD/DqCrrwFjPF+I0tcCJnhmufIbim2LfmIhtyIGE95J0oCi36YEV8gCPIVnDBE85
qF4OqscbrrhqCBr1G1PJhZBhSRmNIbEhKyQvk8xl8biAGSYzDKnG4vZtINqhK2qeBj40N0ZQuHLe
3j3tEtqiD/P8AlFoRHq1buKxHodSWKJFdS3L9TGRsxakwaBWl1PZE/UKdLL7jCM03cZSV4XPT6mV
0hlJSh/gYi+dNFfNFTArXR2oxFGpTEI/WQa0cYqGFsAe/6VGeg5tU3raLzBdp6/X15tI2v1GrOEH
AAQJPoZ2WR8y6kQMeqTRFogv+Z/d80u+0lvvw3uVl0ogWNxZ8DypY9whs2s5dG4snGK0s+u17a5S
ii3xbb9IhGFE8tLhl3RV/OYhAMJYGGxtWup1IfJRaTVV+CKSep0w9484yDI4CxaD3ofl65MNtGlJ
lj0jbQR8igfs0KSHS7wuLTfwqC6jJmb4d4ZpAvA3xkh7stLNGmyZXvcs4X2aT3+eYEoA2kr1BqIu
JsLq6OSpxVdGjQ1hGMSlYNi+yA1ELbs+Sd3BtZkcjc7PC/QG39ZRjcWYrx+piyHElJp4pVtLVaN0
y2eZdOWmax8gpHrxIvdpag5atBuDQ2tICYn813Excic2SvBEH3OmE4fLlaqv5PKHbdZo6AjkeDLA
IgLHBxH+O3/QA1h8z2sITLW1WDe/FjlrUL0DsSkPZA3Be7hPlkWGUvqPWj4WR2cMVClsF/9g2VT3
ch8ZxaIiGt5SHSUqC45NFqK2cJBLtH+cgpctd4rQ8sn46UCxWWF8v+2+gpuEv6y4FS54tLEp2u3f
dKvBb8hM3eMSvUkKm8NNIIVXz2zGIitTFyMO2e3Dp+QTezfhhm/XE0YuPEMwb9AcnhLFWO2vZEaN
EKsR7tdh50Cnl5dvuRFf7js0Ck0FQTRhTnOJ/fJhIk9YrDuvyCbZzkeoBxGK4Zx9jgsI3kgmnkp6
UVULN7M5+euHNDPJAQEnmGNbLTde0PxonePuNTlE11pr56JRKo+x3VcVxMqB311Bo6JAIVdtJzoN
ynJqKF4328WN+kzO3FeIIYP3o6mYex+Gc3mhuf1XMkdD1grlVB4alb811RYLpMecF52X2yndiieE
IF2JsZALu1HuxlFfc1R9ffJOmHRB3zhQcm2uHKI1c3woBkbNcde+/4BlJ46IS+vBkb0gbrO8TDub
FUQS7WZZGrvKe0LxC4Q5/VpEWFkcG/a0crcSEFu3bUP1vs6TsSk64og44uuc2zdFxb+WPGD7a5Of
Iij3khwG+2Bj7MyMYzfmV3R/Wzm6TNOVOUDscxetoTGIoyKpXaGEOtBpB8CeksMe1Jg5PQyGmT+w
HoHa1KBgg0PmRXNg8E+8AtGNSrpEh7FjwG9duvfbTloyby9V+biiI4nKbBJjcjE9J3FRkm66MepU
xEYCQPxHYzbFwhKEOUBpox/6c20edKb2ndEe+AJfUdcKG0Uj59Lj5IwSFdmPe5+wH3eGFv+hPlcu
b8pnBQQAspr+d/4wv+/N/kbiyyROiiwl8CrgENzDkr9c97XSQa2PoWtWnWEQNApdzjPFjlE36dvz
iSlB42DkSsrrAj0v0E4hZQYOH8NA2TDAZa3KvHKeoOGnJU7t1AZayZdLFdWXWXGbJ6UL5MGGMNOr
fM+PNS3iak0S+5rz2CJdg7WgnTKbFV/7mj8oVgSodWr/Kv42hTbtX7Qyt+82mygzFATSvN+eN1zD
CIrpyeGQP6VFo3OQw/Z5rQXlrKM8QF5S1BEyQ7ZBxJJUXalgNhAhQVEhOPpSimiCk+v3Ny7VvXDJ
JAMioH7wXe1HNaICWPE+ZXWV5NgkPCcq0xg+HSCjIWlG4QnwDaA3arGxPipv1h4WmPEyC9Fo1YnH
jj8CynO1q7IDzdguC0JhlYab0e6Ciy4CuWL5Q1EvnNW9ZSgEyjWVafWUjnPp0A0O8SCh02ijkjAo
X6Afr8Dr3AryR+2OlIFVmzNTByx4n0CKBlU0utaaKGLUbFKHkfKSdhRXWlOHi+6DtCqWVNW9wpgR
nLs5jLyUFEf5Cljb+NRZZI+U+d+6PEsqDfgedxJZEwp8Ug+gIEcD5L4y32mynFj+xMbMgpUP65i1
c4mt5MqhcTs4fVE23F7d8RuKq1wRWBXWFr2t/+Hnti8EgZWaqww71PBtrw1q1OKorIhZ8iai39gH
tFmurmyil/AMYXHDIIXOH0wp837arivZWSIghGY7SHZUlfJbX/r20s6kaYwFmFsiC9CUBJvHnY7U
Zi3+GEJrIB2oAp+g8GM2+QZx56AVWlMw4POg44v+bziglI7cq3ZaB1yYiASIuL8RHk1dj7Qi0bNu
UdLFppjCkV7pPGkSjkvhleVht4msmXKf62mrC6a1Cbt58882Fg37a8aDe1+9G6CFAinND66QXSKq
Xm95A5hfQSO94uJkxMiBmcRtiiWKWb48LYDckwNFndmOwrtGqAQT2Rs39XMibTVedk/nIUnpQCIs
uUXzLgY5goOfGlTdxDH7uxymJXLWhFSuj3wMYNZmxO5qwcsfc1qQf+Ai0eMLzpg+d4dW7fem5R31
D4Rzyczs2EmTiuQsTsUfRHK5xRc6SFaPZmS1Qx8NNkd87x5yGpZYtpPw39y/ogu8EJKfVcP8b2CZ
uZ5qfAujvA86rE1g0zaba2ERKFK0BfVcZcE0xJAZ5CRCyHMqc4AFhw8V8IKCbgY8Ghz+BkG/5jZS
/Wk9E5IR/lI1DPBtSquuenZKMPUmnW2nVLHeOQ47hPHpGaH+h+LriKCLXFXPqzG2zavsvfCDJ0J+
oGj8/39Kc3G6cd0XQlwoA9s7oJRKFGVCdJ/ZP/Oioc74ttwrrZt778vFEQqK+QRb0M4IumBWngSS
p6/O0q2ZmF66cR6loL6KI5lxbSOPiOQavvAfkRZdxn/Bn6iXXTYDk/h1JYJdHN4djofV4ct9bg8R
l/luAsLOpNAgmFD6bR8TVghRbEboC8X2DMfN+oKtx9hCLLN3A095+d0gjA+NqC22zBIbfm9dZMct
mcar2kO+vrBRaSzcJLYroS6mKGiVZyIKGvSXVOYINkAbXNfQWvvGnGTzyc11fy1OsQCLWCdn3Neo
aiCpeEk3yL5qvf4mJSTCKS4RvEmKk5TVbzQKALn+UdYDS98xHMzufGY2ImdfqANDwWH0qfeWoy2q
TVbZOuhRQXtuu4c4uY2erYDwQ4VVQ4gAeXGzSgu4ySgVXR868x15jY64crE88KkB7LR5CXVIwRDH
s2R07UOwhi0q7VupGuRBtX22XNRbJdFkbULgOc3nHwBiEtxbRHyzqe2AoeaW/0QQ6KJR/6mPT2Uj
DS4VVmo5TK8oLpgsv0ZD4gDVOiBus9ElsoValt9oEiWybGyOGK1g0Yw0Oou3Ei6abE4ez/ekC/cc
W4/eFvQzfBSzYt8MEejtQD2N83fX/QytEl1VhbrsfMjq5mGt1SckUzK5CencnCWpA5qZDgdpqhPq
l1GI+0Ke/VYqmwzTx0GsVhFdlrvef34qCMqi3+QBQPIv9DtuI/Xenp1R/tjR88Xj4A6coDzxuMwo
GBGe7oTTa4I35f5ZclFBY8MEKaYgBBWKNaqu6g0GHFXi0ucxcnhQ+/Vg0UbvRhXz74qH2RFGFEBq
7ePNKnXz3NhomVT93KnoW9yvCaq841JbdSJQP3tO8QeLH8l3UwYJr9AWKRX795smJ9ASRF9WkxUL
ddg4jxdaYuymIsxrU59e0X/OMNa9cqVioGghtiNbes5eO8rmlv/zhVya75INGe/DbIXORvYQlbuF
NH1qigkDqHtAJJC3W9Mj6BaoknenDYIqSY7QN55UU5ctEuIXa+V1+z69q+20vHExIzyHdf//zoMC
EzJC0v0vdpjsRi3ul1jZS2UfemCixTSkCCteHABUv7JfEyIkykCejN/dSh31BTvilSdZKneEoNaL
X2RWHhXEX10QLLrMNMoJL9JxDu4/pJc/y9IupoXXz7xjg5+1nEEQvuypg5n0vvOC9vS/moWQtF1n
saklaZA9tgs+fUFVYnP6Knq5ELlPnKC0UEwF3IrzVI/2eDl8HHTnotITvYSRovlH8qOl9vuCt9RO
qgmJBlLEYHcWyKDVro0Fijx3p8NhDMds9KnQeLiZBAsehXlJrCYJMCs6iFRs/dwCZqzr4rcJXtfd
EZswzpnRpOK7jM04UwZXN5sy52hgDAsKkPqqFz2A2HHNYMHFXpHvt5l/YhJM0reYMPrPOlx0qfgC
A0jHWB2ROuSJaEou9EU7yC2nYNjX8vyaw1I2dipbjIZicWU3DD4WEZWPN2CXhRcXXGvQPeSbnXz3
Upi5hvnc829iDJTiEHC6n6KFNpolgn8XuggaayGU5/LfSLmlznJdGAro4Qm6BMhrLyLkBdO5Lgea
yB20pRZKhpua7T2Xn0K67z6Fqp9wYghIiF+bD2dzEtbibLKHGDbaF1jRA4XDPYiOfmiTEHVCFGtx
hlDSZXIhHyXapERUeYdAZ4BQzPPYC0Ee9SeGaHCOoJxTIVppwYhKcayPhkY+szdKMNaNGBrHsdIu
cBoQogbRG5hOEAVYIFwV2fAD1ENEaLMj+C1hdlzV6uXb9oG5UXxMSNaWcx2tbJddUr0XYggPJWfq
PEW634QJrXNrnUIPrlK5144pZqB66V7UL1Q2d17xc9U4/ImR0l1Ec6TW0vrlAh67TycFyabOoyQY
TmQ+qIMhG+wMACwvBEOZ08UM78g5IC/J4BjUMe6fp5Oyty1FN/pe/rEXxMCRg4oEWEB/PC2QwI/Z
5FIp59MAwJ6VE8Gh4cuKzEtAYD3TZ1hANMAJbp/PWHoHrH1kQpVTL0Fi5Gx4GuiAFmsqkU2ttPZh
9n/fFxVGO1NwEEzi+h5kSP6WqjnCbj07uZZId5D/3LojkgJP6DTjxTUcHwoUhRCL0JDTXKQlCSg9
ri4Gt5v7kpXDPb2LEDDHHtsT43HQlSw3UdTDmDMUckv53fgBmme/WlMpxtGqdY2TRm3P0vNIsYf+
QwPN0d4A7Ym6c1ZWi1Z+bDwueCrSQ6iJ5nV1RBD2a8Sz6UsmZAk7JmkkFIkh+42LaeNvAMy6sz+d
0vNcoPauDQ4bHBZTLmL/trtrYvuVqXIVdMQB8l6UpvVpha59cSFytREF5v7EMphjMNXNtiiZ5sQ3
snOgB/GFntTQaVrWb4ORsNejgLh35QY4+5Gf8DC3BCc/4zqLYvsMyWcvOPlbA5qD9D+cYfCRised
rFzi7YnkseMV7+BB30waN5+07jX9OMWRES9rsPC6RNLm+A2lhByUdTiLdZ/jemviMAavktJFV71x
RW9m23aN0g1LoWtcwlvExDVkHUsAFRW8YloJhwf5YcUuWT8Pv/LQEbNCWAHWmOKDne78j8fPVdQj
P6jUehknWdyIOfyZKZXX9n56FnxXNkCZyqWcNNM8U+Szb23kXPwOwGN37dYz6A6kj5l5dCgWR9r/
V93l21snhQ54MF2/8TgQYcK0mcMkWdMqb5npOLvKINik3u4wFl0WG/A9UmcFQCMO1pkSHto8Ue9H
WCxLxmxcVn92MElWNdlbqPhTg8D9xx0MSG46xZfAWVsZZjY7aSg4NdnGStk0sihv+yzrf04WwuGY
Dxn2NMCOKsdo9clI7NR4LToOuAx6A3kDGfOkjmbdXqq4KT0GFKPJqV++OYzALnQMaQzCT1n4uhsn
ObyTFmf+bDcNV5HF23KCxl4Tpdxp10o0wgckFHl86UiT0tqE8ohbE8QmiU6LZdD/VDANuVn+VAfJ
Sm+8G1863PEZLEGp2avSQOTBFSU3HZfOyK+DOGo6UG//qUX5lp/YFv7maj39ars9BYORlU68i0K2
EeE0Nh06KKCnRyMof527qZcykDN27cr8s8yoL/ziGmacbDjusXG4/T4PVpasWTaphVQS7tjbevSu
st8+kK8nNMfx3jLFYRmqcxJTs/yXeSQ39EaSujuHW3Sg4zRYk3NXVA6FyJ7V5AVxjjK4aIMw7jBE
JJHd9WlIn7kgRX3cSZLbx/8YWum8ybvnFpsqf8znf/RvJMPuQgcqv/YUZAQkYpDhi4/rotAoEWpC
wFPisD81iYQSfAX2xaE7EPvOs2cA0gnN03iIjvWPWMfIxOdueEPwQymQVzYf5bYlIyZ5vBa1Xi0o
otao/0cjK5nSMOJd8bIVOOR+YDQHwCLWD2k7WVi0j3MHHypaaPMfu9ezM8cb+J/IJSdVVXXdgbQ1
ZtD6dn30XNFetEIO79Ml+pygqGEggNY+cbMuuC0U8N5SO8YfRMu3cTyTwK8OjD3QxZWGtrmVkb0x
523cDa+xID+jmGzxUUn7+uKfeWN6knLxqRngzotSMWPkFx2r5hK42xdU+iZS3uXVpeLP9GMKdW05
jkSt8/MWRPGXcszYjgXfCD7nKAKU4IvYWc8ScYnHlJJzUrNw3OmmNWOMTTbbEsMjQKGzpQoBXjdZ
UqtZ+GUz+9dfiitrZITHkGDFYFGKRJnIQnm5JJ+lMk9jXfiZtPHA75z3HuaMqC6+ae9ARSsYNHsi
gLAdn+0xH5ttDwd0PbgMo2AoKT4j+VBjBNycsuZ4uk5k1TGEQCVMnebHsMrpQGzESly0Grvt+WI0
jKp6bIZblZwFlmVaw12CwQXKq2O4nLQf2A4zC4Ll98cqfww5UqdWXJQJ7RjGlFobRK+G6h8xgC/6
qrIMrTxcN/oOZdIOqr9I/C9cl1q/1MMoHCwcJ/QM4LQsmQEOTeSwg9b0I2c2lETwCmeu+MQ1i4Pv
yZzrDBvUsOIFK7RJU0kLzlujfBa5oGE1q1iC5QX+BEwB7Cy3lV5zsw+4fcLOCYL083fjDQUlkFOR
oB6zBHc8PD6kDdcUD83QElwF8eRC2xKlG1Yi+AAXocLune9hkfa/V27g312p1UjgmHowHrVRLm82
3DKQUSlMvMi+EYx/VCV/GvYDhF8oRXgP0jrsjSDAnXJfb+dolIPotHdosfoqsVJ9pcbFIEZtTGj4
zUFqnZhS7mW/SFx6xYi2ALDY7F8tp4sBOGjVhVwORvsN5Chw5oM+x5p49sGdHtasUiwr6PtgF+9o
otrZ4oHq+hQjvWBxCZCYdFv8fCznYcSA98BM8IghWGdneL4hM/jKKadwEmw9Fw5/nS2VpQA3HiCs
hSyNiy3w3NRyQ4Htqi9yPlOLqCckTvd7mR7jzWMZTO/GxAvRh+8V3aXvxiEyIOgZomtJ14UokYd0
uznLFRXBaqvYa1VeaX8BxXroC0QX1aP1FxwkRpR6CRzoqx62YwgIbzBbye8JdyCurVav+DgZAcwT
V030WIMxVyIcIAR9v5XacHg6XtcGLwbJH5vLOBB99gk4GAsPk8kIbI+xt/5Mk61d+fV72k+b9Lim
ypIRW/k/y4vTkfsgSpYEv4gbS4CVT5fBOdEJlAi9xCCRbxeJxRpTJ8xVlCsN/Q7AGo1GMtCmA4P2
87kGJCqulvPRBSg48D6e/1mUdbujiOCPs6WNGPo9fMxGHlCbde3wBXVvdLKRHfJZCrviOWRwxkse
osOq0zuPoSVg0+s6J/h0ZY6ptzPBMA16g42hBIEIL3jgpzModMcQ8NSulPue6wjtAe4WMm7Llo49
BbuWy9U7hbJhWtoZ++X6topmBH5ewnBJd+AjlZ/QV5yFvHwUv0OcepbYaKwqluF5iDrog38CsT0C
XXWvahW5q769FzM+F2e2cs0eJi/pU0/cqRPVesqPMhlnmL57uJBgj4CbhxWng/W/TEpVLo5/Uk5k
f8bDIPeQ+NI9laseY4oFVXKFRSf6s49KOAgKDYh9F/zbaeMyjqNjhu6ZtImBG7GnW3BJ6bwmJsny
V61P9NUrBTWnoWO9yaBLQC+kmXbGswHm9UkvQY3ShNX/NxDcv/O+5SLwG7Hec00ShXQgxGi2f9xl
SaRXJM9JdG/vwQqv8hNtlAgZFlD+cyo9GFjr5FonPa4/Mtwcc6ZOGlAzxEYFTnonA4H9SPpbkMKP
9V/uWrdJqvyhAmL4Uc7VASFfhn5FkpQMRoXuS63PmM5kDF/Qs2VfdEQYuc+/kOQfIfU161msmIx4
4wECQn/SilMedvuZ59ROFcSF3AU72OqC39ZZQXDWB1Eab6uG3983YlWrtalVVHGdH9Nb6JsroH8D
A9RSdY7DsojuBdQVGMs4n6Mj2MG8OQEAETn2+LhPyd85heuLIXYKvJGcxFGNTySwwhYk/zTpBdbk
qQvya10zs+aVbO0jzWbyeYB+T8Afj+yWMR58i3Q13DK6cSxpaJCL7aI8CKcTf8VFJ8NMeFi1EubG
LtcwVLr1lsvCNIu3eJQUcxpuQkunQ/jXcZPvf8YGa8fQuwBsk8dr+CsPhHYDWf/2NQIqY0NS8PG4
/0WTqmMWfqb2jOoGxXXEBGXxd8+zlUxM5v6n4cNZVXgvJ5uvip8kycHRC1yxYeJs/QAL9JjWk0BL
CUXtn+wh6siyBlcFIIE9yTeN0HHJCWWPyxYGpuD+5fOAPufb9jyZpU2C2lHXZ0jRpPp8Aw+yOH9o
d2JXrHT+aLoF7FPnEJi1ZXg5sKJEmU/e++vK249k1s3ofjeRtFHVaRMSo3rE9Dy5CZmu9G0NIyh3
7XWfTQxTdal+X96UH5d9fgbWSS6shni1pXls5+4Gwn08qVSc6vqYiVv5FbdUpKY8Sx0zWzRir9Tv
+2gEnMZ+zbEPz4ydOqqp2/4HRt195BWTsoaJhtFoYRvfpinnf65gx38b1xFqErcMfdWkzwZ59gwe
D5lHLU8NJpd4NTP4rEiey8dZ+ax/qYYIaxdYGL/waLpWJV5eaVt9oHMl9SzBc/8PoIdy438xlgne
BRDaPN7W4f9nqfZgsCOqdlK8oLkNMdmBTqeefT1kiThuJHXzy0Z5YwOr45BXj1RphmzvWPgH/iq4
KFgbjOXVxONkwK/uUq3FN+6gpc9QBd7vNSXOc27Tq5xGI82hUty9ba+5HFlyWLd/Pv2MFqYVLdBY
RUSnLgLM4teGkcmgFRc1tDvgBxJdXo6lp0L82n+rk6CfIoJhY7VH9rnFmk+h77AYrQfAEvmYhGpP
UIsMhIEFzI9xPOaZ+IoDvkIPf4pHghCdXv/79Bm6A1UMrvvrl6JGDeFv0G8xTvnI1YSPkum/5rHL
qIcRMQ+l9QrTN1vOREqOslD+uHtOZEvNkvWluvE/8EzpofM5byR5HOEbGol3Yy6lApjFwXFmsOTJ
roOAe3e7nUXUWx/JNshyCYN9kIhnaAP4EzB5D8Yy0vPO99E2GDmBvRz7fxu3L5hh5PmSQHtJcXAa
/8lkbFvR1HXJtE0Ud8M2PMx2fMOhgm2UscMASouIeMQqTdl4A3Whc68zvgZfaNySLnqtjRRHxZV3
ocQwV4JCoOv8hImKWJMmm4NuY3yJbBhGclDcnPJlZZ8H2v1SyAoKHuMBS/RynqmoKh9qabCr+msb
Qv7V10D1ebG6TVpkeF2kTptCp3hGyalTy/vlCTTk41xURfMeFAAXjI3e0hWKECDuBSl84tKpx/bG
VRvxGgXgKkCVS806Rxng3HSPqsbsEysyfuhzMVBsW1r+aK0qKvR0K41PCs0MuB2jbWUMBIAPc/XZ
wQ86yDBSNwLaX2BoD+I8N7k1DVWA8SP9H/uhkKyHT1m0AWCDN+p5pDOpaHor3X1Byat55Sh7E3/M
8jiPkg5yGaHpL1xjB15S+I0HdVEQ+I3lgDTMifl2t25JH86NQoNsE5yvSETzxulFOosCN0mGduPf
bWA/tBXOgpbDecO4L3wsl54NO8d6auzprINMqOt07ckRzY9ngnmTZ3l6bEDV44L/46VIJb8PP2T1
llryotnujgQ7MneKH3wMlX0OmPelLz75rCpP1yww7ICpPc5SL3T0JE195gX8d/hXWkHKj4f1le0t
n+At0Bb916BZAxnwgWQvFHohMKKBAAx3D49aEgyw8gYrRlUwTLRksHYXIZSO9bg8+/bPJDuCaY0/
RNfw7uLGiivWgaybMFWdg8B+qpzZFP0ThyFuXoOCU4t92NXNL0PeIQ5Htz8Jo946t77Kyv4ZmEq7
3EN83YOGbVj7byXEBDofUi4Y1XIbdz5Tt4ygzpvQpggq0k864Pnn0tYsiIC/KBihuAFscvz7knpr
nntzKINI7zcRe+blvG4Gx4mwRNLAfMS6GI24RrtWXMb7BmqsrR2MDcoBUVOZSed+G2zA/3ajjxcB
aV2TM/UQjYk7JZBLPy4vXEXkrfwkwXKAVTIWf+EMhkCAy7g+KyLgoJ5c/bQjoCtXyUifGKtFQy9U
RHvkXqiKFQAh941oKIB9F4sFhLIcYfcKvFeSsnqtBpCWhhJ5TVfwq9/iwFW7n77GXCiHT+R6gACl
XNznBydhoQHnJU1dQRyedhXQU2vK3tvFZ8oojT7ORaLyLvbwvtZL7YnSvhDLcAmCkpQ7jfp6+9sE
+wQG0bBhQE/A0vNg2E+VqzrbArszz5zy0P9LBZsT0yNBc8p9l9//aLgpxZeFADME1XM1lT3ESA8a
yEN9p7mbesYKoUZkXD5Wb95KdgcFgiZuToHeXOG1oaIE6v9s7vYytdLjACls82Rr6L19BJh6CGHH
Gc3GbSZa41bkWus/fKYAYEL5GSWIpf9SrBl1MNKjDPBdmxm1vlWczLk4geKOqY+fBl9HsfBElGqq
pDZOL9vvuJcnOaIQC0Xl1wysVCN3PHQ0jjXnS6EOWDs42p6/AqB+wuN74uxMOdt/O2aVraxY6+EW
/NkEtVQ86/9XuaV+LBgKPDeh7t0rHm70tTxws7UuaXeX6YDKrqXoCNqBXRiNtxP5aHpGvinhOyFO
8VSCfYxjFZz4D9TuCVxgx641s26VlVUOtCM/c1ivL5KVqkWaYkGI3F5WXwXuNkJgFiv9VGvteaqy
W3yoWuLoWFWVPlNj9lbF4sgPiXdBYHHCF/6lcZLF2E19uQs1sqiPiBdBLfAaMgj8pXEeflAzmkSn
BMkL4BcJWjMIMbVSChFqsclmaa669msQeiHqOR3Q6dNqAGpHkh2oHLI7fglsCqlvf1orUBvccowd
rpJrhVWrhtELXdGKrc0ESDZ0Gbk/Vti3UEPq4nEixNG1u9fhNYi2ZYEyiPmkO6cgFqC1HDsbBPrx
necDFC2xaO+nZSQtgtiCEvD/P9ggbAA3oirc1fc7iu8yU/ftzUO7Q84xUa7WdmTTfE/2mIvv01As
GAsThX23wl/FfB4VkPmeLd5/ifA8YEcV5xj0DnuIRhPaw/M55khc8HHgRkrnr8igjgEfsu5+NuKP
h+HkPmXVbDs8uvg80A/iBbobzCg3NldDY0RBc5KNcM7L9wtacBoyEoDPxgTfjxZVjTxPOBAYTdcG
ROa0jAA4nlBg0eQY/9Y0AlcKyiPqxqttQ7C3n4Qv4Z6dvWf/Jui0SkJCVPvNQM8LFSDxa2xuhtuD
9Ps/5E1J+KX2i3ljuoFgjw7uDHpUuTj2boS6Ed38UCnDxqkEE/RpGCoUC4483optVOGWngJD8MNm
xyzqFGPvKTISmsLz3LfXQOiP2NM9RJ08iII8gh2Hhkwm+hK1wIjxA7n2gGDf4IlRThjDQrIqQN5C
fmdD/fbNyxdieMt+J6cXFEq76XElgQHp7VsD1F2v8pH4bGMynThrhk1EQ/EAmrEQkG94tuWEwzZt
iCiAslgwj0H2KO4SmnGSdqafUqjFHgIKlwoSXC26VzABvpe9pkSoYYufJOhz818XAYP00PqEBSbJ
TiyU7dJUcgtHsSS8cG1ZxOMWOxO8DaaE/VafKbk+HFBeyypbp/uwqdIyF8yOVn07gXk9ahnt9JjI
Bg3D3SkAwx70JPToqFA+EA60+6CXko9Vu5Lm6Q0EyxjDOIvgh6G3Ag5QM5snOOfz8sw/yDCmByfD
JnXscTHtlmC11pyX6Wfe+hdDALJc3AqQ3G/+9AkKpCQjafA2v8dBXV9lnXfJuTCSXMbhiyK/ziGo
KooMRuPql9vFcvZX+PImtK24NeBrzzHonchl3D2WJiQgaSpjIbjvyRKtjYD2TvxziOPAwuwW4SMq
EcICedIEiHn4xWx9TJBI0EaWQ9s7jIYO78/uI8SZRM0ondJojIFPTaGY4A7Jl+By7+RSpJyPq/cW
93mzOHCOUjTodYLtPnkNjpYpTNDqJeon/HppGGbPA5inVh0xZoyi0lXdmAjovdFGnvwE1Ykw9tcq
o/bQQ3zi3k0w0NV4DLqs0PwcK1H4018x1qrAvEBIP1czVRDQZRILzCF96BvgRPlUxBTx4LlqX3Ec
hVZJFQkvkW8gL4xNepcsiMO0I2Gek+aa9vp/9x6HfuZkcH1bsys80roqSoy9gHSN4zSB7SeuPXi7
PmcGDfC/8851DvflCUn7ilN/3SlSPKw2ROjoIFrfCNGtLed8H34Oa86HWrWM1IdRTUV6pCNncllc
BhEgnpYJVSMdqHIVb1melG3eyjzk5C0BjxUAZjWAfhTjn6eDdy5blFQ1CgmZ00cMEHmYnzvFr5C9
CZzszKWuEMTifrT364ODhDNhe5TuRjBwyiGImLPRFN7R4tnijdGkf69JFpkatytA4t0P85qaHdcy
kVdDD8iDJB/xPD+ex6JbfVh50ecEfVqhS+X3jkNX/uJJC6xJBL/slxjUx5nX/LvVy5cXleksJqHn
EgCDQGmuSx2k3KVgje+30+SWYSwhYexXFIwFiltKWkjRBZf0JBOolynoV4irvp8a7PdP1BW2iB1v
28StHalBpJjqsYkq27Zzz857+Ga0BY+cOQDEoW95M2y3cZpx5r6wM3nu3km5YPvRoQ4dL4xmL3sj
yM3PfGzAZH7sdpEbDS+oLa4oy3o9ajsMvPPB/UZ2yEtlAywDFSj1JuIm7duDVG38ZmdUatCeTIKB
j2Mowgy7qOvaif84Nwv4m3AlXJAfXoDecwCRrKVHpUsAU87moZ9fU8AOWQye30e3g4rGgcnYEe1L
y4S/KZ+0pnJALhulJdUfoKmvVrVWC+lCn3qsHq1xJDL18dPfTfcntlHUg4NBbI0lY+JdhG261B8X
nPq3nG2jGzE/1XmfrRXAZPGEw3Vnf3w30dZfwWhM5rQu6OozJAs458RHRcNsKkuoWITChIQ01FCE
Q2HZLEpSip9cmBLXGwELzOUI/fkwpdGGWc/yaqgB8sygRdfV0HvkSpCJfJAFG6+jY+ZSUFDkDYMj
IWrIjURa8sm2zcskw42iBMeLhzc8s4UaHneV6KcScQEKwF9ALS6w+zC86/S/yCT0FHuVXl+8HUpt
05ZnVD5eJKsaUi76g8rCQNlEMVhiLaloGs00JTHjvhreFvV/kuASirDXKr87SKRLo4GTJLnl/qIR
JSWPa+f/OdKwQuQtkGdGVLGnOSGcXPOoAuscNEQklfSOery8DmPSgbZThlvxss+vCF6rUw3rpSXR
jxYsC/eSajUS76tjjVQX3HUT2HKGK+THXPvBWubqtrnKds2YrVNBwIJ9ZNStIhBtIbCU7ySZgCzz
QtAiTMA6gaNkysuBNTSiiinRO2iEBOYqaS/EVBwdV2wm0k7MQFxIN+CWhx51u7rhURz+pHQCz7sG
dSPNrhHDln/W/jDyCJPg0aPHKCTH8yVJrz8dpcKgYgBWx1FOGquDrJjAr8RNbKub7HwLfFuGevJR
UubaWy2NHhexg+Q33zPzruiqqrda99Z8n3r/GotRgKmW+Z/w6yg1x+YqDiQxbQDCouWEPPZRMBLw
bJ4HuH/uF9HlSRUksA/Wp0ntKnVKOKcSK7Z6put9wjkVsPG9rOWacCBN8oHJjRMnQrpRP+mrmuYA
m/ErUkEK5xTSWfT2d/o19uRqMp3hwhkMJxBhXeIm/6ETvbKCMsaXZLccu0oKflj0UJFgTFoL8w2K
8x4GjS9YW2VPJlwDVm4iY3g+ivO7ehi5TevSQZMN//Vh/KruAdRm+/HmhJW5Isl7SuKiIWoe5VcR
wn0LgnYx5aP0lPKQt0LiD++uvcenKAsluCpLi5CkxgG9ecPpprbhzSVlTVJbrbijUZN0lNxqy122
tRPdIVndkbKcd0NxUQ4Kj+QrzRzbVs+oX2Et3GhQRwWYATpLsdw21RpEhoDM0ruXE4ovT5F5zqvy
sCVmFvU7PLJJvRmLKihI1E7yubAWxzJhHi0mIdJkbE/gbS/bhOcpPPfXoFibT5BLCqxmLjLCHP+d
sw/GamO9GbqYsTXivTza4/dHnN8C7XUd4hg69y4XqH3HNK/yupX8ljDQfDvi5Z+B9hrPqfKNlLad
s/d4OsShy4EHBZrXD8JSs6t+dhCaLUNNwwh6+cxyt1POR37naE4fEkchJepXp7RzqO7RG0JuJFEG
iRT8FP8upuesc/dCG+PEYuhJPEZMFSGJSKcwFpxriwCr36YxsVe0z9323RlMLO4Dlk6ISckOH6QJ
glX67wPOdPUrRhDYcCmempGWZrx3wrvnQRRo4C3LmladQMM+Ur89g92yoIUnRLKz47P55AScZlyc
+V0Y6TrliwGSOy1oqSUpD8IZ49aOsGf3gRfgLqXk35Vm+0SQmzkrrVclL84F6jKC75CGaw1BcqO+
ExoGClzPJ5/AQJRtt2N1rC71P3q85xASQF6hbea/BJh/OiBwmBm3hrxxDWVtQWWJgO1PsE9iXQpE
o3lpGr3MWlgUsuDFoT883WwFtKKm+4ens3Ftc7D3fND1Q9jhH6jEhKEIgAyeZvAfhirxxHkMLP1z
91OhCtuT0hRXDG7R8MLGj+5CW//XQia02ORjCXtSkJfB3dBsdSGdgmzZtHYtqjbdOUOTIczsuuqd
VjiLhLUvhbczEyt/D1+Q9Om5WZQK2y6s6wzAmPAc/jenXxhD3T86Gw9PI3mzRV9UKrAtMsGwouo8
JvPT1/cUIzwhmAUuUlxdS4HY/kmTpHtSGQG1RITIkQJsu9QR2IOVdwfhjkqZs3vNMiMqL6l1W1hD
N3u3udHO7bexxwOJuXzjJbD9wPNHPmlw/pxXLwUVApKSomPMidlELymyAvilCf0NSaXT9ljlS0pM
vAk2xtoQQ7Q9yjP+VqKIjKtvXqT3+FmycQVx5y62Yz0F9X72DIYVJgwzjuUvGl4dQnHDVRDbNNE4
UgjmyAlzUsnxbGT99ckAeU/eyGrA5J3oTLm2QYeTKNjGryOTx4hVY8/xIxlCSXh8L791tC+lQAO1
y23HAa2hFnn+syqvXyA2hFIxB7vWaMoiEMdjw/TcJ/3unQ1KRuMI0ADAlWgrTUe4Td6RtdG5YA3P
D4f5mkTipx1nswXvJml8a53GijRB+ZC61UpSIFc5uV1cRJkQ//65zgzRkYYVT1sdnDx5BdNAPTdL
/oNDOFSvDrbYPQ9rMTOmDVAHs5Gr8/Yh/2ugOdcWCiGgsUSG/JCWCbGawbdGVl4B6hbTvXapgMAc
x1zXWsKfA6dKX3Yude2OKLNhqhRLOADHGNXraHnuNB2XwevQujgCxGjY/M9GwSuGwI/mS5wN/ENB
FvWgTOe9+povGZEEuYe/Ag97QlXnvtXorcSAYtchgjPgKl66FH+8mHF4LzsAw34A8VUURqcmsnZc
2PzHR3JFpvIAcSr3xtDYKTO2Wpx7pmu/vyUS23QGP9xBjqx5zWX88Sx+3rlvo1FObHgCC/hpNwZe
Dpk1/Q+hbj4baOm+qqc+KUoiBaT2pOMyVAf1/CFeMPnZq2anClYqEbNlPtgR6OEW+9msUEvJkTKz
ESsRVlDe+8Vcvrr9hkjasbCca98L5CJE5MhM3awJlNVxuNBsRdIhNwrj6xfIS525gIcMeKH3jY30
+7JNBQB7dmoIZ3/ssfQHCqcErSdDNhV5S7UflFZOxCs/U02NpaljOmugYCtrQqHX4e3IWyjsqgrI
+wo4qPZn2m6HhLDr7lxh/Wn7NaJQDlZPXdZJU4SSwTTGJgICZ1z1Z9c+fhv8XOZAaf46W47zn5aa
r+tg4eLH5pKEGX+ixzBwILntzDfawVS9vWGCl4wYxWvs9kG6B+2ZJrjbKdFXF2GCG2Oo+Fz2MZyL
ETurLM4MDQerITnaxcmjMcV07RRw580CO0UhRmtA+rel5EfXXYmrC1CnQS4JYQb0aqNBdPvByBR9
GWID401PM8Lcfo7/N/6TH9mkaMnbFOECQbkMk2oV0RCcZE5hoU+VX8te/ZxK7Zwk4TufLe6odSNm
D4kOXRgULVqBdxrg/2XIrExogu39HH92o42cOkOQtHD6WLxsWza9lk7iVjpurDnRS1HxCEcpZBW2
2bw+CoSzG4LpS5Xem04F/jG2JZUmdDmk0m5HoZVS901Qd9omcEBnmDJVAlpd8UmAlIp0YCGvBQik
SAQnN5+HQhjAYxrdH3p3+y1oAiLItnKM/t9ajZrjPSV5LxcKW9ZLAeq7QvijMM3dXfPwqKLXUJ4/
RMJjvgxNh00NFNpF78igu6rroO1GLF5Lubdf1Q4GmeReajB5o1wSGadmJOt2C2bulz7noYiR89Pe
44d1jgNKuPJg6pKzbp2FTueh2IHDskIoAZvZXpEPdXlBNNJ+g45H1AyjhEMtFZLJEdiJC3xU22ZL
+MO8QmC4ylS0uKMW2xNulEwGbCYFOSuewVE55hsPhebPVBZK2YdHRVMxMgRJl/YQdQFJTbQVN+pH
RqlxXde7O9qAq2kMyNJi6K3LA8j0J6zP7DZiFkSkzb3KoHooOsv+7zHhKlp0mlu4wVC4RAXtgkYY
QRA26NZpjIpaYyyHWmFBxTVsmMEwK0ryI8aJBawdYKS4wsHnfwgRJm+8AaHtl+4J8RS4gpsGbtkw
FKbc2EmWEsaCRoe3gjX4Dg7VPcGFDVSMaBTpdB6tnEkmKt51T6Lr671KHTceLfXh2ghwAV3lymBn
C5UARr+83CIHy6XnjJxFQUbJxT6sWjKuVTxwOawnxAVdXBPEr4ANpBBJLMoouR/97GDTa808juv2
4PMVWmvGqpsDIJudULrgZ7e2DLtRKuZnVGlGe0U7z0jcGbjeBL8Q6eU/ryJXJ4sl6qe3hxPlfGHB
a+B2hJdLte1J2Yuqyeez9wNZSRtqdqJSBWz0DVDFsvMazb2tSs/X1DQgXlhlJh4K6orG9NOe6cHj
XS9oNHYyltlNSj384fOtoa1UMSmV/xmldu3+VCHGkqtn0hqhGi2xAuTrP2kcNXLXS1k1UKUmoNab
+57b94SKURzGHTSJkd87hMzGoEl5Y1PqtEA0NXYLxgajeeSHXNLRrjZFzYVYSRVRQurbFpnxYq/E
ypMIpZ31kZ1poEcNbmn9ZOvhxcHU9rvtAFUhb7TSeCXrH9zP+ErYWoFQu6CXv4NesuWI1cLILJAO
f7KshlFT4lNgol3aZ887rPCkvj24rwoO84ipJRHn7scvdU/Kit02OEQPkHu1cYm6hiYP9cE09znD
yLFVkHg5Pp4CDN1XZnT5ZkHezGwBi2f4is3MBJuhGP34mUd4V+jPXtW3ws0uf1FLCOdJW2CZwOx3
+dHNJG/C51pwslOdLXVatTOO/vYDqnGAN4sKIgyeqTJbJmJgppD5mQEJGQrXleG+gJ01C3sUBu//
96PDTT3pL9vSRkhZRh9nCxH0lJRK3SQ44GsieNzQTc1ahk6FC0zN+wnu5ZsX7fxwNg6N6aPNrZF1
KK+fuC9aSowQssnAdGNBr6VE0Bzs9eBbuSUH9ByODiwztHms/P6BKqCmgkfKw7uTrWJkL8Ed/e0a
2bI1P+hDqzfI+ZZUvKkuTfPyBUBVTEPs+oXxj2eDBYdqKeYkEqqyBK4RxscZsnTsTmNES7hsdGc/
N5vImZ83UxKQx74QCtspapMsmetCZrbc6AHhn+PYerpnQ3+7eJiYt2rz03mV/iYeX8uUUkZ+o83g
nvROjETZO7g0B1BUyp8Rl+5Ly3ur8LsOLktTt2fOF5v5RqDI+Tr+gcemimXgkTKk3C52QqomCPxh
JaHnACUNhJ9BOSuwDZRN3IiHcAO+Fdvc0C9uZiAE+ndShr0XM4VwZUowZYgERNxM6JyaH6CD4rmb
NvH0v9aNH1v2KXZrpG3r3BBHpry01f4Iz3wBMMwm6I+2frNtCbMpvIobZQJHqv5qNZifhStGZpj4
Gc198N0DlJ7ciN+XRkZvThji+0S0ynWBGqLk8hR0JbMWIS+Z2eur+cdCwbOSlNUBjpBoe2/KQr3s
SEdgLSSWFjBzxZF+/X0Mli7CDw4rnjmDo7YcG5itzEpn4C3lBQIpm/1AlFvBOHvUDB2Tp22U5CEg
VcCu/8hL88kBFLIRk4setjo0chQYE3c/R7C/LzzPTYZWvpAbTw0/xO0jhI8b0kMkgsu8bkYLn20c
uDaIuOrsCrmphL+aKmy0J7a/Wv4dvoknil/Gy7UAbe3CrJkbVACE4THsdaKTwWHJzGytUyq/pK+b
Qa+VIJU9ZnNuuJkOOfeT16jmhf6pGdlYvPT9q9GT5K+KwQFheLqXbvyy1d1j33dmmQkaRd0Z7jkU
YDX4KWT/KR+nQNeUAZ9w/OKP0i8yESlMSYX9UVVlVn577pWMc6geB7q4QcH2tDhcw40FQ6D8Ert3
+v7BLg0QJcLZLD62tQRh+lvcvx8FJPmufMmcXdQLRJIoagZoFKtSA+nVFbm8606tMp+wWro2cgwT
DbntY26V9ABagY5HNQdFdHnMDoDs75xgsusYQ4YDuR/HAO37RZWqv978GKqYOLEB1vtL2OTnDuzs
MQfzFAkyTgJszfpSvrx9JVmxv41jTkEiwI46OC8bNFsgiSHIugW2BZgnc6Lj9SzWqKKm3KG5WMu4
+IwFt1jbJmmhLLTmhQL0htMpR0SKdg8ts0EQ/Ej21/N9p3LLIpIKTSSWEO/qPrF00wX4YBJ8eB5L
b1h/AGIITx4Fmx2hmhQWSIsNhtwnVaxqeB9VVysG/rMMGnNS+1WXeyqqrpeN1OcdQ39rwdYvBkbm
E2R2Uhe6bOzm2ekwhn3yAz03PQzxpD4lw5ZQaVJeVkf9YGxkjBZd6hIq02khQdMmDCydVh1LvBJJ
shmcNk94b3f8UG2QUzPemb5SuD7TAKcR0hwszJhF+EUl0EjbPMew3RhLgiTjiKFvGF6hbP6As19T
0kNckix2xgWk9jbEsaiPwtyCTdDIVN91K+a3PwDWRYlMra1yykAy8rVGrS/14QTGMGVkhCSSJePz
w6/HILRg8XmP8ehE3v16IQ6hSGdLubmfXpYWLBTws8vckl7ymdJQBpelyh23v1mVJdLLIKhEj0BN
iUjSVlWHhd6kymZaB7/flaf44VUDT8m5OOpDq5lo7KxaojemjFXIQPAAIQA35YclkNOYkxwBwlyT
JQiyxt8swEBoyEFqHrL1QQxs26A27dxUmRRJk9zaX3y3WHj+yAdBlF+roiaC8LK9BiYrFAaGurE4
Fx+zXKry7nzZJkTXFYTK+R9ECnGZkFS545Wocn7zSMqsfFYbk4zmsgSS9FlCmtLEaov1IEMtz6uw
J1c2OUSKcPi0SANxWGCN3PXD4zXgcOedibJmR1sw4dCtI76ugS6hwfdWN591aBbqb02qKrDMxWBO
4LSud4i1g25zDi/LORZM59+6osN1jA7YTvZUTKsq2wdWsNqhJZcsaQPyCjTOpPYV1G4KljN60Lkg
7FRLhJfHCyVf0icbFYe/yuE7K2wq2pi0ZEQbOUQETJDeQRaY9K5ptTsFBGrnbwXQjDrRaY2z6cmK
ysfSEJQTrIkO9iPhC/nMQI5I3LWXEOfiJox/iTnzZ49D8M7dproH/8FCMfF9fAX+K/YxMPNZDkCA
uj+YvCfXUVupvc0H1ZM139h+FGdGCTaLc3/ydTmJHQvr6T+au88klNQWTXTzgE1jJlRTimg4ujDN
0KsykLG64BwhmcNTbvzSDe62z8esRpUaIN7eAQFOi95oC5XMjuOgaQ/J0qNCN0vqt3fo6NWthSLZ
QbthBOqWLVsj6nxDZLBt0ln752gI8YLWdWc3l4MjKHxjVXf7K/+OqJTFJiWGhcJSQs87OigsIjU5
1gioxnilU6VEdSMuMNzss3EB0glTmlFF8oNBxoITFYWnoYktnsMndsgFejrdE+OVfCNXMGato8mM
Yf3s1SmlyPS1pp46nF9HP0VK4sBFKaVy9VIdbOS71jfeXSg8D1RfPFo9NCwc4PVspzzovhkdt8iV
UXhPpR/NP7aZn2oegs5qVqev43zjb4LRvgFppJxqUGet6yOn2KlFx0QSwL5uomcRNScOU/kOCUdU
PTEoGQ9UCqBeG0rp50+z5LB4fh8lxKyPS7gV8jvQI8Wz55aIXQb/ssBvUoclt42PKUqWaRoIeszO
eEdU7RX0Cdywxv7wwx6Qb3zkpk8KsamJr/hE7JmogbjjkHiNf0j7Z2DqOG+qAUB+BNPnDnuY46M4
ggiK6+0xfqVg97oRlvp+zmd/CviGKLzGM+e6yJnpJtrg5g/Wdo95cmAAAvg4NOv9s/wfksNSRDr1
5/XVFcEg0LVnMykFlJIiYVJJrEcfAu2LTRyNjxv6d8Z7hlxvZMQZLd/S+JIGfiVFHYgnlGytK+0B
b0N2e46TrU8f0mc67/TQ2PzPVud2zm30/WPlwzCxYvqlMZx/7cGMsIfRTlhKx1lSm/NAz38qB649
Oev3N9SCCx8wxs24QblzPPLf4VQ0snjShUya5mABIm9IYWHV1D2dioxYmKROwVqFaoQ5mbCh45tM
KJW+OhL+AphLdWgJ9eVoas+4z0HB4UgCd8dZ4c98vtib7eZ45FEw/R1niGnsvsgcEC9fAD/9PHGR
sqnQ9qfmLQPH1dcbS90d40OH9qOURZBTnrBfwDJHQqur/D4BGkQn1FPiAHcdQc3YVPcvrEqGQIK5
WJ2qmsKkqDtKM3tDCcNiFVdPOb5ZIPTDhnKYmRZQJ0jRsQR3bDQoF2zxC6H3s4hLG3pUZlsjsfvr
lABOuUadBCcvZck0iuc2VcfwaYpTy0xHbDC7G8O1YffTNNtYjjXptMRcqD+eAQfP2rPCdEh674iv
PmIAdcgyaqHep5Vu71tbTBgWpcX/E9H5mP580vhTmdy46yKWTSlp0C3blejllWzpwX4meXh6j9O8
w90HjcIinQo3r7SLS1dHqtAEMjDH90qf80Fi8NP/HHRvVshrHM3jgKo/uEzCqCypwdCc7AhNCI2u
4aq6wCY3uXvycOs++IJswhM3nIBTLAEDrFyCVF3qZbLBzRZNsf0e9JLmpN5CJgFCHYXSZsfoUgMi
Olf6Ab7IKcc2lmub9LAsZk5rb0DzL9VEKYUsi77P6Agawp1qNuEbSFaJkjPhDOXpjWWRKivs8srA
2o/QEVJDGJ8HOcR1QvAJevb4WadY8dASondia0VFNzxqig5j1ECJ1xoRTGzCYWQN29eyaNSAOcjv
vv5DC1jyd9T2uuHzcU6B2X3PlXFvKqYgKTyDH4n0RvLHbwXknqLRH+kbIkSNpYXD9BNB6ptkZ38H
RB+O4+FYDOjgjNJELzs3S7kyahDg//2sxJykZn+x2ehKjE350NY1Ucv/yj73D176yR99i1whv2La
SlZ0C7PCkcqibObFHD9jKMCjYfufB65Ae5ybsNr/KqMFr0CVL69vzPJXBfu5NyfEn5UdBuyXQEJO
N+mf9UIVqu5AMisUZsMBsF3CbFYrQOv9utY1rq/EyuhEnbQoOqfY0XhOTYcmgqG2XGzuLN/og/f2
ENl8gjxkSiN68gowZwxFBEsLqmvOjEnsLAQiNyQrqrwwgHjf3ETm9iUxbtlPROhj7JB48at5J72D
kneXrYGyZcybpwDPQDwF0LC8YZMLOLKSoNbSrTe84TFsCpfzIQYW86iZi/rbCrrsHMyh7Gd8aZSZ
ak7G988Xr3DftHdOrskAPyvk5BD7nKZ9APt486OMRE2MbTDoTlEIg2mmqt0T1jFiwqiqB2r3pDvc
DXnFiI3EXqV2h9XIZYnI4T+c8hfyW75sEaSQ0rXEqYIiBJoG6MzhKkEeXwwcLW6q0/Pf7BfWxsqS
1ZzJ5q7r9aRWZ1/Qxzd8UPt/igENIiXDNuso0d+L5Ut/IKJsN5LNi1mzOOq11Ai9zXHElsMu3T6f
30krn8wLzIJsi0SyfGNa6KEkD6SkCumWPBRUc7n5+Bs9qIbarjU1djPseOL6wurueet7oocGIyiU
r1hSQBobs32g91t9TWLVi+VMvp0bdJK6L9oUgDtuWJrq3epf5Ud95iq9yPVqT1Eqj1HWyd+n93Cr
/RkS9u4PpEn3f5Vka3/244pUJATgYKBNSQkJjpL4zFt0Xl8sxWxzXgJzmEjC9GABng+imwyEiSKr
5A1W9wUL2o43Qp7O7RX2JzhoBCTRnlNLeij5t3NPcnTNe9clSh+3m27ft9cstTm7JsNX7SGgcA9s
ynUguN5hRnJqIZ4msWLmqWXyx69SWnF4DzeXs0t7TGVRUoSKd+8VHmqxGeoBTcMQwW2BCTLGodY0
Xk0bgjzDJ8UHK32gHS1DcemQh19dHH2FS6wBurT9phvdV1ano9CAlHrlheWmDCydNrcMaDMLmdR6
yyhptXFHZNCc8xzmPnlrTSYXR/IKiy9Xy4YgSw8eoN8+1rBM3/BcjvQ3RaV9PRRRfstZQmn+C++T
RgRc3kSjYeyIAWR9Who2re2UX4FGVA8gDpmM+okc2KSFEbE4gtyCMojvQMTY20OqYfHzLYyBF2kj
eMq/o0VQ0++cmFsIv9XBbwahVh70p02EieDYjHBF9v3d3vr0RGZh5pkqkHqj7Z3AZdA1e4J0s8iL
mXwM9wsW5ndmWegUeRXjCpTiaRgDsrSZay2zp/ON0ICG2E44nL9inPG+hjwu3AOpxCMaIpYKMs1h
V6Mxdq5y+41B90IW25v6ViiZo967EfNBRTNiTdhQyPSNgpk62F7LiR9mh7GSO0CEa8LBYp6tdYDQ
kmT3GrwCE5JhVCa+5yxcfj2GuhIuUP4iviV+2IdxAS9w9OQTWJNNUN2l1IwDVGLyIKLL6/Qe1Gyh
FBqckaTbSX2pXYC3ZBPW3LoBhN5/LY4faaCQS39iNAi4EKG1CIlOVQ9JiYS7bWbi1M0Qe9w5WtEv
XEXh8dvyoQ82INk9LhojQFqj02ZY+FS5Ih90zZ3ikx1S4KMkFw1s1rMwet+mHBNaTtsvVOBRazT3
zSVt9v5DJ0Hy3CzSD8Bq70hZqs1o6tbP3DFATOxgOfjnmb1iw+xaMBbl8lu3U5E5QE0MtYOApmiK
hnkDqNQxecFNmW+4RVpcujNO6LQ1sLKS5SlVvr4hFF6HHtRJH+T88ZcjEW5/QMQnwsQxEDHVLIb+
bVi5Ak+VM4irMeMrtddpB6cXIAvGDIM+B3uG2pJ6f6cL7/abR1leZvK0ndcMsphwsF1IY2mfn9eA
mUHSmhaYy68jlHo0yMZfHWaQz/4YT8U0ikGDy3XsCacdzcIwYLyiLdhghAdE8CPbKo3nHSZo60Y7
5kxwwqevCOJBVt58PmRcoX269DQaM8AxCUUXJlg9mD6qEEU2vE6G5Kys/CQDxTxkPPtQ8Pla0XAp
9YY4lhSfDOTM3Pje1Q3jEwLalKzYQE1vVn42rIxiSfkakxs5NTIRiD7U7eJPj61kLd+xglZi//XR
7JR5jxy3nYKWsQF7nDQMyASxh6eIHMKdIbVvjzGZcYoGxB4ahxVCbgLNbpXPChnFXmJRBfsVfwhM
TqimCr3niftZPgOiSPTeBFBVo3oTn8tx7mRj+8TY6CBM7ucgS+NSI4fH4BXr0vYdmifwMOum+8Y5
w7T4ioDSWbdi1nRt1WwVXE3Qep7p4rGznYat9A2y3gtrRmYuBDw7WWI+Kg66fw5G6rpYEIzB5Mkn
hm+49TxzbfVddgBGkAIwudzsi+ClKvQEzkvtWHIDjMbMNjGXyYGknaq4ZgqEFj69x9wYJhwKTgZh
2lVR/tNt1ss5CixNdAoCFnbV+4eRzKdKfIZmOh2wxvg2ruKcYHgnR4TIL58MloGO/RNSJ9HHE6xH
9PwXMRDb5S4nrGhrqC6ishZcsNXKACHeqYkN0lnd1L5zA0tITCwFT8sAVDeKsi4zAPNKFZREX2ea
vEwFU52pB0eOGSgSvBoO/cX3dYVX51kzctq27kU+AYfzU+qlQRfgVs0KeODiTIQykC2p62lMMpeF
ufrwd7WSNy91/JtOOIdq6zjFOl0ZPGlfJZqr3b4V2JjMYI279Y4EX2WqAonWqkcQ31sBxb1bNK4P
F0JoPC8Bv3BUKxmQiW9eraVlcDzVscFQB1Z6cBWXiY7NepmDm54txXtTNdMF/PF8L7phbWWeyaDi
s7xOvEp3xlm9dQTxrSVm+l2lcmbimirxd7fRWrNH56ARYwXBJxhTGOWi6p1gVnXs66dvc4rvaUzH
aXQrQUXXLzjopQKEeIfZMzYlj9XPtp4x9K877Xy+kwvhgM/CEovGI6kXcg1EUm0ouUNt8f30dNam
5DJLDBy8qFr1KnWF0AeV+Ko9u6mQEGX4niYMTx6WfvnsPBxyQpNEtxn5hPR2UCkCK/nwOCWvceah
yk3+iCvFwVbC3TF+VpQ3nPa+m98SCj9ebD5A5kT3plc1SSJU+ztvK/+/mpbOFhaJ1AidCEeDQZ3w
eY5VCB8sc5xotaYMlrfkUHrcVU2XD6ODoE07QZF/VjrhzezVd5laH+9/cCP06hMM9ATzeWYi11aG
/IezbeKjf6X6st3eI9YTOYB2hj9jIfsLX2+y+vFL9HxPQx/fPfIY7XlO7MpPVpoiVBlzyz8lpUcB
KZGMHJoAjEkc8uW+pxApEBi2OHvZmCtZK2IuWvbV7gvdTVhPeHOinZeaN1IEQ5II+pIxi6Mkwb75
qQDWwwIb5F0Ou5Utk3riQGWA0+Fj/7UB8t+XnukK8EbZTDcTyEuckJCALjMRuUx4kKo0e5i9aKYo
xagguG40syHQpxA1nym8nfqUvk2GQ8AnMagnGJ67VkCda1MrjUNRed/J1EWbZGQvqWp7FlXnrwSW
w0mr31dwej6vK4Kb+5tMy8QMiCipewPbgEWcT4RIKKsgYwW7aKjuwI8bV5HptHW/aRfx2NL+eu53
pgnvFcnh1N8kP7CkQBbuMEgiPJMo3dPYI/jPmcqZsik1OeK5m7GR6LjUCCMW9qUhxxDSEPeljL1e
n747GSNWjesr2G7+yeCt+LxgTBs6O0PXCwbPMLU7oTRVIKAQCQpXzg4Ag9Y/UH5gqvd14nTIQSWR
vqbD5NUm7OJq9CJqDAsYXyXPaMPNBtHeD3Di2nis9fwxbkSYl3Wgx0tGZSoL07yAFJcGHI6uJ/vz
pT0q+0lvSoD2UVjs14Wvv2duu5cHXgDKRSOkq0sf1UOfnWzq4URqC20U80i8ozGApuxnCbsSrnfW
PjiMtAA7HZvBjzp47CpnguSO+3/bHzgjfp4jhsMyvDYFPQwODXhPqtH5fcrkXWoGnvZbp8dRAvUt
C86zyv8aSp+hya7m6gSrbZ69YnpUMJ/tYm9LGNhORt+Afy5cJom63SzdjuqutnrQxsOzFu3fqymd
O/w93eXwuM/hgVeFiePplEAcy4NV9Pct8TVUcG73wuaRLhUQRpwd73g6LSAkzr1nP2vrDZH8FsLm
slk3omjJAuMYYhJny6ENIVoKsMGly5m/uBBRiNnEg7Xz93ukw2hc4LT2Ckw2ZcFDx7WTPHwl43oD
Db9uVgRQLJxoEH9xIaMX3+djSDzCu71NlPrZC+0TxICtjbtUc6TSqbNG61nCYinJ3zl2BYOcwKLF
W9strSinh2FQ3MwvkvVawQHwFMAe0fWqDS6M4ruNc/cDakeZYTdJENtgaE3HMG7tTHwAODzorGl3
9Hhv2HOEy24SWKww9R6Y1YX/sO50gMeXHkgxOh0RW6fXQ2rnUi6zqyQEcTRR1qq9olzy9uhW7PyR
guRBPn5TMje8CqGJIqGxqT5pkSFm5/gM2xDhYCdufuGHer36PPivx6rtPN3fVNmfHFy5JVI+CqU8
GtixaGgiMyS95JvXkezfX5JMlH2GgLO5ltKbUF1c9cRpC+j4z2+OjahnbKb5ltUPHKE6+GCvnE6w
uBPKOpAmVKg7vuWwURKZr5JtG0jPGr1QUbhzRh6/OiUCKag+HEi2BvWl6Dx5VAxQJsIWSZIqflMq
Rgra3uezU/RV/s2ZrP1WMZ2Q5vvla5IxIisX9zE9AylT826ATq+sQNUuXNHACBDXE7H1oTAlUw1T
vyTF5e7rbEiho5JcQ9G255nmTtCWH4KfUyjCmsVW24yZEAVGD1w0IIiLfKAElrT9i+l9b0kETQRa
F0pIqLL/vaGOvBS7+pafVKRTsTyZnggIT4WBxXo5oilG5qVTVvDSHMliljj1XuFqCvZPu5CF0EvI
vwFGeXEYWaC1o5NV4a5zG8epSWSrGp8xUWqXZKjiarsBKI2361mmNqkZxuKoByJthurv5O7EawnL
bqZSPxAWzvaoGZPo2mWrGgBCkhl8XMJ0bfwSyf+uZY+qZ5tq9mLSsfjq3V3qWE5AJlHIYJbzNu8j
GyU3sDJsIq+jGnrK0dv8Tg03CIkxSVV53+hhBILHpIUf1yl8PbXK7p2sHdKfbw8uK0Pa/HsgwMtd
7P3IkJt3B9wWqZJQxrFJcrsq19VKFFAkKME9w2XalJlIwGFFoQUl31pDaCSghGNx4OeyTKxtdw8d
RlG1lTrUE099TsdEzzXSUXnVy1IKHBBaqUeOYQXoDU1z3vhEJVX+Mdc3eAHs0LYGIs7XSj/mPqMA
bzkTrIVNIWvhj1DZzwig58r6bcWqH+i0IZ3aRwASNOQoyi95yB+/Hdyw8Ewe61Tjl1ZPI3/N1Kjp
yeD3nTtk1PXdjFSqZMPOfsQBGEj83Kt6IXbI5ClYl0guFDx7xdJm59/gAW9osFHnBjr12/IqPwYS
9sz/0HrwUkd1vwQpvtTT8RMFWtBL8SoW7DniMWeJDvVWbM5n2YZn6YSou+IfXW5cr/FuN8ctmtvb
QvRGmD9SgFbSxXE42e41g9aHTnSB4Un+r64dvS0eZyJou95CkFjvqgRdmpqDhERhTP0pGfCPnchI
j8XCs5cHZkQNmmf6I2dS6NX+hqpBbVk7fWEqCZFUGWZHzZt0RjeiNB6irJ9kgEfS15zLY5wHa21N
sUf0MJ7iSfn5B4wZIl7pR282zvs3PYjov+zTTHcrU+qcmUeXx/iREEvqxUmiIqUBMT3v1l4k71iL
fGNBsIjWTCzUgslBZUJG7bkuIQvCst677rqv6UCvvDLt7pDJqyCecDpwXArOMnPfB1F2mjGmT8jr
WJHRRMob4uwsNLpK6Cfkvr7PxPyJY/2Zo28GHw6UT1tYhei7T1vyDkx9wJ1KN+q+VWDae9IvAkZ9
yvM+D456W2d9PCe0F3mnZrIcr3dupkshixk6tDiF2L6QuSqfkm4Off+KA+jhQvi/EJNZt9FyvbnA
wW+ca2nAhlv//Bx6X88iloqD9KuRcom5d76Dkhjwgm11bRyBYOW3xR6Qe9y28caBlBZnbtzLZAWA
hTmlJ8E40irMgQlrp8XfDM7kbRBB2V7wR7NhdaHJLI2OvmdAx7LbfnrsXM/UswAUiFuGAC5Tbdlc
VbIO3KUTS9utrYkg7FdCv5lY6dKB3L58PyOjtTwl1uhs58efhQ7qeqnGNnpY7hqzsnaiEMdw7UoA
WOlIlieENJeQlKC4XKZjEGYjy2Jd0RcdCWndZ5sOABVzCsELvf9QioNQ8niwvwFf3alJxbVWckHP
vj+HOAA9XxvG5K95e7m8XBH1PuKMaR3NfqlEZTDNvXeBiFe9TOKjI3xIGXbfX7enciTANSwhUYCk
CjjYGEUhp2Ob/BEFqFWLFTho7xqvrkt4aCrRdNVfYGycs8X33Ij3KXHAGorIh3nfskBCa+QbYZA2
5yNek1vl7KvgeisY0506vO19+F0qoq3+OBQuTeLTgmlHK+FyKdusuxqaPirA5LalgtaMSwQ7PYQu
Yldd92tS9Z7wm2yS/r55NyH2qF9Q2hoewBx0+hd1pvPRUAWeUB8x/d4k+z700cp3s89RUJruEh6S
Pi3DC98KarseTjC/YGXT08cKBBICMUom7K5Toa1JQm/t6sDGYMuK7iesdf0Hy5YiXrZAg+8uL2g0
QrYQgEGoPPNq48RQXSzYi08FC+pDeYsPIaxhcRi1nhbVw0vtLS+M41gBT6/uvgwXW0eh5zjWxC1R
0FpuSZrSBB9oUMYg8FT2daQam30GhCFrMnYAvqnep40RN98+2JjuyXXVwYHh+lnblsv0taBI6pZj
02ZNb10sU0/bxZyFmno3N6pqakqicHh+13omH96bcLhkrIB0gqmeGRhFIVprJzdwUQUMV6bddyG4
yDiXEJo7oVN3UlnhG42mMyTV7DxYDZA1qYARBDrUV0mJpZJmAI7fBFfSmOwXbVqYwtc8+cw6atKK
Mkdl2Uu7r5L5XNWLORiVQyiRl1V96whkOVKtPedMYnC4NWFz79ALAdAf2blX+KCtn9g6xm0sIjqj
CAobgAJt4b3GZAxS/MOBXi4pCHkDmCHAb0VejcK2bIdcOZyakacIVWdU6VGmlEJf83k4QBkncyti
7QUm4XdPTX5JZwX4AOOZvW7IrdCMgoCLfTVGOA9mFlobSlc7SaNIM6xCHuDPR0H8F2xSNzWL2z3Q
/2ne964Otua9aqPdU3tqznitq6hsGvCqBq9mpf9cnG+7CWKrFXnYxiRb2VVmieSPXox0Yc5LWImT
XYsqGXan25KwIoR7J5LJu30AKRdQMPxUHXS6LtdBXNRHPSCBYedyY0nbRBDlsKvEMK6iKikyln/U
qd27Xc9Y48oOqZd6kMcsvoL9bMHk9T6Op/hpK9rZfptnAxAmLeqrbZaKjT0MH61Y8hB6jsgWwp1Z
U1WkHk9/bMNjqF58RonB9sKskdNo4wd56ddUwOPwbCsex5RlZ17T/X4So39rbkgls80HKwqjUfxk
DW2Ddl1BEplGKN34RlSEOU2iJYqnaW5WqJs2nBe9Igy7aywqNPAhwF9oFqztzs1j+LGCT3Se06Pq
Jk4u/U+dHMyXl+364zXL6a96ZeBOcjv8Obvtx0lRWROfZ1aG9bGEYTD8TLX2ZT61Up8t9nQB9B8Q
4NQNS4BenATD4TjjKJkUYphHLoEivfOpvYhQnqpzi0ula1rdX4uxuSTic2lGnSaxsOm30g5pi2zE
+1E595iNYTjqHVdZFtVg0c+ejwpjsQODfnAU209o6qXH6n8lZXyynTI4Iiw9PG6sJZdqMDHspOsl
v7GwX2Q2PI+sN22+zXW4vTdpSUCa+qIStail++LyMV8vvJw4JKIlDAaGVygX2Q+hMdyIU3r0LxV0
xhfmx/R2M/IiRNCPGYCQmp/iB1lNXhrr82ZuApHCIyp17W+4X7by/w8U95i1Yux7aGKMVFo+EJPt
GfuyIkUVJNPO5aOsiVUqG+ilPo75pFziVay6s6vA/w3XgoCfPdidLKrCC5dosLi/IWrESlaMbBbD
k8FdmPGGlC7wUxF6dMR1qyc12JQaePsXse7zrD5AFSyEYT8+1Q/nll+SLlXRMO8qIw7EukrHlope
g+AYq6bFPT/SRBxMf0fxO7cWD7g9czOTgNjymtNhvrRP85MEPTpXQQyHdUy5C2T64oE0D23qJGgf
X4E1LrZNhWTs9Pu4XVmIgFWSgXzFWQCmc9EOWkS6uLJ+XnBCvWhSmrwfA1GRV6Uud/fjOgq17fsL
OA+8gMM2PF/XjfRBEkM+vgLEgl29NQF3Z5rULM3A9EPnnBRc6hZXgpduvyQMUxwuBi9a4qBln8B2
lZFnfVqbvsczla6isdKjEqKKWMgSmHPNLeLeb3GreN5kehe8ot5lOyuT5OsGehM7wBQxhWWvQDAC
Le0ttwDwEkD9PG7J13YHtzJnpz7PLFCRShwOWiWb7Ot+RoDMwAnH5MlmCFLMW+C+sUcoECIHOCmb
FpiSKT3ecWlQyF+5A+KG5zTVzoAip+8rnFB5mznsRFoGkjCCPJvL6w4NTa04uMQvma6dXIiQNPNI
HnlKayBFtTdINbNZHG4kG8DvYX/UCwViovaqdzulQfS4uHIw1+Q1eboX7MgwzJlKfst2koA3pVcW
tcWLKkfvq7J74J3ng8W12Z90woJCH+qujeUdSUAPlMekNr+47aow5Cx+DjICY2m1ikT/5ONEM7Ef
j/iMcdvk0LuCMSI5UQbW3Ff+ipUMclBy3alyDggifC1zQJ04cWKJFeqp2YibgGTiFl2W18GSPfcA
4Iq8k67rU2RbgyJXyAOfHZ6IwAX1NENSa1y4iflcd6UTeBMhXupYJmk7RZEuZslPGmvf534ynSzS
+azvcRWGYYHSWASB4Ehnj92WYYN78HcIwd+q4F0rAa1n0RzKxBfqbnTVa8xRSKphPQj/xLb8S0WK
v8BVyOKiyDhF1F1wbYVGF9wBJr+OM8+cLgZ6WT226bT9p/ryDDTOseML9NH8mSj8Iyzqb9y4VFrx
t4QS6kVSi2EOaMksWWqdgmhw8pO6nDXJReQph4cerH2W04nA4Uqpf+YAshj7GEizpGblCKi0G98N
Co5q4HeNFiaqSTxHxj6WwKclJo6F/OsXfV3bWuPJd3KiE7cg6HVApFe1RbCallh8/0iBXbRfEnV0
B3nJofV8GLlAcUSlgACVr47XXyaA+BqNwRHcPJUpBXBZr6LGoWuOqom+EfDCV4C0khZSwxuBA3wK
9sLmH5mR8YGyBt0/wx+I9+aZijYpsRMLMvXFWcdw+t0OHfpjCPxpugpEC1VY9f++YLjfCszEEWKW
R1qCbYb92lDzh86+8ylmkcbZxJackdwed8H4kRDz2qUNIT2V0ONG/CrrJVUnTW3rPyRPZSIe5KbH
HA6HH07WaYnSgUKfpzlSfPUWon7bZDBlJZ73y8yD5OuQM2MxPT6IpKtmV0zXtY8lPMDu1XMJUAKi
zRZh43sMCE1vnorzBO1BrJ5a3qPwgCfW4y1uJtd2A7uQK6TNRsKFArd//IwP9m66sN3NJ+ZssTvV
kBQFqZrBDcbao+/sm/F8+AQgWaDBmGRJTwetySc5n+MO20zRsfJHREAYttdi6NZq7zpQ4/QCTMvW
KYaGiJRi1bpXc1UagQFCmImc2yAzghvDS254S2iX4Eb9IUkvIfZvfAzHBRcnEnie+n4blyuGuP6K
BOd5e8tDsF9DKcW2PKenEi7d+O8Oxjck/sGBa0424fXVv4XXKvsQGERae7afNRP6fksEbZ1en9yH
NHwdSrGPSgqBsPsnSFK43E8jMRTkvVVEkvhw9bkdnl0+KNJhnV9F60X4Q9w676hSSJzSsX/grhtm
Fu0CgzvOcyvjSYckMiPIk650EMq56hHL24wxzotfZl9sj73IV0XDyvIsxlvNfac5pGVU89MYcNgV
V1Lgmzid546E98F7HPuKhUAuncEs0hjp/SAvvOiOXZaPY4/fzIjXUVwkQsVsLv28TaaxMYr2RaNk
3E40TEQKx6GIwPmtBbsRhdvgDiKcBckVsrPGTjWH5DqqHjPOsb32CzWWsUqJgfKB/LyJGRQfOpkT
AqxEa6feXMIajhrorgZXCRiZKvt3BVDxnBIpC2fk+mUkau4O9NqZFXp6y7xpFlC5NXGaRXMEdMkn
bfvIir+j1axm4F1Yor3d+DkMw/jTBENtBFeT3eFPwn5shkxq3O3JboXeBtmxQX9fpoc1IO+QSSTN
kyfLHgiyg/3+skCJ0vmjucE8kFGZ60NfJ8cTfry6ZESp5MtYw/8nS3E0SHsbaMvpzuMU96k5aTe8
IQUmYWAng0W6dkaLqwBjOyW20n4KBMyaxueZHU24QfxRPH6CQGhJLb6GtdmNLEEF/EFsoHlGcp3b
FwzMAyaK47jGZVQsyTDZEqLI8TCbkH1fA2vUdpbxF/aXj95ZBvAxrtx9Olc00oDWaX9twyMt0Cm8
CVsDbtXHGMKmWfGBE53p/daxJwPv27ClrzBCRVhh0tY5ypJKTK9UKEbOLdMu/wWhQ7bQD/t81Afk
CcO0AirfadnCqquasGH2rLFT/1x4dMNFNjy2IPf11iBDxLoAJ2Q5hcxfXyygkkQpk0fnPGJmmONA
wsviRvd4DHojl3Cek1QvlB/ZWy1AN+CXXkvAx5hVENHHBZkg5JuCodEPMjwZIampOwk/Qs7Yobkj
Q0SnRjvU257CU+o6upO7PLDcDgw6tgDmhpvXYx5vkVmoP0Euab7Okwayw/IGTFArgPZ8VK1WesYT
A/X5YTjp22ZNPMU58nBJyutvMKba+2vsZRxcW9lOaDZWltwNFvVC+c1UsxL9Boikg6tOZ1QPacqC
VU/zi93oC6XXOYZpMGxUh5ZiwKvgrGpjiHkb3Qhz0rioU050sjbcev5FY6tRQS5+G8UoyaCjQOw+
Di0pFD6sbcF6zBTXDBsVvYkMgyKTow3do2JP3uKx99TUQZ5wsS5WMeX0X2ZcLgvYInBddoAm6Miu
JL5/3OwLflcvZ1EvL8v0GEFF+6dcJQR++GmypfVY0bddQHG544WaipRiA5zXQvOhCt8WvEYtBu+f
Qji0vUBqjOcvWRt8WFwFCKCsTIq3p83EXmKj2h1FbkS/M9+f9D2nKZ8fVOHCzrseAYkxet1FeJ6U
emJydwryNnXWVupbXYzNF8NmoEzxR4jS6di3MpZyf8UlqkKnlwBWNtfCxqUQxVssAwksDTva7mlB
YiLYaU2ZSMfg0spG4+zxB5SNkaUMfeRa4o1GK0E7DQssyR6IsO2HsvbVcFkZpUyyrp0ibuZVxQSk
pOODdNKq+juANhiFyrkxNmI9K+o4nygMzdyODxQ2TKv+x+hjufz8kw9Qy4d1vmcHhMoMMSxP3iDN
jevw3N32V8hDYcGMz1mXtrEZxYT86zP9RoDzgNYPraV6gzsmtdyxLSqi+WBkwtLq9Du7yRVE7c72
eRvg5mHeINnojvDD3cscD/A1PNR6IBwIMHLXjhQFW0WPDhThcKuSC+kVUyyTqQUxPG2Tb3pVo0uD
XNRMVParMaDWQ7Tpwj0m/pSRE69FHCcA4VJp/rcOEP8YvurhKYxq4lXDDui2MMse0A14fUMauJs7
oA26albx8XCxJICRAVkLhl4ZTHaK/uWLiAjV3P6n7S2aRHZdlhQmrgf6uGp3fEXjxjMEQlUcQ7hR
aKiC79VFkLfjR69KGmwi1AxeWjBA8d26K9iLfhf48Kk9klp1HrEBBTa2+TTCW5LBMvg6qs1zi2RD
ZNXpEUQcC5vozwVuhSU7DUzHYrux6e4JkQce86Y1KmTts+hKGXtGWfXgky5Gs/tIkgawXKDkqzdF
znDYv0qmxtWWE2bp2ZfyvlshsgSek5CADh1ZpE4GJpCT/SsIrEU/GyPdYtwK5v9hGjEU/TvKD0Gf
Sdndbc4BizEO6pwsTiXKGY8gAA2hBN++HqWmMV6XS6p9yrnI1VmZwkJ2ceb1pmugjeDqIfg8kxS7
du1HMtOrFYIj2FxSUIrn4ZXhi538IbSv15PhK0+jbhAqBcVkMHOY1MzY34QN2b/QIq1RfJVb66X5
lquB8yWGYL4ZZ4j68QL7TqcjrhNEy1VFcb1QyRTBucd4Ts3o+2EI8+SiGiw/WKB6rIRgADDTBczD
3WVnqChumf+upVpvmX2WyqzOd6DxBH+9Cnmkrmq7FyF5VaeR8Wstsx/UOc+3ZiYjWs6QBVfKlpp4
8o5seSRsh4sCPcHdB1HzUGRnYh8VWz91X5GaomrvdSxLpvVzC9LsmME2CAO770/YQYsPD+WcpgAE
WcVSayyosmDle56EboHSvKk03LtT1rGrABJse/WV2YOp1/6aZjRJRcjUSS/1mp1dbElS7Z+YT6uh
CcKv3+qVB4mQTlJf50jFi1M3SK3hnG8C5+v8eiGfnWasem5qwGkschvphK7FF1sY8NZDOc+kNIb8
LKrJvEWtMCziC51KfT7gXel9pS8bdF2TqENuu92NYKLTCST9kO4yZHoT2tF0Q11KAp5AgYhnMeUB
ttFTfc23BdGhI6M8rkSe7yGS/oXL/FzbX+AbTWDU+j0Iif0gEwjheNrzBWFzU9kS/D6PIL5aJbOA
riDuzuF8jC4QCi1BUYgp+Z5y5bu7DrozjKC96B+4WRzHBz9yWf0hzYiyWLue5j1dfkDf+rjlTQkK
GDw1QpmO7hY929oSc2kz5teIhKUSJllSkN+C9SIDsSO52lMmEH+tCp/E5dLqRA+fZsitC4ReKiTt
6H1Slo31eyVkK8IovfR/QxLxWms73TyNSyktO4Cs+1Kf5+C8NouKGw7Hw+6xnX7gJphIJJ3rSAnd
Bdcarp+pPli9Pbw45KvBihOOM7SV+pyJbeMm+Q2OnCXqVPIWhLEn6+ESdjwHgAaRE0JmLAk/894T
359s+WDBbEsfPF7eSSX/leiacpa0h/q6HOr4/25n98md/8URuqJcpvdJXJuCu8//f7rWJvZfVwtg
Sjdo8Mq//2bVUjdRCYW20ghtaBgECfqxOQVhkDk08yTDk3bJyEO0L6uGw8Y1TW8fTxq0l+4+AkAF
bliBY65VEULwJ2/xLO93vyVpAGxF07A1h0xKo6MDI5JA0CLC2bQHvktnA9Fmc+zEuOfkFKVs20aM
XSl0ZdSs9d9l6GvLBHnbb8lXa6tsVuXvCpfe/9xTc+7RutQukaP0U8UqPOjvIBLWXal5Chu0Dnqr
IwtCKRHPUulQeBunmU2lFSAXV8DyKxAXE1YH0oKGsuxm75Kood8JGQrA/CYzJpIIfR0t1Cizdsh2
EOtEqXrEufnchk1nSOr6mhAK+lxGOQ/szekcBFdAo4O5g9lYKfMN7oJ64umYAy+15O7Z82sPLgCh
WFzSYWUg9p/Fn5UXsujXP6ks4MMvRDV6qCWeDp+33N3IJtYosEMg06zguxviUk8XkxNFHag1g5xX
78k8LHLxVRiH6Kd8OZ9DmuQEIcIYmJq2IJv7MxGJJ9uXO4Es8XyatKk2ZVIcpL8XlHHiUGz04QwJ
kL9MyjpNerXyEQ+ENPgJC/mnBFUTBz58wZwffYrB8I+Ej7N/xugML/gOjuwdVMCPlb6vF39UlzTH
k10OOpkgeVde0rvs9LqP7CD+q0PKAFpy8BChISmhcIWFWE0UmV+oXbDqFlRDWem/oicu+HdMuXyQ
DTkobv9lwqCOoThtaJIOB6CUEhNxAEXN4GgzkO1sD7whdxo2S2mLHudB2VH58C/4XR7c+ZMk5tRE
GKs6y9vUXvuV7YcALI9M75SmD5mmvjjnzeyvdHnb+3vOthSoI2Q/itZEc7Pxkla+1HvBlzGAAlUt
3lSTrntoT4XgkesgH6fwrI/K7DzC5q8HIX89kPZTemO0bAF/Wz0/33VbM7goS6xtZxTcD2y3suih
uUlMkO+qOdX41OvD+O1vabobCg2axOuHIpVaZ+QSvsNdoGyOXf2ll6Wx1W64lmBmpeSCbR2/7O+/
UBKybkSOysxRkys42QPsjD86sLfEbtgUwibaE3IaVwBBN+Uf7ObIYaycqRvRdUUvXq0A9WrSPVDA
bOSoCpZNuS9W8be5T+8wHmlGwlNVbvqpHyL+GEYQt0JVAcz2B4wxOLKF/+Q39ZmScs4qEnR/IQvN
bjq3JpzabpBW+zG7Tuby3buJ/CdVDoWSU8UUO1+5f7HwIZ9ssRp5kTbtyv559dRxqFmdL6Ca89MP
DMxMpL5P75eaJPPbhUvcy0l2l2sgcB5a17i0UnyDeu46AskV3f4RIIxR+ukB/xRmPnHEOzKSxqbl
3h/gShufNggCCE8XSH+1zxhbrwnyvQ+pjBxiKzSVhdR3p0YQOqKB654fibuhH87A90xq8eX4Ck+j
crCFt8auVsXqvH1uNXcsprgwaujJD72VCOrE7+4rFo+mKaBcrtJY/QivPbHIeov365zQ+I3xO+y+
+IaUv5PDyfSwfM5fxPY7sK+/+8SkEt1Ar/Akmm/rxQN+ZJb0oWN50cRippepf8M8V8XHyaUW0zw+
gJ9mRSV5OgRVRUD5cf3W8zJRehIXJZAsFO5N9wrQZHEbunPTR1vmC0byG8SOL5ase0hsGSknBeSA
T0igRFI7dTQWuAuwcN97Pl2h0dSKDfVcJR9JSuI4wadFTkOhMOxItZHgw9y1tSYG3haekt62Txb2
vOUk+Dmy4e+yRbfz4nmTh4YltdUEKZiLr7mh7aJajV3ukYVOOYl/3FrlWs2+0GSdM7DuTuxcOt4+
piZ66Mde/2ctWa+FApIjDjTlgox3yY4jvUn5rCnx1lFfQRfmcAYClTWoADS/XXd3M2cQA3jImwkW
sGZW5yQWZI01/sefbZ9zHifqeK6evn6HW+IHyKG0Y0XdqT6rRwPFYMi2H9kzoE+/qee/Gol97yyu
UVBNuZ8dhsjvQRw9cVV4ikFL40WXX64giKmBhT8utn22PCH2gNbzpQDiIQf/zC1x0npym5Ni+j6L
poLmWnCU4hRt6alwQ7ctgEsQAtYJe1s9fFlteMfTJojAHl/JMPo8FDK77Z2pUzTuqWwnEs54y5in
r/ycpqBnF8+/RCtKTrFd+TTjZAINcVDqXFDYlwkGIFu9FVvJzDsrGL0Fkg+bctUdnDlR1XPPkkVa
RzLMzn8LFYa3VbTEusSH3FoAI3NjWoW9iltcKHZaj5wjRe7v5/e9268Oc/RbsmSm2U76kmSoo3TP
ypwoa9pTogomxX42Uxdl2DykOoh4f1uca0UJEiVEyBc4c1XD00pcO4xhfHpfD4jkMp7WNx0RTP5Y
OtiRmi/8vJ1J8L6KNbf1rxtZQwcC1kJnrYP1tYttAsYODbh/e5ZS3C9ePjrqm/AzBuJTEyluZd+Q
PFLPBFTasBJa2v5kwQNtlzCWJglR9z59zEysh/pbzpqgNp1UavGdsQzQbn9tMyQGjuer29GTeCK6
i+RmGqLofl4Isw3B9aNT9Z6pIoqrRHailz+kc7fpl/QY8YlHmBgAYSX/A7Tn+DlN65SxrnMAzePA
iNqedGbQvpsW8yq8ih0bQ2ZXh8UszCuEu5lefqSLXxn+aJSTHjHY/ZorswmT/VLE1qFG1c4VSiwD
KtE/xPsDVzM++nDNY1h7xA02AU64MP2fYZFC5+mZjg7NLvly/O7hwjn+64jFZLSvs28OkLRCXkcK
xsVDY3c4mXzSWSpvFz2wKPzzRkSPxJQSlXM2DBqOSGvwG66ySpFkcDgp+ciyO663/cKY5CmODXUJ
s41iCtRv94/v7PHFmo675zyMwIww7bsR60vu1+/f3TzeANJSWOeJyK2Aorh/upIkk2Fj1U8KkAsb
qbupRWhc2B93vIhjDtMIjEkT1VrMZoxq6QS65IqrARalxe1iAVhzXQ5TwZ0W5w8P8YbKb9elPvwe
kSZ2X4h9HE6Ry5A+3NAfpyUdNFQ+u2upHzUwn6Dn+uZWN+4Ba1AxeGU9AUjF2K+YQ1bzrVHikYoY
CUxO9fpVrpVcl1cl1yzwWQgN1mjCIzVA7fovb3x5I9dlcMdM+fTirJsOwvirUw3zFJ6K4yzd1YGM
Mpog+B5h3DUzVxwThRC+mxHXIZdYMjK7OB/ZFHG6cM8jVIcxsW4Lu2WyWS29F+xkvoW8256CpjfC
kirfoUPKmTaP5YaXZxS71bSheOpeAcGTIN5y8XaBO6kcywkm8bd6vPFqurswJ2lPhMY/mvdfso41
5xGKm3ACoSUgNlllIzrb9zEmuycSy0rqJ4ZAlBDAfZanbxVXIaqDtoJhtlTnVPbxdza7MWuKFDWM
d1e3kkS5xinu3+oWXCMPDUg6Pk2OTZp0aqcdZTTVlbr/0NHFnkTwt0gkk95WhjeHf8lGRyqH0Dcx
Aw9Hw709BMTB/vLHVzbeXGb3GSVe1SEYVmuH3tAgbc5c6dxWDyFIvOkNdmU/X18ApCyVHkPsmxWE
FFPw23uGgd+W8Lesnzjxr0qQDmAewSAD5Wo0FcWuZajZ7X/6LSPmUJI7ScfLL91+JfHEVGIToPxx
dTM5zI1jN3lBetV7aAdBoK1XbxXrHv2Anm+fjNe41cuUpu7ceDSHH7HWkS/8yfnGsvcol+VT8QNz
jkFsFluME95oiw3WnEs4YdZ9omrzGjhaBlmEkCN3VqSF5oTuHj+3szJN0x38DdydXtGafufunoAw
SnU3wAqZWKDbh718rKxZRFvW1zTmtXkJygap6ffYMantas+iZR6TuU/UxGBJp7bsh7DFjvTpfE7D
F5pW4yMR+tSTIYCUlH0GW8XaAeWTXEzfO5L1GWXFL+am//1xVfdwsyyxuGX0xRnweKNpztEPgioY
4GYS7IhLQx7X8kc38NdgeNGNMbJZWpc94T3nt2pgwcF0xoZy2jybrzTcp5xATS4NbRI+RdVAOaOQ
KOJLgr2qYHuJMZSLdoG9iscOHGwaH4oRgARcPjefQDQxwung7a/10PweCW0CQZ786NXwaFXeV9VC
9zdSadEf3zgWXF/ba0j0TZ/X+pfDCidryMAu9jO33GY0Mz4/jRRJph2ODHjQbA76mSPdsYGPSXwM
XhMJO5ewOU/mUV59Cxovvfbo9NDf/LlQ95ifgqtdccXtFmzh8LjW7tMZicxyxgfuMcRwRD33TPV+
3rvMn7qHkxer9Z5H+GwvyYmAZFIrIhlvkgJmxuVUeHKYfDFixbYFRiBgkzncw+97mLrHuUVPscIH
dccB7O04vGrlQQPg97TFW7Llf1jhLdkyTuocrSbheWseFs1xo6t/cK6P/ag1dKSBQSM3jGByVjLW
ieovMNseZOMHD/1T2SAnSA1NJlPAMQaWVgBEHMGFYeI8Q9bEjjUQYGoOLA1UHZSqd30cVn+Q65PT
Zxlg33Ed2jW4/sHonBQnqMjOoqtu4jkyiwFeIxwdWoxOrKF9Vw4+LL+ACjqOc2vHPtyeL9tL0TP2
HIYVTqjRt8w4wuYxmyzE4909gc8vP/dK8dtDjD2hMMW1jWzFi4bsTYgioHG7Y4q0Y1HtXU0hr7fP
Bs73oLlTtkvH7jZazZ+XZigv8BZyv4vFn1uXiIq3zWTnjfiCMeV219w+5VPm0Dr0HArSfZ1IDZzP
ft101hi+pZ9Uua9K2iuA/9IXCkAT4FnTVMYvrkipzypSpi3i40J6mOine44fL4Dt2xMoJOKiRvXN
XZK6zkre+BF4kLtWqV15+EkTlQuvsmRrxAVrDM0+PK98ridMiTtgEP5PQn71jJG3DanW0/VEE3Q7
Ei1JVmLz3OaZc/d6b08C7SHIBg4VukS354u8NYIVAmjh4IhdFCir1NMFOPvIo0D2xr4AC/69+qLl
0OpHsuETOoN6okXtqxcy5I4D6zJOztFXZ8TqfCUl9OXvdTVaoQ1i2fNCY1OrZyEwrI0pTmoQN6nc
tWvLGQSZ+E7fi2D4AXPVExtjRrPbbSj1a5Fyua3X/zAXs5dXeHiMzXXE3Zi0ExAD1gS1B4I52kT5
HqreoaQf/f3zuxackaWXzTs05XCCm7SvA3gfaBpk4oShneMs9/mVR35aiQ1ULuUZlryCzPx+XjrC
OdZEpLyeyuxBDrJ3G3BF1qm4odiahTigO7BjFOxd30V303SySgkrr9G6VLaTx0t/p5q7/xH750rl
c7rxhv0TPnlorSNaLWC/sIM9Gxdnil01kcS0yoj1wqhrfrPrVAIT+PmSV3ilb4hrdHWBinXnph4O
eKZkOghnfNnX/mpE3bx+3MLUhdpwfF/V30wqq5to1a0TAykNVa7yD0XWiNzzBot7CTciMw/fa24d
LkHyP8e4QI6+9bGIfjc+HHmjL8gNd7DpEpuhf2AMxEkcvS2n8txzmWMIaSH6e7Gyo0LTm7gt5fxB
vptXXp1kK9Chmh5HEYAO1KQBWeWkAjssNtRQH4Bvdr+jCIZUrnmk1tZMOLXs7bk9+BE5FSvwVCAu
UYbLBlpyc/4zzE7+oPDMkB+hjUbVaW1FNZwgdvhfJBbD3QsFBhxtaNmP5Qai5WE7yGxonD79FbXU
o6PgQWQ6DIIbptdP5RbQob+K9Nx5AQaenV9nnKEpPO3ra3XvWiqwdThfXVSiSNDokGlUpE2DrVg0
LFLvwIgqSNSQZJhI6uBMFb3NhIVmePW1jjEfbto9AiIdGCjWvj9bVzTK+HdCxjCuBJ63YArdjJVS
WnrlwliZ+w7qo2XiPrsPqi+Hc+ywhTgbRWWImc/4nIEwIb3kBvTtxjrebNNHErQ0Lfa3XnzVrYKU
jAd7X7ptZL/nWiZqVE+lYwZXZ1JWuRU9J+v0HYtrIUAZHUZImn38rQrSDlVd4UhdmcAm5Ds00Qq+
C2A9mlkfdUhnwS1sXGDHkEj69svG3Npn3p19+aUPlvjgtZxJp0uHlzjnOYuAZqYslcZjnzGpNmFC
kP96/4iKt6oy1QTJPyzlQAd+ZTGc+NM5Q2npFU3zeoVM7rpB0s3xc9zigO9MhWnR6TpEoeMvaKgS
p6Wz98TegdlSVrnp0e/Qxpe9Y/bqqhOMo8ikkRshEOpVdg8uOqy6WBrHCcWe65aquZVZPFN4KvgX
wDd4Cljs4oa9haAH1Hj6j1FSr5fympk05NiWtG/iaZ3UD9gEh2QBtb8dvB3O8HBQB7xr0Z8Kye/N
MdJsUVHjJUIbJlrvrEmDOHxOOuLUTgUoe8ns9DQu7mpV2RbWG90HXIiiJ1yOotQz6SKSgV+wNE7b
3hJ4ksXY9TbVqwUpMqRADTXrfGFrsd1ikBwhARepe8w7A0OGF7QNehwS6woZvJJkH5x09jOnI1B6
2PnXZOrQxw2jn5lhqyKbVENKwtYEspcyccUiDYYCZusdt0g3gXOo/zpcKkA16WRc8MmgfJPduL/u
dGpaRD7RRkAE7BgfMYPdwCmHaaBdUzFPReZKGzMvo5E3neHuUmUmK38TEPu9XFys86YJ/DnwJIqa
7T8PCWAsAyr6p+dT1tSU4R58M3LcfBI2dVfF3B0WLKcT6KbQXY2ix6ghn7wqcITNzVHpBDdAp9Bp
ZgRRvnjwk8F6ss+x+XPs5Ga60dJwaZUHxLufg2KasX1xgQMvZwqDLgvHw0ANbO6Tf9V8cvL6xNSZ
MoWQeMkymV1RHZOLLxD8WvY1VbWZcMDLTVrqt0rjwubfVbZEJL5l7qzchUGZIOAw2/jvvjTDKRmY
dCyIclQF7dYXKrEk6tw/W88n340zTyD3Nx+w7DFZBtg5vtyM4WaenF8fNZL8QXmrf0u4xtA+7eei
gJqyXdtxuzLQlg2xzNe9MA+PFmKls+ndULavIaFGOZtx2Fo9VZH/KgdVTm46DcmFK28RSfvXJaMl
5IlqCVKSR4egns0U8KqoQzG9NRHVCO/QKvIuPktmL0kpbxyRdoDs4YHg5S6TCIrh28wNbRaHDfWd
iiir7aUJgU8zSvWHZT6qAdpxLB6sKIMjAR2VArq5Glh1vmBrajN8QLhM5VXHzCt6HwAsYoWkYrxD
f2mDQTcFg6zmNPxz8ejc9EyhXM/Auxi4035242et4/s1xEr5vQEmCqtznlzG+gpu/q/a3YwElWCe
nw23pW/1kxKx3z7UOq4ZZqqoF2iF7DhjxKs/TMcFdqd8PDHtghA/U+NyQ6V7LvfeHXRs0+Nx9BGx
H8VslGDdiQ+zd+PPacrE45FgsDT2q3KhIlofw5ejJIUWqWCRFqxvBD0cNN1LAzWjZlvX5sNYqgTI
nogZ+xlh5GfFdcCirT3J2L2nLio5/OODkcYpyITDUgXRWx0ApxPJ98PlEUA/3TLEiP5N4Lx++XjB
AxmZiHwEPtyD7CX8w26ApzVpcrRlH0FW4Kdr6n67doYLVHeclzSXO2oxQBoRoDNACV/qeA7LdfFt
iJuJdYWxJ6l/2f3b3l3acWv9Z/COunluEkn5uXsLnlkFddkXqRWPRLvTZgZ0BR47N94SxBLXthGp
hmRGokYolQ4qM+FMU3D5R8ZDhchU2FSPpY/6fJuwCbws2cWJi3E0IyHBl1qPh4Q8PdocNcSBSj4T
XVaeUXWRgURoVwMnONTpT5cVPCYcfGpqp1a13eMYJEYdEU5792GqFDqxZ5EYnBVp/AFM/tkh8zH/
JA2puFHkPPFZ7xvqBcxnVDe47yxZ/MElLSWlRE533U5etRkYUsb950+rVfIDMa8Bze/qc3rYcDvW
ZANgMRi1JDfvfWXlGxez+iOh2oAqA0/8DT/KyRqdrcQ6E2xyBMv5ialLRNYyM5DlyHK5Pk8iP1l+
dURrgXILruRUJw6v49htB2tR45/v3Lo+ohICaouRqQ+rQVrEhQNMgD+mm0FtTiwXJlJBgenULYTP
qhIwasXwicEKo3T2zw+zXhbEVvVzmDTczlL1/9uC3LxEQVxx2KNwdBGRo3goONrLOWjyA4GD3xwD
Fjd0w4E9+4RoIx4ghyHGsYp7SQ/jAg72aVYST4nRQbCzcvYIRbNynRW+aOsYMJUfz1zOs9/i1s12
CT3ExR7LSxc+hDaBj5oT5yhnNVZFhYtrMwQXa+cEgC3TZkBMRYbWj4fGT9K+LvJFADTOSxiqB/ks
WdCLJ/BLFbc6u4YMjO884SMfHfkIqE0lZke9vCiYG4oBa+WV935K9k3iQbHmviKohdtUybwT2+gF
e61xv9mnnFIthrGk5F78hp+FElF9uPkA1zHfrDaivAwsVy1dCf3oT/L2+fEEpPq5PbWRnaR9K6rJ
Mt0L+ckOHS6wR2SComkUQwFZ+bf1aR2SwCZifcw5r26S/ymj4cMjPrSipgA2EhVenlhMmVOz22PZ
RbgCiI2M6AMQWE/22CAOnWBZioNxMvf4ygBQSuQd5ciDjljfagdp2zSMveCY2KMp6RxEBbc7AMa4
HgNvSTMnBdSEYRTbbWgsTA4WK2RIaZhy6LfeOoOZN/LHQWJavTvaz4OqzcnZ7kRrqv+j1rD51uzi
hFvjQBFEJmk0J2RdR913gigWG7eJYuCTTmvT3faz9Kc0f9Uc59Px+M00QKQqI8tVCz1K3CgD8Amb
T/esMCd4p5nVWXJZNmWSBp14D6nTGfRw28MCbEwSavBqUtdiz28dlsjYuFgYjlw9OrVVsv65FMzN
OHMIfUats5HRZquF7Y4PAG1+SLXfWRWeh4DrBI83aD81OwMcAj1aBMMgvKxjZn/Htistn0JxjMis
kQPrBPKgswZXFFsw+uhhfrE+UOUl1NlRuepahbm3bKCRKN2RgUcCBJpFRKgGbixUmhUCmWgLYa9y
qup/3ipuF31R5xfSREI2UsHDXLfOo36tVnolKaoUMSlVXKT2SzD1MEc/BjzP8ooVNA56A6ZCXZtO
IXv/rM6QHRrKT/De1RrRTybPc9oemVDZ6d7uY2HNIbQO8Z142BbwHSctZWCVNMY4kye0P5WSmHb6
ZLQ3XFyzah2mqqcXRObOUnNBa5VKEkooO/MUOngo1rtv43zWn2vxc3AeiDfVgSq60ThPmD5DPUMF
qE3GpfnQ9Ob1Dg4mIvsDd39FDYx/PF2JRdRFmfWZ888PhhmDfamceGEzK7pJ0lvfHekiRp7lVxuu
kqBmpRjniPfuqLbVsJL6Pz8K8vHuFgeQL52la3Nrl2b1O+tc8HcP7m01RXEJPMMwUCgty9o5iCKF
krrBMop0af/j4Df+t2mepW+0e1HEBEvRYTRvn7KrlSoRGF9q418sPt4vaLXIiKYThGG490loGIIX
vQ3Y4MbmtFfG6qDp9f4vWSQGQ7jhKOatcCAuUNw8D/cw4aU+ebUW6lVTXKYSIWZhkrIFMsIjwOaJ
WwC8QfZmHtXVa6qVUd/FZ8M2JnDCjpKs9f5suxdjbWSst0xZ1ittxNQZ5IUEIhG5QNvbCw2TehQn
kJ2Obrx9MNDLfIs3qbP3zgbLDCiFKXNLcZSZuvIqS/Afp/hD3gOO5opO9TtGlliZCS573+oUQxQL
lpmFYsbmiyQilBFp4rYP6ntqDAddBhWIftsXaI/oi/PLKpwbDz5fB9Uz4gr+9oiiaZBGs48XwCMc
HGpnrPshfNXILLXd68DKMQvETBuLUi1qTce4NoeFMZ2fF4HyJkmJvaaRraco+XCz/YLq4MRvr16+
1fh8l8hFm4LDfpiVr5YprrL80IvFmVy2+doKZujg27oBG6fy0RGV7LfPt2+2gzwyF3bgExELKmpx
6Et7nOPtyhQO8jmvntxbfkCynyDwMFGZTJHAWx2N7GeW5E9M60Pa3YWE477j+nsshzmavtVjT0cg
0YpqFycQK74pRAGS0HVkKFduKQTOjkzg4Umk/FQFQIp4tSetAYEeR+O+tBpWi0paEmMHqi5NFYwt
XayH4wJketohMSKTgNxkYDFpnntlROmEsA1s0HXVUH/MOgaZLubgbRJolNcTz2LXaCZk3/AfMRL+
CqCRPUAp2qbToYykkP5Xx0K7HbTiBsStKqJ613U1gtS7IIY6OW4dECGDFoLGx2anfXJOAq92YIRR
jUlR9B2sslej0lmgeHXOjjUNmIYJuYbInPW2S+x2MZmQ30sjVWCx+D75LVGAtR+e4QBbnzmfktC1
F6Tesg3mpm4uNgl0D5TPsPzjvPORT//SBAwFuFyRm1eVcrV0OmHtJLfD+TorWbHei5dm0H0brtZg
4KWdOIf/Hdp2mNVcN9+spjv9XF14NbPwl47Ytyy3wrI+wnFqBa7/ZFfpAtTsrri2mJdMgdEG+vFf
eL5iY0rvGOBGhV/kr/0AlWLeWDYg+kdcfeWICXCjNwV4yFaob6qkHm2d66ovfuJLzM/U+nCNU6FH
FvTFDT9VSHKB4kaPhgX9y+kzjiudr87FnvlbmmClFebLpIIJzPcxNJnvAw173Yo8kDt/pl6k0aXs
2A1izvXoxP9ilt3mmfyCyGUrNKAdiwI9YUJVldLj9KieKnaaiPUrfkoawuWeq++fy+SYfcIezpCV
OH+e0g8Ju/RIJOHozxMv9oETG3snlmNAuzuodEGABdljAiyF/ZdMya4srdFHf2RXUppE/p6XAvHJ
NpQlCd709gq5NM+IBG/ynOaDEDMdhUOBJchECmZVk+6Y/vADB80F1ZIoyIEe91MyJXeOkIDQNC7D
YBNb5V2B1lREZ6nBsOGfHRihTy3zLfl4GVQy3ZH1GI5qQJ9paCkzxr0GD8mIjfQqP4uVh4U4264z
evlt+mt4EaS8GwQ2Y4nQYm0qNrsVPPisUTVgB6xyc/XYoFqXknJHbhGxcMsY5eOtmBn7Hap76f/c
aUTDiJW9F3zm/PNeVrqwco1cre5YewjMtgJpxo6txMKvETqxH9T1BlOGGTsgt7JjJOD+/D+PV2NL
2aHgG87qtLPOueYPQxenq8euWpvqcMP9IZev48Hi6NT1gv/OIHPNBWvOnDPZvUIafB5a3hI96zUd
lqbhoXte3SVAu7qQrCrLz6U72UO04GXbZOX5JBZs8BbC6tgrlLmn8vBGpCQlaQpeGweCmvxDW/4Z
PtYrtBVR3cbBodkY2gA29jiniq/Ii7cO5FjMhb5TGfWRKsfMx6adw4MBNpyfNhSRgBNq+KbLxfS2
8uFo/YVC+u7+4K8YlsmlAD6xNRT+m6kDtHUbjQMidcE0eWI8gKpM5kWNnP8k1GpV5TnHBd/GBG1I
VC/l8rwz9AETsYwe7jQVeHHN0XIJaMXLhq5dIWvjqjp/F4elwE8m2vxBdNRl55FZa3uV188/98xn
PLAIG70r81QXONohniH1M/RSyEVnn3A1N0cKlhPf2B8kjIyuCgfwJ+dbXK0JtPPd2T/SLCzLwc+X
L5UEbaWn0gBDwtLLUe8p5kWCfUvnDg2hIrimRQG2YQ3YlRVV8gNCEAzjo8B7Du5rjZ22367hDeAE
Qg0rcWFpWp1Kt6Zk0V2HD/A0ApdGFEK2fkBJGxU5nt81d5NMdoD9gXMnDefWNZsYH2c0FarxouCF
80rIqwURvTxdzFyr4JfqZVKa0Pr8Tck6GH7KK/kpyvYQN2Lp6CbPyQegYIcw+gB3IX59omL7nqjJ
t6hG5DTBZWFc6miRqd3j3utIf3EdKfhbrNQqN4Ndcp8e2acRcdYdZLQ5Nb2JsNHx0ha1H+TUu20X
Ni+4ahZN5lrxtbZBQbQg7fikZFtgUaHDjkqsiVSuQrnfaN1RS6poYBHGwReqZn6MKMWCapF0pl+E
h+Xm0VWosh4yVdl9OmgYV5Ygx+GKacngLJ2qE37W86czJ3Z7NaXxgaRV/JVV5y0kfZrkmUpTCAVP
b5SVwjsK6UBr6dgCMHK0hW8WUUEsYqL91Z2JejC7RddWAv6kitx0XeKW8ipWi7oisYIf8l7a+CFD
VPSmda4RlKW2GsZN7oV/gqY72JeL2pXtNVy5SLqT9ShegatfpDgCLDI3omrNaITg2UovRKjr7/rl
M8hbDX7cDy173GTgais1dFQKMxisAkXWtJLbkCUaWs4M/zxu9gCWwMIxGlJGqXt2XjDqqgYjAXoy
RbdY/VdG6xkoTnZPIFwgT6p8JZL9H3MKfhk3yLHzQhOBerhjlYv8pIcOHOwkKzajktXoaTOHnzf9
gZa9vYCSLRPZcJQcxdiXOuQWyHBnGupoozWuavBLxl44J5J4AXwN8Gn1lVRU2zwzgelCc/3288sr
e2mInwt9dp3mGIQl3nTJvwOKCAASA/h7JCbHPZw/NchUHvcqRbBePHD9LoeONdjL3vYzk+gA0Zgc
S3Qf6uZKz4pr+yYQL4sPWHji1k0hnGNK5g7YBeL+b+oFaa/9skSFGZXdnhUcD7keIisuoOhtDsib
P/DYzfsQfowsxX/IFpHUmf8nYpqFIzQueRWupIE6entjnsMLwChSy0KYVNV6M4tQ0pqBPnVR9lAf
5nWFSp6V7feQRJlP73cv9w6HW6bNy1q6rSqnoXsLkBRB2uC5/zMh2dVdJmjs+gTLMRwui3az6M4p
kE1/NmVgUUcnf8ZzgNMc8aDgRTV6vUMTAEtm2iERwF89Fmk/lvWgdYY4sZJf86n3yYwXFK5G1vbv
VBvQee8fH9NUhilaF5zo8cUPTTbjNNfavluqwcj3QX6YAbZTRj7bIVYNpNwqnvPBQT+7GjjV40ep
MDzmiZoyCN4ViltIeKqVJcwI1hv4Ee/Ozgv8Z0fqz9x7NqPissS4/kZ1y+cOemuL3FQrXAIVMxa9
IUgzBate+Orjkaa7bABbdRmHmk4/xm6ORPjK3hYpaALIym8d9VY1o9mQppfUnzcI/bzSxMe41AG7
QoQO/X14CnvU81+UiaILpbkje/doyhyT+iemv1cZNnkwLKlfwaRqzCXDmdMSkFDn4weEg4+Xkt4I
hpB2/4RnwHtMoHIoD+kJN3DiARC013vtud0S7492ZWKnh91jWE0bx2V4diO7QKNX0lAdhYCXLlQH
d0gBdCvL2cXnP5HTa3Nt9XVuwgX8+oS6OTJuf20qi9QMWApROEmu/BZEsUZF7Kncj+4ovZuN93TS
SF+AV/VNaviINmkyoi0hLVbj24TnGNweOA3cAATNTTWrK1ieuVp0wYImJb2hmmpwY6bBaqevxyRR
J99Zoa9HJoaVXFIrmZthw4BdtTmAgC+bGR4YdkM7MlBdCycrOv7nPobXPXj9B/YMkx5eDgyNtvop
Hk0QRFYrzMmCvRFbitzg/6K7uSNeQ2ugAkBYZrhFbptuDS4MEA44Mo8aJ/O8j23Be85ZYSfhfh6W
G2+nVMareWrMhtW+wmycontCvIv4auLoWmTc22JJNryglFcIizP+gFsryUAp8a/PMj6mvSVlLntJ
NHRO+EF1VaHVPz1Cbt5Z2yysWP5r+Mi4s0JlXwft4xlHCF4gn8E2GjrxjfnayUiWVljvBm0f4o0/
cDqIJhW3PCk25w9DiGkJXgZeKiVxP7q6m6bg9uC6e3PXL0U4J88HOLHj0n5d1z/ZlHpjlWmA3vE5
O044kE/YvEkqjT3gU7b6abJZ9XmjzgKa39L8z6QynzBAkT80puqLakxm0bIkfvOzQ+1vn5f6h1FF
+5r02+khKNX05+bwCVzho4EkZyZ/kDpSwQ+piuqRD6EG9rJyBxrZO+I1lsiHxGF2/hCW4bX9jcjN
3mfhbb/BahSsWpFOfoqhYhlnLDOtqMzy8mbVfaSOEeaF7JlF4Dhz1Xhvx/9cbKvSGpr4a6ci5pUw
dnq7o6r0afJWEgWV88Z9lm2xFDoYORPqKPuPTQgbiNF+pohV7y9Ypcw/niJamJ3Ze5oH44IhSaSV
jklJMnYPXLw2BSWNOC1BjjA8LSxah1nebrxgDSnZZGQJFze3+gVL7xcOA1caH171ELS7CcgaUYmS
mg9tLuZ9h9aPAd1JO9xCCFawazFWuOr+o9aCrIXVurpMVsze1K2hnJ0NXSHA9aiYskQqpi84v7H5
KODNLwLnM1vwqc/j5MO/zPWxnDmHrSxOM51G6cvjannzmudVvKivIdcV/9NpnjRUHBHB+5fBVJvl
SV8NCPbAGLx9N4Ld6zw+ZNdKJmFSKAN6vVwYsy/3vtS/Q89imhur5zesqHaQPy+/BAbtZRYW/IG8
KxvJd4uKuGUQwG/y8kUwPgjGtQ77Ntf5aT+Uybr/8C8+xkVdC9oAT3ioMuY7Fe6clclKhDUmgYj5
p444u7pD6Bj1iaiMG/dVGQjfsUQEo36w5dQddAh8JaJoPrwyiIh3ON6PX3XqXDMxJkkeyg295wJS
INvlJK/jMCcodPXAnnO9UMbWfbQE+UxSsZSR/Yn5nYuDvcG7FX/sxqj/tWx460+cYwRxKXgnsMO4
i2Zsho7LgkAarjYRLxHFwDZ+7d2kzY7/PcaYkxyp3/cyUjcV/EvcWlxs7gVGlLc+a/msLdjzCp39
ba9DX8ygIjIXGOJyVewsNc503Uy95da5kuv2Cn3FTqSwkxkanQ6+AxYSeBs+leWACzCh/W/NkGwN
1LLL7JD8p5XaALh6+oUvdpScmkaoiIDJyxoivIVKoIz4QWECoclhivBTdKDzMGwefACNrXP83ZrO
XZGqb8v6/5QkfQcTdbDZVjJPkUosNQf5PX4r2a84EcPI/DgKvEU67k6XUPP0yBxqRXQcVmogSut1
DP40aLkDVe0XN4cQZDccuAfDhHQ3/U7HVlPfC0uNrZOZqi87rbGYr8M6xDgEqC8GnBhiSZhO6nM3
DXrMSzitXSf4ypJqkBEte7oAYY28C8+mOE2dxXAjKBAde6URqD8CFGHkTTZyET92WrX6TRZ6QBkQ
OAlFUUXF/7ap+Y0Y1yYLrgOetcdypzUWyUP/vHvtQ9UQvtJ3YZE+lo6mtzy51BlM/hQy/AqJPltC
h3mgvS9iERh2yN3SwXQIAPlwcmVNRUv8GcdFtlIFJgRjUPBux7D/kYYXjpChHfJk035W7IhaA4aZ
iwDq17AtJV2TqHxUm2j9xY7h8qYDhjuK/hxeTDfLT3wKAX4Udw3TxizcB5q+nQ+fx75d4MxlPfgl
6EuiUehrkWGx1fhkcn/QcQ7OFMtKw7orrmITPtZa30Q+TN+KiRIwcKI04NMLCMdsodXlpATAMdsX
GNG6ALdPLqthg2OXF8ZSfazq6ABjQwQUaagmbgDqyQHXMFthMM6e1Fn5qUPamP5caGxVU/0/TAao
VQdWzpz2UrC7EsvzGGVG4KEfM3fis415rbk2n7McgvEfa0vE8k/tk7NzJ1pCjs0gudyCq9msR0jy
90NBiLge/eWKEOGlpRKCCDPxyUrX5RQs9pN6dZPjU4pCN3Ryk5DHxabkLS0E+J3kN10xh6xhFA+7
zKmL44eIBOsVPYM/AH/N2NX4bsSMbpl+Hf0kZ0gks5bjyieoL/qVTi1kbxfP3xSWPgkXZLlbl74m
yevSWstKCroGu8F1fH8WIBrUzOvo1WEubrpl7vCPXKoZNDW3xNRpKGL001uLgEqdwKKekhNpnY9Y
sbg8qu3UF6HUDaGJVS6/rboiuInW7wjGRoyvl4mn3ZmIiGIHWH9Jj+ExkKILCtkvInLdFKv+jKN1
6SUXCTYx+iAcqsqXxWRS551Xq4of/0W93lKKhEdNgtFTqnNR9xed/7vIx8PryEvxSSp2f1SXtNOZ
CtjP8r3GCjolHbqrpR49CUmkKFFuycpfIri6IJ3Wjppu8fAixaGWX42JWyoywzhO0SAkiOGQoGuM
DNJ8fGruxBCHn+bmMLP94NAprLMkK5DgEY0Ir9lco3FZhGk06sDbGlWxC7/iAqhBzfbsZQ8QWId9
21Uv5eDxzIm3PsDBzRQhvNsHP7t18KrIOaEzImV+EyJwiUF0y1cJAzny4gip1xcW1jLUUeqB3wtn
cNGLwlsb/bMmbcF2htnOvKDrUvtVcLXHrB3BXYZL0hybWctbS2mhhIJk6ue3z9m60QnKbxdhlkjC
QMdvOX7O5b2fv8bijTSxDvNwxu2uqJxYh3X6Czh0O8I0JH4qvVpvTKUJ5tJf9PzJ72UG5gMbns/4
5AzuXX0Kz68eRniyDlmSwMGw9DZ4NQKvEtHOwQm5fCRZLV42OhpUHPHQllp8thRpr+RYDh+1A/Rn
OtgQThOyH1kC0i0gUH9FoLmlLwjNm/R6XFxIbWaVFMd92GPbCldIH4rl6GWuQyRsqTa7yFc6IsK8
Ygcjq1AoDmp6PLw9Hhr8H/fzdDk3I628LrKtbm3WrmBmEeMmP4gpm4bXWoxj8XxfYt+r70DoCcyO
NNxKz3M5LjA2f7buUIqF9TH/zLeMLMfiqONj9vtKcEQ7kVPEBVHipoI8JWvhtHushU2kEkO7DiR1
Q6gJ4bRcTs2bEb/tFIIBh5zbFTrBzMj3+Wo4qnBhusnIQFEevp7WPh7qYz5L9o+dHqhfTyoinY4a
RHsDJOc3GoOSqjmEC3ncJtPP1RTIIBOw3IHUJmSy443jsoPEkUrYmVi4sCCp322c8ETKTi0+XXij
os6UhSFX98ZiNc3UwGM3RA3oKho61nFaBsFP1QdD/vFR2QXRJXAaZLWS+1vxO/AtuJGyygO2iE77
9f+6+atEL5nKBMIfL0WmCP7wC4HTop6BWFHjmWG179a7irWoEhhLWImoH49t+VzZCzT8k5lqoJEB
X+SQCmKMVwf7LkDeujLWzxCSGCZKlzTAG4j7spheu7sIAxVttct5e3UgZHQ/TIpwDOXxabJ3/IUw
A1DEjAjhKtmiRwORe4d0pGgf304atWG1o7cuF7GRw9LmdrdyRl3kq9Pef/wWlUVZX4h8tJbR3JoE
H+1KLf1cwplsNCtq6qdnIFsFUa2mg0GWeLpo3QRJrdacWkE6AG3ZjtqMmJF1MbakQ5+aF5Xd9pyf
OvC89VTNmetX1eoVjvLL8qHNtllkWUc0BB9nfbyQtD11A4jVfnTiqQC1cSrnT3LjVjE23KaA8al3
8HWyKBnNUxLichF39TqxKDmPnhFNGFVaMtUAiT1zbVji3I6K8gtguuyb8uLOI64kRs1MJdEYe4U6
I/JXwy35286pjkuAiZ7vTOljD6EKJTGvOLyS1Hij5KFOZ/cyCrOmHuL0mE167L7+qLR0iYP1EEKl
KPxLbC4xy2GzOdj2zYfX3XMJtzJf8W6gR9nJdn8TZrwazd2P6YjrY8M9EWeSsQgMjZWxFQVcjrtn
ZUsh9Z93//rjAoaj3oFlDr9K2BAd3oQIyFmja33Uz7e0FuWbv/2R05rhY2ymdbflTKGgRPT7tyh4
zoSDfycwegX1YOhlBRolQEUldCnuDdY55o0bQ5wjilYjNKcKtbfa4vU3ETRUIv82DuM7iNMKjL4X
jZ/M5e78mfD0l6jmBRrsM+q9Ij+pE3sNk9MFs8QqVvnXdQhh1ZMR7pJklJ4Zct7JyeeHpVp7Ld8h
pJrJmuwC8gpT7MGjNtcN6/6jbmG9e67VK5mWZJzd9rK7Bib1gCSUvfaE4lD/psFJYmtXmhCoysXz
BI/HAZWwKeX9JCmaGxhCNm4shokxih7Pt5izkVjVQqCYjrw04bF9UF9cE4upBhYTboLMPI9WQPnM
8vw24Q5ZXSPaUGk8pt/rAmaI9ikXxmjThqycYsXSqIM3wPxgqlnrocuf8YyG43xrzoSyGdmLH3DJ
a0BUbIMIahXjRxAU77ub5knd++Uj21/CS69PZNWzRasuw4eKpO5zXT0sCuQ6ycyszinCjV4CioMA
VlwgyLuCyA3VD+EPg0C1Fdu7BxLgVVPfqCZ6t9evus+tR0R+lnq8bnLn0PINFxKFc1CEWKlEVsMX
5XibaOCfuAXkCW265fY1gkuXsjZ9/KR2Knc+zFhNlIqyVuW1tq3EkY24zV0MSc2oOrEypXHnRudl
70xmre+Gb6/4qp1HIDyNQ7g4yn3FORszjrGorU17VANVmV2wjmRiR9yUzXVsS23uQTljSpZ0lzSX
lYgZOlGX0vDF9XloK+g2Gk9OhXAFARvvq5qH0YMcSx9yuGKLQPyLOLTybOJ9Qom/NFAveokdyRv7
pysWYbkUS+bPYlQmZjR08AHwagB4g/FH6fa6cpQgas+uP+lOwlNzTjU2D8QrydaKSiHtb2sJdKn8
SEMe96VDJ6OVQMcty0Vo1ALKIUzO3laZ8IlHZPfy5Kl0pv7miHITFe/IB+MwmBC8kv2WYBSDgpR9
47pnNXenl/+GDEVUQuaxQ2F3zsVy6/3hzYcVWDT6tm9fTs2Aw/ZMHz/6YX2K4vcPODFDcpptrHp7
wmwMsY7cXqf+8BW78r9h5oJYKNbfFswl68yRIi7GZRjkLYgRQj2ZvOzzLUha+65cn1WTKf0h/am7
ed6U2y+NpONbBrrw7O0ffJKdBYDM4CfajKqsbaTEhxC+25eWP7CLUzXmOWed5XeZayP2/lCKxDXj
CzVz+C+zqGXP+E9JAhW4yZkqz3O2aAaHsKjqZVzDM4FmGCqtPSA769mGXlstuXRzaVnyd1gF9mbo
dbfRC4/f4Gi9c+Bs0YDUqVAFPsf41ocPI6Zf27DcSstOgiZtdO2z65aaHYuFHiOpqi3caDhr9ZkC
kWIoX1RyhpoF8IR8Xm1UmGH8csC9/IRQEFezhEy34zXQYeUkrMUKU2MrfetgsDWFK0gy5wRKygUJ
HR6yUh09cxQDpB2iI5ZUPV5Mlo/UvpU83Vqpmp+r904bC+5d3lzKQanu8TkiMAHvm2gakB7B1EBt
aLxjpugqOgMgoJxm1mdt3g5FtJTv7e4SkQAX9vDUFAY2V2tvY+J66R8MphHywcqleKfX3P1zjops
WybvIiNJ/Z/MQ8+f46D6HF2tf3qwiS0Auc/rGCL4Bzf1qCyqoAF3TKcOulUgnz9LWc8GGlVe3Ug7
JTPmTTX39wN7I7QhfrvQnEaTp4qde8RIUD/ywNfwqL5+sR7+xNH6zddO0zgyhzX0rTw9PeDzqMiG
PJZgSdCVN61xO0BDGhttqQEC4Eu9a/d3HveZszIHbvYp8YVrP8E3K7grzgCOIpQwfK5LbOU/yqdN
J6b8bLlvCUqAJX2uDBn+5yrz4aaBbhVNvVhZGfxwU9tbLFyxHF3icqc3lTov0JPugr9Xg7/ZQGdW
6aEVgWLmn8UZvkwR0tzDVumzSlhXRCjFDRwOnsrLk702i6FWW/IZoCqGVGTTDK5cjzCOMGTr4Pid
tD+1tKZ0EOvS21y/a+6JSs/b0fHLcgPgKLQXZeemyzC+0OGEASmQgN3Rt0BsuG5zfSdvwGnjbg/U
bx7dXB9W7bBls9gvlI56HmeuJfh7iWiYcHTucC97XlcqrCsiAn+E+p9XXXGx5T7Xl1xt78diqH6m
V8fhe25JE5xeuI0GPIA8zHixJhwzlA1N0U4XvjT+bq+zITDL47QKpCX3WC0ufShSW9ZoRSsnzZXb
3YmgjMU9p5fx3ywfFUR4z9B0O8TyBnmLif2FButVmOX6oAlUMkJLl2ZCeQjJwY2yOyuODo4dG4Yi
b9M1zJIxpf4B4BIALRbPAe2KNjpuy0ANKx+gFlIWQ570b0ipfYCr6Q4zfvWJhCtBt0F3YYNZvPYM
TGEV1xs4dE46SK8nKvPEI+5MHGQgpWBkJYbQ0a0QApD95qaAyH4XJZ0/DxUZKZ+LieHSthXz+Unl
yu1e6ARLlkIF8bAySjdptJ1zfsBoL2/eouEXlVtVvUp5J2jsuSf3C+H/4U9tnSkib8+eGpu831mn
qRqCZ7EhGqK9cDbuDDa40uyu6aN5VlbF7nF4xcyigFx5JPsu98moTSYjKE9lgj29+bMa3D5F2ELM
4VmodQm4FJWgFV5LJH76y5Hj5xBJDOmgwi1z8xCh6x8sBhGWriiQUNVmcTdNz6dDg9sirfwDp4ZE
DtDSE769ibxPYmXeTqBFGGic0UnTcVaDsLmT5H5jErJUqnukltX3ALwzNnoYN4+ceMsm7WJw9ooi
D0v5JppiobPzdI0Dgq0Il79EDzBuZmVt7ymcdbsm/g3Hhn7f6V0biBrQweM72GDNYip6atxFlZw8
jMGHCsW1LoR+hwJlvjgrMV6E6+SoKimwKBuf64yejMPwvjMgk5sI0hOAlOykVu43MNpXQfuzRl4D
cToDq6MfXIReowyN0fba+HaNsQkewYr8PGPiacGpO1jTf0N+1zAzNPKkhxuiRQt8E+FBNKYXUJ2X
EiV4lgoYqfIF938TBqU+I82h/s/IAeKnfbkT5bsOBVfMo8mGMzUUnNkDZjU8sRj3U4o1QlHaCn0B
pQDkqvaW/4mzPxPGnoD1bY0aS/8Sfj+LmR489YzCnHqSOrXxA4KCPN7ciWDx+y3KHHVCujOw+OjC
1Oe1176mhZ7HXIN+2/BbaASltNBY9ks5byY4c8MOLVyqTS7ehpW7GhM4I1zfDOCIBG+6JF7KKfGY
zRMsiy3mvu0AxFdbNGh+P143vH5uE1HcNtKO0mxYjOXyOE/WB5giGhgXDoEx5uJvYgh1y0rOT/pC
qjBB+Kr0QNNaYhB0sunabnXba3XgTf9bQRcme9DO1Vk5xgxiZtO0IuhjMnquw87P5vnNXTxKiN0o
KPtTOpBYeSZtweQucQxvj4iwFLR5PGX7cPgSPTLaFR6SuLNo4RV5DzOR8Md9uXa+DjLxKgmAPc+O
6a5AeAKfHg83sVrgCPQ4YQ2jkf0BonngLVFoo/5sAF6fGezfIGd7cFYy0S4SMS87+ju7EgcIuYJH
fxkEbHbgA52l/FzTEGIyV8J2HlWKUhGsdrj+o0ZVuI1b4eSUtpMVvPoMwQlfbs1t37jmmEvse0N3
YQW4x7QY68AtGuiRi0zLIMMnznv+HsJHL1yQvPIntIsPcYRkXDuV8YbphEffOo7iTH+z/JKX0IBP
1sYSvaFA8RPxzDpExfr2Q+4DNPFP4sGqjTzGFnOFOUo+s4x3wWsyPoVl+d5kBX5434UOXjtc4Edo
6cRvUeJM+OqcX9mDf+ex0h7Q5XHb5jyXMydfd0Ee1hQsQ584Yn/hpcH1vTZg5llzMYEdRUKkHGQA
w2jPcRiiVke8NQHw+QHXrQkAw33GIpb5qU3/BNXs3N9W8POu4K+JGXAVunuqw4ziyrfI83VZ3b5c
FaVIVArsUAZEY4wvRV2EjH5Boc7IFgNuJg9OY+BVDEdch4YPzv6yDPWM+1/tv9AI77CIoJajs0L9
TsUZYebtgpt+EksL0XpfzmwQo3ttIe3OoU711E1N3EfXGmpB7ONY3BZerU6lwWE7EkSdEqm248Sd
o4KVZSOTqkg+c5FwNGeD7CYqQnx8u4SomxBvcUhSUya3tUJRz3aSF/ksIOGocqc9S5qoAV4jc0tQ
Oc8CmVhDZaZ+itAWsSwwzTeeTMAwnC8nY1y0JTlQ1hDMzEhrIdvHCCa4GfhDx/dIrMgBSL9ZyMF0
O8rLWWQXR4Dep75JkX9oRmHgAq/22+DBBXFi6v4SVl8SiYejkhp/4R0ZLodMS9MqUOSuIuKV2cQa
Ptldfft0Ci6z8Lg3bKVJDC4rA9qK+DCvjPMHCeQhEyTLceymqa3C4unm8QUvJxGDb2TfUiN2BBzG
LPPdGgAspVLn5vz/L+I0p6oYEa1Jy61mwJPCNT4mWfOeK3ouVsI4VT+MVJB66bqEDGZ9frcprfPc
o3P/i5K9fU3wQcRUgOphPvQkVo4krYY9GVu68FyeRECZd4z8mz7M7Z4PPKMMkYGty3sxXCGPkh3G
BV5YFtb/7aS2APX5TI5AyuSkSL6XJiMeUN1uZo1pYgfC+EpSpOVwQcxqQo9woa1Tnf5vdXbXYtu4
8K5DR3nvVST+NjCi3/bskTy8WwhmGTB8nn9OAnDhb2MERAXwosvwzh4BE4w+BVocGOrKxcf8XGtm
faYK5VSe8FMXuwtLTpe6dGZ05svhK6zL78vrixOuq6fgv0BhZxmSJMNJIEK2pPE4QgxUINwXwk3U
FOipCGuzMJAIF6jokOrLIR5jJMXz66FR/+ZfMu8ryIF8upGMv+1w4Ncmt43eBANO4LLZY3fHATHk
LMKTyJozDI7pcCr0eqjCOPC+Kzez43FfKcvkzM5Nc/MLxz3wGJ6/hjcDb6t/zmbDXWJJ45rKxJc/
h34Gy4Fd1mWP2HgHL8LilAwv9L5+95q81D5u4J3pQNZLfx8pqvhuA15sq0FkahCCbACkGsBHqBVU
1jFIgZPA4dkttikMykw1HynUx3/p6ItLSsV7Mkv8gxmLu3l+Q8wnbJh5y3bprOLTk+aDA9seFdXK
O2/hH59Z/rkwjc1FBDOW6wM8nH9PV/oG/3jdCjletbay/awjQuITJBJtjUdsd15lRefg5U+ez/wR
ZoyJ7nwgRvFsQVhx493l2dlU9lVmiqur/CHxzo+4sZfysNW9dsvRanQ2IxhlYtDWOFU+e2FSINc7
86/GoDDKiq6vkyt+NDpG/3kth2lC3+a1fXTgML+niacnkCCT88OHPcp/r/obUAezx8Cj80vjHKQN
x1yI9qQGxswFUaOJmbEfRZFL8eyNbZVcMlNpnMFLCkV+p6wWtL6TErdM6OJbXWKrSka0fhf50T8+
P/XOBWosDSK/Le+01GCy4cSW1C0BNv9TUaIuZ43Mb7aeYSNQWN4UuHbRjRHBjRK76qCON4+8PUen
2KSh6KLRtzd8Si72AFYTjxxMY+vC1Ry+r+jJlSvg4XJLLV6yZq3v7ERoYtl0qPyzNRGrx6tRreGA
uUEeG3AgnDITULgI2roFeFrDno2hPd4wpDvbB7brcWChsSkKX2W2Bf94aUqwohyYgn2WSl/+BxJx
U/Mw2msknLzddOpOQrjqOJsjasOlnEmYZVQprbamoyOrzNjzT42n+ilPktccxuXWe1wTtVZqmw4f
HTVIt+uxdfhyxiNXHGWOX5e03QF+m2DprMVKs8fcWbqttmvia+2G+vLONg9bpwp5OqO5hkgtzSX+
gGdZYfn2DgjH6F71Cu8Y3mrpb7Yc0647UOOpUPkzkZ3ywOrTLC+pei7pQadKFgozet+RLopayU7d
JiZlcCoRXH24t5MU8teIqvE/VBNajkhNfqO54w7BKx0zszjhMHeLd4fV6BcbckpMGOTVVmxoKWb5
ZFMkvB8PhJL54XN3g8wGEpRzlXi8jKcaPvCZlMcRDI/rHNqLc3cazhXlJO7OWSK41hNvh/02TAcU
bs/ZhqD8v4ad9z0xFS4rUnOhOFobl/IjUqt/vWUIuoOmqkWJn4ihiUaKCDFTRx/tSt7vZJEUxjRo
iynR02rTGK9xKKBp6Mp9QRlUThdzrDXRzdw3rSpnFzSZjCcx42ZMXNwbq5HvKUExVqTRUskxJgJu
UfIkNrWNyRIWVNtNkma2zQQYNP8uvWoPHptYYMZFRK+h3dGcTfx8lp1n4tf5UMnWhbJ0ztGrFoR/
kXo6sRntoJppfheJ3bUrNb0KWZWrt/WcLmL4HSLzvxwVdQSzg/tiATPBRB1mlGNtvQ5WSpiQrS9x
xQdZRzLZeilPeVowdkrNnGOxzhR012cv99xEeenJp2aF65yPjqabuRlJamD8x2Q+Oovh4M7bxvy5
1kt8lkS4pKdXdPwm7WdpphabI95oOdiaDm1xcIzvNpziH5wwuhtFpA68WwU+jPk7nzGOp9Gp4p3s
KfiPTASAOeD0ZVeZkGpPCtiqNM71U/jh0X6JEZoIlfBNMCFtCZewyxStQtS5urip72f1biFrB8Ll
Ohaec8qTuuqb9gifmoFgrfY9DNe6OhsbRjd3++ZuVA30vOSYtIg5YZPNLErkugNJ6PF+etqsz/Ui
FvlGHwwGyVh2RNUm4d9Unon9wsMBCzuLagJDue6VG9/UOslGdTIK/Ja3qpBiASg3YsgTYSjuPngi
K0tt7fu0Uf+SjPTLmyPqjXYL2T6tZQYvdNCEqZKs/vug32HTrGU6nVAlvVS2M7a7pCSy7dxxTshr
zc3d4++En6sHvE1icYaWL4f+S+aAoQUw3O2Ht3tOv9ZaYi78wELiaet/aQpm9vIO+pHmU8vrXl1a
0GfsyJfIpOxXy4bCbFvAxRhGJUH4ARSvwE3PHWYLDIp2QzLLxuAt+zo9DXT1q2ByzynvJXtRJXx0
svuOeODFvJ7f9EFmz5XdQsIdoKrZuT4ymTuigZOdBdk+oBzSqGS1GidaX3DtKc2LADYwLMKCE2CG
6M+WboZUsldw72tR4WO1wBYjTe18KA+M6l7cKWkRgqSA08Ul8WPdKLQgTZFGB5SYcszkYbB+qjMS
Z3SuoGWuXXO9BTh3s8PFeX0I6S1b1ZeX5FT0+P6ve89OHfgLE61ix8k8HTqmHf4OajR1VnO3IenM
+flo1Lf9TYBQcNTc91HJofaQeon3bUcFTPpqOnwree4l3Y/W/OUeHs1OUSapNgTLAdguAYQ9BQo4
vYcM2VMCN6xFqqSaP/Uc7lT8lpZ8CzxlLmLe6QGaxofzk/ZBp/5B3E+hDfwGqCFtBKaiBCUKFzv5
qBQtzrYyIhnUTaKpVS6ZDugVW/Qt8T9NP5JK0JJR76o/mHi7o15PHXEmcHLix9PwF3m3xh2pPzRV
mFaQt0ChL0OnraztjPQ7xdUbeYlW6NX+P6lmSRo6B5dVatyc5FAVkfepNUkLgDJKvG1vXnocg+D/
7kLRUMBReB/RG/LISin+BNW6j3sfGereITdDZEDSnsbdW33z3Ug6vC1QOyABBRpnogRW+yVyi5Ef
AqAocjVE/f0VW+wdkP7giAdjlv6bNKOWfeEcC2aBGf7IyP0+Cqf5XoiK/vJI9KI/w3rtJJ+hoiyJ
Wc63dIY3Wr/MS0WD+YehjKyPc3QC7sWrjuXNt+RJ/l/RjzjB9TaH1XnaGoBiCKh+8qEdJM2d0dEL
yseoHt7mTTNhIV/T4jxcl5Sgv+w5Cd9eIMi25XNUmeSqkXdIsfEp/w6HVZx4eXfv2i4dUuScpCWo
sBxHvhYjWAWfZQaPfZr0bMnUbW8Zjla97WzQgB7XIILruulzPLjhQ7JBejbqPwhzVaZ4wCILyjE+
LIBO3F7L3wRpfuytLdL/lsIQT0KJjfH6etNFLAb1P+djnCM6/sIM3I4L8d5Iazcdh9pWHp3U2GrV
BNeYhb5OWJ5go/mvmrzGFRT5OtclQ2qBIgfhLnFroZ0GmkCVHZEMvsRMR9SJsjwmxsOzNHU5uh0D
dANmQ5zIiSJZkT5flfqSwk2vXD3LZwIo5MSPLjx+8dHraKTe0z0VynFUHMaHQDNR7O0tIN4f0mzs
jnmdCq5dZPiMM6Swifa6VvZ0Etro7y2yui2U2tiZbyPfebymi6FqHYapdYa+OYvRwICD2RccvdA6
m+AkhhHbZYObofH7RyjKKGEo3/z51C/viG1W+dXLWP/DaA9ykw47wlDUa5UulaHj2VJKRa7I0tgj
m2bn8Vpy5GvV/3nxeKiQxkYEscOCKNPOF0X7fq5t+B2tqQaJjTfA3ZSa9swsILnsp9RlPZKxqYVK
M1DMxG1bUGD5sQbz22ZRngmJSFZo/u4/kAkFETOVetp5bYDhnLWT6QawxJJo/eQxNlQUI2mtRjJd
m2AKu5M0rORj26W2rZUWViNYc4VHcemvFgjZyjKiGXmvdLkyIcmFauANhloa4fFgr33G4IRIAT3F
kWPlSEgrs9nHrR1hF5Ys13k+aMQlQvLhROLjnWzISksADW4pORzjRjUngY9TjGsV9xK0j136u2QT
agODIRy43vXZtMqj848xK3P8TBELhg9KDb23bBEQ4Ko+llXXv6kVdd7UP8JlTm2WoPNX+4Kla4Bf
O16IF4iJsn5wfc8LntsPab68kK1cCdDENVwXpcPh9iLgn4RBxBSkxLgYSAKe0Tgcr7pVyic5ViLA
VsbAkwwYFdPSQ7Aa7C7pia618E9lMOD/5tja8mmfuPUD/WP7s1jrZ5Kt7iAFkJmc3vJldYCT4gZo
7kgZnsz1UKPZBOvpdZlC+tZZFUN1a08qGqg3SDxlKD9+PM4BNuulZwVPT4M93yJFr3/K5OJUHOTs
7yg99WZ68HoJmQ2SUkWLj6gPDOolQOosOs7aifIezxiyTOsgoI9mZ6fzD+zvrfIrZfv/ISLS1YQo
hAkiMSQpWeboc7sgD5ZE4a+ocR+4S/5iOdSd3PblcoDVg1FbpFZWtw39is5zMM/O8zbF2W1srfRH
JqFZWZuxy9TbZ+ZIz2EiJmpBFxWXGmucm9IYtfX3J2VIMY1pc+j0sjvHL29koKdRXTCv/L0XbL/K
AgxwxmZbVIZKL4UNXB77Xgbg6JY9l/9dFUQaOLZQRjxOlZRLBCDmDt6UOW2JkVmfWrgln/UIGTgu
FwtkJn3UDXXfCg8hS6VTSbVzNT+nyQJcNT5vuAKRffW0OJmg2U1nglygoUgjCR+Ih4XtCLH1DdsY
+MKqOLd/VqRKdqJRlQ84tu+55RVmzSSUn/nRMRZjZ7FqLac62sO55SEvkzS4sNU12JIUt5XQMo5w
AZnDk3cqq7sAM68QdBDZEY/EiJkbS5OtiBFO4MM/vPNDBVl3l6vuI5FDHakmEpI6osKXcH73vkrE
wiQUm6F6KeFxQioWRFHsM/JUmjrKlPrsA3a3/Vqdq8Lldfn8Tj6qqPmXtS7BsQoUqad4tMAS/vsz
1UuxDBDXvt5iR3M/ZplUeTIhYY1t+D+ox4pF3xNLr+31w+XuklOtS3t3FGpkOGdzj55K9SPqThSY
GoCriIXun8vsP3mEpAdm/KEkeUo54M050KAZVQU4nglT2Atxd8q5djZtETh4WrpNF1ltGPdPK0wX
bxiZngiQYJRClzA9eM1NGYlL6KcHGVZO24zi+OMoni64GttuSt1/jLk939W7t6SeItWkBc2CfXeh
lFMDYZnvunf77fK3hWMJkzaOJmuMNpOD7oCYfOqdLsycyokb6HQT59ocunXJ/3RViaIJP/2cr70N
aE0fUCyo0LyoWDdgU32MKFbXPUso186ELq4KsOZuupiCZYhyAGWHjvNfR/QKctg9Awy5bXQYjTuk
UCgNKVR7mSsJ+TQx7fuX3AXSk6YFOidSPa7bv52QFd2mOIjmwICAtkW2s7t3qTQJVO4EBpaONFHn
Pn6zjQsgPsYwhcZXpjDgqa7BnDycvgNbXb2zCMnAf3GLpq5Jv7OwumrchC9J8U3X1nZPewMl6eT5
DpFFk2du5SfjN/c9+EmWtdftNsX0c5Rjs7HlpC2elphWVMq3s7g/IprwfwiXzY2goOzvXCjChTzh
4lG3kYyb74k4blJ+uxr5/faVTXnNS5JEs+I9aTlRp8SlsnpbSZOzBVp78qJTEQX+QZ9aKyFx6sUx
6Iv5L29j+AioaYvdJdvalxijTqJYzU6sYUnM285+yALNs1xfweV/boOt7VjYjLMJBiKhVCM41Mlb
o9GLyhpA+uEExmzlKsQ4kXJcGSFQE0hfvHwtgZWze0o2r/tfnXQQk77mj/SQpyyufwt+SHm6Twrm
M/RRAX3zQUDQsqRdj1vs+N6Hk50MVmV7aclxOspMpW5T6ecJeZKaWbAXevRGKOt0Iowpq/AViUH2
A10H6T6Bit/NZ4023kYNYWEoNdbpFfcsHdtYqTGDiCOytfVgqS0fK8h/Wl6qzVzVV1hZbgI+Verm
2j95MLoj4Nksz6PPkvbqRdzcoDxq9SceNS3V79z+xuZcGqyOXnUNfUprEAN5zdUJH2R3/OKJzJkr
NG93egkEt7kLByRCP6+lEgdy07M2zt2YKxKhV0tj5Vj9tdNHN8qW6ClqSwjOZ4NO4cFStD1OJuEr
+fSIQZ8vbV+q78V1eAkir6J8JEgEnGhJCTqJYoSs7XlQpXEFoOiN64wsaRB4mpOQvz/yTI+nykhw
sz3+qn9qOG3H06E5gmfgRRQFsP+m4Dk95+y51DQbBm8LFyRXoRccWuPQDhkEDZMLV2oY1KVYfOrl
cTsVRYRAS1PeEPFJKZQyq/Mm8uNA02mj4w6vt02J5dtGpsCstLmG19Bq9HJDT1EmkZmroeB+IXQo
Tzdt5OPKwsUcJgAxzyU2RX+UuHJ7IQc8QQRi3Xuhs+WrkQw85FLJ2YM+5YyoMg1ukP1RWtUQRqrj
insSKKVRIrEBK9kTxQUX04/01pv8O8CJmPEUU5o1Bmqx+eRgtreIrbjdNmqRAfJ0RA7b64DKf1dP
mAE93Le8dQ/KWyAv6QkXNRjKIL1g1G/UoZTSrp9gkxRFUyke6/3jsMcFP2T8OGyyUie2D9edof9/
giK4H5OZzFc5QUoPj/1FNqWtpIHEhp3FU9/AViAPSOyQwIb+s3rEWymnIHWZx0DMQ77Ld2HV/IvA
LOI6gP3c6nEbsAxtp1q3xNT2L9w40dHi6z//V5n2Z1m56m5skS358Gox4UQUHoH6FMbISo5orvXy
MlxCIuqs60XA3cYlYSPJIVZiiozqq5mjg1KazehiwBGb0QoDV+FQ5sBgGezP81yWylW/kZq1532L
coGeZSqWPEUvoLD68Nnb/QhYnlhgGjIgNV6UKm5RmpBJnnvZD6nn2uoOOeUX+jXKU2znAl4qMJZQ
0qwTVah4VDJ4v6ghbtAJWJ5i3sh/j0dPZexT/e5PWwV2N9ZZy3UqSvvCdUg/KEf6+GPazvqxPIOZ
07R2y6XwACIW/SG16jj6VOoWsqB4rJWXlVHXuYknkWk/OqBSDTLJ/WC+0WwYdkSIofUbDidPJhmQ
TokimU9oouhW2td2N7NlGhqWLPqO823fdSDJ9/K+fw7P1sWCSzfbW3LZLzSj7TR+tei7BhBuY+gM
rHW8hFk0yVT+Pb103S5zpQvaobWq/irnOS7cy5hfKzyJigQ2pSkdLpF3pcCW5GxPk2OIsH/z//mr
PYbg/zCk8u0jVM/K/hew0SU3enVuTkM5y2L3XUPxl7w8DXvsA8SL6x2BhRcFId4ea2VwwGzWEjNw
zZxqcrSANlDdwpUOqYvyXuXV1i0KS9TcplndwlTo6j8EgxLP7MnrNB13StDYdbxC9htuo6KmVLUU
J7jx8D/TtePbXe9JMDfTp3IuLUzIMprcCgAZHwPXHmhG/jzNCHcO++gV9TL6eZhG/mklPhQMjjWv
87zXMuipYA7bxrANvN8vaOR5IbWH8RoCA549G96gMKQLWBqMVTOdfJHU7bxr+MNQwQlW8LlCU+St
edyz6gddI4S3wVS4/qGMZwuvT95qaw6oWLZW0ZxlPrUua+LJZssdqggnfmDJPjTl1zWN3BcUKyND
KQz0IrS/3Y5eyR9Zry6dSVngXrPdsUecnN+7e2QVjtbtP3H/HGX7NP77wjY0zZyk1KyB38N6pFq7
C1YXAJBjj2BnHiixoCz4lt+j2+rz2DY1rlNoTR2tTWL5gkG7cFqBiKpGY82p0NE8HXElmHeX4LjW
9QAqrLi2VXZ1wn7PmqqeeEUkoo5hGlp5I14hMic/bRb30eb2DI5ugsKlyPBy+HK66VZN3/mI5mhn
YwxqcYZoaQxY+Jyy1Qu/NMCLMU1Nk7ibirIyiXZ2O4BAvpC5AzoTf+KFwrUgaayZPJcMep2gls/j
IfPhg0FF2uiHDo4f8ehQybxT4sTzm5mKiRiAEW1zfpMS36rDUGW+ZB/9Rsm6+siMQDjuJv2Rj1Dn
YvP7DYgohPcaTl/We1jAtxVmrnClnwf7nnH/eD/l4ptihtZsuYlklchf4j/RyQF1sXxqMpbrXCSB
mHrVWeBF+wC3OtJbwft8hSnN4+9uWsIS3gi35W0/xvDG8Q9VAECBnaCvgjphvGpmc8ByUHNcADmQ
yDtxyFJKC4pX/IanUOo6uGPXH8LmNaWxM/DxbDaQKsKG6AQMxA0nTAuliHJNXWw/8zWUJoQ0TWtN
NbbJR8oQpE8wj9kSOYliQtYOxJCwKFa5jOHvNl9D0t06x1g0oxo5CIJvoqR/fBhn8CTDq5EXy8ss
LvbVLXHA70ecwgDB3JHnXvG/KlbVES8f4tLhNnPPdwYu5aE18lfGY+hhdoo3zAEPQ/V94tjvPY//
eUgABSPom6uYdqaVqq7kRAw5sxWJDttZfTA+EkKXbicpLUSp6RwpTRk43Mn+7sd1jkjJHMT+5U+n
F20XpEzHLpWfd+jh9daawLt0xB7rauLKxW2HllYE7i947yL6+tsCFWsExNw4EUV6Un1ZPz4RyTPb
SO/PQxi0pe4JgR+9jISNZIT+K3odxmlcuLJBb1PQSVQj8WJu/HFsKpgRkqDD/cUhXcENEZInURBK
S7lAoqZ9UUU9Lsh2UZoLw55AL+26E/2S3s6eCu0B8p60j+ZhBYeDHV2Svkky4BQde0+Y36EALpJf
PID42UFNHs/sMDIslRl9olk1DwXWUnG1UUsd2zYE3+YKVK83BpxiEAykTulLHEqcqF9CXUYUg2Dr
RAdTR2PbVlNYU7fGeWUeyBKLStGNpKJ3wf5rO5D7+fUYKje/2b+HORjBz4v8/onzJqAmwGupMrym
PUh3DQueRdKc+C5Uxbk7ObmXHGh19lwt2nkPOIo2HoroJ08KgFgJhZg3fQwASO+VH9MoZHNjgoT/
pOfPAMB7p6X8MiAZmf9/ZLBTPMuXgkparcNijxde0+68B2W0ftH01Y5OKzUOCiEgyXx3DsWGlmkx
e86stnVbNV9vUdB3Xcy7EnL2Ldaa8IUCvn75kbmKdvAWi0qpr8Qt4ct+F8XVOISUCbdDi5vngq9E
kw/XV4g8nndiWTMB1DKD3d4hKT+KJK9JBMBlYnTqMFOZP158kVqF/4ee68bZwEkHIhTLl2L88hXz
HstMEOVZUqHfmbGegom/tOM2WjPwhb0CsH9FwXe4Z/ozoiXBUk6jeBdSD9EsvfYr8gbkOBaHWyjM
ujSmPMwDL4g4m0OAuGaRZfDd1XGCqqRNA7pgxNMaqNQcHy2VqyDN1/4VhNZlSdmU0HCWNgX+rfUL
rfu7uRjgwYVrQyth9siyqmKw/KYCxWEAKhDrbiVtVt9l9zvGBWe9RIl9Us3OmmcT7AH+iaRyV8ev
lRcOol1i2qiU9FTlN954V7nd4C6U0xvX4N3K34x0xT0gcG/Dbd0CMfJVqiE/cyWjYfZJA5LTDbn9
AKewOjM4FzFStXK/9XjPTjhIrv68FrNfBd8kUosm7lXtGTK7VFyX+HbQTa4hiLxG7x3hRbexHbsS
m3u5CBeFdu/hcOAwemJnSTzorghuYsZbMjRQeL1UtftHL8wNvpqz5Kt9rBQOOJBsYV5Gg53CC6Z7
hCCmtI/kzdxvpMe7K7fvS4pPDuBhqdotLR+EDqagGnRYgyLeTQK94xU8K6oMkaB5Y+QbqC6KHWSK
4yZMnm4ZljRCHA1LD8tU1+6upgLh9xpCyZ+AXO0/0F7aklsG0bNfMLiI7YggMhD4IT4dfip6DEG2
/yOVETXAAwwA3LutXGPpv/XisUe2rLrHioB8QejEzs6wEwem1IPwnFJN0+LJf7ZaVfT/thO4qfC2
v1sfLZ6+lZszJ623YIBfyjoFSrZkhT5Kk94UW48r2h/RGiEyZsxj0ReZO5/lqQ3K9FQ1yIxVYL/G
pUKLz9jWCyA3xzP7z/QnT2u4sz47QItCscid89AXGVqOdFVKXhPEwwysq3uD/iMpK8tKTdQdSeXr
JclLh/0d2MukerkFwP9ysXRHbyCY/CyEYRDfb/7Y9Zr4vWbusGMRLRj9yq8vvAkDnWJchx3NvRn9
K988p1TTILofHblXUfU29vFcwfhLwQj6S6xMS9LuoUNv2X5BePz4t6BPzBjfKxqM0f8WAvOSZedN
vtvZPnsHHP9O7KmAKsmQK8m5yeQK7KEHcGAKFD4ASVI5fym853t4SVG5PlNXxd+SiKBcHcgc5ysn
8KxlFDrkZc+LuNVmAt9ayHCVhzxiGe6vDy+/s8QNUtdd5vdIT5SwmrTuCjpVXp+/nBtZwA+tqtIp
Aw722nCM4AxCj9O+ZHGvHQP/QOVQnL+XZU4nBeCQQblocXUV2oMmyahuXx/BjMC0UJwC1cIPOawX
n5CxnyOR83TmsrrGIg2DXbxQ2LvW2ZGM7UQqaIe/DLrG+hoHsEib4OegtLVQZL3E4ieXo7JAF+4K
ZC4j/8CTVTy5VOEflCJ2XCPVaDOacPO+kb28MmwtLGhDM22P9AomPLgVGRcjd0ErmkKdKPVl/YQj
iMTGm1XTXnh2I1/MxnvPK97wWCl6ZPmryQA7kL1KXsRjYP4WjwM6FC4ixuUEgqnEm4J50GZZXLES
1LEs5980mTWlJ4rHO6AkJ2y+3swRK0uafZjbM2PkvqvGoEeR7uti9mpEbUz3NePm6ES/sXUezAxi
QJhibTtxf4UGPxiIt722DuykdvuAfdOKFK7w5Dd1QVvWTVdWuC0LqoytbLLpsQvYMk12b+R7aUsZ
9sB52oBIsHub17+NnAjWElZ8wMpMiyLdreijcTBOD6OmW3eQ+EVhTiCj/0kirzR50KLM0u7fak68
vswOBvgd5hJ6/hHCIT1dymXeDwjLlPh1UXLVcZ0A0X7O0D5zVW8JnPa7Cn1Q/TN1rEC9YiXKYg/L
TQIcZy9KV/2DZfCndcLfZo39/17SIXS84G9Ascv6wwjZvSUed6KgoN3m1EyMnTr8sEpgcw6n2gwC
jjgVCFVr1j0aLzDvvJMMpYq4SwAWpX39RniGE+mASyP6NABAt9vKeE2EWigdKRnc+d1NABWYEb+p
dvu4DPmsXzWgP4hf0MFCIX4ZCQjGfNDVdlaH1EpdGevgZQr9OGs5x68EQHuhb4zDNFW/3s3p8wg8
Bvii7d9TYeF90HnuvDmz6K9tclcPQjutWHyR1/SKkh5cT+xcVsyQ4LwfZFvlqGkBO2ZVgDp4fmxJ
AJFR6yRSmcEwvLUx+CTTwEQ0VeOKN0wd8F2kWO762LNn2rKW/5BjSadn7TEsp4ws8EIiFr4AmGM+
YVxJDSczqZ9n/CJiJdrAeoZq1frCTVshtBH8c23wwPslWgX4YFnnjGnTv6Z6rNgtz2D6a35h930L
0fWMgAgt/YUwxYmc7m84/Q1dFq0+43RZoRAjUkR97SWXNIX5YWYNubq7AuBx2HBYxc+0CTaoMzqR
U0/zzMCELRdy5Zq8mWaigDsJteyuCfYUu7QaSDepZ8q6X7OUFkn7+w1GqbNsFEXuhbsKw+VL3wfn
spKY3turQ773ixZ9UbXc5IEazyW7TKv92AVK/IW9xvdpeFliG+eZvsqAWhD5Xc/D/tjzn9pr5dFX
cRu56ENH+6R10yfmhG+je+KKrG8aSmyrThLZ8w/lla1NjFQOnGJq8UJqHAlDgqyzIBNImeF1jHsD
XYh9OCjTwZWhBkoX8+OXDIjgZHl9GJpCx2zTxe4dwN/xFkfOVAdoXuFlBkvqyMErphFgNemcc/IM
QzSMB+R1KdR2sYGMhOq1D3CpyZ2VfR66QdgAbH2vRqcA10bTLwBfka0RRuyzLjCwbHvHoRLVwARU
M7Iq/1VguV/Wm+6ZRn13i6T9Gyr5YV9ToSGxsp9375wF7nyb03IYHRG/hJBVYXsxvqyQgC0CKDUE
HOhKfzTWQXuUe38D4RHkpVSy1CDZG+L/I0QwLwkC7n126KK2arC2i+PiDnxFEiW+pQKIBrAMdGs6
O5IpKiel51DrlIVw35Rh6ENq+wV//Vt9LeycMrWmAOE5GH3JpYF/sUClA81s3UgGDFHPL4wPZazo
/CGVE68KaW2zpmVyJxzoxa58EmrLj5mlAK8iLhrp4mZoJOc/qEN+D7AJxARf8sZjO2pq9pAnS2AO
ArPbQaoBDJW2jtN8i7Qi0gQnCNcxVVFdhrtZK5O85B2y+H7LmlJT4R7lzwyeqFfa0GX2FHHHT8we
tdbZ33J0a4W2a3crf/+7S5INtXqqBeGiYooBfIqN79BclYU9NI6vkUQ8LYTuUVL0QFpZo+PjFki6
511MTMwfAQ8/XKutlawZ0Ai57R7OvfKmbMBGl9mRZPP72HCYf5scloPnckabqcSgz6JBrO8GbsiH
BipBkRxRp2uSfhcvX8whfqXAo2p3OooLfihc9hSIQcdTktmTTQCFrcndWvDAJoO613jGXcBmvUVR
VpmTdQwZx0C7X8wYEnsr7OIAauBnMydPjnzOJFoKAzKugrl78egNYMPYYJAutUkkmanTyJo1k0EA
ZLQX+T4SurQECjUNWBAQ3OQ+y6ehecghX9yISyr9tqWBlinePa2xVUAU1muCBALvR1+mT+8HlOje
oXGBAbG6XWVpg5FqcyGK2LC0PM2maL0XTPsqdiSKkPbGuyZEpz8vPpeG7LnfnWbfge03+fahMEP9
44a8+/IGjvJI3xFeuuWXYBSVk5zNB8lWsvn6Ak8TclvyU5KOmdaKJ8OBPEcFG1WAtjP/cKrTWLfX
kPpeqsTTTvzMlrKR6bqGSQD3Hf4sf46BW5x+VoBqoLmF82QP0Pju9Qr8AnZ2mzMEC7n9jazkJMEt
ZZCWQBffPaVBdoaMJRfaKR88O+Ntm8/RvKA5V/KZjz3Xw4nJhsbwn97+C5AIGTyvAtTTgYL08Eb0
KFs/VGEhsLCCQAeTZG6Jlg1OXYtCm+b+xaFYh8m3ahRbNYCqX7cc6KSA/+gNfAR3BcKcCDl/aDZ9
MxasK4VoDkfE3lNcj8d8K+YysQ/wts7VLdVlQ4mJdYkeTI6hY48mrirvim0gFQuizp1XGDYOVM2P
toVxahDm0s0RfXnf8xJ+oXqCB6cj/lUmpQ0UQnboWKlAZUZ0ifC7ng7M+xcx6Y5QMtthE8nBQhkl
5JSqVJFUtWbZ9+KtM5vokUs25NwtJqYiaAvBo41qdnW8oi6UWCt7HJpE2X9Cjc2Wtp+LSWrpM2w2
dHVaiXRKDRd/kr6Nj/PscdxGZEo2xe/604x1QF+qNYFzYgbfx8pU+6bUwJJ2+FVgSQmIVdJFaLt+
lKXxlewIELtoN3kTGZ9pvACs7ljFNO2D8ejMSdMzRPchGRufxMMWgqdvMOKluK6/W+5ObfC92p1G
tn/psxldEgTQlxHxtkY6+rfU0KSTpeMW0UMUY3FL6uoZe6P2aDNZUYQ6zWQ45hhhKotBR0SByZNE
7M24tOGKrxvpfcnLweD0lozUoENSoJRGN6CXSdY8RAqnTkuxdTFRSo8liixgnhiYyXfVzJ3Tjojk
oZgsn2RoO2h0BXDVCBAzdvknxY2HOC8TKqQ6f3wF0649NczRWK39O1iBhvAuvk1EtbX7zaacoL8t
54FkA7AfmiDBf5CrHhBpYbEUBKhd9apvRwPpn44HKS5NEr21fn7817IVVKtqX7ONRI1LOTYac92l
UCVwbbDM2IjDgdI48Eg9NBBI+WCf08NWRX/IJAc1uCtEtYp1RnJziymqMcum4aMUoaaudRpY0M/l
t53Ct+s/ktZT79vFdF4Io/zPZ93lw03QzA4oOnS6P3yFuLtAYscsDnQ83nnaer4PsSA4GbJLe5P6
DKZ61pD9k7GoPcEz7YnfdZWLa+QUQhmC3j6nUg1O99hO3FQkfifcDXL/TWc6tUqDgtO8VekrPVF7
LDpyq0yOc4SwYjw/2Yac7ho0puX9gA4ARlBW3z2lcXN0J+f0N4Ht6tdTocdZk4/wHvA6mXHFaDTi
z9S8+Ca8lHlwdY71foYPbUFs3krwRhlrmNG69zZfWNLrwwHjimI89Y/HlJ8j43K2kZpldsyGbe14
TIUPqQ/gW5WbKwekWvD/FwXBE8N8noD9x0uQxbB1AU3LQGiKkvxJKVBKVwMPEEeISHfERwEbhXf8
JPjlH5qyljqfMel/SGnk7oQk05mM2RC3rlq24drW3MSIXzw8qITmUgVRRWuba86eR47J3Depgl9A
sarXecS1tNR75B8r+DPdL5oz7lhPmt9gpR2hOXDo3KeAQFmzRllTt8zo+OAQCEBbwJfFGfMkSYpr
C4NBSnsF2kMNI4jQ8QqN33czRGgR7HyKwt7Oe+PCUt4biaBynE6LPkE77ktOXiTKhXDjVlhR1Jvr
tIfXjXq2gWEMTf3MyMmv75JxKEm9nyryeLGwG+DL8x9CiWkiTDaGHroKEwUfOe+a7eImK18hmBKK
yvHhbyBYiNBOISdQJvYRYFpsz1JiHm4d3E/KGpqMRez57sBI790Mb+9F/SB/mNMqgThpKGKYLRTP
6ra2DTf6tvVztBrkTKn+2JXHQSu1XTXKmfkayKI0Cq884lfz0NTkDY9wCC5ckKbLrWXwdpr5rm2O
Jrko3KbyI07Bd6zps2/YSWR4O9hq5q6UPPThEzxFcvbLMhidpMGOmhk/dlqj+lGu7OKTOEjk4NZd
Na3WuyKHW7Pq62KYFsKJDFrDf/KFEQUcomaQmrR+s6ZDWxjYhW1I5D/VbgyZA6WezQyULj1yAbB5
K8mwC5/U4Kz+V3p0iYekmIHpNxz7yEgFhEjTuw72+SqINZo5YPi7ZR7cSb5pkcNaYF2qPX5pSR1J
2pdOPrCJd6c/oZTmkLWw8Zr0C9nmaargMwf4LX7oktBUCrEhoYUeqgDzXigGdzbsLFf5ghAJEjyf
5B/DOEcirsLmKXRD1pXLx6kDFgMyZ8EL8pLVpnqOv32upAT9AN6VEmf5uThaM+Gq66ipKxmna/Vw
7O0dFIxI9e/DnHaOfOSvOtgM5rXhlPXb6i6pbiFq96TkyS111ISCjOxxWcyp4wvZpXz5pJx5hIju
vB91Tu0Zj6VgQnR3Yjbt/U/pRZ0LKtXjHkWPm9Pi+tXC6El5Y+sW2hZ+K7gRRVE4KTloHQHcqC3b
HCBeB3twJxbp95C2ef0nuARkSHwv494+xHsTEsnByjEhYmKXVHPU/wB6sAvi4XUaYKMGWL6b8Ey2
GrLSVpY8YEsZv+uH4XpoHjLl5Mw49FruYS0eKMIXqTgMcTQcgq3bndIHuAHYiYgXk/vJjOrcGQVm
xVjuMuKCkCoiNXzvRcAAqcmJjLAGOdOesD6x45wuCSHk7Oyw8bsDS4BVdJ9Wxbx3pbXN+jwy+9JK
RD9+LRFgiSSrG4VaCZqkys7V6+rVnKq+9EhvZPu9jDAfoBkfMD8XmLRo9C8rgvRvtm1Siadh6T5K
Z2bS4iQALsXs8NGji0uylgq4EZDZXIYWnwX3X+9pRiwe/haDIT7xOG41AM+OezWhO/1/MFqPqoHo
akmQV0fpQp9PeTmN3Jf/F+OZ7Dk+b6lb1O4fCEAz2rY7bYjhU6p5v6zEGuz6VRFWLKkpuisQEnLp
9TTJmt1Sz3z/qkLbWrxHdaw38onV2Gmmo12xb98bwYnv4BY/ZdJ+m3YSZotv4liNP6D87v7LOaxN
LQZpiPdf4/xj2ysQh018gUh5A3Csxx2pYILBOCwjlte9Yz6dprbbzt/4Tvv4l1tQb/oCxiQVYnAJ
hPvajaIT9w6vnBq851wnwi9WY23vPg/OWSu7O41xWj4g4bO5WHzPBhaiNAxr2JYC0XOB4PySbViW
1EYyLbwxA4Abhbbz7YQVca6RyZB3ClzuhlxtgdY8SkyC4ltEN4+9FZNtK/3cR5UkOyEhMZKINDVm
WNZP4e52TPyByF9rDzHlnbfY1ztQLvVD/yvAzVTQYXyTr3wOY8jJxrnCrMmI1ojvDgErlfg3T9+K
4P9IY5l0TG3h4G9Vn4ZGPlVKADHf1EUoMOuGg4JQfPyBOrkvZV1czUryYhsALwVb4DmWBg2Uo8qa
LnIL8iRjWayOxpUVVzx/7NXr5DcDtMhsI9/L3j59T3wd5I+pv5yKzgq3iPitsftz1dzOCpbZO2+j
cIbgdN8HuykEi+26LjOsGjE6djR4b6x/rHdhfP7RsjBMstxN5+EqZs79n7tzogCsQxjzUEwyN4CK
DdQ2BS/sfitFgvIQcE023qVoEn6PnXEPh53i5suRkhi+mqzpwSwRcrCQpI+nDdm9pG3Gl1T6Vzqw
dI6vrMPv6JLY9hXGicbJTgUsEH+1zVTqVCcRmFn+NkigJAstbKSQyDAAvm/J4rK+fX51tNlJEy9z
LKT6+Mcjq9nEMLc7nPNyb/D1LX0hFEwkHu+nYHMtXn5HCDksJzVQFzhdRjFi5N73PGCoRJM2gbSg
hqrVR9VgyaFnY8dwdgon+JnzaNW/SUGu/18nfAT1J3WI0iCMeCwZz55rC8X7q4//sCSAcCkipO6N
MLwns/6KCw3hfs7AVRmqRKfirajEF2kKJREc8S0OtBESzmuqSi3fBtDNHgBKCoHAHZ2f9Q913OzK
d/bFmzjGn7Yy14glCIGHxo/nqHV6nj9+AYMmlpQ5xNNnIaD5fKXfIKwUioukG5YNFTWOEQWBDM1E
kuw23si5OAlajmqK9Ui/ShHiEl3qaJCTe7c/K6rr6GRmc5B0CH5UO0N3mTvZi1GBiRVjcOd0c/N9
AnC6xpwiBgNQYZxXZAtMA8RDVAtBGkcBU4cGCrqLQPl72pfIm+twhcE/0pP1IF8m8kkL2x5gzTnf
D6dmKb8s/PGrxOYJa+csks3IiJY/J7yFLuYGiL3QR8qK5O8/2k3cWY0Jan1USv5pCciUtF9noNUc
BP8xLDNGHPAjUdeDTPuUZ4DLuANYPN1WEH5YBRsyo7tvdCJM50MnbnusyC9Dit9pmylgfNRN0RLh
q00Tb3wugZDSiVYQiZYSY5y6hjb7t0AhgZ6dg7iS8UOpV3XvGYfCbgbvBYHKQo3UFxGRUK+3g7K7
aEHcz3W5cX/NapSRT0YoUb6SWWyvKTyh+MU/wJHi/Xin/BzSFMvQk48ugZVDAOVgsw32SkT8LL2m
0+G/zL83dRoK6RlN0RFV7TIqFQbjtRPMTa2U7TRTZUnUmWONtk/TSQ7e76gJg3cR3MMu7siOjeyA
rmxE/cMYgbu30Sss+ivLYrruKrYK78DoOSA8z/yT++dOGCypdXXV7c/wn/KRBVWAulpjNviAUHPI
10PBFQxxUZcKfZW3sCLSL2gV5cuR82n6cwLq/R57hmkm5iAq4Nw2N3DskAxMKBisSqEtMfNs8aLZ
37j6z7FgTTAw4UgAv3Fma7XK9fuS1mS1cZcHGTfPbIALcZqOuTEZsmfKhWZcipTEHlPtjO390HhV
WNMsBSaYopCov06ifuX/w8XC9vo01MeOQK79XSOqfO9lkqp8TJey2DSR3/H5sAtnNBHZuCx3SBc0
QVj2Kai205PTtmDxeP0+zSGqNm9WcvV+6Idc6vzHBb4T0e6TEGI1feWKTA2arq+5Bl6WAszKujsd
ie/tj08RZF+e2hYomqziP8STx4fVvmH7JtjSl1yOZON1vhgNl9SH2KXN4O+UZMGlOQPU7mTAw2BY
qTsORH/k8JqZNH55U23UgUaXO7BuRa1rB7OQr4IqN1EnJlj0wTJbVIKvpybGP/PYbv+F7sB9Sfyd
FvFVfn2Wv/Hm2TFIjG+9rq+RektzMGBdWUPmHYpTI782IpOczrpRcFonFIrquvheS1MfkIGquWVp
b7cUKNKtup5MQM4cVpwr+xSWcmpM3BvuhlcwdBt+GwBKcYFk/gjA4h6VQedIGqUE1cUCDyBldLol
2S2T0aChJ79H9pgAQB0rmP00pX6YdQqj+lXxuqAk7OzcezHZ4Ts++IbjAnju03Indli1DJJKCmFN
PWXlUM3Z7U2N75MZPcqPKhYqoeAeOPYJwjasqW7WhS1QAN9Zil43TNTM4JjbdVvHlcFbpFgaiwwV
4u2r9BIfWvUDe3+ZVEbQQAAidAGkCVd/qGo33n4zMdx5TjfivZuq93FPOtLSyKhaaDtj8722ySqq
jqyQy+8AhPlvRkqmPmxmUNXrvnsNBMg7F0GCzgrTm+dy4hYtONVwFote+IFqU6YYwiiZQxVfgv6k
1TB47fBIddGQwhqN+Jew1y8gqER4dm+OvhAdlxS/KrlwXq6PTwXg0KTE0HYXRjt1C4msDxG+FNuN
Qaqw0AO+Gd2gz/0kGO+pWsMVwjR3kKjaFQIU/g1uSdvG24HZZ4dtcap4Zh9LAm28LMiXOeZWPnkU
KsF1Xr+ZMRTo8U30rTYH3cRR3eaM10yB9slSgul+QGJ7lRNDu3t+iFHTFChYwDjA/WzWSHj79mp/
v0JZUmJZde3mAvKqto76eExZG2yr65wCRjvA1/FMDAiR/cVnyj9rJlteymVCttSneBTWU+l5Ptum
alwh/wH9ed2BLgfW53mw2i7GmZNi2BfdexbwEPUNRI8rQWlWlH6Q2NXi9hdOGq46TikC4YfnxcTa
//TWvqSzgjeKTuLn1SDRDbuDJa+XfnIZVVK+TBzAvXvVz9LeL4PcS2UjfWzcGL8kzu8UQYLGVDJK
yqwSbayYaEsYBq4n2+T+CAnAGz8KZsZi775AL57Ieq9HLzR5HINhmw5VvZ0q1aCmahL0TtXRVzAm
6t6JfVRBw/H5DCW0E6OgG8uadRi6rI0qCMFjq5On2DlwayU5r5QRmjmTr2F/HNHBmATgR4n2q2gD
oWwaCP6hkQsV/23hZX0MkCGQBCa0gFwC7VK2hmFb8rozFSSQl9QMXGfa5vsGxSUHWNTes8LKGSbl
s16EL8yOQ3RUePC8W+2coH4syGLd7FpnSemaLjSxFdzmPIXQAUzIOdmLhcB7oQT/piOz2/EARouJ
FTnM3izw/5FdfVxAJqYauupkwkSLvpHg1MxIXbRVbtpDYt+1AEGssoU5WbVLkUt3Ee9I4dgXtiGY
sr5UTSgK3uxO0GPvl0uljN+pKHbgSvrKW4In8MAMAQcuhMkm4przBN/Vq3bhz8G5Y69KpC20m9Cm
WaFionXj+I5Y3+KlC2uuoQs1xOyWUBt+xweCwUlCDGvkaMvkXG3yU42IOcCWC8FU0PLwG9s53fuS
zPnhDDvPW86rJHJF6BJA+tiUrKZtxV2HS9ndpYE7rrFk3MDjE3oYFkuxakC+itxfkx9+RA+OW6YL
WI5xk3QAlK8KB8eveSMZ957cyBLC+re07IbIVeWNVRKNISEj7FKP8x5B0u97Qhl0bu6aiNg542up
0cXxLFRZs5dZkEXgIsIsojKei3tx2RbtXFhIrLZv0cN3159/YKY/zyEDykd0Tabq3NZXZvtL9BS3
WfCcDHTDQowNInj3e0mMpd4XdBiJDjA6dsh7Kdo7p+vYbWx1DVp7XG63r765rZFfL0AIW3J7rAsw
S3zaAihtdAySQVJ4obPzt2VpM5DTFVOMlCinMq8IzvlhRGHcxymgZibNZMpk+IMuWx8tis24j3/r
6VOr06nytCDaE83fUOR4s9XKoYUqM5aY53Jz7pwIcLS1XOriU83YsoG5lySak56c4i/30Ftkulh9
gbaQXiBd/s7hUNxCXGqYI9Jsb5ANOkkpsG29P3ZxDMYowhUHuZXHHTYULYQDzT6p7L+tfdXEpMAa
M/kQJm5JvUMoh9XgKc2lkStbESXB1Jvk+XSyfbgkxLVJ+SXcIe/UtJLlwlcWrpJXU+4NqyfNLaYJ
C/uYzCbeBH0D1SvD907HU3cfJsbdt8nAY23a1OPyX1TZyrx7rk0QwOE9kMFK4O4s4cs+3H/zS9pK
Zuw+P4q7WbafVUGFRh+UaZDyjjwHNgs16p+bRKCYwdwE6l36VOYxZPsBICChFnG6xyRfgxxy+OGj
14ljkLIDCswmRk06tkiBs5LaRnh4hmt5yoZvdxaFr+j/bUEPh5stj+fmI4+fLScJoqHMuvroQ9N0
yCzXOL9qNNoyB/eVLOmUz1zuuDbGYJgwP6mtiilVPIqcRnI6kWu0HcTNrJmLaj2zoKD41H5FNb8A
pxwFEuyshS2fyIfEIzKbF8z23wq4mB0u5qX/tXYZltiu1iKAU3FkIijV7D3CIsnwy8S4qa5QtHP3
28gOtljrQN/HjV5xG5dXYQjO8nQgEbX9tYlswICwacWEQgJA75KF39/jwzg5+nTXHVx6MkF38TLE
XTJoMIV4mJbzytI9FoG5KTJDkLkUObI21QDZTa9ymDtcufjIc53sKxNXsLOIbkbGuwUc9Es/YtaF
MX03H020sBmU9xTlUebIvUw53P+EBspQabixWbuFzr4G74TJw7saeLslsun8tqUVZ+180JH6uC7k
BTtFEc6yBM9u/rJ4nRNJouIzzd/mgNj1gcwCei+dqAI+5E60I1x6Xfxl6cVppJBTCW0sBIHBg1af
9bQQREW561GSuqHKoo9IGceYeAISJZTFg/t0QCt6mq397c+4GBBVeWCFP7kqZ43wNiPdqKca6630
Fdk1R/uX4n1FA2gaB2dGRiKvs/+3epi2Deo0Bv5Qjkuv+KIgwkUqyzuUSRINmhQMUkIFWFhYOu0d
jOBjDXaYSARyUpPsax6xkmXCClODR5TxLuH1dVaM5SPaBJE5QFN3Ms/6HjJdB9VB03hZbgdVNcT5
XsjLBpak0F6sMHRIEo8upcI1wwcjbEoiot46L9qTVI/HeHHlkHnPYhELeXAsYLFotVTvxgPEglri
O0O21YJHTaldoGypkeGXKF0oCdyFgNQmzRhEJboXPdWx1bTy2v50sb6lFxB1XS1vVoU4DsN2pofW
jmx4OJZQEEO0+xSybONLEKvf/iivp7srRwrze4ALdZZCrHmhVsnyBiQ7fO4zvhHzB/xabZiQakfm
JQpsWsELHWnHBnsAcxtwDj05MIrs86IQD2WmlMIjNzseEnrnkepSvNr5k7tjP4AzVibziQc7sSLV
0bKVejmu3iemWXKT9bEdCEenzmV9msNwSVa0DPXsNEADoB0CzJFfqRufFmq4Mozq/I8ymkdyd8V4
R0kSAwyxFOkDz0RjRJ8MS5FUn1mIG3u5PvYN5fRoS2H95PBAfcewU51YEwJlDAZORIse9cW09x8e
xmK5qmbekHhxb7Y/axavWsqcI4gDGtMb/vjf1oXYA0BEHzG0WuwuFmhHq5UY/WMRTSE1uP5/ZRC3
oUlkcUB4+sYmV2yb8bSiGkpIio1F5NxVBXzTpMOhNNlycDrqLo4NU0EtcyN0WCRcZhgJOITTk4J3
33oRpvJApNYQuOY+gOZWJtz/pjOMF6bCavUs5IgmJjFZRqC6jOYL1uV31qOHNdmqNiiIPXbfgtA5
BBZYbGIvKu6kzGsGwL/aA1j0kQdzG/Y4weASmjmLEWrsxFXWVcEubb0cFebOb8KTiEj8EQvwtoHt
Rg9Cc5qNLertpFgh3JnZb0yDRrklfrwSqmyijb4M00deECayfR56um4ZtBET1T+ljRyGpin2U6ii
codwxpDbr63gK3L2ewneIowPFL9k/njC5yDoDY+anXFTixzXxUjQ+ZbtrJ0v+PpP64qe1+hymavu
/M0idaJi1Ph0tO9pADRzSI/ZDC4EJtcw+mdc4RkyXHN3zOuI+35EMHRofNU4idHEeCJvNHKUuSlc
72TSFiq5yJsyxwvR+I95VFi6xKHjfMg+5JT19TJTCEJBu3Yk9bswXJkyTMn0KmF0ehxq0f8WO3IY
zPjB8mRFNpYxO7Yi57tBJYWJ5eH8RZxr1LA/Yhov4doRkD1SleaYqdjBb+Fro0ofAa2Gad9Fc+ko
OQRzouwFadYUE46YcH3UTmQTb8c8zHmP853GPMIiuP4KreDaq+CHCG4QUZF41Hpryuo0pz8RgCwS
dLhZ7Uenkq4kSj8NozXBCeJGXPEGVwWfTxUE254FP2zF2GZuoRr6UAKqsSFD3/KxEGlFgs7WLVn3
n1GIWuk8vZOHlaHgLepFa5c4H8lh66bOcWdekC2KcjQEguFk4LDYgkLaoYFL0IR6hOFie5PcAkXz
rSHfqIu4tMZ4O4N76Wy7Zywnb1sqVlh6FTHV5W9qg9MayiQ4shurimERnHADaXV/U8Uz08kePC0g
G+hjpoRIPAqs/ZSlEXonFG//MzmrZ6vZJTk1urONWc9Jm3gEphzG4GhLBPItjXlJ8RQr7StIkKG7
dlWOwnAOpHVd5lWwExUSLOdlRQASsom15ntvdmpXKFvLiK0ZlvVrJ8tJg+T8XrcCyAsmOBDa1b+q
oZt6TTdh6+3ljonr5ffDQOdzBbVi1TItDHCQn9QKv6+eoieVVTJnIi5zb6j/J/e5lVTNulaMwQGH
NObHnY+4jA6SFyN9VQVAX5+/a6FBjWF3njsf7a8TQ1J58e2Mpz5ti1z5csHN6sbYsti5zdbGRas1
5To9MNbMyY3D+SBIeepEq9i7Um4uS+enM7BF7BIlhXqruP79g5r2+sXxpJnw7bUttmUvYLjuEqML
5DJVLSy4gpSNi9L6yN/JLEsx7qJDIGE4TImb33bDOsQvdzyNRQK9Egwogy5xGTfLHOzK0xWcL3VY
GUOaxLLGWMMoIFilSr0kmx4V1+DJwMzHCx9cW6gLxjH/JJrhilLVaa0DteSjJb4BmSW/rE6492Fc
Hv79/7uucljzYMJNDSmsVVPvHGp5w4DKF42glg2APyLRkNscl9IHo7CUK7ZmSsZU4+yF+2VMfw6q
FLLiSO3sc/gTAlpSE7W547g1//PajdnBy2G7aPy05EZffqGqGzmxJncqKbYpjG2d0t7Ltjigxv25
VBdhcmpo8zkU62I7b8Uv2WSEbBOp1oD1mOA4aakNPk9VrL6tgTGTRZhnl3/lntz1x1FcOe6tTcK4
x5FkF8sRcqEJPjBxQNQUOtYc1HPVFQZTSV/o12mtzsV0C2hukE+2Za8Fe38WyR1MIexIYNj1tXAu
B8FejGM32HURDh2bJbpHNACf+CE9CVGGEExNYz1Wgkqo+H6WBjRVh3a/hw8gT6begmShLWkhL5r6
0+3589mBGlGw0EIz1LuHoWXvKiFDtmptYWfFCXlC5C7XYDFZHNYhUDsFipTk1z4N7gM3abvQPEi9
vHqjb04Wg5TYCxlhp4hsdPg6i6JxYFT7D9ECRhxvr+0+jFH3LUx/dQOs6u3pCNrFM2zwq0NWiEfp
A6cdDxkNwCXHn1U+x5oz2w4oY4Dg/hx18UafTzph1ddwSAH9wSKHgbiAuIDCDm0ityFKAZpe0G8W
ZoZKmVooyF7bnXyMNzdZL+/2xXxu3bKqIe3Q7yKGCkZNO2VT31pgJJiABPv5XIQku1FZv1tAspfS
qmmLFW69iFO65X158NxGGldquTWnOsMZXCQagwhYN37iY9NJCuPomzN0JKspvpAVno50NRUb9t97
R5sdB6xrk2pXGNhGjub03BSbXEP8PFb2927zrtovJk28C0wUiPeYiRBJaM557l4XFn1X2tLzlhuX
pZ2CDwcIKWmJpXzRoP3KD83BOel8gr9kwp41BkWV9Z5uzKyZFOZ7FeAWieUikmx+Ezyb8WhpGUyu
5g6h05FNWo4RcVUe0RieS1xkdbM0BeOFWVsA6730/x34jvIQa6h1oaOvUMC2K5WSv5rv0Ywy8r1i
qn8JU4V1H6Nj7I2QtoN3gZH6akPAIrQaKGHuBxAMnv82VvKUhFalbEf1802+W3AM51oNRwqplKLE
miZQECJ+fieIhAH0DtUYlbGWwHqIf8SmJK/avqeoYA/E9oBB72wi6muJ8b4GnyxMTUsrscFhci/d
Hbscr8Au7PcCehotT5hsWiCMiXWHeyMFpnrF4Jt0eLnaE0co86xSLxYPXHzteEQheJQGvDaqJeTw
WYPz+yfY9BOIR0f3Jpt0VmUO6beKkpiICWrAw0z0mAdjx/g+0WxdciNJbLCZUwwtCAXwSZYMJla/
2S/A0GWxdBst6tYbQg6Sg5zyNTlq0Seo72p2XSPisdFi8SZTDZwjn3NE2M78knWWVaFmzDpPaNzg
kp6LabK2LzmBXuOqqsK01PSIP5AJM212hapkxe2kmw9UfdICSY6w2tmOn8yLTzOPxbfjBBClLpF2
0n0Apc+7R/CkQ1YR3uA0YSeBvF8qMyttbLb283irm6/6G0fN1o/mB2++mTGYi27Nrq/qwtb10w4S
9rOvLE1qVpiGEYJfb7C5ADrsk+7qyDsLwwJcmmJr8bhJxCCwH8bDCX1Bw4xdp3DgHKkeWYQR65RY
RHt16fQ4RT8QyVMZLt07OUGMqsRBtiE6h4lxsNYphSwOa/s/mJXOG4vvrk2T/Nusq9CMv8p+hqfK
MEcXfireza/pi6/742nU3+wRErlVWQdaVe/YpDalXIjit5HHLYfQvjK9DNVuwDGakUKo1nC9TDhZ
yqR0f0MWgjRYPzgZG7TB1FxTJUV9SoQD/x930aSTYaJR2ULeyrMrgnAYDS6YaypntYwmF4ov03QN
9E7FcswMXRUFyP4V5FzIqcJL7EunNCzzN6qLMosVGCqWrHpuEo8HRxRqmQMJ98DRxLUcFF6Qpho2
nRndS+em7ANs0BEODCrxwTLbf89TUhE82eK53jQ/OkkdfYK1g3D/EZsKoOdyHKL5svE3kvGxONJz
haN8bCPa+/BfjayQ8AeUUnPuWX/X0uZ8otHqsCoWREE1nLnOm75NUi2A6qrX1ZnBm2dpDo6/Vg0X
5r0W4cSuklLC3s80Nu3nPzM1qBtsbKWzj2veKEsAjR7/gCTFfWS0Pcx7wFq2sNTs8Mzc7MreaiJO
lsOghzdl9KWAO2G9dHMrvc1NWN2CbCMViw6M3xCLRkMhcpkMVeVMEQOOSTlYtb7MChcUNIzBNqGF
BQCHz77HGSxJmGLpx7r9HCG4kj8Cp/oC9oof6QdyKHt+bzVOBsW+wGZSdFMphPR2BARfSMigFgWm
zHX7nq9aFnxb/heYqnU/fDotajcE+RlVzvDuhRTE97h0rn+HtH+hOT8EeYo85l+kb3OZsIKWcVyh
No1NeEoqFnOov5aBYnU7LxkFBoebNwBwPGiqlkp+8biHV/x6PV2Kg56QRwzOhJ/luAbHK5srWPME
hVDA4fTcQjjiVjgYsvh65/pfObIMXDZ25zIGoNFnkAuh1yd7IwQq8kt5VcabBgisNKORAwRdSIH7
Kezlbm6U2eU1W5e32UPMvjzTBe05AUae36BO9DnXdqoQlROPezCUivo9SXClbaWYpqbW4/ieXAZd
uK/kZIzlJ1P8BfqG/NIV1VhTIHQh1bdNSWd+/okDKctWeBa/eAAr/txlDQH36NGnDJMYsiutxXas
BDuHk4eLOVb95Rk+tHSmgvyMgViozJ6FuLr6YcNSg+pTWHgDGeX2vGPByAJi9d0VDc2nsM2MCY1Q
1Q3BDUQYxb0OvK6haUBFoWKkVAMBy4MR3i6lFXaaeqNcN9V5sVrW7Ct16jErNJQYZaCl8ephO54m
qEkDxNwiCZEnKwY3mlKzN4dWoEy+Rkx86nK1Fjs7YsNebCa9rapIAeLEEfpdVmokeLDBCq/i/YNb
Ja7OLK+BoJYBNiPn6P+rTsbeEDqGQmf6F3Veau2F0oOW9I75aF1kWkosZO2kmX10B1tzTEwRFbDv
beDmdv0R2adPq16LslQx4hDVMc1Iyt263gtPYkJj2IUiGSQP1Uh/yyNBjHs+WiG8/CHVG6cNtZ/C
KppLVAcD9HOm4nlzgDLUpJ9ove95DvO0FmlpXNGLD+ZWgqHfMfN/uCPoN+OmEHbQy1BqdbbOcDUD
Vc4uxQpM+0xj7GD81VTArOsz4Cdmtws4NSKSMzYmr5QkxBrDyYccIat0ug+WZua2nlX5MUke1LAo
yRIWbm8LWyWptxUkRzLDo2dxFOW/JgbUhl1SDF1mHrKqFu7CmK6v9FIfXYttcX1XIEJa572OUaon
8dUTy40QEQxObzBxBoK7qrvolGH1smMEGTXGMZ1D6kwbW+7aM1kEvwD2fmt8wDgM9ceidaeLWCLr
yu0fFW8XmfB93xuFJ9L1Vz1L9Y4WReqGuP8N4fdHgr1V2FG/tyShSffUdDeE+7h0Oe5O+UZDTIWi
CygWtl5QUa4/gdyxIXszclL8lOl4NxzDz0VYai8Tsy6tAFuxLzhkdfGRMVE6HKT2gmVBl109mttu
vcT0e3wclcobTQeL9yC/bLwSfwGYHwZhkIk7v9s+mvdlV+Vz+Yk+49bYHGrNdSN6vBR4U+MgVZhB
l75V05v9YOkl/UVGN9MPmO7ZuzNdkuUajilVRHVOVNrTkZOZS1NhvHVIAeQoPmR/BYEf41jVs4eo
jV7vxYo4VdhT1etj1XDTfkgsGxEpVaigBnVGd4PEm5Iwuo/enw//YiP0XzzXBSP7KgZjTKLWEfL9
4X52Bn1iI7Krg5cNOgyZJaQjZ3d3pXIAlgl+YcnC459wNLvfJhz42/g9fmFa9lZTkvt/u43rQQWh
molgLU0zaEii/62pjdoAcRZGJdGK72CeRThMoQCv+vn08sLhdGZp1BtQfWZTZO9AO9E2tPQYdkl9
IF9riDe/EnOAYIA3McUzJIDDFMFuhyiEEiviSD/UAoqFsI7vbE6lTjGdytSRUOqxqkIimWvxVtzg
ceCcvgV1g5CFb+nYYF+1LjU+SMip3mE7znSCcA4VGTSzMtx7s5FVioyvElJtwZOjkTIoup4vybIr
ev1exTobBLBzmgAR/DePZAF7LCAp9UcGSzF/hdl1LdM4dGqMZfeRnvSnddc+CZVkvUbByudboTHk
USjNiWBrxXxGBfs99mC5FmmCNHAHd4CDcggYDmiJAwh0XqGHATUuISkqdrgSrTick6sFw2a057k/
e8Rb53fFjCWRHf/NM9DRSdklMcPFi+0NCPxAV5pEiXv+yO2ovsmibZVYyMPWozIjT/00zlcvgSfD
CoZ0VPQ8B743xu8aFg4HBZwroGrod64O6wTtEuLKBogb+dfYThk/y4kYTvO/H9HAOs47Z+w/b7lc
+I0f8c3QrwMTbqsmvneXqA7ZFkg4O9eNYDJjXV9KgoAkEpc+Z0OOJR8YVX9aaWIyvZDWILa4D9co
pU6YfqsTUiuIw0qEfQXVhR0tXx/czi+gk+MUPQw/RUr7Mj8juv4dD3f+49wQ3PgrFIhaMg2CX3TS
K06P/LACP5jRdneRU1bgGfgR9vUzAOxUb778KTZlV2Ay1HUjqJER28Y12RsSkUmSIjDY44O+Lqdh
6lMek/w/D/xuMugwBfDy4iuUqVVvu54w1za2aYTZIVx9jkJ2c19clfmDRk1ExMgV9zrDgH0aw6ot
RwyiZSdR9spEmQ1pk04Y9E3JeLMZ4if+vcKUeh4elzqtCpzx+PN0+RZcolxYuEe+4DnzASLvn50e
8qGtGY+Pte5v4LbIwat6Bwti1A0lav7p89CMZvNPgy+JgQZt5TXO3CXdjLYZWYdwyAIjacYdVJ09
82uebdJdc680mZwHglQ++8DyxCl2B3hoV5HCEjrLRK46rjGvNpjS5GKW2ooejNurBTA5B/p4XS9C
gXnU+UeGHOmcjb5NPC0tT8/yNpyBXpnLnPt7/rjFlx93g6ylzAT5yPCyEDAgi/az5MO8U2MYAsbD
HIIUWAFZSJzbt0Zcv/wp5LRrOTtTwAIakxXAc9EWmP/9AHH3YwMHqpDusTqqqQGmyCf7w+Y9gjOx
Q7L+sxXik7pI0llx6VZ5h9TulX4y67kD1gjbJdgilBiw2cczWHZKtlJ2i9ZU+yLVHVHweIvImtkC
6rRrQl9AMcrG3YJKNQmnucbxOEH+SiQwPfyZcWRs0ypGkGHv0ky/defoGi1kMhzYr7FdY8URTo2x
HorLaCR9Nw9CZOPttOYtgu+oIMAxXkiHA/4Qjec9gOX0NJX7SbXBFI8BjJDHEi+9qcvg876u+g+V
7Fvj+3+mU7H4s51Qv9/DXXXQuyfEt/dZO4sJ9FpRnqMMUk5JMOTjGn2vUVjyoExJDJjOUB0FFVrf
DsgMzGrznBXG9Ob6vP51geTZgsexaphncGOPQeo325uK/LXNHDAAzImsvRMFsrA5pyEFbEBbu2HS
y2oVOASNO5/rM0abMGNbEcIpgtzpBDjyElrTsdFCkl2pG1uBiiHpYpYQEAot4D18iQ4SnBNlEkpL
EuBE8cZxoYXXeJHyautwuEvwBkq2fYLp96t4lcyxynpbLNNLfq8uVZD+3IR+a3nZaIC/GcBlFBSr
JtnCJtOqPnsj8kP3aS84EqtKX8DtXdnzgRP12f/Hw8OvuXEEZviZ2eZzWhnaifMp5fUfQl8tIKyF
d0mqkAla5T8pVFVGmUFp0jU0wYERmrtkkwA42jNNlWEkhODDkk8eEk8XGQ5BCIO/GYDn1Jfe0bEZ
n9noiGWrY9nH/LyAcQ7E3Ns/+K91j5uI8IpmAbh0N0LS2UgszVyB06f4WUr3FcJuq3EFL5BSlUhs
IpCnX9/LOpJXQFNk4WCNFoxenkjxxuxcOCYeiobh9qOegdrmfDACGjpFP1/fEWANDn1XyGJVgRM5
f9Zgp5t9Nv0fYrvXezHad4iXsREpKy70u5kfl16yzfRBbGa390Ao0r0/6BgXmfjPcIna9KtV/hnb
kr5i5X+g/vK5aM7GKjvXefVoxAKdqC/zCA0NDwfwRPTPPtvHHbGasmrRoG9wbzMpCu9XOv7fGW+P
WbtuJxt3eFMr2VyU8Uob4uH392ba1I0eom5dy/2NkTdd5gKzvn8vmh2rBmwF50uSyZalI2Dr3YAD
fspvhU3mKq6CZ6juZW5AXZurVE7cBJr/ncsvrI7OMp516Yjyk5WBxvHMkPQV+OlNDLKGB42bCgJz
Mu9lCrUKiARP1RkPZR4zLaHYb+1ZSi5hlPeodfvmiQiESM2jTZXb6CM66CgFeSvl2NDCiyF7z89H
3shVmzvsgj1Vn3rXo22wDYDWG3tilH0/Fh+NeezenDNCwDWpzUwloe3FQxBygs8XYAU6JVKndGJW
dViravs+grOPI7w71feSgKH05K3Lm0Avn6V1hZA24SboerfusQ5QJLt4wD755QreHdfpAJMWotNT
6FwEcUuJV9rDQ2nKFFqDHLXrfeoL7TP8PRlUJp9CnCIL8X+J3/V8Nu6mvt+hYs+vUEGzVXXGtnbu
TTNqxv05XepE5+iJy0zSw4s2dg8Igh1DOpBhyJ148CdPDI06XILZXuYvSavqZYBxA0+79sSv19sg
WMgeqRwh4zlOKq38CJLxQ3Hc2PSXVcA0RJa76P2MBCxnXDNxz7U/DZbDplqfai8TEsT9KAOOkTCd
kt3+efme3a/9nFh03n8QJdnokvnVHj4ERtG27r3LXPHHSAdf9KQza0PcdUJYCqOUFzDjpV7beLlU
qVvWkFmsfBCzpzWwjCwQ8kZhBMEIqrvmmiavLF3681p4Plet4EB9bYgzBybDU8BYl1GfePxANSJ1
hFr3kRQhF0b6ReQ38IlVXAiZioMAa7wFXhdvKSFBGJKN7xrVDvMubbOTvgWTx6dPiT0SE05vRA/4
iXWpIKXMgZ7hXSkupGmgeLDe4/Nswdio3E1uhlmkIvdZ6yS8SnWWh/kyqMVVflc4bipQEaCo6U3d
x1KTdpWYLitsc4juwr5qHqllTJeYQknWzCv1RmbWintSEX/Z2W8lwK3fmvV00J2ahr9dOPOpnhD4
HogVszv+rCJV6KPcLP+dystDSFX5qjNq4/BIOt1MGOCATnXOQW2kAyJH5XCKTm4vk2Llq1j8AZbS
tv3KwaCDYqY2ZmUpEbfNQ9Pkg1NutwDgxbRTPo6s16PtX+wxntkp855/UGA5kLFrwgYqZ92CRIwu
lUlc39BMxOZjTRjdTdzAPQqW/U98qS6qpKwLz/nL9g90r+YsSKXKdcYClFv7Rj9nW/6zTAeSXxqu
DYX0U94Bnn50ZlnY+3tH7rWAwQA/eD5CmWZKVq8oEKvyA/WJFik2Zz6jcDx75DoPkQiHVm+q947J
C8tB0+BfIWFkbbYm/wTgdKzr/COKeS4iyCI39l/uPOxZCNstQ3DzhwjUvaitY89Ttyg/xoPl0s+N
vyLdeyOQLgUD6+M2k1UaLylEUAvTFjYxUN1eVwytIwfogpxgPAr34HUO7H+at+UCWnbuuZ3T1AR8
9Qe+1AwPsfdvV+X0yNg5/RX5v3FIktIEaioU73Mc6A9OqTGUUOlepZ3Ci1ZpAUwq7uB5fBDJSIwT
fRtPCo856AAGstU6foS9aSUz2kYvOCPd6/MI3gQoJ9kkRUtN4Yk4/TYZr+bx7vKh40tNTki2571+
Dn8cws9DanZTFU9kQHKzWr122ztmFAxZSJKtLGFOU/GrJ0VgsD5m2qEM3pSH43AYO0R+zAGFvSJU
FVn9Jlj1ORTm92q/OXyM++k1af6xvXBdlndUqPwDKKgYaGk6qmMHhRH3PN8PvxopTO4m9Qaq/gX8
S2nFocTBa9/Taok6ik9+lWCZFQl3qufwbAtqPS4FzdP8KUEOtwjdTWBeljZwgsQiy0BLrvpndu77
7CtWOdBORNigUCiV8Rg9se5HJQqRnXxusOcqyLF5pAmiLPGN/4dpAX2PBjQWFRdqCqVfvoH/z/DH
rQdnuszpjvEz0eIidbtAimx864Sl8FalH2Ex+J5/pLFCE1aDLEwQRDogBtepdauEJJM01r+K9Jnb
Jeclu55roF8R5cd3bRv+vlFME6SqXW19CgsF8oSqxI8huTm+e+kD/Zu9YVaHGEEHAZxhv52GMQ6b
1AVcddfZHb3Z1oat/OZQi5nNlNQT1tDIbX+IHR22miepwxCvU7jmWdQlUuvrR+jFKz2H/uPh2eDZ
Aotq5WPAGQm2zie+Rsu3tSJ1rorQvROsrtM5QoNN/fwu2WoyCWoMk2Pn4iYlXF1wN6PeW0yqOsPo
lWVkOKCY6/2zuCoDI5Xxd33VAQ0oO53DlKCZAJvfGTzRy20Yx+QmWVwKVf6jLCnk41Knge15Ckq5
KfIpKFbsy1Ix7z1KdxwTrmCOW6bus894bW9k3PN9ABMMn6w3l/bwzbrlj/fOAbuGsyWZWCyFyu63
+k3m3XHTH5wTeLwHLSW3Ce5GcuR92bV5kbpMiaD4AKy0Ny/X+ySB4Pc6+RLOHojHz15COZGPYr/E
CqTbMZbRwhiVxqCgh+ntDzXZHoljmt9SLWEOSH5ht8/YF3wjGgTaf4a0+sYj1P14rZrXpxoaMHK/
PH0Uz4xwzQUqP+TGhtqP+SfOCC1NJYmGZvhMURLBPv1FXWFek9bWeCwr43vwdfYlMgt7u5UrukcT
iYbIj7nfl88GfVyUecPcuj5CroXw10VdoXk7H4U77e/yS3F+hDexWoFiSc2MKhl4kW3FOIQHxfOk
zeVM1wJ6Qm4bseFJsti8LG/FIpXum0gF/GuUDfNanct7ZB5PNJC3M4WcZUXngQT24cQIidvzZBl5
HviwRhtQQUEsTGAzE3DWzDQM+a05c6q5ry9Mdo6afCXGTw1sxDi5LvxH/t370w0kzqFHwd0w4OHP
D8GQJlSmnvzyOVDEkjBmvU8f/tgPNrKkNj1he3Oje4R2pl/8aeqPZ7XN+c5WM9F0LC4VLDSv9oln
9v1p/tNjf+kRD8vXFJJu/A2QWgkrusO2bO5q238JDxQGqZRCFgwH307YVoJ8qpmybRS/AkK5aqCa
QpcuImHAO6kFiiQxM1bWDK5NKcEEIZ4Nc0ym7olZE5Un9R92+SDTOfa0PAjN4Y60/K0JGsa5TpwA
clV2stK1wO4wzyH/5CpyQoY+wC/kTW/pUiQV7zqK6uTShfJhrMtsfYlY/0T5oUnrpdT/F6Zzyzsz
TAtOzxkpClbCIuxaB0pGa0RtwuFkU2zRtv0C/ES2LL7X3ZUvLYPnoBHQEFkrhCSOdVGiQwhW+GXZ
OPCPhAXavbi6VSUDc7JmF4C2+LB1dT6WEaw1OyXw65fQD/TFJxUdIFdX9BemFhcvtTsqOgc9j0sz
5yBMR9IO2bu16nNw8XFMxHQOOJVXL6sJTPy/DdKdvEy3WKke4AgSNFCoMNDRdyNM1mTnAbo0Ruij
iOIl6gUyHfOGSUC6JgsVykxtuch/5VLi6xpC4NaIavYhzV+T7pnPRig/2iIoR/scYsBu+OVzQFNC
f0NI9HW/jywWOZqkPm2eIC24QUWI24NV555Tl0n6FIE0iLme0b5NVwyu0pKq2mKvdBFG0gawQFvn
LCP9dL33tVlagFmvZlY/4FhUOTaV4jbvDcAi4F9mUguCaBPhdZSqQx9Iit/3+8q7XKut1hmRpNP5
fYyBsf1sIgls3vZGRqXPc9eB666CF8lnnCC3PQVsWbsA2XI2wiXKvv7TaksS8Y7sQYPmKezD3+ye
GwNFTovL98Z404KdtqSi1KVXxsjX+SOpIwD1fdGJGQ3SmQLqyLN0IEpePPnE53HEp1+/0uyx3Pjz
SaTi7ChSM/px+/PyhwvuoZtJ3Utwd4FpyvCsqxrpXuW2BjzGfUXKm6ZcCZTarckD5XscyOEIFQbT
DHgycdM5JDklDXZN3kDddTti/GemSl34N/hB+pV5cZf7os3pRXo7Ydy0Wr4bNzNOGpMJ7yfDUqA8
QmhHhcqQrGTdqgafCpe4kP0VT/9tupxFoSivOJHqu4p/CDm2dnubcNhjJWPvt2azvYXDXM61Y8eW
DP+3YEdrquZ/pFsUg8CdDl6wjpSMLjPp63pKpzQ/TE0L2dQrW6gXs4LeBtgzvT2gKsHOY5DryPQJ
B3/ENmiJXSxkQE30uc7QjZcYYdkox6erPpJria9jISjv714RqQsHDzfxY+U0Hm0b3VpGDQlwb3vC
sXqroNh85ox9+loaWmEnPtfthRdVjYB7C3RaPpNH84l2RWVzqnL1xb4Am2OuxmC2WTx0lbHGfoml
pg1MUtP6R41SESg06O4nK8ieJrCWTZYmwVysHHPb18+ZxBtO6dIogGQo8jekx74KgaFk8pgCrJ4n
y0aumb+B9Q9nff7rswLkO2gLMK2n7gUvxPNzyfVBliBYsRJ61uaqCBlvpJWvOBs8qNwXgHOOKO2A
nMjsvQ0dnj3470pZ+X/fRJ1YtH/HjPb9lT9/uoBGJuGxNj3ZlIuWC72kVIMGdzW86uizaqXeVxeW
2G03clUWIcsguD3ZrQCUa0++L04VyGmL9/5pAX81hKtekCQ76P6zbJDzyPAbETZggU8SC2KPxVPp
M8xoEzp5Z+tRAvVcFPs69AJe2Y6wxYPZ/hZX15ibW338/lBZfWrLSfHyQW8xssN6PYl1/Uy3WL7i
+bGCy1nMsVF3OieIWsuKhbZ/fT0VFhwRj/8zkZ5cfzwtXzojr1dxp95bq8MwTjzHUs7kdi/Hlm3L
aXtb/p2i9mmgFD14u+XwxJH930lKYMk9rZYx35Tnehw1BY7leHLm7L31alTzu0a0pXLxz7A7uXbC
1Fem0/0/zXZTzQKL1WqNMqhFlwSUc88l4QxzYd6EJnmbFW9KwTspOeSSRTeeYorDQ0IC6t8N1drB
vnf5y/48hY8ryRwGf752p1chR+USWzAYqc7U0boYPb4lb2QUK2cTA32q6bTICrOc9/4gPBSbHyir
Ub4aOg47ZGeMdzMQHowBVLveQV9NUxStrmDWLDB1s8q06vTjNn/R4dhmEtgNT4L1KpBxRBSuzi91
K+DcSg2/wW02D/9V47LgPwOVU+5R3dICVgeNkUUEky7EytF4xDhIfc1v/OtaBM8EMEtimwFWfSxM
rfcIlj7lb41P4kgJw5DM3/iNJjpwxP1+ajG3eaX9cIjaWsNfjJq4lZLZYIVPY3ViUaVJKkEC7+Pr
399prSQt4glipTlUOkYoZODu4jY4fgPuFZyuNVds4SwfbM1kGQT5mlPLzIxiJc5q/peLhIBK46hZ
6/3URO42M/ufHYlUaQE0y7wZk6JKZyym7AGuFygYyL/iAD5jBDORAvw6SCmUA/oNFEB6eu1jKbik
dNppucYBS66kZC33qCUkr78UOe8o643sH2BjPVI8EvUfFJkNs5OSD9/mDA5LDzoS7hG+uM23tnso
qwO93w5PHOQXDv9cZr7S7IM8v8wM7gQ/XWh+pvNMVleZpnVDbuD3hkDR/xGGkLlztmsq5GsubmMZ
Nn4HLU+UTV6eIoTm8Mebcvw6CkK8lXwKBxcu/0fBfD9YnaDwtUGzJUBPCEpaEfH1+0sEjBjIvvF3
6qP9S/WweD5xIFAS1e4iV6tvpJ3P/AVqVAu+5/QUbgl+Ij/S7Ncsy6ZwPOWqxgrKAW+Im+DrOK7H
K9RdeD+ZKW+p/J6UtRN6QtEf9vJaleJdxD4rZ4wfF2jpT5y5+VdYImkQUzdCIhkXP51jcTduz9av
dQI6s2pvVcjkR/0INyfu152CGlKFw6V2tcNNnrsjYOHrytV6Ym+dS17XF+lqb4rR7SpQTIvhw7N+
tZ5ezbhgGeaEPudIBlAJKZrlTOvRBlGHtapevRilLbrb2df5NSaUYr9oRFYKSqtRUJVljKxGbt4q
yBQOZkOEtOh3G3AhV8yidGJE0NwTLpyavGBjz9gXu8wHQdd2qlaPQYs6ioE53fkIHL61nLgVQDvl
MojT5ZgrKbnY++naHzMyUENpwEj0U7FuddPvWvs0dkhwina83iflnkmZQoBG1Y+VWaX7U3HL4WtC
rexOhQrCywBCd6nAf6bLRa5O8eBAqLFWoBJlYQhnuIGy93EE4EJU/HNZjNQVCSx33hp/U97OY5JF
IJ51jL7p/cgAKvGfcFAV6XXEFyk66VqvEJp0b5opjQqbsuX/P7dcU+Lg2vYVbKh088rR8GF9Nlug
0nq/habjYd1puRbM6PKEOZkyy3VThv7yD/hvXj2g1O8U3tFAKEvhu5W5PtcIZnoKpU/CkhYxJ6nb
3Nb/+oXApTZDdxmPz5EsGhVXbrFLPwg18vkI7bX7gtf4GimG8unl+nghhOGl/7HcfyW4UNTy2yM3
816htunuf9jAFa9+tmkeiz8ZxjWMv3fqv3rt0ClJPSelzp7OtmyWQ5i+QPZQjhkTbtf2we0i/A4U
A7QUItXJ3CrckPz9JVjh3f2hgbHxsShULSEwC3kW467R2/SaYXPXBuSwsRKlZBMiIucOAfkVilBx
sVRq5kjdQit6giAfXIjtVcSb5OmDuaap1vC9kwsXXqA/aRJzVbBrrzOr097vSSWGOcvTy6KL6W69
zfeOzTnIyqjIpPdEFu0L5wDsjFGZEyeLnBsrKeg0m+Yp/t++hpdC6Xh/wAojd9wK8AN2lY1Z+Wm6
RIbwUPoklkOjGVIU2rXPePyjL/8TaGkkQVGhgP30v5yApGCQ+vc4FH9G9MGJQ7AtGVskvZv0Pq5E
VObm16zRj0ZkWpy3fMf4wfFEUnQ+OCptQXM7mXq3TdrUWFGeZSBvzTi7TE707zRg+O2pgiSx+M8r
LGzzXjUrKB8cC6L76Ex/bme9qGJRJmR3q7tDkvV/KLvgUXjqT/Q4tlS8hOHhc1OJ1IPpTYlfYuzD
nQhKLHAgG+j+9cPkL0jSjheBLsxtkUi9VOw6ypOVcEvZ02x5kaH3Cwkbdg1/qMbOVEN12y/1Madh
cuA7IVpuF14G7oBvLX+H72QbCaDh6FpoEMMTDSR3GIUqONKlrVqKdI9FX63gODAYuQINwII+F2MB
nJ1hgvbJnAyYNLCDpgK1vw+SLAYf5C37EFK1+IOsWVOZ7rwsIIynAgirurH9Zx/vQBHuXhimq1CB
Kw5KYRJ4Jh8GTijvsUaQ4lLzKEBjIkqbjLOOMEbPmu0RX4TTKJgnnW3E9+hsCSxq9FWNrlgFKBXO
8hapHqDPDqOFNxVB49Y6RgbxN4aynTdwLcMgqNL3FttlgzE6bewhsva4IEc+5GuIv6J1Mk5iy7XK
8lPMwoSbYq+L+/5+npVroAZdkNBNIOjPIkwkXhX//K39EZ5hVyotEKMK61hGNzoiy04nm4H4cUNJ
hNUxrdYUBteOJod+DMTCm5+LViHQLAXD8nE+4jnO1Z4vrykstY6e4rnKXNboI2kRpgy2XytCMfjg
jM0JCxUdo82YPm9efXBgcmyBEVyTO/jOAmWRU+PfNINxWmG0v/hz08HhHQvC8rA+qEJIkKKFO56l
hZm4BeZZR/bhyqhN3qptNIZrPQlMEUMzkkewVxmsVlAIaSLk8bIP99iOAvuKdLUQPKNhngjexaMR
ZYYMhG02nCMSYOaeS1b0vy5OEL+gvkY7dUqkuH3bDb9ohc5ctY8x8A7WH2hT5o6U6V2gyk45TBUP
DW9Ui4RgAUnYWDJY6NrzyBy0Qbaa0b8LVkgTeptr0QTEoM7d7uHANkbJ7CZ1rBh9kazFmrupwxKK
QeGiRVaRSfjCK6q76jjdZ98lJyg3dO+wEUZDXrwX1Us8R0gRDsnRgk7Pzq21geMJVtBkzpYqxFI+
wVggo/jRTfAGl5f3BDdGE0j/WqbxxTLKZ7SeBrdjxW5GQlya8koVzx/aG3zp0pF/MguVU8iLzrQh
9OnMZKUmyg9XNFDl4g7tlhj8pYPeUM46d6O2Tx+q5ipWfyBTrODuRf+QzSOyVvBGohk6WXw1LMD8
2pG4UyR2MhHrOY9oI1CgBkIkbYLGgUnF0eV2FuZXeXpUMMbEu6j/rUdArxSaj7tVjj8lGIHFKJjq
N9vcGtM6uCQQebh0/38YRVEy8BnXvefwVbvXA8NiTLD5XaM//OA64GAWEz1B+IED6keTyqioLo63
zU9s1hiWoUgwMhJehlJ+xyfvqWPAuWnNWf6PMZ/t73CxbQQxOFsxXQLfRr/3TDKuQDBTnSdVOh18
7UBCTHm56eitpQlNzQOAwg2n3twMHcRke0pS0nzLz0W0JtLUaDAQ5d176pX/ionA0w52Rv43Kkjr
AG9gQMJrJ1nJoUDcmXYjQjaLKVn55Ot3n02UtSce4cpzCTgrrixxLzZdrMDSgRsMvfs/ytyNhtdW
tI1A7FAJGG9Nk6M8MHuHPqUOIsE1sfVcJvTZMfhfViZ8aQ9sczOPVcN+ijRkNaklJuwT8V52ughq
mKtxcN/4B9einAUcbeQM01R/kx5RW/cTmFQDoaTJzC7knAo1wtPYm0uGoVD2z3sVn6aBxtkk/V8O
uMUwHxOn5Ghbq+PXMrQMx755peIAQwsltJvl1nqjNTWBbSoK1G+PeDAGnyQr4sbjZCVicQ6tqrU/
vGkT/j57IN2e5RD5K18Zyu1sp/ixBxo8iJfTdfVGER+/jVDJT9rSA57rR6zKRY7j7rsz/Fm5HPtM
tWhCwFEt9TiOrecu446TEN71lU7KhI+HOiziJAXz0bCnsG4lbEn4tmns93PjENLf5SI4dT1YpLW0
0AxpGujEGKO3wm2OdUKx9XULC77IW65dg0UrUIWSM+fALIAJMgpwCT7MlOmUuIxN8ktjHuFZuM9F
8iBRmHufHLes3YehHHJJAJpqlUhq78e3WijJK3gfFR0wXDcGEGVn05lFN4n7TdK6npNTykAuHSr9
0SRvib3qnxUl12i6ufSSsMNJ9721B/REulAxgyQAhg5qfLHgceQzbeb2xz7EVQoyaNca6jFrT8Yz
TWxRuPkxoMHqdfGfDMqvp4IgIiBe+G8KGVC/OLZi//61A+8w3l1/V1krHxxYY02AlDyScILD48Ry
P/BpPOO9CZCemrWz/Zi+oGHqe0RiRqcRDWFHUxoQGQdpadRygxXdd16U73Qc2mO3XDiWwLXhxkFn
cMH+CmH4bkzpZcD8nGxn0pHKvv6bFcRqFALkTOjMzdiccYTIbcK8+ik9M13Wbgv6rRB6ZQBCFZY2
5g+Lxk9XYzOE1/miz43n9FwPH3o21rJnkpJbvT34sDyKWAv23waUrlGMwaN3HjkfBRviwEOmzLq1
vDZ79y0qzzCeXcWQqCQpCOJZSjcgyukzBuOPTJHrHRWWJV0vkt9DcBRzQqYcu6Qsj27wbEJ0M7Lo
pkVtC4vuGPXGLa1LW+8SrNyABzMVSazhFN8lbF8iBrS5hqDNHeDcm7MrpCwEMAfreCSacAKV4Wt8
YaRmr6ZG/DO21bpjvit2NUhBEbhFKqnrAH2KKzbc3XBeHde6C4YSg4tLydl4TlB4O8Z+D6WOTbDo
V5vaWsURE1FAVN4cq5fyWDoQBGakdIDutZpuMhecuMUxcnAoaZ/4rXjnFZJIBmpGe/8c6xMD1a1i
FrNGcGcvQXp0LXhWqxrJhjn+NePvXsXdvHL9QF/biqrD68bpZcNvaJvoz0Vycmk5EshrZbsTsD+I
KmCS6OczunkPxvlsxNGUtgF8QxkvVfaQaJcknUjYw4cH6ufbbkZwg2eeP7Om8VIPPR2B/f7LZ2o1
8qOBAJMgqXyoOyGWt11xYWBAdldRx/6o0iE2ueZW1ES2kk7HXRY4kOH4ThjUMMw5MzxrrtWZKDyB
Psx2hMvBVVP6+Jy0TWbNPGowpyDeKChg9Gz8SxwYVJ2R9iDjmFXjFRBqg2K4x53q7wwg98BZIxmj
4le6hoU4i/9R4C4MHeam/wJcaT6Yn1GUwixYhcqJ8H10jUqrKUnwJeRmThdYI6/ZCIVKqrOlQp8k
dJy/HBw0vZUH503/MnSO7NpYl6fN02Ddm/E9/Yh5XSN3tngRcZ5Mk5Dx+RmOrwK07pg6ua/6rO80
QWX/urkiOJg75hmXFi30a3fso5CeimUhgrcW5XsZQizc8fMmxbXzvmK56kJ75IbpTsPS8kX7QMvy
QTR3YG6BuqzlFj+9KDyKfUYUbxRSul3+qFTGqMLGsNjTue0Zs361bGsNf4fN3PXd5OQdP/LuH1U/
GGMymlP5u2Kop7IOGqqyEfbEqnb8RZ1t6WSns9RUprisjUZZw5uLS2GFBCDZNx3ArtqVVpr9w9mF
Ltr6s8JiAiRYGcIMQfEI0Wg6SXCgk/Vhvu33pmxD13HqGxzoskzO9zI8LcjRMDAkKP2d5kvBiIc3
mftbjrudv+IkjNFNjIS/an/Bdjf7GQI0NV9LklYZ/I7yDUvZCS0BCuvKXfr0Pf6MZUtfQOxtS3RN
ymel0xBNaI3ZDyytX4cm8EywxP0c/5J4fODKFTT2XBuhQXAU40iST7WQ5pu7ZZ311A2VUoJ1IMNk
Sf501/1udnK02Bkli2FJH5wQKKGGQwjltLZZ1pcrouq08abUW8LdjUVDhEc4uLumQUfZeuHThyrj
xWeiKFAs7kUMTd/sIiXE5D5Mrswp01H9lOXVPFoeB4KBWwhztAmLc5V4E0dkK/apOY7aLo+iZ2EV
ng9fJs9nJPoqmOakcowTnubP//wTc1/NfXQCPscAWDPuRy1dUqfXFadRJI1oaodtnNtgEF41aNbW
/49pkH3t7s87FtRGneDWQCx0ZLie25iiDrhlmbCbZOBNq+F9pmEKXRMPVBB74v1Pge0ULqcT/GVX
c+rdXAXnf1QhQK3J8UPWiMmoFoknyJb/KXgYukydAa8O3FSfn31qd2fprG3ojubEThAOnS6T/eou
sKQkHOmzPlnVbBh4mda2FqWuqOI/SwtsHra5RyyM4h3E2q7xHc8ZzwJQmtGL2JMIJdhCmW5A7NZN
hFBzhP9MmpyDYDoSxrceQ8p0ZkRVmRr7iWEqP9PFgM9RTo0XLpblrNwNBs3qDpz0bz4rG23dX3sr
FNEt4wlSVdF8AN3l7FgeGwMLCExeukz51gg1hf8Z0BAQVBZifZHyv5lk/E3bQnALbEDIljRO6Wzl
CPoudE+uH1z1H7DndB1uDyBLHamDlzZaAgaWOcV29zDRjtNwzhZYWCiBky7gruCq9Y5fVWT48vKm
dKd0ATcMFM7llsKJUhv1+ICZBFQaMNt3LYGdFkPFTMg+gWEMRktTWQFbfzeH2ig9gI2soVzSzFpA
YPE0licElSCISThbpX3xfJqjxNDSvHtySKSvXdzw5MJ2paHtsn57jMO8vhi/eRBM4raVoE3Z5+YA
cSyyV3Tb2u8WFn4Cz4RwBzOld0+M6Rb+RzlNMQfPT5OX4KyNMtVjD8mxXj7SNdhYvGT4HpU8o02x
SnRQXf11RbNpRjB031TegtdqZeGgpJkcbCF6oB23wus7dbfOyxygbQc32KjiXnp9KZMWZriwRqn7
Pquox4POeu3wJzY0ll/iprkw87/S1Ym4oX1lmhwc6/5IHUpnvd+3054N4vwrMgDIWnMqn5gEJcl3
xXGT2Y4/DNpHn4hOaxrnf+f0kwOrY1ebpUp5FES+vykyxCXUHJnRchd/gef/FGQoNrUKYpjZkuk+
A3yyWFVMpqdoDddtjdE3AGnW6e/n9P6a8fSzO5fNJ0RXV1onkVx3AN0cSkvF2dwuN92KCQaS2zLr
TS3EpMQG4MuvWDwQHqkySqlxthM5efzvQgG3emMmsXmcDyLmhfiL17DifQdA3amZdQIsvnReEPbo
TcIHpqRjEWpM4Gk8dvJZEJb6aXptOMj5wbbEsQVuwJB09W6L7WwbjP8pF9ThYfoHJuD9JRo2xfx6
yZ3e5a+46+BQ4OgF8652IxoChFs/DwIf/HWLeIZCtvCbalyCgNA6GJeTkFpPg7GAToC3+pH2Yogq
ywaP24zh0uZexZpYu+jFF7ly5hkj4ylnxIiwXuZnSWxbzqXpKj2h1vtyHjHKy0OFW9uYOm3+bEdp
PBqc06GuoI+q30OQ7oMIvN3YwXyBGTIQdm2qZl7wZt6sVp7eAs8uhq+1LSwvSsU4/bz/ucwOixj0
BZ4+Tld0vXjjtXeEfqaPCLUTSXPz/Kia+03dgFqcSyzp+UIjYemYQrQJlkxAo9TAT4kKNUrgqFEs
uO54lyhDso7s8XFekvjD+fx0OChgMqakvnUD8rk5V6Ko1fPQOUw/DgP+0WegZfxUzeJYM5Nqxmeu
QndaYOt7H9suZ1OBDU3LyxaEZX1ctMw7tBUxHrSUuZF9v78M4HiwsRavU9g2WMOkewcU/hsw/MDi
qsaRyF4BcB5Lms5cifDUdYLqe/NraThJpoomGg630AY7GeIfKXscY4ZNGRL70KXC24uP7oi/S/k6
NgZqHSuZAIZf8buj4f67jrAW7/Dw0Y9kL+i0OVRq0iH6Ywr7uhISaL8XJeD8XATBSUS8PaUp6y27
nPn4QLon52rSTa8opnM4JpAXUJw5rBHB/NaDjyeTqog5eGhAWmZOGNWF2aYSprD6+8hbBegChtxl
+zknM41mnlzaRltfinha64/MEL5c+TpCZl3S9pBaW+YhVl5TnG99S25v08m65x0UY0CzWJSN+fjN
EjZazMbzVtlkkCB/WY9CqKdwItDv3wRD5ku2HdNKnfyhNd94Ce/sUGp+kneJcI4VtZU8KtY55xpD
YpN3uvGqWre3W5F6y3ziE6FCCzavN2h0DOm/9d19mVONoNSSpAQaa+jD3EPcYABvmLDT42pKpJuS
D1EMEu1yu0paV1TW9exK31RPMEH6M4o5urLvk2WenL1xioLBweAogB/uf7Fmb9Zk5FTwJAAYIJb1
TlJYvjxBeppdDMhho2AnxIJisbxggO2L3AGORU7FaKiORK5fd6PvHHwiVAVKgcyRlVzW6CfFfCEL
YUWNdc3XnJmCOXWZybZQeY+PUjyCywrBLlW2WuL9snF6wdzU9E+/BDoVaNkyDu+njSDrlngIgB0J
cGCQrtGIgq/evN3/QUq7BwDeqRV4/tpw2HJuwDQp9sOquvaa/2rqIf498aycyVgfPJmO22/LJxPf
tqt4LCUqJ0R4SwyJDjqo1dZFKlP+JOEh+GH+m5XUpTWkNhLpCa0enraNpOW57dz4L0IUhsyctoNu
TVvNINDd3DB/Tiwv8UeSJZVXvXnwiqz/U0PW9IG/rD/SjlAJN29uFlyU6/w9IGZUgbLHkgl3mIzR
b+ppFim4l0s9QWSgHZBhP/m6zIkqPHmCD536ez/GjMmWZVqofaR6Kdu1JMVqlmS31xvFet4NAbiT
Hu36lLQ3WutJ9zbfU6YcVT7TDLNseiox++Xj8Q/UMXuTq0pSSClc672yXIM2XkFqT2K4pA+q07TN
+6gCjeMLYOTEfXdZzRAodLe3vrEqpS+IGi/6zVavkdlKY3VL7oL1PGi8zxi/6qod479jpbaq2n0U
Q0yEWwTxJEW4nojbr1g+a6sWM/W/nKakgHHFBp0I2VCbfVRmDD5bu+m27opAaJPk2jlm9d/SCO5X
zEJea+Cz6UTY2JpjVr7OwmNv8ec3C2ASY9flrlBTVC7LvK8exVNhtoqZ0jyqd3xBXaCJGy3yTuWW
tGGjest1kL9LGRkZMnmGkQWA5GkLIEv6iCXgFSLkPHjuP66hg3hix61XgQGFV09hbX+BvzeS91o3
a1GdO3TfPw14+k+ZTIjBRDCU9cEvwjtmZ+iW3fdf0VEFXLiO4qNBjgbXS6bfEbQ4nmNtfegiG8/E
XEX5Fpu3FImpQ4W2VOzg5IoqahUeJilg1iY4UjZWf/dlBUePT7vtoWjLZESls0LcJ7GjwnLGIwfZ
Sz+pvEBC0pYXE+y/bHK7mm8AMoNcpeQOEeoGx5i+lppS7hL1+TbqkanI16Ns4WyJAFvy13zuAFuI
NjCrzujvNk+EBzObLes+PSRdMrN/pE6sYOC7gFCBh33C623ciOyBcyZAG7LKIK12FCVIB1yaSm+s
0pS4uD1Yi1gcNn9E998zYXDS4gWR4Zj4BIAAZ0iwwN4/jsfqIPP30MQF4mE5MKVbS6qoHrpz0JGY
pn6vPqefgmdkPofd/83/cq4atWTCj35G8P0CjRREEyod5zCEf0honzcnhq3gv6ihVzariX0pubO8
sgy/mH3dJCJ6k+oqOvTEcQz7+ngcMXlZTznSFyQK+6ZnwE0nOdv0WyR1V74SgJUPgA63VsOYGNvJ
zLcVfpe3SsPR6VUV5wOP6VoBGWWMP/2QE38mB39NXaWVRi9jiIk2AQxJ120KYS1Xp0uNrMQuW0OL
MP1ANEJRrD5JON+6/gRKWzZOzR3kETCbnLtbWjFO+5EtvCQOA1SBMdeelHrlXE7dFcVtD8bd5IH5
2kz5Z8YJQ4fI5DqPxAmbQuzLpUM8YysLj+YWXrVZYwNY+akkW0z893IDmYudiI2VgUa+y9/2eSMv
u/MNCKVU1Ok+QT1jt+0ZtPghjteUrV2xNZKIanaSBr3s8Qzx6LddX6QsWQ6K5uTBCUnSXI4Kh+XK
sFcoW6GPk50V0Co9VMvWuZV3LFKXZYzeYbDoW9NP/bn/42ju/NBK65kBfnmA0JscomJJHevb2Mdc
j6XCzagunVNaC3PeKsahfM0v4aD4bxYPUj90TZNJXVwRBYWwcqlUVn2PRxrKdRzkxtEgeXoiPxmQ
IR5cAglIxLcjRiFozO/zcsGmU4muOKxcmsTeJTmYKKxCXkZSbhYh3IyZ8TYNR4tgq6vBfYSraGtz
vnhqD63LIxFf47Hjqf5EY2tRIhTj0bDv0pUP5BIRYw/M4GyGqdM7k8CXZl26wWvTUBPJW8H/p442
g6+a3hGNt1Z5hnFJfogh7cEBuX6ZIWDTtRr08JgBzfkEb7YYHTsBbox+9UKhoBBEVESIshT885+o
l82jjgyogsStCxnCmilB36mKODNU20lq1sReFqz9qcX//kwtA60cNd5pdZVezqWnvwbVj2t3LWlh
D2BRco/9+qmU6bPrIgQPm41l+qMxwkk3k6EKMiZab/Z2EX0LN084z1TR4jEdDzh16pR7g5ywMES3
JzBQStfilFuYoASwfEWWQMDUvmJDcIw+8ZKPvZlLPS/zghwRl3/37ARnAXjmWUDK3jl7e2GIoY8/
HPpOgvFgBKV9+SBSfYGLaxPoXPZj6niaynX6/0wD3lH4FnDUFnL7D4kmpRCdrCI7R5iV6KBvI8uZ
bfkX3mxbsE7HfzWtUg+FzltOT/bHmGAdGrIXG5Uvo4APH13Cqx/nnrGi2jqDyT5xs8bc+RQfV33i
UOO9Zij28QUatprgRypJ9qFTkP3nYBfPav+b4pGxBMZpAvrMl1gAiWXdA75duWOu9eMoYtMPXGJe
cCC0fUrASgPntAT32OML72k5BkXjTVB6yDfP5tR6dEwnTYeWANHxYJJTTOKVJR8u30HgYuP5WJbt
rP4OEWlLghJBkNOcxJCSJNHTJSHG+Tpv6DztzuECup2i5nL1yMkbZDf8qiBxfTqAQi5V4xbE/M/Q
+EGdKjnH2JiJsw5OAnlBS6NQSk+iPbiov+OBCR3keW5RHUOxcrq5TUF/O/H515CcYqe7jAYFUJjf
oOikd7yCCCda1yGnGpQuc4knlUMSyIOhvY+qtUZ1oxeukZyM2LuxUk4z4NTLPb1g5fw4zEH9sgY3
uGn8ULc2AIJA3OnIhXXYhkyR4NudP9sIFFCrSeLl77lpDsSW/yeCVkf+IAzJPD/IZ3dKnKg9j+ac
ft/iW/vNCY2w005Y/ZPGLCg3+VIAOaxHBe2ZEy0cGbA5qWer+nHd0AweBqj9So4IkcjF3qn6Clum
60kcRHYasAL+9fPBQHICltNLxkeP6hg5bMOkfLYoQESYbq+VOly9Z99+DwWYRYjIngFUtYbYKBDi
Td0oZTqd9LjfiHdjDfVJwWuZZ01kL8fyHrwXZNbKC1cP5S2qQC46DqFq/BMz1b5+LKA7D3yj82u5
xi0PeP5miKR3yAd1GlZnGwAAW1uOHMoaYhxC0AAUs3KL2xjV60xJn2EIZtUdxjSWnRHMw7J+D2yj
UoIno5VLVKDCcTda34gJsSB0tZvuD9JbNheFoxRsW/mKZjAYtemc2QaxENjuUDPJ2y5dX3rEHsMi
qfGkgf1kz1VjX/dnALn13XfqpwEt7y63fE4KvhTM0AduS1VFAuzbb50MEflcs+6tPWp6w2+hKxYW
zSsGmqo+eKRoXbKMC0T6KMEBrv63RRDGRNcAsp/K7Vz5A+mIdUtmTC9QQhV67/xhHU8d3PQIqCKe
JqnJUGn3b5z7Oh0FAw3CYvWgYFNx1Bc7jiThvNoquJIqNw00CE8kz6L7YkVe6eEdKDqLCRcN8HzX
T6KCo8YmevbuvhAInLrmSf1JEB5ffJPqaKUIwIie/7DWiXxqn1eYTik7ktMNZmC2uM8JENEmYPF7
a0yNvYtCQw1mDOHi37XaxlP2xUbx7NhPg4BMfFCuGbqibJZFPLOw+vuJS4apPLTwlGes+tCxk+xj
e8anxTiOykn/9mxsJJuIC46EY8LK9ysjiPmHUSs1Mpq8WRX+hbjRZ/70wYwery2diK6tFxRa2Drn
yhsmO7jvBn+fSVIoh5HGUaq/ppF4ODfF9uzwMLHpEmiCi9DYoC1PLOMddXAQWyX3Kg3JNxjy1M7r
zqsoXa8yGTBYTKAkcT7Nt4PSbeqjUjf1RKx9ew+XY5JQVEXEpfgtQgF9opk0DrQYpXFrm+sreqZ3
Nvpoc/a2p5dlbIskrCOtWVGQSPS06LSFkC4FTvN5xzToSHPcMqtBsYaSx6o7JotKO8EfPSoJZM5w
g+0gGYGjBCCl67csADGa+Y+Ezdz9uLW09d4KSaaXrmB+gSwYtKeO2Yk+JZ0yOdEvYWxXfMI9vDsu
ch/w1O5Dc3RONH8bgT3VJUUO1nlRq2cW9wpuPb0e235PQuS3bJ/iKV116Fl/DbMMpXDMySmyr8ii
tXKWVLDXjBXLcmZ4b+LmXaxvGA8r7fHZdhGQGissrMpH7WurHiyA07Ov7o0aa0tyHX2G506f4+8O
Q6TaH8WvaNdlTpaWL/M2YjuaiI+csC5CC4WeaZfhGgCRnFTXzZ95mknKKApjkvp9vT5scGgA8Pi1
p+zFDXykTDfjXl8jhPz3iCmxVNwvmHoRKwDTH6fMBjo8qEq111/wuiAcDhj+npteU5gvUv1WF8nL
/HOV439WrWIfGAZu9V28Ls2Rn3o2j5srZJfOhvHCzln5IS2i1J5t8pQfM3P1tvqsZqscODPKDqsF
xpzcEER7LLSZKcrItcgEu1TRyJe4+AGlvMyMFM4Wnzx9bxxJyZgKx+/OSm3gENr8HmcuqreS/CWU
QPxOAyX8fTrEiGWlQmvF4UvYJhKEaWtioNgM9VfjSSS2/Xd0DRy8jugoaXaVNX5L8aT95ZwIrdlZ
pQzSouYH01DFS0uNy5wThKDlgat/jr1zf2PFOIp3IgOqLt+RwOO7nknhauQeNbu2v4073svuC0Ta
WmUHKkijA6JcqqCQ8IMmAVVlhb81C+wrqjagiKp7T/G2Er45aFVbgaWWXiGWBrQ1XZ0z0sCDL47O
2ugiFRvz6PQ8aeM1CluIR2L7vguX/v8Fqej1HR14MbVMpRI3aK3CVWLvZU3sGYTX8qkA5HvsCgAp
aKTBpKHYa+b9Pn0OmN8e0s2fMcVN7mC9kebbuFOUWz0q/X/dyfaKELmeJlVT7UtzyxMkQb7RSolS
/mMwcuqChbUw61qrYyoddKuM7OmMeZ0SDwAhYvjl8DcTj1FdEOnu4mflwT72U47gLhWbGC5slDxh
yzPSPaOz8eT+brSkNQITiEsyNjbjDnz1xLsdgEACZONN2kDtZsf38yAZXX+9VigR42LV6xwUTieK
xSEUh1d28Ylja0vkuOzafvN8pImwCUXvkay07+5N1Bu8D9vn1B7TJ1GvK//C+jx2mVNG24RjnoJg
hWVZqWV7cKsYJV7XSQrtYkJmpL232nPpEFo3DvBd0hUqnXUe+WgC9/RwTXwdDQrNkCSVWQLtdmn6
1xc7XboX2cj104q1HQNsPF3HDDPe7T3z+3kD0S3XkcoaWmz9m780SWqN48yLu/PeosUYRVSXgl19
IOGgMnuxaSQjc8tfQInBBm+EyIJVWgC8WZjuumKXO1hFRyHNY0FDm3vZPZoDG39p74slPMKFrpbu
antgWWgWzZ1my6EYf4VePPZFkrK6IeggbQBj1zuA+kkul2cdwKQWBxRpDcnfkYKFumFI17k9RoEd
4ge+JU7lkEVum8eTBmFy7YT6aNHSFqBmS1mPa6KSgKVKPSY0ZdRmCZ4uZ5GrKc2UTlbf2Q2Hd1ID
OGpLgxhA3Ja/cB7GwOcDGryjyyOznm2fB457dtM0nNSRAWirJmdOZRaGfKxLIdWKB+OWsSafOcz8
nrpq/mXZSVl0IUYvNNAd2cnNaNzo0mqpGuTZf2d0WwUADkxrR6flTLEzErtHV76kXg/WBNmPvsDj
iugHa4jejBpC17mKp8ogWdlCyMVPpDQtlWyU2Z2/l21yOrFFTLs1ks1W6HL1Rfdp3h2oFmwOch3w
XQXltYWyephuNguhd6U2aZsXS+W9TjbqiUNm2pUoZEnRgKLovFKHPGomFWBp2f4j1OLgE8f0hdtK
tdJEaJJe+B4ULq07a4qx82pMejCJ9GuwkRC4dWAuNUEy9a5Gac3IK9tVragC94aFtPb1YnltNwSi
MFdsgtnEbhGgNoyQ/Esj3hMywAk+uZKOUZn6V7Wsz9cKtmUdeSJhbfBSf0zI238Fkz8WrqZXIFa3
orkRs8Up1NQPSd6let1hLpAO4dyEBvtVuWIVPnIgc0htYw6ULYVR7o6KHNTP/GDJyqV5uTeyjOka
fSHZmCgQj6ed81IHcda9RPVIRQWv+KlN8HYxGb3PspXUcQ7beNLIaB1lIYQh4tlzsp23r6NUBMBR
T/pChGVUI7uaO5vfKYGowJPd3IRi8VSHwN6Hn4ABF0tsBSpm4EpwTX92bWcMLnSiFNYJaQMsNkB/
ADOupUY3GZ05JAOE+iQLi3768eBdyohanX3JxUSURph6jjxyR+xrk5Xn1Y5lTgvOFKHugoxd++2+
j1na60TGVcm6CS5AwIWA6cm66ctzMq6UgFoCHKVHWqdI+kAYTVIGmEMH6H0uRqyWC5/pORNeiDGI
EGdca0Z3Wneq/LUEgAAxgHPYSK6MUEo7wx8S1Mf45505RSHcFl4hLqr0e3SaVyUeC+vpbQUpMb68
o4gfOctctoDHnn9nsUQDurYLf/lWYI0hUqBur2PAvEJj1hZrfpfAuz+TICggP9YcPY2Ed396L4+5
gPrU7W6taXow01j0RigSxOSpxx192JtIUvyxvmYI9RUbfqZKxXcXa9yW5r+Tkpny5j2FErEeD4Rt
BXYBcjlmBdF8D4W8t4xKu5cPykQLpawwLVRodTJdcF0Me/2N/R5Mi+YKAZcbkCvk7/eidK6dHnqE
8f1V3yf3Ys4qGL9kqDv5Y57QU1GVJylc+0kyrUTFEYCphKYzm00j4P6AdC9QF7vJ8CatxFdyZKwQ
vOK2/P9KvqI3ZRvadfD3YEllhouIV/a6DCIjxuZbMk3xGl2uffgPtI5DgpCQr+7tCswUFcYaDu3g
1QjTian2JWWhdJ0I3/3McWjWdY6ZiJWwrFAya5GR+jQUKZN7FfClIBLp2hTujISWu1VE899Saiyp
uPxPH7PMAMZ0l4bfFYClskE78YxkxhlFdYfcBniATdXAX23VlEdzzlcKnXeH24/z9xF7Mawo/o2c
7AWuKHjD53PLh3ca+3VbfMuz62oI2Ar/J3+XYKGay2PBIfCaro4wZFtrgA2TxGw0JLXgyrm5qm1A
uXguPLZ2OIFr1ZNC8KTg3xA7/FlFFLiy0rZyoEl24jTwIL6GObUCTt5SIfxm0Z1z8MChMvdAh+Mj
+xkuq9gWfBsII0naQU0kk/W25/Y8Amo2i+hMbu5p+5+C+J4yq2qo/f2jq9bk4Qz/ncT2jb9DxFsw
h+qvuedzKSn8sOm07LNKTTcD9fdGo3/EjosRR8PnltOIJkemKevbQNK+kvg95jRCLGinh0LbYwTx
YioBiD0kEqt0C5YP+XsaO6Cmkexx4HWIv2COz4euX/xIgWKL8EDBLlEBJumpwiL64rfLE7a9eTeO
kkPSp7And1kk65LBw2EXFAgz50FAtucKobyVSydUX2Kf40SFAySyCnvS5KgCzWU9iSOk8gqv3yjx
w+6dtWWTFo11p0L6YdWPcCTm2ICas8v6tObdvmTeVNLUxVeouResQ+V2ygeGE5AKH2KHXwMspvRM
juNlBAmV+boI8qPlFmFx3yYsHFtrcuDhFmJ+ClsBLojujFPBgjBHthEg5ITjoxSNS7oZg1HnaTW+
jj9d9jSui9bU2t1HROqofixhe17DI1FBhL+cfvoT32SvLKuPaK+CzkphHzQ2fL/JcU26OCTLxC2I
PccijAY4cQsga3iNx+YsRDjwIqt13K3Rq5mnWa7JM+nTww5axJUuuIWHeOCVD4G8hWezD5tjdTb+
FIKasY6kluho4Fb4o+LIGGawq+INcm399kuFwsFRAYOB0lYGFQE3gyTARUPMRPpLuP0CwxQH5KXz
X0nyBI4KMtOeSxe7MPpRefYyjDd65G9FXjTW7pf9NamoEGh1wQg/u8s6G8q1enaW+15ACvUa6FiK
VPTbUA5w8D13U7fNSz8xCGkUvf3GQzqvXe3wMnOeDPTNCoZtK5rToOYRzr8UN20lWyaMS0BinbkR
87A5o/Wu8kPC5vFyfzjZCkSmX/qo766/Nm8t9UFp+KMqx+RsmdLDthFYj6BdW1NNTmqzkFRE6M+e
bdseat6adibcnx7HaKrXaztmKRZBNe1tmEgP2dEpuO4Kndi0LTCzxtFazL7UktbiQ1lo5RqhUQUw
HqvgetggfW32rhkSqBW5cpD1XpwHqcm6yDFpzX+TcKHc7A+YU4Xrsk6KIJpC8aBvKayvmQw+px+Y
w7vxqczd0XQzbQnF2CCt/Au9y6QMZX3JS6lx0G1c2dlq0uRZicdK/c9uYrtJtPGGreVW72c+CsWq
cDfEB3i4szhxUhw6LT8tS+aK8DzyFOFXp8ror29oqDNYOh3r/e7Zp7o86vmhwsrMIRtU/KPnDVaX
GbtokoSEkanHGVcW2spaJw858/ydjDLIJz5oIMFivXDzVHaO597KODTy9mFokqTiLPb0IjgNATNi
KROBbFYGWSUud3RMTNs9PQzmXyoSzj/COF4cl4tOvHjeKZZlbq78rq8MMrdtNV3glPyPvSyLx2cg
aRlCBikkrlMWstbjaMf3FMq4fvcG0K0dguGkkHIPIy7JRL/TWs/kOKmk7w9qsofypf7Doh9+jHe9
xlRSLdSLQiBf6H/ea7tV8FieDAsvETauFc+MQKy47b4InX9oxxyzv/+/rz62F425lyaMu2Tpbyet
FC5DtUIa75rtgSXeWMRY7QoW1leYD7xS7NHz2xpWbFXOPsJxJCc0V0ctAKlG4pm5wgE18ahU3YQp
sNJF1toze2c0eQLG60aGHjQB4caBYD4eBnAicAuX0Uc+Q4Y3SfJy53PhpxW6IVffs9XcEU8jeyJh
j9P65GSQgHI2xA4zdPH/YU16d5Wic70QTXQPPvKMNtMSp/8ofELsIi0HHMDhVU3JEsZYH9GdPHBe
sagrd+xI5GlnViXsrjYrSvAS6WPUyVNhtGRg916Ni4sQuLycAFSxg9CTm0d5nFErVGW3VxqsUywx
jX6wgcmZ0XtAIAbveKh1pKCe5DGQCFdz2kVVwAyAB/SgUv0CbHWgo1BfNvD5H9YLN+tnLovUeCjj
HijgFI0lU2z+DU2uMK/hsYVFY/Bv3X9Ipg8P2GezAK1xV0lKUd/xSUyS+ooBfmdNlS6gz37mJYqz
cDS/ImCceGeo/NuoBEEuXN/8bYcQ4IQu8wFYiu21TCrUBZ3Xm/FoPZdmikjsj1dIAEKfCqQm0bSx
+D/+TuUe0D1FkwetQYK+XqsyULS0tBSyunl5yNwoGq8s60WzixH6uvdiLBXudtQP9/ELASUb1x3n
iPlfVgHkdmARcKJAdyr2+bhfaUlSJ1DSBbSg5RXXDjRfTSxeKzY7PXBiixIpUErYJpck5wJNO8gT
c4ab/KrENbf+66b9Hc2K66KJO26lEsSqAZOBXE7yq2IoP3VTFzC9BDNTnX5XTd3RkmPMfqDSXLv3
fGNkAZspC/44HpujRv2AlaZHVqeD8cwTRxNIzx0rjgfMsW0iUXB5BWyPrBGKFn5ls7Qjhp1nJtVk
TZb+apEtAKkB/eGxemeOdYBPQ/ehN+NpiJfoVDYZdevIz0tiKyO2B/LJQ9I8LlJkTcq05A4UhWG3
vt0Bo7YYe4EvERAwOqV4C2q/2gcjdyw5k6KltihEafNxYl7L3fBpBLVCTskD0XwmCzEjiRhkhw5Z
rWfrNMNt6lgOV29StYOiCnuYMN0eF3GCW24qcpLE4iIijFfnLRl77Sez27MJj1xKUzkvl1TqDALi
GtF26m3JBmPuyvQtLvzfUIvs/cZPStUmKPzQ3OHr3kA5I+U2hR0uX+ypC1xFh2nkFqte47MXh43m
26Zc1orzfoIEGLQLP3A8IuM/ocfAyCnvRyCYbiECag6miEW/G86o8a8IMV3aS0AKrVzYzV6LzYhr
S6Rkob/7gvzWG18FUbdIewJBfHJqZfBtN4J8ejq1eWTq4ovmzs/u2MpbAiQspWE8r2FTqm+LiZuH
HCBFqMNxqdj1JcR6Gu1tD4uZzubAGb9B665ecYxMLU1N3ca8xF6qIF02RdNTFQCaF0eSk6Rmf+Am
+nsgAuH62m6QmslbYnzKGg5npP6knpNujhGV0gIrjy8LuMjhiCGs/QAcIEb1axQztbzrK56oYtQz
7Ayo6a35+Lkaa65FmdnOHGTudfMeDJgGSc01QaXi5n9xkxiE4m+V7v3vzXa+hWpmIba4C4i85h6w
m3j0DijnbZPh9XgLrifD3ov/FK0zc7PiiAzlk0TPADijSs/IXZ8lnO1/6HGYG1zc/yNu83LSc0C1
pNOvrXh41fCXg/Qa9JYsy4tPKu5kCmILr0vVx6voO3HyBLaW8Q1/PV1wJv+C7KpL3RmZMz9ZabWQ
xW1PXQcrgDti6sSfCfHHfaPjkqSQ2AYoXs1+XNWla/M3ZtxDL8m4De0KHfcqT44RJRU+ZPp0R8Uk
fGF0a5hAYQzldUW1fpazEiTvJBESSPf2s0l0jRIZZQpJXWjcQ7S1fr4qLyvviOWgzimEkuqoKWrS
owz+nzbhWlzVxc2UCFdzT5VtWqkYjv8Z6vewhV0fJVVqCKl4S3MMtb28uaUtw/xRPWhsTRes3250
JVgowCGUzBUD3zyyCFgeAfoF27wnDnC8AeyRYXZNBZ6KAB5S1BT97rQgEr40EpXieCRaXpvCAYuP
P+1C/O/LmQsBEZnYsrjTsuTUUlKCPH3vUXtTKIDi6BwLwfDKBP0f7iWKQwSSTBaIEHAwmA85jJEU
Nez6+F5b1h4sC0bv+OVE5uQ+wR9Wa2fadbAPSkA6JubrY28u5EZ3j3hQHW1yaptxWJ+ONZfTzIHT
7XqcnyEtxwPck5nl/Q5+gXD9xkPyYP54NcDw6TYZ9j+ZGblJ7LCHyLv6g+hCwAk80iUlqJUHJZz2
Cpl5ooBhfXkaSOgWntLOnIEPZbqiBIP2dubKV1uSsiAmbHw/jDjRHJpFYu70yLxE3B/gM5pUwwM9
SZxpgJ1Ha8yqKm1UFNfgz0XywV6THv2I+RuZ5/cczVG/3zu97dSIbgrKWCCU4H2ewRGFnG3Wb5PC
ze6aYGWJLfAebrLG7Q7fKOTcBBKA55LdhTAIITS2ChnNBQ8fOMXj1766i5jMRlbGHGJRbiVVasp7
VXw0zkzWqjcOLG6S8vO8xR/dJ1xRsLgKAD02eEoZRuFh2FCZaFlkXYDx3D3YWEjRc9PbojDh6PiJ
0/T0o+gTFxq1G99fjl9zBW9rGd8h6zRg00zLc0iaWZg9xitQMorc7nmvoJjbySdD9XTvnxtM4yi4
3lGzJss/+Ik4/lmLBLwUvG4guay+ewOoyD78ftvssWhbiUbAbf+lr1blZxIBTIclKsewkAYOpU45
7abiQMfC5AorkMnY+bVNo9wkEx0VWq+W0v//tS+GCuDq7zM0CPSdEk9MnLis30hWVG2heBlWXD14
K7lI/Ra6E+iJWctcNsvKtVDpSqYdi4NMDbFC9M5ym87CaG4OvhUi5pl1Xa093h4uaeZdL3syh0v6
HukCiYf4UXb/bMlZmZMlH+40B3KX65LIVAVBSXcjZj2hlsv9fWmoIEozoLnh/kRGz44WXFwih4ae
H8Uzv1EEQoLF4rUYaYpn7BIu9ag19fXAKk1HYzErsofi+v4M1ZIKMQ6wmSZU/lQAJe1n+loGKsZ6
jQ+XERJqXvAkrKHTRVzo+iLCmeblYk0DojaeZ9SWNfBJxb6wnhn5NVrDUhXq45ZXIGOJ2f/F8ZBO
qj01C0ziecVxP2acucf6pTWx0RnTeOFmwq5L3T2M11d4tQV41MDXkh4xAXkCcFAzIjQyioe8Kgan
TG4zlly3n87pnLmtldoWOpknsYzg/VU3qvH3uArUHdTzcSFiEbqahnla++tlWy4hzzLn1OyQVNv5
dbGG1q8tgrVg5xtLhI8zqfKDpX9nORkFWJCZI5EZBumoCLtlta0++jWgkCo9f2XKL2H3jyEQ6mEK
cd4fLcPR54aDD1OrePq82YHIntr5p6uGdm/5kdr2wXJyss2PmpKqhnm7YDmp+pcxXZKG6PimCHus
oRE9Ts/0gL3+3lUEJ/r0qTUZLgXkp8gcVSjEPS+SokT8wkq+KkEwrYXaZroiMb14WChu6u2MLoEO
mOrtN7+TPzesVOK6lfawGzwcSYOT7T0UgwnyqoXaShD4m+3AcRFNYBmX2uufYLPWJaILkLY7V7uQ
qkPO/VVlyhWNLz3woYj3MdbncP6EToC2PzMIk9fz6bo/eJ0EJn2p4vujkuApfHUjn02uu1jjVOYr
2+x1p2ej0K7hHWunALfC4ipyeWJL5fJ5AzANPGQJULYr4NtITBB4ZExa7sD5VO+wii4wYyejjlwR
qNsP2Sx13jOdbcot2+4ALfZm9TWPmsI4t/UmytUwZAnEloU8LdTstXpRUQWtOpuonWC+gBqoXpkp
GCEYeAv83gzsfypbHP3Dvb212VRdr2AnVfjx8k0STv84YURU58UrXmc4n6sr+Z/3qTMSi+0HjuUB
yl3Z4EjbjGeWG1FkjdVLfLlIaoAzyDn0nyCtd/9M8LFkntUDilZrhaMhgcJIWs7+K5ExfP4YxDMg
Gd6HgH4SFdj6feaM/r/fTdLlbBvVpOU0CARACtEgruXbxzD1AgihnsUUy7jF7ehv/HA1ao3QUuK2
xeCtp0PP9uXOVH9zLFtbM3/3wujMN7Mx//h6Mo8I87JsQqu44KFBh+Lerx0V4pc5CE9LUAYHOgPV
PXzyAxGehzaRgDpUYaUOP0cn63GUO//cmVFTK9XnwHzGR4oG8LHIj5j2SiRqCkpSLqVV1YZF1P6X
/b8hHpg055H3z6EFrs9ADbc9jCXC869N+9+G6ZasloVvW6l80CX6F8QIQf5JALrEFjP5XqGWf1As
mHQ2n0FvNLoEs3ORgoQgyZfuKRBz9PiMiiV/nlWMja7piym9dspAdPlEMsVXPz/u3wH7sJ+W67HI
PHLz71bouJ2+EXJU3Wks76K9NLSGjHyT8qM0fOh7Z4jMZraqsmh4TywuzFIDDaDMV3cUpNgfOULw
3SBrrwaPNIoaozgb91qjzbwtZfkUlYf4x+nyLfTByy/gN/KaVAC3QXcy2IsSOyI8eC0EpGhwKDaA
4UVjTRkYL0PMgeLVXOk30slmP75ZLzA1lBFEqP4KzuxLYApRIU11rLqxTAjd4UzNLYkV8Vb70l5q
4p1Kym8811Mc4yIzyW/HVSyNP/RDKlCzs/+zAb+8NXmIi6ZPFe89guvBrlk7zPkJSKcR7POJZ7fh
mp3hjMjZS+kW/w3Vy0E1UzjqGi1yHjK6pINnZs8st2RS6xYRV1OZXs1fH09nrCecp2P7ZuGsBjln
9EBBgYqtuJCsq8TzMkaHiCkaTedSYXYJ74yNVCVh5nkaMa8JOc2kumpnODnMvJUafUX/GOmZ4JJc
1C12YgoAKINwHOP1l9X//7ioz3dZEx8cTuXWSJZV1wSpuUsXhew86FEKcfXufJgV5OAlWd8pjbuG
dL2OHUJxXlbq4ATUb5fNFxVs/FtG5rRr1i9q4ZmcIYw5S2KoXX5eXJ74/wz7IpOedbAZQHNPIEzB
hjgfhJ1rHlMv1PBRsDMwwaWcIGTDI4jnaG29lPsz2vpG1mPDtOxHRj/QVOnQhw7Q9MyZSmuVWjqg
CjcJ9/RyHWyW8trmFzmM00+4NVa0OTfW7J0sKqd24mwKQ/I+VWqF5KGvuyMMJwiQQ/+BYjC8Kv2z
0WA7lxTunuR192MOjuqehTz5S1n/fVhq/SisS2JHmUnS6UaHVAZOa/PdWiLPXuxHfPz9UVHPeTi9
021RKqP3LMwwpfkFg+lloEwZT3I0g2vTFnhQfnpPlG7kBa6na66U+sCQH5wc1v/4SQD4rC/e9PvC
miZ6HQyiFGD+fHxqb+0JNnnOAOJ6KUE1oGn3DSw5F0JqHzrZODU5kSHKnOK2aC7A6ZIMU6yt+sRX
Jv3qvG4Qh+xJtpeI44K3zr/mjByzOyy/C+p465XiRGNxY/Vu7JqNu5RLoAD8n+LobgAJAAuYuHmo
nI0jiNMtb7P9Oig/ByYlcQ65zRlAZmHt2cQeRkwr79tiH/Ct+f75jA5cOi2V4dByiWef66cqENtL
0bszIkkhCzMGPaZTMVuqoQVrA0/lQWSDDBxSf4OTWmirZVryIU0PV5Fodg01gCRJr8Bn2NII73cc
U1go0lqMHk9WzKHzdkCToxwlLVmvw8XMxjR3YwV6IwGIM0mEKiZY5el7nH295uX2jZ2W9vvczu6k
lmRRNwIMd94hg6sK0Oa5lcdpgXvNASdJaa0zqxXBzuJhs28BJUxos+BT14QXEtO4JIkIxP87Nj5h
w5vPO969D3N2X4YBuDWDCMv6N9NZU7h048VSvtCL1mVSBplLnmitrqzMaJ0J4v8Vv+F9dbv31yxm
Hmli0wM4qgMnYgYadbMiQrWpBSuzpSC1yBVncwFFHmlM0bVi0cvnLDHxC/diQfu/eaw5G00ZCQ9k
ta72z0ax72BajLqd+DWfSA7vn8Qs/YmZdYeomImGS3/Qh3tSafjMiq1ghdF8a+1Zm8MgV5eAr0wQ
cqamfoBJxeJjgTPxdyXm82jsZaaFUnV2RlENP0OCMthlQLiUppJTFpWd07f86zRfd0M/+JcFkRsZ
+tW9uKpNSjyrN3enqKXgwV6otcbSxHJhUb3f/M22L48x13MyyZ2Gwjn4eQoEvA35SxYtwCi1MAhu
KsBxUKHTjShliC7JU7Vxnrk+oHh2DHE8PB04WqoKp5IBtHatSoRnMnuw1pwvU0h+0rKZ/2BuZzcz
nt2yMoy+L6SW/yZxcSAUPdX1v4mxDIYYs98FTALmZT7MO3ilZL+6vBPVbkBv/DFS0DKba6RlOPZx
Um8Iha23o4PAtVtYXwTIhKGP9ZHhBkp5JZYi4EKhCteVpixIgCDFWLbD7N8pt0DBMNFsoEcotKFV
pZtOUd53HMtjpFWf2H5onigxpMayIe+9cz2dUNGahUjsyQ454969V+XO3U7BpJCT9a4DWYq2+Up7
8Psn1VTFiOi6EGPmzux80yL3df7VQvthnSVlryWiHsuqkDP/tzk85s65Ca+7vneJAOwe8b/ESioO
+Du4d+m3vhLM2Gkk5S63zfwwQayH54zA7wWA9OqV1KMBsKrgUgdxhcMgvyI+uy5bTZu2L5BjarkF
CAdGpofeEGsboEvMChXW01ZiWM+SgL65L+wm8UEXuGt02WmHW3PB5y7a9UxMul9/7u4tLW8qndsa
K6EqomW4BuETct7MJwGZyhovA0IZHGl8HPuCbFWW7iTiXpxWVLOAaxr4CFAxTCgELyrNx+cVIKRA
A4g3sUbGo5+6KfqGs46I5Gneo4s6hzsxm1/VE7+ZUeaRCTfOZju0ufZAG2HcCvLkWlzuG7PaMaBu
zGDn7sWiLVfky4T97JdL/Ue8Eam4ungwCzHb+1e22wq4aQROduu3DKjx+3Ru7PWoOQZ6Hh5RbmMS
JTAHT3g8UTigpF5d7nX4zPCmheekLayNeoNJwTxMNw2hGWM2feRbUeiT9zSYaGmj8q7wx87q2j/x
BUSdwu/Xiu7TDa9zgQ3pfh6X6Gfu3end34hqw1BDae4oG1NoWvvF5VEHH0nSMCklQ6TsZnXq70p9
lWZI5mD534xBWsFtYD2stwkK/ORJXCvLyK/cHSaZJLfNZTy+gAYG4kwrRWKQkGDebAcv3ydRBnKX
xxw+0lW8bIyM553bvwGg8AySxXC4QIUzQx4qDCRqRh8vyfwWwW2AG5IOptS8A+/taK7L/m415OAo
8MMjjJ96spITJuQnIs6+go7pmqEOdj86V2AWGZmiRUGc+V/3Pqf8yyffDQ/om74N0+D+/171p3aV
cz7QgdwdMI7UuTVwqz9MdM5IFbFURVGAdhJvsHkuGVMYns8F4nRGm1qDqVknuVgU9hDXWg/htAua
Er9/szDwWMUM+B4m2rNOrnMlpDHXLdzbDbKbjJ+9nPzX/7mHi300+dNwbWcBtRBfQLmCq66yIvCU
0qUZ9bNlpZAe/zcJdbmeGovnOLgJ7U6Hww/r8cfe56UEvBypFSGk6wZetI/3VoT2C9t7+Wvo0rEu
2QvnCw+s+GGvJe3NYQt3ka+fmpZkR2CU/Xhg30DAetV8XfW5Z0gkLePYzVJ1sIo+pyuskO7XcRRs
DD2s/HzVj0cnbHenuUrk0Kq3NuOyhmm73uVv8xUr9falGZ480+35gKgAyW62uVDTzV2FfTeyRyHq
5/i7rvbOEMqhDW1ByiJ/UkAYchtEZkNFdaNOhe/ePnjn2y181KVluVDixbZnb2FRlRDGYNpfWg0O
kAqZngtjmFWzbC31eKeKnBgsqDTHHg6tDzEi3B9UjcqV+lepQFIAXAc/bmkBkjtthuyyrvhjlf6s
4Sf6YPtTgYOXJKtzPrT812JXZsGO1SBihQwyZFSiN4Hm/XhLbM1MvKqet5o9SemH5Co+gB052YAh
5BCgM0dxCbcqGbmhYJkn4QafCGTO5awNiyNSd+aLmIFr+gqnAcN+0lPAAlxmZ9x+z6FnuWHksfWp
yyoh52E3WKrYSHR6dO9VYpxH6H4dyjRSsjy43fUk44N628LG99rteHJYay+BVpdAu3xEGNBwVHgg
X2sM8xiApGUMLeY4h+Rc0Of/7s/an9hNIzCtcTmNh8OENSS4fJUM7ZwzFl876dNC24VleFnxl4Up
466xcZx/zrFMoivEafEw+H7MU6551tD53B7eKVHnqLRaNW8KyHBxzlQ+k8kXe9rQB3DtfQSxZVfr
ukt3FCipMLNuVay2XsIY34vXrZenicwgZKmpu1MNIPBnOmatIxHuK94VTzRbzzlM+3Z4ydK6XfZh
tZf5+Dw/SaVKbvma3/GsFqjGVCzrKT0N8/MuWfV0Go6vnwSAF3WGFDVjPBva2uqLqPZvzKV+PBYB
s6GaMZlXKoeZwcJiBbJgOdzWGw4QQZLAvCgx31DW72AHgoFtCFl4Kg0UY41NaRHO1A7A16Co1HP+
ieq/GzJivFXs0hPHponFoV57XXgkV7V0xs4WEJNW8F7rjzFRhzMPY0mWL0g4pj5rYjEa9ZZSxRf6
OXRFeQxx5g5GSvcu2R8dcBGFcMBdwMyOlYUDwd8Dui+D0RAL0ptjCoGo3sEBKMY30trb34R3uIAi
D7jxGBk8wHUHc3n21REGwp0XNCCVFsfkLdVDjY8mnrhYXfftAGz+I3Q+E5RMPC24/3Kf4fruKZxT
TiPv1O8UqUEt8s4CLoqU5ZQrtZgEfeU88YO//KksEURbkE7fZH1xVDm9U2Gbrl5CJtP4rwXGoeTI
vWoYCIDL7foib8qwSnJUXIKQ0B1gyjF9dqfIt2yhJV0PgqSAIQzXt7OIQroXFfIxzzLEOpJF/H9z
ZjNEimMd0taj8TQRyTs41f8EAoQY9OaSEXBNzh9G6xthfGhpkJHua+4Fx3aSQEfQfNpsNIXVoNMP
3u/XRJzbY5wGtxx3M1ZXQrOFUVG1IDA9TDAZYb8YFLV9j6/p+/4tMBlSaE+g6Ht4Yh28yJmexgtA
KxKtOicqsdU4sRPsiBCNJsj3fpopEqCFW9BbkKIJlaN6GeVXPyXoc68kMqqOtWKFpJDwhjEFWue5
iKE7beLbkXW5vtAV6TLftrQuYUCEL2zIxZdvScZz67d1kr/obKig9mb6/JbzABiOM2uxfMeeps6e
EQoFIASm+PfZvGByV6Rq9XcxyslAZ2A41BxeNNzJIHBoLRQttw5oGmKMEg40wMfMcadmBVUPXNRk
E9YH9YVlsl9Day3IT5jw1AQ9RBUyV7LMSEEHmWmka+SMqyUm3LaTujxCMmh7nMmu/eIVGX4yUCFo
DfRWMo9UqL/oVoObNsegRRCzRY5jtSTrlJHP24utu5b33CA3R2uRLY1QAWrbBewPBNCJumBCryAE
a/OEk/tMy+YixIqp4FrMwk8ce4PF6/tT8MWef9qz9HWNr8gbG+W7mD5zAe6rj8TTbmPa7uHfC/Cb
hShYeRxspyM8im9quvKLEbuGDS8uSbAWIsEyLaQ2fZx5/4bRnIq0tZys7+Z4yeojn2qTnyE+CUC6
k1YsSlT825XC/FTuf50v0hWt7DzccGYcRUE2b7ky62wc3zKveLBj2tQmm65sh/sEOTEHRAvXGxDE
YuKiHUvied9lJzhTcD0J4bQoU4c0FAcPQY/UJYoISYVxPUBzpEVznseMyJbQE0IsI1C6XfnoIKJE
sFThrns6nUDiZMTsyXxN4GsvV2olgbG9ta37fxeKl0gbn7PTyk6Rqc7c5CKP2YUd8xKmR3Ipt785
ipq/Cm5vcq30Dwpq3s2mwnVvvH+jQvfonibRmXeE+2pi65g7EsTgVdSjwlYgbYhXHfD8/QUvpjZY
VHMn+efDOPABK1/zNxvk9tPrMTNnjWoKLQCEd7aRe+9piQr9ET0GuyNzuOi5BWl32dEVuBs3s5em
3IMmmuRA1P6q3qRMHYHM9UA5JyK9u1Ue7W48mbjaE/6DF0L437OVfkkGCW3VM7ypNr6jAP2P3/N4
6xHH2Q5kueFwrK+Bif2QPD4TmPySjIFDgrnLtl1WTIygtxlzTm/Ktmgat/ALwI7CyzIhMNQzQZHZ
4AZdkI40C7RhWz5RFnogfj8J3NWE2Fj4n+JpJmXqZ1a5P9zuBbvCoUbH81o+WGl1v8rJuJsRN7pZ
i2wRgHPpFmFQBXcHrES3mAOLLpj+m3LG4p/4QYJELg6s108DZQ4E1D2BYqEsthPiYBzZ4yJJgprY
YqTgO9JRiaGu5r1tpkowf8EfgbYIcITz5LYYUtb+QQHDeuZ72pw/C4Ktj+HkfxjSXfaCmEX6RuWK
DU1fL776CXewR2p0bF8leP/KGVV/nW7Eqye7Msiup4wePkRQYDgNSOtLbDjAb1811tq9StUIihHc
q9kjQmUqx39tec6S8J/m8XU0xXiAGvZSjEiESRMmNbA0nrNNDmoo9jBWfVDIF70WQ3zp+l7MQ/OK
cHJ2kScYicO4Onuo/JybQVXXQxdNvNaJgH4Urb/uiVpopxPlpKEnsD9JjHMd1RjF0GFY010C1jGI
8AYZAz0e7a3qNUJK7f7aqWjGQyjOT1YAq1zBIG4xGqNmW7WHhfv0imnselJAuLWD9DAXh4NTsU2F
6WvOhCFyX1H5U7jvPJQtuy08z/O6llur98jYJMzxzNBgrUE3Lq8L4H2OdNhfURA+fdNPYu0wEn7B
2j7q9+l8VVJ//pQ325jxhQgwf52U1NltaWc484wr9lrbmE4uaFWK1HHJ0hCveb+2ptuQCgP9HhhW
WKdobZLYRxH89zdcLgio14xMyIl1Sz9t4C/R+gzg3Ey5SFlkDX59ox7m3Ow570ALLjE5dd7l48CW
BGS0fGEKe9qb2Xw7I4TM4DuwFdtk1lwY4CaFdg9csKzoc18Tf3VSx5rVHmM7KYIzqC5xo4ViEwJS
U2LpoRuyI7MnXfy+2IYS4P3wFQN3XekZJMGXRdiyM8sXyl0Ls3P2P2UFub7HPdxrt6WCgG0qJN9Z
2aEbhFij2Z44XvGP/KFP3pEGRhus2VQhXRoLhjssVWGieR3swY5VE+XOLds10fZ487Sv1YKrWFpS
Q0xhRvV5VCaptjqofhXh3NYj1D6p624nAi5SusZU5gIO2fm4nTa7w61NGIwqG3d4mg5MfpH5/HBO
dC8FJp/vGmIaV/lAyx/9pAKHtu+ZOMWQBlhgkb727OLHUtfRCcFl6Jl46WZGA+ODuTUfLNyggrpG
pd+5w8IIs18R0smdK195cHQWVtdky2PeU2CUwqFZTmfuqMBeE90P+X9qTQGrdTPjy2/n6bb/xz94
EPxBeaGqE72etkvQqPVG68f8qS5wfoQaEU/5jTvF2cDDYoOcEasnI/8cAKlN0VxZjF7Yg6wUx20T
sKwm0dCV3gYfbE87lDypGoqjSyYPRbKMS73bqaYVYlRnHdTayOozzSipckdcccoF+hWWKsmDGCQR
C9zCUDXV725nFY8h6x5WRV/7hQfiErWl2i5kUr5rFqro9NQgJsAd9zNDJhNqN7v47nn+jai0BYMW
kK8yJzpXdO/6W7Q09T7R3sb1Zy9kbDlpJfJG7RNHgL6ISQCMCYj2nT9ByUeRc4/xywaEXZIYEYO3
z8o/1uxKx6+HNPDGRTrRHNlE/dtWKcD7hyVfUTGYl3XUL3OhGAWa8l165QEigAOI8bRPmiNXvt6c
twsCfebCxvNireWDSxlRGkItl9eZDBkwo5v7imGMqGY5npbDXYuIXn0kiea3yRTlExKGW6D+DASC
j8xplpv263ymGDxFU7T18OzgWJbZhY2wMv/8Sumwj9R1wf9VhrXnG52yqwlRSJmiP8xioNULMC1r
1srXt3KN5/TGuEXqFeRI5rVuCHBhzn5b0zm8/xpQRoDbjQH8n8jwXCbNhvuPjWdTC2cTO1U0d9H3
Lq0fDVHH8VEk/8l70KtwEhv7hUAxFXCrvM+QXHVZCIgobFmoNojrFF2BfRgHjGcu7/Dj/7YpxLgN
GYsXN1hqiQH0zm3OW2VCXK2YiXQau+vkyUIcsZlfW4DZ3Gq5mkil8Lr7z3dnv4SmtBDsAI4FAchy
RXaw0M5VbW3APKwCa4jIY+CSJb32YDbtsn+iieyRRjPE82G8HJg+QXhUwVJVc2pLGE2cz1J4NARD
c4m2OrsCO2j8cry7siO3Hi1irXj5u+RNXTiCKiAQo3HKdlfrak/NSWbF6NJCnS1EXPAKj6z+7X8C
ddUOTRUUBN3DWHRuEvyiapEFrcXzSwEw7YKAFd7Imq/2nTrKn57emO09fenQR7GuqExT77ZQAy3M
3R38SXB5NfSRK2SnCR597uFlkBG/ve7ZxHuS09waudxNFWd8ha99meeMRMMXe+p8zopCp/GlzP52
uX4keLhJmC+ZSBGpEHkjzQxSTkLiwlg1Az30xK2XdIYAquFS0fDOnEja3HYaAn9N9yDpgFkYQtkX
Mq68LyTXrkCgzzoDgs6KbvVxF+3hJZY/Tp0AspR6fjH06dmckhj8IOg+Kh8SxO7Smw3UhHaAzgbl
5x6utA6DUJCvxfgmIUzvODw8NS646XNuOpxEompqXB4+jlxRLun3d4M/7PQVsxbBIkKLEGEk5PH+
bI/u0mWe5k9llII6VCTqs0XXQjXTeQOf2CKKd/fo8YTNn0xgYpYTe7yfzfg1eXzDz5Pxgm0d2YKL
k4IbdmAq7/CStT/PmxxsqlU5I00ug2EVdVFiaU9SQDTyhy/IdFlRAIyRI6aSo5pFIXBNbC+UIxJe
w+CV3AMg30PwcVA6ZpeqY4cQugUReZg7cT9MOv4ELZU+2JbtoxKB7PoqyLP3aupgot9TPpx0SnAh
j1wUKVvXMT2RgkKORP0sWE3fM5X84+sCGihmHRiwm90BYE0JXwDPPUBtqEG8vgQ9yz3dRAD3CNYB
q88kwAiWAwdYAajb/IB9rGD/DhUki5VgtXbxZ3hqSBVgkYRRoUvmF1raGwvusetiOgYyQSXTgcZa
MzO9g445RNo1a79NbHvljhbAQWjLRN2G8MJytkH+n/9JGPRGaGMTEKhhkseBnqIDk5edDuJLRPsU
jNRz/oxK5blfaj+75enCQoaTs7NCBTmGCpEIDJLdJpXOsOzTukQUXpFaXvuRlEIYoDJ1dVCVTOMV
gYUjJII+PZs3uow1xbUC+Zln3ftZiXEeVJNxzlxeEOmFxbzrLdqdRo0z9H3ShQTVqel1rk5+r00s
useozn1Upb9KkUzuHik7hLLy46L2XwXviQNv3QbbmC0LpkV+EhY0+kLuHORsbYm/bvxqeMG9rjxl
TPZcILHZxM26L3JdJX27q6gEf3aCAGv3D4jXvNHvQUrDIpLeHQC43ejV9Uw0ZXJEXVcorQBAuq/b
M/1BlOqcRRBHScroH62aj5SZJbgSjNRFvmWgopCHO97mNn6imujcLHXY0Lwa1snuZkSkrEKnokyE
n+YdeZkVgSvybTeQZZ4GTKRip+Tq2OXaKAz9XxrLAG2c4raVtK2NME9ltROSVg5abZRqi803iU66
n5/U6lM0mzk6gTlXFM2mFVNMRN0nGmvcpFA/VSFIeWuNTA46d9FBaor7JAAMxesl4FcostMqo09M
IexahXLcWvAT4Wwmj1ZB2zqEXZzomGHsz0gxumn9x0qg4UgHckD3zCJ+i4SdbsuFqiQKKff+oLav
XtWUZuC8Cv8WR42VWfZKdZmbI25WD6Fo9R0rILF5OAjohGc3d/WkZ55KkYmjVNAmPWH2agFAZ7cC
4S9SicuTb1CiXPkAYyoE5X4QDF9PDoTBus4tpb/DeHtZGrMgPuSIVQdDXmWYDWtph5x6mjuSZ/Ba
fg8zlCqOM2IdzvvX/kYehEDy3gr3iTif0zcaf6dHfnhoDseigu2anKyVnPwxa8fKCJFO3HhaxJGr
vMkl3lSHjpsFH+YF8ujezKAiX030lHWdpULdD6IEbRYNq8Ve1lHBfZsKfrlb6VW8Ats+9mMv62Zr
apcuu22HyPonQGPCfdD9nePN6TJKO5yktNzMlaUDZatrVPhQU5NdzJfvyADCjjGTwn1Mltp9dEnC
QuDIrV3Z3md63VEL0MqF3k5e8WtLD/NFsM1/MBcC7JICFzT5C9rDJx/v+lK+F1VwlAU+H9HEtvSF
GWeg3gmzy8h+Fuwc7lD/zORepsQNvUm68jOuTmR2z8wuQzXCt8g5KUeXFowwe39TmNs4XnLDsj76
zLGIu7M6ys4zfo8XN0FVrZMTaoUGDHkHuqHU2FyMDb4ZYxNT7bmVo9VjnUow5HlhuhssjHKG8S2W
Mo8Ukk9H2gjiZxYH9CqpfmUyHAIACeMD5ijuHAHOwqXd+JITKhlcN3q5AF0hx9IygJuLbiLi/ijv
3NsNXLRECnOv0DRVY7YfzbwFUy5bVqDrefy9CdtN8WwqejKS8vMGOhyxEBKti52DIOZ3PsGSF1/S
9NW3ERb0j3jcUhHeDkW+iZUPOSDP34HCOkKbuAg09Yh7xyMIgkcUM93Zasn4Due5wF191adHqDwb
ks+zYicu+J5M1jXkoN/X5MZW3sJOrTbjmIin1HV4YjC0YVcYfXLXR85s5CtSlRstMUulGP/+dRwd
Sj5cLfjyhdd8Lii2zxc0HYNRwmm8O1T0cMYGWAvrOZKGS/WnYYOfrA+Jb/cy4prOF2uNganvpGfp
xPF75I/i40Ec+e1S1qEQC68uMsS/ZTAh0JBaYLZq3mcrUBxaBraBb51oeHuKo7Nt/fUDT5jdogoi
iMVg2qPM48k44N6LrW7+2HI46BjOdBdRsWwv/2OJfWPjXYArnfZMRGF5v+hHpftTcDLafb1NGmsH
FpSb1nwKmo99A98hn5aOrY9tnISbuJIhDSr9DkPGwBcwr3LRWDK93fwekaZJF14xfdIfDeigby7z
+bYKEL6+9Mdxrhhts68KZVui/6H7wZHbd8NVBot7cYM5LxgDxcRwhgOe8KOVMb119co5JMt1bCcK
IkecYRv1qoZqOEpzmJEynfS78H9VH5FnBObBu+ICSsPqmTrkgcmO/IxQLLUFWC3z7AYdGVAvgRSY
lz8ofvIQltIHRmFL9mKUX2+yIlopAMlFTBAQU9fvabFgHjgCQqauwWthD7avSkVKtFASLEvjGZqr
+Vn/+q62skVN9KBYNqQ179zk16FvA4ltghEC59rZbH4YH6JlgeiX5vPcCB2EQQl2WpwBAVpxpvZ5
IE8u0+KlXYpYbksTGbnMmDDTCjcOoj2ie49QFvbLrYYJswQYhpgfGQJSmgftvFt3UvEEO0W1Gs1c
ldRVHj7jfzpzT6kVFcIe0h3LoIj1BMC8csWaLJkmicOydfwLrdDhTB7Q+MIo8Iq2QcWp95kZhzCa
Pk6v+ByFAf+kTc92YYAIgIr/KSUH3uWT8ijS4v09xesTqpJ+yvL8bD4zVWiXUvxnVhgF8PASOZPQ
XyPJSPDOm9+dgGqWwjdySm6+zRiYQQc6dZaPxkRkcakpxMj+I+tqNHVxEOV+QdLy94QGvtG1Fd4I
Mn09+JgkBWosKCrC0iGb3c0Gb1xwKJ18mbTkyYrSS4aBE3Y5Ov6EYJoIvN1OTqDKoVAbhBtT1R84
ZknZy8BTj0suVZRqJjWQhYLpuuvpB0c3WYQIMQt9Xv4QpzLUEAHIUoUEfQ8t8KwGXZxHxFbfx2lK
90Im0OjQC1fUFReRy1FQxIKLJrimdkis4tKXqUEFvCHqh36tWr0UcHQd1pLOfl/HZTQYA2zkZOry
FINlAL7ARgh4782CuLvWpSVPPq2yPfH9p4JA3JGYrBPek8roRNbS4EOjdFriTAqBa7a9jxEDM2ND
O806pI9MDpc3K00jQNmON/LTELpfKaTUhBiyDbOAOdu1CFoVcIhkU8ONofy+4iZH4EhJg22K8Lc8
0QU1c7UdKJz2RChLIIHQKGMedYaOwajOd1BiIqybb4oyQ/63qYf4cthlPoaV/KUAMCPRI3Gjtt/3
1tevtSNwna98gjDhN0bE9ulPpAmIwnbKPvPFSNPpGWywGbJrzkDi5hrywZdUDtp5EAdU7U6iVP2J
r/AUjmc6eUI/DFUBGtZRxFJgPsM7MlcSyyroSEaatjLCVBRokW4wG82hsuzUL4v2dJW87QJL6phu
hgFCxLkPxtF43Q1Wy00y+VdRfmDRKcG+9Wa+fAb1nsDADi5L82t1HiLOxyKRY4t87M3IA6mOMCwF
VJc/vLjXFpDPeLc1BLR2kZdSPeIdHlIoZjVN9rlC21j+OUqxeaOLzaPMy6wcUN5txGzkg53RQ2L6
zTdqPNboGrbbBDMvmZEkLuq/PTUgJUEK8lt1K+mwvrzS+QXGaCf0H52FPdvfXk+RtEIAPp8QzHxy
IahuLo/eVzU6OiSkoUZyOjbLYCgCPJ1RmZTu0UZeTWRNeUn+tXOePlaoqZbeEPXLNh9aDDITPfdE
YCjw0Ipx7un6yji4a7zdPd43c91T0hEJCg291b1ndbu823qKOpr4WQWq/Bao7o6cp5sXEj9/sHut
6TzDfWifSWnSRNp/pPLTlP6XsxhzQwht7bdiXN1/njglwoC+c35TZ/E1XbVSzuViUDd30x4ARq15
QGBoJnMUDxlDUN/G7ZLh88//iglHjT6V7prMdMRKvN8RfNY02EqsbCQCjlt8i2DfYO1sDaa6hbXM
agEcuGWF30TJCVAv4bhb3Rfw6/DUnkIUEwYJ0/rwb3tJFCsF9rGVauYl4d3ySbDxpRHO8F168Lrx
RLyXFmEXweLNl99fNHAw3VKJPaQ6+X/9OYtvtVwTI8BDQ3wIojk3e+cTBuwNdR2awTECsEVGvPCD
nkKAHCqKy3Eh2Fz9orCf/bpdGrZksNxzTbiLAsazmGxZqrTJbP1AeqbxSvlibdhbGJtE9QhBiiPC
Xxr/4ZixNyYsAmwitBtqu2hvq12ZiLuj0Ob/f9dGlWAbMW/OOS/RyKa9yid5sqh8wPz8NcFcasBz
Nwq/6zTAJiShsrIMGYEZp1ChlcwScLh4/0VQYOnDvTUzW8mEZAnrqwsR8SVibs4Ye/wmnq+fCLZb
Ub+ZRweL6VvpkmBeqxCu4qKPYmpUQcudBUTuQQenkHpLkkVAoYg8L78T34KQyLuU7IJ5JvA4pecv
6THqgPMkSkdYF+omuN6lNAy9OJyEChL0zVGktBvQQNagOEnB+nhWr72j0buMcB2HhjNZ/bb7Ubet
RoOeXYODADw8luTB2yjiicUrq1kuvNsubKULlwFQOfQv91MJ/F+Mnq5ECHcaeBoIGb+9U292ppaZ
amcdZQ7T+tSnEmQK5vYE2FGhhaPwibWkPP/ss2XlEllbJm0DBCyQDitoD+Ft9oUJHIb1bWciOWxn
r2HAidCKLygLiru3+73T6L2LB39DOGeWtmTRfEb5sN4TP9TsY15cXDTK0YIrKcruhNXYO3OulJKN
M3N5ewq1kA8eq2ZcSeLrvXQn4LzfUE42pI7BH4nYlHYx57BKLAg5aiwN3jzo07uxyj8aNyeKKUKA
6Ims+Z+IDYXn0942vNQEHo3zJWAZbc3wdSr9uFbrQh4stNCXYE7BJbq6m8Z+Dg1VKWREH9UoF6lx
Ye9A+sGP586DrJfdihoSR1fHSMYLzOiwbhhJRLgB2aTc5L1SmsZZzc5okKS0eASsPW/nXwiGxouN
MdBouK6OUXEBpoj8rXEx88nA3hs3nHGlf++JslwdAqfYlQluvwEZGSmxIwfzFvxL4MbeXKGOWJCQ
nKPkacTghKEl/VgJUg5jmhl1iYgMZ05CuYyZKy/mOYB3m64Lee8aQhky5vWvdYVuDz6rsev2kgDy
JHC3fps6ZIe7lb57btKisIWatVXHNLGXOf3/vXXIkSy9YRL5qiT8fNdyWXO9RUFGUWXrMDanJGOQ
LISWZ+WLfXy4Kv+f7ozy6T4TOOVB7Mw9OVG5vGFzamogN9qGieeaM4ZfpONdZFx3tZ6kgYgYFIOX
MSiPbwhbf3uEBKgdal7wOWukD5TWxbmcof6SHjRrWwUtN7e10sFBEQWvukjv/jgtZrt5cQ7pTe88
glqo5KAKG8bYxLg5cgqBYEsQPs8D67uVY+4/nIRrvwg6PyxvzYh38V9+1vw4VIaPhuGAGFEn15br
xN7AZ1IOAkP0cPEYSJDiq/YABXCXAGxEDI8QGbar1Fbrcp2bmFtK+A2uxKLOt7VtYS+QUnl4+oUS
6seG2eC4exIs45c/cWSVzTU++i7Fv4IN9X8I9v7zvwa2O2yVeoPBnRF6Pm/TgfjfK+6eeqlte3km
MHVoGz4G0sQsN+lMzw+y14IdXAAhra4iYl2HWJWDZVXprMC9BHzaVQ4G03OSXYL3b0V2o3cEKDrh
Z1VMzZuBrUDRG27m6PI6dAwk4sdTk+9Rr6KoJVLZn2LLhoxOqk/i2pkftQtvbRkF3uwEHthjDsYm
rEWAy24UahfqVEfUqor710rMPE9LDJ2qqqBoPbrODNDi4aKNWiIa9ntX9llcPoP5AIdoiH4MeTGx
PISx4VFIRMIwgFxKKF8cbyamqP+dNTKE57bcPRAKA+evJMEF5pAqVM4nCRGSq6k4sXMHsEoLqOyC
/sHi1Qb5k60QCzJlP0BrsW+icSfNQPZGkSS+Fqwcn2CT5LcTWVnEWhTzGwZFdiEpFCmPRQ8B3zsJ
//i5UceVn0EnzGFQ1R+qy043wiJs6Zo/kug3R6Nx1z+6nb7/HwxUZemt/1FqY5HwvbRAjxBwuldr
2xYMCzz8DC6YJZfk9s6C6Y91+Uxic4zdK8UZdne1mC2ZgGea/X/93tDACsMjUV9TN8/Dpx5SsuBS
oc+pXrHsbr0z3uelJSV2OP+fg/e/1rL7PZKc2ET6P83z/NPHGCnwB1vheh/2DqJ0ILscqgPmcsiz
Lz+/DMEq6g9dUApFDqkVy2qNf+GbvzNtzXyIcoV6LhlP/+7Lz8IWYkDzy624K9ajm5sRWLsaL3nY
wwa4R6kiXPhqpvhHyYpa11q6wrV1M5YT4IgFxOOjqw5APJNeFvAKNtnxIu3iMgOs6oUp5b9zNF8O
MzsmZwJg2OlSQBAliJgRQ3St2wGGoSCYj+CBTU5iCsYz8v2v7WxX2m9TGuLPSbPD26o8vWDs+4JN
MmfjL+o3qTU529XpxkRVzpwehC3sfNrZ39faFZW372xUdIgUzmEe0xwLFwV82J68puOJBJwKf4I4
EiRkA6YK9nIps47m4snRo4p7kp1gilyn0n+U9N7mqHPQ+g7QUQ9eQVN0epI0Tm4h+RAqmo5tbfiY
zDOqyNvRknwBcmNdNhjoZZ0fF2aWjkUPvqyw+bbHtAFzjXtzrFjsWBnY4CQajLhLQYaPJnI9/Y/Q
dR9uM0r5N3Wb55IURm8SOPLjkQNMyqTFMkvpBpzybnedjnCyza3gRw2LVUUkEXiwWWdJwoPBAMnC
HWwFveXvxJ2Fb/xHjpnAk5j4lLOMkR1nG0HV95fLO7PzAmwut3Y3xI/jfo7bM8VnQTL5m+lLy0uh
HXnVBq5p2N0McBW3JjVGdFYxeibJA3U4mtj8NDer42j41FlAMe7oWL2VVff0HiA+IbHdLr3Nc1CD
MgFLcwa9ronY6ECplS32UuMV1vjuwpfWhVs2RWXqIPstKYtzc+Yak29UX/IENQOHG9G3dcRmP8X8
5tjBKp0GKnIJsR+/J+Ybh+JC20uwMYuWsnaLOL5hlvbKHP9oqYEo2r7Ye7V/XWAOfRgH/iIXy2ST
LL86njRYvsG1yY4MxD2OLJ3krbifrBvdAUhIfzdTD5//GRuG8uYIAvGHQ2cuczJCSGhfN+Zgo0uw
VOIbb95Hj8hq2pyhZX1w+0NpfbWvENDZhqBE/q1ABLBuIromZ8NYGVDgd4ZBOjKxbhjtwi9pOvT1
L9We2Vs8uohX5KU++FGDhaWPhAYZhw4pIqhwfpXoprJvfmKhuERcdH4lW0gbw1EIF+aEkqyzfwFP
Q+C0tQoS0s7F6jvkKbNX5fl2Vpi7h3hu7FzgT2ISMJ/MV7EIlip/um9eQ+6OxLL0//xwcv/IzPTE
QT6I0BjctHEBCtG9q8hMJbj8iMVkcwgtMKIJKLqBGeuRKWl5RpXmY/fLPsZ30nc3mWjJd/ZM1ijA
t3W2BlnsUMa8fdPh+Yejntu5MIAAODqjtnzxbwgetW+kOe770Vb0X9sub07gpzXHzV1E3PlbiZJx
cyDteq3HdnR5+J+B2dJAoUxTu9VFT1vtUofvWzPiIniiq59OBdduRuifOt/GoicWRf423gMSVBJm
Q1RGEaaZUbRs55a2GBtMxBjvyblWcCGsbnz5ttgYhwu+UnrVG53BhG1pN+LMJeoiTkTJicacDIJ7
/STKkqhj1VBS1Br/IHoszpbernHXxNXVYgmKfwIk2hClVM75hetAA5H3fjf1yRj8CPFaGyVEYkYG
dgkn5TeSA9yvplHXIQfnLdtI9A4wOk9xSFh5R73CCxWmAOUzD7vqXNR88MCdo7/zr+xJ0oXqWy+o
mkUeWpGDaH/g8k/L1FvQ7GCBpPgLdDK8fQmK2SPWkAiIpBJXAI6L0FC9W18FzRfNyYTtHZCOmyc+
UpvIgW1F/6Hc5VVfkHT+NE2h4KVnODAvIQ+QZ/mvbMpUiPpdgTf7V+h2BTD+6UdQqMhxqzVHTbLs
EKWFWbDUSnPLbYh8CIHDiBFRGeevdZ61/zRyCFwc6eCrlqt6x+yOrUGOVVrmPdd+nPo5hnK2QEax
KqtqD0ZwItjTN5yWybobNmxIzqBfMYpGcTetPb49JwwGq0kZOQyrsI3UkN3NxTUSNUBj+3GWw9UG
7L2p5sQrplT948Td/xC3+PjhNlqhTk3u7k5/uSNuuaZ1WPLvihGat5Id5ayC7IF52CVFFe1rL5iJ
7Q2YsWwiUYKFJ3HXNtsXVsoVyP9HofE0PEUsibpLA/twOibW/JY54oxU5Yz3hmsbLbiBHMCb+ASz
CbhjOEGB6vDTD3PtfQmIJdHnZjqZBweB1X6jCCWZfPlq7f1CqF63NBnHw5VM8jEpjvSGW5TCk9gL
YNDdk4VUD6h6wSso0oOuLS5yOKQkqW5jeBkX1FumsXYV3OpRWy++qLE3xoP51nEIfNa0o5IbcBBY
GRAlKT299qIRwoLf/WBQLfq59h1NdNmDz1LB3xu+CcD9P9WL5VVR5mvL7CjZrooN0+JCWv/hl2Yh
J7+yHego7xmSibyqMsG7Za+eHalGxGXPbJ9PNILLk0Nu4Bv1J51pWNtHZV6umYpUHRBwkG/KEjXe
5nRsVf2Y4DThy9K/GPoI/injEFEPNvBs4O3lMpP9wZi1W3Od45oFdYlw/ykGQCL5Hw0A7bfsc0D6
LuW5tjgDSV60fO/KHiAHPZeKQXfsnwGYrspyWGzoxMrKrVMxS9gclG9uNQfHg75TuQkYb+KxYIhX
66ye4z61XV6kXAA09/rv2wlbR9pfqVI7tRkeMxGBdMleJe0mc1S3WBOVWBJwcGePzgg/UQk3WXKq
Ra0a1cxOsgoEZ2o0CDqv1qdpZcfWZ7xT0wdcxmhEMjnH6+V9qzLG4Hl2l+GpF8Xc7U5RRLa4dVT2
O4/refnkkJoIlLXImEf17TFUQEs40srw7j/vryD4fRt/sJ1ZPfsw21bqQtOXIWEL3hhdIEMWYYgp
YPyhRD4qw64W6ZUPH4NnW5CPLZQ4kGnh102tNFZW34NZ0fuQiQegZ/b8ST6KWlFiUiGXrP6bTtmN
IrmmE6ywfmkBh/ndmQ/Tq0T3Nm1RHPxM0GExk4wh7A6VewDFx4wXEvdD+TrK/yHlNEZAnBN1Hns7
iJU5UOIAnvx6RRlRjHDbW1YuWhbKa5i8X/eA1MsDFEhQq1n+UtMy8oG0w/jqXD6zeCwSMi9swYls
wg5jQ0S9qulEmxWBdf6aXAY7Op7dD4FArf+guzpj3W1be0Tzn8DefVGN/P8DbLR0XbXxSCLe28q+
PsAHkIaKI2N13gKm89Mo0P7QUwti/WvxQf+SBdhAOWnuVFMbpG1sGTp+wqSUjxp7hy3C4R7EDqEP
QQRZTmeq+fV+4cNtWjvWPQ6pdXAGugL5UR1gY3EHDJ6oel6LRKP9aSdZZgn8M/CCcU88OlH/e01s
LQi2LdPMyvmaWsRPo0m4xyHRt1AtBfLY4aDW020JmuZ46U8jtLa3TLBLsK0/YmvIkZrH0r/mVPz0
A79splnWhxUDjGPNNWAFIqmy8hVVvQf6985LtTW4mgYPIDJtWXWyHXU2V53PUcG5SgiQK9Xr3jFH
OGBKw8jXFNvVZmNjcWW+yj9viXFn2h2T7gnOOqsHlZtVVMU+DG2vkmUSn/8to4Jipl4uV9EEJp8l
WEMmKuUWMfpfyFs0BsuvnCofcGsKdiGSIO2mHKtWCZ9rjBzmmNO0tIIL2Xd3JE8a/I1PJtbiYXN1
tftCk8kZnalxBZxdMPYGsZhJRN1ye4DFD1fwY7XQkR2GrV9rxANxCM/DzLk0rbrT7mxfVBx6PDtI
Rl79cH44tJBuiNmMsHdT1AONYLjCvc6JfRS4BpkOd/aiR3orvIqIj51WgfiiUf78/Oxu8KXKpoml
G391Lox4vVqEsrk4rTUTkC/FMfbrbgUU8GZzFRtpYc+eRNUKutTng/qJVmYzYHcKeZcs6Dtd6wzy
UHGPinwpdswD8Qubk7LGbQnMSbRDdL+i8kHuN6AItZLKtZGl+WMEoNNvmVVYqj+tQ/ojJLkPX7Ac
59exhYR4JZkFOcjHTMubwp91Qf0x1JBLqlGZoj/OIHGgyoGR6Dv1wE5XxexXBxjxZgFzsm7huf7L
cGPUxsXe4wc2D9Vtp66KYUdGHPFkl77UMyXHdLAeXz6o6XAQvXHaeWZKcLyNUK8nx51ffXMkDe9t
Lo9u+RlOdHYF2cc3tl1B/t96zxRHghNnbUZTCdV0pju4CH7txTgQGmawg+MUQcM9vDPpiVJ3UtL1
qN7oF1OJYwUeDvYisNyxxmvSY4j0Ewc1YGFDoXHuHV5DtClOpju0DCophlpS9HpERA5MHviRLx0y
1Ng242KPYw2hwD5yC7pTc9jteqTuKRYnITpZylP+npNLoQC8v3WALnDZNau/vZzBYQazdF/d4T6s
nxMxTIItg84Bob6kV/L+DTOpajTZQZs81J4bACYkF4zkZSxii2pqEJrhiGncIGPKzWHPFUKcFBh5
upDdUxhB1ftn09ththyrB3jRQviHg4Fhw23aTU+J8ZHLiB6nHYknUpTc24dOMAxOj/wBO6TIcx8y
Ysuzr4FJGkG5f0BXl7sRmUczk+OXCB//m/cKrJwif4I8HXuep89f3Ol8V9PhW3z0RlXqWrGXUNii
Xam3UuNPcgH7d5wZNURrcwgTkR6xi1VOjH/a9Tl+/3ZO43WyObmeytp1tdFwnXdmeggXYJ3UvjH+
iDMp9DCaYoYSiEiLLO0tQUFXt+Ov8lSEBJW+/C/23tqHF688Mbz9hr3EgD3Qf/qfB2GBuWiFz096
RhdpoRBq+NGSjXscTsj+5tINQk6MJGWKns5Wu5K/aEVdUcOEgD/Pw7FEvE6B68OBxNyPet14YEvE
KLa3YnnXuUtv0zXmKAWkkqYHnxY3p/rG6A+EHSDymouUAsYPxkcQUrwjrFbhdpLlzYVvlHpcNVc2
1h80fmlGGNKuIe6t6M25dXa8HYFOxe8qWm7ECZvnEJe+Zxk70oJ/Pgu+LjSOwvNj1W1E+vwlIzw6
1GzZmIIiEK/jbh2A7IFELRm5WX7XbwN0c8ZWglObwcr7oaPSNBDIsS+CFnpfF08h930tOp3fBPpB
oa89x9i7XQErF84V/PA0dC3F0u8FCm8SQIMVMvM1K4F6UIOdQTa22xQ2X2su1qsLARW99tEIc8U9
ouGcZLqLWEELBQatJsPjHD/acTC8LqHBsyypdrBdPnvJmAMLtPIIJ1w8cLwTzBDP7ASfKOmxUypM
V8ieAjw9hPNntrMtn5w/92TA3y4tOTc4BzO/SUrvClR8HppAXIqh4ZvVOMKZb+attHob92fI545z
SyQj2oog0RJkWylswuW93vDDvPAcrYs48w/qXZ6qkxw9dEetlF4VDqS2z/TGMqNLoZtJrrngs92s
R2m9kAkP1c75hLL6vGM6lmkYrQOfBvtQ9UWHSqti+5DL5cyvO1qnNpjXBtJL3fqVcbhYxgJC9Sjc
oDuZo5zZFzinAzuBrG/g+330rRsdSXtd8V7aC6Q6prjCSmYd4+zwSPOi4KhQREMJIG6by1/eDJ3E
CuJn9VLMqP4xzlQSJdrLRDEIQUSg++IQPHKIx59kx7xysUR43ex/vfYJHO0n+snEvNOB0YHuFepL
82dXFfp3HUjCgI7wMQ2c33cezg4b9XEo8TGi14EoymqLnHaEz0tGDafsIS7RN5/mASS5yOujq0Y2
+B5Fp/Vln2Dj5RMpRCIqpj0iqEzav7DATiFzKa+POUrLcE1TsWybX4U2Vz6iEPUrzw4BbOeqAwyd
Tx65y3yfiRVKuYij4ipsvHCVhIOUcFzi/4XZXEVkYvtSnX0Uq/mQI6zn6VvtldXZ6QHHepBX6F/2
kzl/orphMdQBkC28oJjQSHwDcyg7WSVm2/H2WQc+AMjLcZubonfrKZAhwPFJC5TrftfKicw/Vz/F
+DMhtqUPSlG4a8G3J3nj8y3WdSrgPKtE1bc6mHvyfbZW/KjCJv1Vn//Bf6WkkHRjdF4rmEx8NQOr
bPr0vZ5YLMcLQ2t73DGc/96sIoFIdPGF0U55aZkfpu+DTRrf+pZHxtUKia1FXqaTlOkoNb86kw1r
bMcLPiuWFcLNAfcZ81r/yqQwfg6XhdGakLCOVWykn1lEou6Ywyl4ci/CBofxDwFep8QE0sntzP+U
b0q7cbLw7esPb/6SKD4UOyKE8ATigT6sjQYVQ/6afmfpx5MLtbu+easDEUkiKdmMWpYi1nWDlYQe
1H0eU0FQlcaijWh2R32zVyj+XXv8P69i5Sv9awHtw8zdIGF/Pm8dS73WLEcqCYP2r5LlwRYJj6gT
nuVAwKAZoDpnhbSJJw/wJPpMq7rs2mNOR0w5pg1Ze0i/Qu9UEgjkVvKQCRcOj5cTAAbJ9kwJfkIH
J04534jiZofaMMi+4+7nyCKFCe/yRV5/vq354+KRHdAvQu/tn0UwRPqvNZPtpf91kmzKJGFoZP1i
m/ENklm7Q/OsVapdBNgnphVe7+UtCKEGU/gXv7ETiv17hLyPhSTXwfCHM/yYA6l+rfzOYujOj9ag
bqlZfZ8rWe4D5YpMftEvcOHr0q6+Swp5/WW+7OGmgjmoAgczgrmAXzdtue8IRNUjWlNvQGDWY3VY
Dcn9i1b0maH/60yhj4xMnhC+yd9TNYDurlG579LFzj6Asg1xUHet2UI51ZH558T7jmZya4UL9uI8
QWPwEqvkWxUHJvgznOqw7+N51/LNhOhjZ/xSFPNQ5tWw6ZEM7G6F6HE9TTQ+Xsf0mtqKU20HU7Z1
0KNWs4K//Vx2SWspbQTmQjmTW5D/CHiCDHUyiqupvAmS5TlLoPEJcEn/zJQvvSpjdOgg4Nl0CBzv
dw3HJgGsGo3NRHnbGMS9GJDpoNO2tvbE/DMTGJM1b+tIhFI4HpsBgxG4HQGei7LmhB4jVCfu/qXi
SW0oL7ovQEojj6jnqfQHe8Px1U7jzjdbQssBC9WxYBDpz/zV5cQfRO7vB1bysDuYNk1cmxaibqUl
c3YCF01tfic6e0ft2Dmzsawu3vC2wARZbP63RSf63o4np8iADcXQeHxB/0VZDAPj27WnQCOBaphs
nxWOEYS4TyUzL4xJsk6NK9BS/xkFG8yHI1hyeMRqVXLIcf8Kv39jy6goC+3txHLLqqShTyBdttC/
atpv1dP016Xka7RhuBlvXAYmfwMvAfvw7WTNikE++A1x2vQ2LCHDlUBhAp+LdbTqp+/YPPXK7FfX
fGyKgyl0J1Xfb47Rz6DhiWoI9rWYOP9T4ygvnpPy0Yufzl7rVJwvBoqgszMOo/FcraEX1g2g9dQ+
ZlMu1AKuwzmeVG+J4W45fuNPJib/C2Vub8D2qCAggblcnnfO/ADQvR3dLOMhRUSmCr3z//tL7bAb
QuzwwRDuxzgOM99naw/+3HSyMR1QJx5L3YzC+cd0Ob+yRcDE1Wl41diLDAPNSVQNVb+4g1s61dKS
By9Jk9TQO8Mh2HS8JDf0GWxhv5HjHOVlwahqVLvWFkhxUKO6nJLIkunKXhIQPxaBHaa8q3ws4BwD
1Vf+RMOuChAawYwvs8zjsKlMZKx0jj+IqQPsJuz9LLPYCYWqSkv7PC4qVTdaEuVfzRU8gc9pjrAb
CbCYPUe/ci8AXp2gZWfQPI2oF3Z9N+Ro4QQDT0VN665xgcX2qS7jsGEe7/NjAZ9Fot/LrNsGhijD
SJPaBnQ8BbMuTDWR97s8p6vZaul7Fzj6jLbHhI9BBca3A3uC7N5t22Kt0z9RlM7Yj27GhMmgebkP
/RqDRTTIoElx38EuU3/6I4s7pV5i8PvAJi5nQ6w0HwqNeqlswBmKVw9MVTwCC+1B53M1Rfuv+S0H
+uCJQkYAuAAhWwuV4LNauUEifSe3sO4/Ccy0e1OcGBdjbgARgzQsTklfU77uTXmDQb5JkbYllKLk
FFXQ4Q6goxryYhPDQlgud7o4zw1CqHXbnG5uuWjANlrOXLloel3gqbKOu/6jV4Ck9IlSeF7V1A8t
z/1w5ekNsMmiQ2G+ktT6Y7xXSJ9lNyc/BIOb9cXNzExbeAeequIHX70siovqbyTDkcT/QNNbe14d
zpdLzScpd0g1O69EHT+0OjRB5JK+1zbm0nX/xHpCDeN9Lm0+MTsTsPZDkRycNoJ2PNGIkPGKIgPJ
BCT1rUXdW8sb9VSps09L4QeeF2fcHHl5ehww36WEPc1HKjR5/g4Vvmni3vat6nBzTuaoLXZNwO08
9+mYf1UVCYnPwSJjJJtrq20YeObULRRBpZJRdRXiNuZiwiQdgR3B9a/uuJF6t7UnRKAp4iRmrU8K
s8ZAVjRVX/XG5pQaLJfp7+SnLwxv+nTzsACzxkh5fAYcmkamG7bUb3JGa4pOUtO9JmQM89Crg7vs
NCw2QJWgHcCfkvXC2rD1b7W3T4WNzuD16wtm5nDe7xLJgOXy8GV9JyVZraGxtcKtg6ti0zzT3WZf
SEKvyINYZOZ/FWEmpyT8C6icpZgnOWOX4V0/+n8VDq3VFFGLFMauxFpyWQmo3i4o/OsPwusYHasG
tJwTNq86tmWKaDeNB12Prrog9Ab3mhvzXYx2NZ5sztMSNLoTu57QJQpsTVYUE4OmxTsD4Xt6p+nN
4GJaxnyKjnHrHAg+dLrfnMRb83Ga4Md+m1t+gsjRMD2MDO9uiZi0NXVfu2bsicV5tXVKw3172qtp
EpccvoASurwpvDe+Rb5+/PQCtfGF+7rHdWZBrVHCBz16K46aD7IkDF7xVCZxYuS53QAYG6bsNe4W
MjE/n5zbzLqkkOxjZQnnNIAx81qbe3lECT3hCS6UmB1sAS7nHduZqPihQ15Vn0iSq24HxJX9KSDg
sCn7W344Sx0EXdP1F6aDFLPuwnxyoZOqz7URKTg4x3Xcj5k5AzESL9fMaUafAKMYd/7LMCKjQc7h
lAXMcbFp+oOedby4qFil1qLFCp61R04R8Bmy7tscvp28zrsypXqyLpXPB688U/oq7opaCSzz04bv
E6IAv9MYiolWd77Azj+sAhN7EYtplf9VsWVGfnGKwZiBFk7jLfoihyjrRGst3h0md670U52NOh1m
wxtP+cQNKa7aDUapaAiy+g9gQ5peI20KDf32LRRu+T+Coswr2s+VO3z1SY2A1p49xSCt9SxCDct4
YuKOHRQvkODxDg240QeJdkz2Z6gZ0x+ASouDLoHROiJyEhrSinecTcqREZaN2KKWswCktflwqKOy
I9GdDHB5rIORoMAUbJkgI7FCmcWmvBOKkGA7XY5AUEfIM+KUkbe7d+2GoOYe2wekLSvKFM4q3byO
Ycw1mWOIqBPvGYcPsp6xDmN+BMkGWTaWSvYD4hvnf5m6f/0TZDAVIKud+g10bNvcnERIbRb1rsGO
cVK0j7DDf9C2hPkVGPVEEYHDkXN7PMhPCpgrO2SckoV2nhdNBtpTqmr33amQ2AgQyQFiIsxD78wR
/2FyHajneeVjADIAGbmXMiPJv+SdR3HoYl6j80CWCnzUzPDsFaSErx0OoIbhsZIcA4uCjBydB8mE
PZKy71ft5yCwYwAqEe2TTL7SccH1SqLLIc9n4i0cK0bKZhQHhwkhfS6HYA9W2WC40xwde5Khck/w
/ORWFg40n5dhTlB7zT+RoRln1IRftF7DICv2gjSXKdFZV9R/a8pl0CLAwkC62+1JyflPvCEQAljM
lAldfXWY2wMlDJrOlzOvLj62fVSN5A2XeEmezuvgcY5fiIeVgytV23tFqYM7a4GF0nzKNmCIXtL2
FWTLJZlhaINV6OAZteAa6s3kRuxlS16Aj+KcZkx83KZYVR6mGfMbiA7MTE/g70MuZ4uwd5h1yvdj
MG5PRxYdAbJnXKk5SF30kc5xmE72sD90VQk0W1MOT+T5Edgj9UpJ1DduvNvl5p2/VxWq/Qd9sbKR
RFYkRac2xGFyVM2MxgcSCnkDL1ZKsn/jZMw4EGOpi5l9Fj5RZcA64T57rHYp9PViSJLdquWYsaFM
etk7wx/rj/4x04OWzd2h3TqfnilF4D1hXvDgJOinpO/7GdlOs6wayvkI1u7akcl7DlQhw+eFtis4
Q0u2awePMVAjpsu+f75JiIE8NLlttevSljN201bDjVACe2gX0rP312KDZSEHCObjhBW9JlvNV7o5
Lh2OYayDz6+tWJLsgREoINE8efChLiR5o5RVIpXI5Md9pmo4o7I/x0KtpbMKBEHOO0/+38tHiXZa
H5aDaAVg5vzaYf6vW4lrlTaJVeLNfKMSxejFoltzgvHYg2vnfMMhmrLecdNxEFkuz8huBnAvkKpI
yVXE9NKLewbDajglaZMiEz/BOYscI138FwbD4NvThEFQT1cp0S1TeeSpA+aCmaeDlNGsWqaCmK2d
ZhbD35nESoaNeVb19ZgMZh3/lB9mpdQY8KnIWeVzM1JcD9tPROEMES9M95vF8/JtXlDCvuiTU9hp
6dEnOuQxYq1eZdLptF+kX6VfayFvJRkP6nm1cRluhxEcPkm0WlU7djwYRq8dqWLksZFk0QEDigbP
VBV2ESYyCvUIJLxuTmchBwoAnwcNITZMc40Fp5SpNXB8p85lBCCOtfraoV5KZU8lZeL0ozAZiqSI
evvDh2Pcaid176vJEP/G8OBpHKKO9HkOVOVUB6Gdz5KCzCm72D5YlAJcMOtbi/GwLM1OTxjHWcIH
PKqx0RIXc3A2W/JYEvcEcLyC56WzTvV0aCbeTP2p5olEJe3ikNHxxlwLmm/9ZOsfGueNxJ0PGV9W
0PG9Ar1HyY8Qft2r9Epqf/U2LOYTPi2x6rikQt6utm+TvGdArTAmtrRDR8JhvtwRP3tHm2hy22mV
o33HOgc/U6CM3Ts7bqg6MoACEGORUUMHmjmA1oswanu3T/eugSpcFZ7hOUqKVMaBw4g9uj/0A7Ai
B0uvdu5Kqw3G8IkDuXdPeV6oXrsTySYWPttyjEWOfJF5/M0UZXfAsxekpJ6loq8bMxURk/BPmZVn
No+Q+ZrN3UXGt10yns5EH1HElYR7Mk3TKwo/n7248F02dfMAxQJufMer7mg6PYaF2PECAdkClxDB
ZgKNn80DMPKG76fei15mhKPenoNBZnyHLkT1vLaFC4AeCQxOTOOYkchYjMWZqhRqvvBKd6KbrL9d
VetnEcdXux8JrIXp1B4bugdO3V38omf0uvnGz3cHj3WSzNnfkxpaM0cwqoa+Nz43Xu9KjMQZsGcw
mktcNukZxvU1IL/3H39FYg/7EFHykh57ZREWvbNih7KUgUTIT6grj0GYqUCNJGI+XfwG1FdV7Fk/
6mzrnM/1rMv9hgdxhhj/1UQ17fx4i1Ck17ternBNrS5TnMb4ql6N0vIGRIK37IPeCdof61vCAhEz
9HSy3cM0NEUJ79a7XTL0UmwuqZG0LChRa/sfR5PuhPS75TfKKmM/1ZoHiY6zq0LDZmEsdjkbVzkJ
omD+oBQ+7aDNKFX3ttZ2YntJVqOskebsUjouR4JCUQV8Sa/4gcaJ0O8aSuog7bSJFZb+3vrVjOVe
o6u2P08JqVJEfQhxVSDMMwu6Tc4XxeRhAR6WU/BftXocEMsFJ1mt+fvGCA5R/WHKXroZVUMVU2wp
O4BLcRD8Lr39uZBdgDpHufbjc9jNYgS3ao/FeuENOFdO9dBMFM3NH4fi+8rBPFTQoDFxSoc077hD
37iLIp2PnMeG8tMxzweN5Y/z6ME+aKu59dlzHOVzKvD3a91N4Tqd6S436RFXnMUhXfY7fLl95TUB
ciafwivT2IhRazmTBb7hEwQVG3AbGRSdJ3/VC1URMCjPzyxdGN+YlshvtkMMcNV4ty0lvAf1OFOJ
hQQuxyXNx3DIrT3XxN+2ZlkqUsIEQcrgCls70vAik62QmUr2swHtQkD7tkT3NhHuaBxnnFqyiT4Q
7pjAqaQ0WyicEdW9rKl9/p+SsLzKGPxzx+It+eQPz17DIL8WcMBsv72vE7ZW/8CVxavIXLf2F74d
euUfd5KfTULla6TNp4ppfbsu2RjQwhXsOPc1giyA1csXxcKAq5Me6X5RZwoIzJcyiF+7drjhqvWn
LHbqGCwQRXn8moqyzxQtR7ZZ6WxFFCBmuHImJ+StqgXOLPHO3ualCREzW6chiZvFerWS8/uSPiBk
TsFUYzrFNCB/UoSFemLc58p3AQLepdlVrhnUHiQYtQZZ/x08jbY1/tMWcYBI0eKBq56kWPAp7kcq
pu/zAQJOVrxn1DFSNUla7TPHXKJ8lNXD89IKikkiotrZhIJozkSd+qg/CBUo9T9T30SvVuwVmQFg
YE1cdueHucG7IiUKkb6UKeUJeENUqMavomLF/Qcu16nnrC2HLr9RJlZpKgJ2e0kLIFxWh4CFSnHt
t/EFVs5bpTp2tR2o74PzaYwTT3Baku2+UaBbogsZQxdg2snv2pbc52BmlrbosXJpksSQKsNCLECZ
Q9iJvHdDP0UF+JsZTCUrU9+nX0mQpIakShRQb3izwWUH/2BdR1dy9m100IRAIKC1v3aUHT7bV8Wh
aj0SOrW5ecDwJFe9OJlk0QZSTvxNcOrb96Qc5DbZgbgdI9+f/u0zWjkTYLASPllU3hd9y1DBfLx0
/WB5q9EZkUgM2EsKdLZU/eBQJW3QHVWfYhZWdQR8P2O20hEv3A2Ff4/9KKjwJZ44HH5NpqAZiYQl
hlkY7dcyD+ow4R3fg7anKD8Kip4IxieKLFUOqif+TxOjD2mVVaw/nVaHkrM6E6wOCwigqBO4SfS0
qVe0lQiWm6JD/eVSGPJConfZm478l4IHmydXsj6pq+nFYCMbLKM3d3OrRG+Gg+S3qyiIbcd/xViA
3WkhkAr24QF3tWI4k3PPyneQ3y3ZcBtoYtaq6l5DNB4dgeU+k3QqBg9dp/qnN1H6xRCPl3ZSF4L4
E1rB0eKrGOJqHdDuvHqgaYowzn+9zxZB2STmhMDpyOweKHuSMvqIugTyKt3DIe1uJmAoY3Ue9F+k
yO8lIofZLCS3KvxUQ0Lm3i/vonLJYN3v48y35ndOuFTxWhbk/9NxluSDN63Dh8KhTkpcxRCt56R1
zzORM0rfjRsbyTbNNIx/7T+YVtS0GAO/UMKZPKKugtHT9JVmyp17LhnJbBUNnKQcHDGL5GGo5EvN
ZwbusY0ZKMnXHKOi7vLgXR9YFE/4f9VXedOki5YEVTc/D1JlEPgBwfTOXsON2xobxgCpD3FHJLbg
W6+ZrROPro7yNo3oVX9fAd7iXAZ0aC06mF2J6kRrL2g+Vf0qYWPyXFFiI54Onk6oCxCJo31Lkbuw
QCHqy8q1IHoOCl4jhbnY426hZQ3DNHRjc3zOrx+0pcramXy2tYlp3Kkvi5SDTOXYk3qcjB0fW0Rp
YrbKb528W8G/D3G1ADm8CwQB/jqKu231gC7EoFyU1eOjOkysdP3fud7JZNtQCyuSIC3huSVjq/AC
CuSTxa6ohfScD9ZhP39sDApuk68/Em7SUw4iNGu35xzcw6puSJCzQkUDTbfbBCN3u2Lz53+X1PKG
IWe03gfRsoNm0h3ZSFkrpt+qJFPKdwcr3Afr5nGhlIBW4lphgzpELj9sfPgnEbEBuhcWNsYalyOe
21KgRepqSjbMuEyPBOwKofi/0N8YG0Nt6zB09cm+uli22s9pSk80KxEPiobaJU4L0KWmrNkwbjXT
tGS4WGJESwM+Rwop+Evs8ARVwGQr0qRJ6DmmC/oEqO67cX5Wigc9yZ0OYfY61Kk1fvf57tlKdAiH
TolYsAIxkKijLSmw94Hc0h1DNTpo6/M7SZdQKxqE2ahpeC1d+ZA2vHFzXjLMTf8coXpxzlwYsAvI
maUra8i6XGW49JgU1k6PS4GX4ZQ8+oWLGwS0wxEdxfAvH6V3SJiHjimvb42WefjBGaSmGHgbpLPt
1HhgNNOECL60AQKkPM9BLsW01bzOPOQVKpt23xHs3kJy36iNzchRNo5jjfGGqM8RtqZDCTdEtz0j
TH60EC1tS74k+mMk18g6TENtbWA86/vFJhsYhbk1/w5Ph7ujrJZOAn3czkq/M9ERxTdAk9b6g5Gq
6ouUXiMoLnlpA1GBgrz5/xnuLlSeM0sbK6OSwapWZtJxa4JCx3wSPu0eA56JFUIHl23UEVzHYgwc
yotjDvqp/kCiIYJKr/UIS9nJYDdEH6+cFpT61fwzBaNQacIwKSHJf+62lbpZe4cjMzuPj1ip4PPw
nq6bhaAicdpgOcJ6fuZhbyMitPIeCIEW1KvNUzq/RDlkhQB1wsjTKWnle1iocCvnesTNmYmWaUyy
DMwa5tsTO11LXoYBU1b+su5Y5zGyfT36bmdtl7U/Kq8eeCSG/T1xqbb75WM2hm0qO85Jx5Q7W3e4
h4BIEzqjpoveYoM8lCYFQzrb++rfy26hXWXCTDAvBKltpYf+L8SnBUYKdG+56qkK83YW7HaBzbk6
SPpbLLVU8m3H+mTu+3ho5MHo6DFX7/IMc2R2n6OVzzQ3wLNnLl8pIFTaCC5b2lbpjR081k9YEyRG
gw1lMTpPqM44mRbvpL46Q6QkMshfwFI3t92hRCVwYlw50vJzuhLmi77Gc+t+DLl0OKH7bVy1kVaW
Iy/D0PBeaAjd/kW5VgUlleqEqQWpDtWgUsMZrS9mZY5LfOhdZrimPDfhfshwB2z8ksIHkkpkuSsH
kmN7sUgLqf6eeaF3ZsSxpZ4YytzD63NP1lFSYjm1ToGTWv9i9u3xftwie4mJJLJvk2QD0I5WR2iI
tUYt7mlkrsmLaO3j56P0J6ve51T5wnUQzsc1XR9wAqdUEK+JMw+8udVMJjzQE2jhjotaYP5PRDb+
QOte0a/Ag0LpxbBAru5Mv3Auqpnp3USp0fjaMCVpD+LeveJDASp+SScNKnQ6BxONRfXME74hZ2kQ
EY/+OHlHAfJm11cMKJlf+byYMNtfSx73N5sxiLU44lppMSdISE7GNNbE6gzzLmzQVO0yRu1jX6i2
3cBMGshoHenL5Iey7yPYJ6AW42sUratfKgdhxgDpbmiSZkX5/bbwUF90FOH9l9r8YSzi6GU0XoOf
WONNYcu3LzTfaf7OWigOswmXiJD+gyE/y7FxBsMKsuIKtlCpOrHIGh7yKXX1lKlUr2e3LUE9WXkt
xHU+ShTOUL35pL+THJGVFpoOAlqpyLW5ztE+yAYZzik/beDBLQAtbgUSAuaMx/E5VgzDxz02GZA6
VVo4DXOzwBbDoN1A3k368bEV8g4rO+Ifp2NfHgQhY3eSd7p1wRydQQFHVVOmS2leJLtLTWyf9poU
Io4Q42kI9kRWcXf/iFtQCwm3H7KyUghzxfdqXPWwDjZvPF/P05ZBl0IdkJ0EfHzYQrhfU/ES5iG2
TU8E/YmP0HaLPhEUjQcmjorXUZo9Y2Vn4CMpJumPgOZah3GYYZ4D5S0jnoKH/gaCxz5OmAFGr8+B
WXzdND7ja5mTL3ZHNJg/CvGAvNumuVdB0J8yPDXGmTd2DLp2sQTBwiCDtXiZwZEwE8sWfvvxCQO9
mS3WfW+5ZQreUnh/RDBc+SKSFUW2/ZFkXx+r6nhfRcf+WTnloVFIhNAx+8U/aAu6D3kCB1RUy6ze
FiqZmcqYPk1c5ODyfeMnP1P3G4DC4AhbluY1z4IAGMnZZzQRYyjjlXpLhIuEf2EfM7AyKlarlPwA
m5PCyvnHapLZD9V61UoOl4GSg7654Ezb0t/6WgzwwbdmYdugBnmZb4k/auaPiX3f6XEfz77OnovE
ipIfKN3GLCXERcauscdMrafHQ09v9n2luBl3iRNpG7+ZpWySp6TcgmWi5rscVY1hHPsmEq/62AfN
RDR4gFPybE5ti6aRHgJ4JaPfpguDVba/AZe9mpXessJgDmUTgQlYp8b1rpVnQ8JfLaQI6vXiVbep
rnqhspmmdg3ODUkFhbC74/Ji5wEIU+wIs+F0N8VVo5kT3UCbuOXIrANPy4S08bHn/1AP1ufpyOtJ
IJNGMRqQCxnUv/KRYy2jl8NYcNudTi5i70Ytr6HbRH2oS42mpgbsbM69Xe7HOocK6424nDE/RRgH
E+xQcLZMxqMEPNrHRfiu5BU2C0N+4hivdGY+aoPOUrTga8xlb3/AAY3bvnI7R8gt2Snk9w1nQgGT
NlIiAUrkZESfVk1phfCQDrMKlKHwZeCehkzohO4wP/9r/bUUWnB1+W2ZMGj1yxgRpoWhsKDpgdp5
tgyzwAVT0ILNqPfJJXyCdOjOAcQ/eNjMbZYVkf/62oUJnwiBg4rKEIGmk1G3s50iGYV4PWSIJoxE
y+boRErKtfH6neKh/7Vn+hkwSakQobd4WpwrqsSmkPKIZS0cPkONiR4VQuVsmfRZhRH+8DvWHYjG
SPw+IAr+WAPO7ffXs5OqzuptXxKLA+XCAP4kuHYgdlWDji0AQMmufZdy2xoMB2N9MlQm1sr+6dpl
EYmootQX5osZ9nYqU56HAj7vnk6EtOOAcFrs7GbO9My9KT92unnkdOEuvbhn0GsS5Es/D5UqBexU
1Z89bTwKkRi4LOjCsKXvanMFUXM1n86o7iFYY50JKtMGzfGQ3LmpBgjfI5eOdsVFWNOk6sLBCSfw
Vv7AlgZrdKjuoIUUEbfaAaFqBxEgLBYIatinTYejIwYjf/YGS3m7WatJJwk/V0rkEAh937GLps0m
fE/TuN5zF6VBQ5wAYHa1QK/JP7I53KoHgwFx9iiKXBlXDoBwEKHsOsqAEus6LYPr/oTFKrDTOVx0
c5Yr9Zrketx/tCT2CApR+7OPAbQ6VJq8eIPrqP+f+H/PBN2qfZ6dK3wwMvBNO04Sp6Dfq8TVYK16
ijxGFVup0N9RIzC6Pl6f9Xv+Hn5JAsrqbTK3gjHsPJrDY+kCpcrwGq1j0HFsDsk+fOYyHMxQiTha
St+l49ZX/GwuagS7fQSzU0l+TleAY6N/wxeq9+HhznkCTHFPrFwnmzOvyY+/Bxnubus8F33y6hNp
kx5P1MkB6VQ69Sdg/QyKDSMZfgAIxcvjz/1xQVq81s5Qb8SCgZKsZ9Kqm7aNOTMPPCf+Jsb2TVw+
y0bkYgrtYw3ZRfFlnpV5k9z9+oHMxusjRxplTAQwVs99QVaYdBVqyq2TD9JUIMYhpLQoJBMHVe2i
oEZNm477hyNUoW0gCGfDBu96d6U4k4IPxsPoH3OWY781TrEvH/MUgUyWWaU4bSvgekORumbv9IES
WL9hJD+XbrX+b4HQgrOUIIR466d2lFshN8eoVxAsBbYdg1ilSP7VXp3i4iO9nWf9zslEJ9yGTcRx
pKWqLsBOMbvODveIVzPD3Ox62mMN2zGZheS1fU19l2uhczVbIptiKwGczvV46yY5ENzgSxtZC3pP
R578F2ONBtztBUxd5ewSbdb0SyjuZL9fBqRWVlZS5f777Gwtj062EzCBOmJgwpPmpg7vt5tBLDIv
uTEsG5pBF9PC+CdR7KLJBeS/zhK28g7TLxqoadT9YtsGloj3qvdH6RWEFyWzmPj9iZ26tykEfpUc
bAeRCTZToCn2mAe6WkmPQrVwUqkst181e9+SwK+VjX3KAqXA2/z5S3L4UHgVTtcGr7zzPrpuVoxu
DmUhTJksl09tQAYXYwAK/rk2IoW0q26BPcR5SDS+V1pcZeRvCR7c5q8Ozh3tcJ8Q05EAskC7EYDL
nluosrPKonG/i1FhF3+mQkG4CWWgYSjs87lpyXHDxkcd1oS7AnlifrK5wMjEi1ISkZr/D1km9HgK
0KLoDRiSvZBLrfwrdIwZYGVZ9pwTcYlybkYxwWFaQi/diOi4Z1wEtR2mIdrXpLlqA5LrS9RuKbi9
XtC3K6M6TfeU81e+fR+kOCMkZI30j3UC8FTeynW84eidh35qlrjeGIAAsUpczVsP8gyIyVTzkgU/
/Bu2Gjl8/GNLUEpCWWTk3WFm1+q4+12Iz6ZZllqNgmYbXjmZ6dyVfyxlkH5k/2Fcs3xKnWy1TKws
a3xRhJZ8PZsuwq/fe6VLHWpx5Po4rGcVm8A57OjegW00EquR6oro4HDePyE2mECEzWL5+i5ar1fX
w+DQ2GfOJA0qGG9Qbe3J8u0HcL1DUElgP3OrtGwEWrTmDZuobdUecBnqpw0+TZbplXU6JKM3WOvC
TcH5PrUNpIp3eaf73RLqanJnQTfWuqHAVVnRd/QqXinvLbvZ/PD7k6A/bQEr4laQs8HQZgRkCewO
AqsGPnJ2y+5BlwkIjglmR5RI69JpbrRmV+E7cdS9Nzsj0ZL/bo94OYw/M6sVNWD1FjlXMnDbI8up
ULKG/FpjgoqRA49fHB5mNFgfwxV8aluo/BXh5bgLWuH064+WBRoJr9iaEah3jntwNlZY6sY5BpUn
GqnGTTLxnidgAuSO/SyeMjc20Vqt8swmHilpZaUnsm2H1ITsRjLOt8sS8vD6fp+QaLyqRcwNkds/
5vokg/7Qac4HHeOHx5UxQbzuGxkVuZp4/lFaIqSWGSeKaP7oYGwlLq7EpU/CmPgPtVMN5X/Ko31r
LmFIN3H6Yl9m6AEeqd5KKdNeKi/MsK27nNsJLG4KhtE8KEtKZhKcZ6fXB3zUyPy5IEXjkpZyKzt0
aRVbFUxg5iW8SxIJsBg5S+wKDOeGLw5fU0gxEvEoTmO9XpDi639YKhlWsucYXrhoQZy9pELj42kn
ek7+8bEwxfnDYXCApyKpIOQ4XJMBm6Yof6LX0U2p2rzzrAi66hn7luddM7fF4uUv24qvT/52Vecj
IlwDNkafm+wdGwHDpRFowGE+vGkRoudxbp5ATLR/mMC9DjithLGS+gOQ+TD+4ktvgLSh7TYhQvnV
dGglou82zFcWxZh2TDO7ez5V3TjwXU/6BraYcqeDvWcJmly+gFE06alMW9jwpZpML6pHUtzgcszs
QI8SorWGZUAcZ6edou88ZCEkYi5NxhzbntMtTIyocdkwdUU2G9qtr0oelSCaB9wUAgfzNRpPLEFH
4en7HOF6a9Tufs01tKxISiWK9QmiCzYYorSWvpaFbobruFYS1O1JNDQoMqdHDH5Tn8pHx6+KlKUc
o0N6/TL1tqdnjjNiFjjJOk7t/FsG2fDr+qDpIZ+1KNYQI3+4sHgHXsFibkYlR7GEi5J7tV4mpR/3
gdlWgXucUB5PcXcHSDFCV/sBVpGnGys4Ty97x6nBkNDCLCUC25IvjgF10U4Acca0m7ti2DIvpkZA
PCf3k/6IJtIzeNBtRMSCjsztXztIpRVCByXqB+XVJGr7yCrBV8vOXIp77lFepvfjQS7W/yJ3KhK1
X62XKHjktH786TeIMordX5pnjxcIX73r/3mkF7Ga6aj7qLUwUZjrLhVsGOZjhTetiT3YnJtpXuxV
ODRIPudmCpMgioYqMb+eFo83aMKd0MzJQ5xM4KH8nOPjpEqEIn8kY0Ykf/9WjfK3QVFScWPseZWQ
Nw1VBVqAAcWOuB7ecYi1uSp7st7WzDBcL/mskUpttShgDs/eaU+4JD/GbVywckiHTR96Chz2gP8p
uKNIkgd1OOZyvJAu2OELgDA1Z/gRg7o2INPEV/p7foG4zkpvNdtRJbN6VNYuiwMDjkRg7y1DJ3FC
HGrhxJdLtIXZ5FoOjgMU1jzTdFqPxcJfUIgEEfoPNS7LNTDgXmjQoJwN4FhnTzP1RvQiF7+bB6ks
w234aNs03xz73LoYRzhvGqlMrn/gSwuRtUOa1u7s82YBm6YAmQsccIZJAZUQp+3fDkuWBI8ECRl6
hWhP8+rPnBxxkok5izsn2souJgGH+ne0WA0/bNufYQBJjQ6o1+XLEQ3rZCtOP64DEBsAfJymprjv
atjU0BfthQMICTi1uXaIiv9uEgoQuRvTSXBC+u9GqynhHqJt9d8xaGwWVPZdOh8c5dyuJ7wLHOik
qk8InV0Gv6Bmf+y07oDJ6X+/IFQsZ7wrWe5fxPeDcUzvJY7K16ZXhVOP9DRFqsDekr/5/QoPWGqe
3e8QKvv+pG1GZH4eUIXCHqqlnBCKzpIoK4Wa7xJ/iumAB7epnIYK9lNBsXL2ERcVPEP179lB0sfZ
axB5xgwdWIKpdtTEvxrGL7N4AEo2thRzNgu+3WDFNomzTWhG80u4TXDfKBD7E2kUYzX4Flcs/QOV
5w/pqzPKNOdOhMpucR2xILFGHP9WpAZhRm6cGByUa8p+z4ZncmpF/LOCUxeHnRnBGCEv/MQA1L0A
wFTzVHUX6BEd6NIPsbzVvskW+elIkhfc21Y4FhhjfTEW6Q4c7qlvosFGRbUeOjTVXigPNTJ0Afgo
38EtVF9nEC/DqCbtRVYnMZOgwgVgA+wK7LNVLla9Ejw6tm6r5FVwaTsTEBu5OQe1B7V2cc7g6+Y9
aecPC4sTFyoe1h+tX2Tfs5B69cd3/H4hJz+nXqZjrY8yM/e1UHFVSwPhOU6h7vtpIZyeFDjgCdB9
cEveYz51ycXLlnE4mOWiQUugX+XYhKvKOhtUVYoa3PlLR2+QOYh+M9yNkPfiWJpCOY3o70cwzuu9
SUINE1/5tmDbL2VWaEy/uONc5iA5Iu6H3xKDEaG4hOAFJ+enJ5IFzC49Sfz47mr0YC+xjQyL/tkS
fM6fmJNz0fOJrax1VV/ubgyo7DP2+VXg8MGEETVpoCpdTSBzL7LLS4uzThJnWUDaT0Kf7XW8jFcK
Tpv2NZviOBpbr6GAf6z1UEhlfbRNAGbmr0Fr17fR4dWY8vmdJVcxJ2I5FNWSgwmj41S34GISe7PB
lOwuXlzjXQDXd80d4Pq6LFUXPztQTFvSGyD04zT0/qh2PaC69Y0Rak6kh0v/c3DGMkaEzRZj/s2e
jXgO3ml9wCe3JfAAqiUO2cabZZc/J6yyxsseZ/kBuwn9ILoY6PX2GL4rqbkq+GY8n7bnLfaDAIP1
yvf9Y+SDcoGOov6Dy72kzMxf5OL7gOZlYx5TsPVsQ5jRdCu9Aqs0gVFx/Qs/Uk8Q4xhJMclHyqEq
giyXqk0cahvEO1CV8kXkhymp7MEp4SLmTTsVUvzDaATeDQTSvPPOkGAOTMDgPZ1hYH+KfE/pRSD4
8zZN2HwCc6OX3DsBALV8KOEg5o8Cicpqy7QGu6Sqw6wAJqR/E3yJByeox30RN5xVypSJ7CPSZ1R3
+DoUGU8OEHCe8HQENic4Sv/tUqVZToF6g1mATt/hpD06AZLlC3zCf2H55KgGFVfOJcX7gxNQRgLd
W9cM1ews/5tnG7gXTzYJnF3qIKmpvE+1uHIuweasDuZa4oltjXnhPixc68XwDF/SqmkRSBrUqqqs
DuryiiO1uGGJQk+gamMeyio0ngeRglLiLBIPNH/evL8dWX4zUvHPzK8sqMMpjCYWgHnrmAjZURFr
fz1+ljuBBn5+ONNGXJtJRotvuj5/g946OZysIp7JAQGvZVEonoSXa4CLmvAwj/VnzpHrfaYWjR1Z
EXQAi/GCjqswpGaRCjwDY3M/G4rgnVxNo4/aeBWOxekajhmdYOZ/1BhcQ00E8edc7tTW7n+SAFEH
2Cer6qrPYA9KrehsYNZweQuPJ4OfBjsGbFYwxjuLbvo2qCpCySJYKjnAD6LaQEuIecfIX6AM2sqd
tAHi+cb0JX8qnySgN76TfV4qKMpBbonb3kvR10JgQq/Q87ez1wyNWjsOtBvrmKCHQlEdnKTwoGeR
/KOqU4lCAkf0dL6HtcIbHQdGaqpGYCvIjee+5IGoS0cbe51LjcYdlEHxPLiluqKHICM6Gs5D/nEA
pIPaGq7XX1VUGRjyuxtrGTThulJb/xowD34Ja9IcSn8TAhVVOY3pAgLBB5SjKNsOreaON6rXPmUC
V680rvBDU5qP0C1EBy6Zu+0PukTrIhZpbIj3C3Worhh45TmDdseQlWoGmib/FdTGIvjMGCBEJAPG
r45zXSiEF2Rqv/a7fHftGZQtxpq/xf8b5qS+aKM3gX4XlEJ1a35UrYu/x5yiFSRBMsaS2rXVY72G
Stc1TfyU3So16zmlg+25dygDk1KmgE6zlkTi/HqrQYf/cmSUvtmiEk4VP+LwQpZtUKfJCJzT33q+
imYrG3PMDykVSwAEcxLR0+e/7iL5H61hg8J226ZdKIoT9Kf/pGL+agy2lsJO6nISdRhxj/7qCEhG
UT8dzOcZ28SRQ3UDwSpc7rBb9f42sW+nT6GG4htxCQCCGmBAt6TlUoqKiJw+gmgpeCfUMzX0GZwD
F/H79MP3LzTT4dIUIIJ3JraOMNlNm0xNwLut8QAZRJ543nlFVUorBstVBB3VEXS4nF/ObHLWn7bm
6UeXavLaaEx6aiIXPWBmMmDv2mmyhrO2k0pw8C8+yCOB6gF1h6cb3CNY85rE9CTm1frL0ah3xX72
utdrJ5F9xv7qId5bf3Nc8GxL4cNXxrGuG/trKMArdlNykjN2A4GTUiVmJY7pIi4dkl+BMXGzSKGb
qgdVc6shX9b2QfANaaQzYb3hz1W8JN3CpBOLjhfojS/ig7eAeQtdAomTvaEBRUzno//IFMMKK1fJ
8nX8LstK1Y0pO4cPtNB2K222rb2YpS1wojQfwknXrnxrP0nGRqofb5TUGM7BygDhRqV1uZinrWpi
eOVGNXHy8JkzHK5O399ydctultw9nWTakCBkbkabaWE6ujWLAckov+XGUneKtamKTYvt5YH6ufXa
HkgrjFiNhRWeGJmDMa78pJbxXT/8fD0ieSDzFCIk9Mxj7NEekJrq2SHQqqXy0/nRmPkj6FSZmRbS
TllsA0orlRlzbnxgaCMFrtVKG26VUtlcn27I29lr2NuJK9ASeDDDymcYdbHllGJGs1r7lElm/5XT
Gzvv4ES+PDBS79CwKXnFQLiD6quMoi0OeCwS73IzwqYznxAtNmWAyDiERUxn1X923anNzhyFDlsT
baV2qjw8BK8mJhckWMxLdNZbBJkDqBkUL0d4q940GJn1k8HZm/aLTjupKktO4a/51t3o76152PqR
a01NIMeT5Lmy51Zmg0f9lGdaYpCzET3kDkZu3ruCkSrzJrWI7dDXbecQefYqA+3XtastVZ29w8He
ktYinWsxX9qFBDxypQan4C36sCFWqMNoVrsQHUTSqmzVuZn0U48kwGsF1DABDHAxoV8Fl6jnIAxK
UcAW0wP3W3lMmOFE1zWpOOeeHkKZ5uIsMhhegCdLDsz011Gu1aa+YXSnGz5P3L4wJVK6Iv9MFtSN
eeKNtd+5by1ZUd8Jrr0qP0+s+KRquZv/XUzQ3k0ptjsY7zaq27UGqQkR7ps8MGOf8Mau++bMYps7
Ij2vekpvCJX7GwIhoOz6l8JjDYWS/1N8ot5oosXu7h2Pgqq4cXsj9LM2nsSZud4Pm/5zbsWSVFpw
qG9qks3K9vd5eXp3wq0euzLd09NszpXazByDj5FAqmfrtOKVe498tnRLsWaNaw9j7YpgdrlxE4gp
NNKl3wZ19Z4WbPnAeC+VpHw3QQ+iTY0nmt5uHcNWEZ19bLs72Riq9739tyvEBelX+MULCL6S6Blr
JpvNQ+KrQ5wPZe5uNTSOb8ZOL0tohwgx1hywurbig1EiG3VhUZzfyG5Qnu7zyznCAtPWZmVZxVpb
wZMdrVyax2zTgRuSxumau4TJ0bw7dkFIN0MNE5sY2mBFV0B0hP0Mn0opPd4zq+FVrz2Z3A3u4ZWm
iOmeaI28pNoz5SL0kvcwUcE85XBj0BVhwr1FTJhQPHdsGEDmmhS7j+Vg87u7AXyou2VTrqoU2m5f
wx1VD7SxIcsgn1djXhDCEG5GP5aXJPQ3C9h1HmDwvmktN5mY5srxKrPxf7fK2M0LgL/vjSNupiKb
waHOpOz1fyl1SmuFSJsPmCWA9BqPoFAES/ciI3VCWIGJNEqlAQJU1p6xiJR0B/H83iQkyFP3NseY
wvW+iyG4YB3DjMTwfxGahpyrV0vqlCuq8/Gqbe6gybYQM7UjiDOl+tfsOOAVCT3tept2Xa2scG1G
Z9tmiQ9OHCdPyc9W4zV6L8X/Wae0S627gTWkBlT5LEgiyo0qhEVkOU3c1Gn2W+cVoH5YZiFgouRO
FFbnCFW7kzz5eTWZn0oV1Hz9AImfuoZB1SsDrqmGqYHqEDpm/HQv+5KTJ1BHidGOHEFCH8f/kYsV
XoNFAM8TLKEcvYui/nkbubqMsDyOBlTyd3WnI2US40YVS9lE5I6Z/+Xr1fUPfxOoSdtC9HURt1zc
9a53vktv3PSCKhrAungL2tybK5cz2WdchHbunXnhsDYmV9QbayYwkHfIQkstRhfvZBUz5pIhShN4
qlJMeSivVH7uk34Rv3lZlKa5jLjm38kOKGYnhvvnKHR2321momQ0DKbgbgi5hg/cHzixOX0alvWa
KfRuiptm03KHrzYzP78pn9O5vRVrN5/ZYaqiKhJsaQ95ex1jyIVyAs/ik9Ycdea5j8FrjmdqXelb
y0pmHRBxSZnscOOinj99ZxMB5ADkDMiBo5OmTWR75SibxJgPV3XU6ngZG5mkJXN9JLRs9KpNcLCL
0bq5hNl18aSXfo0bkcU4w5fKOX1AKaxE9+jFcAiO+y5OrPL3YyU9r2/rgtdGXYXaCG3Z141AZo2Y
qPUpTbfIK6wFYuxSWifC3pQuVCGQfPnkAhNnDwRKKpsHCqtbLlr1BMFerq4R9WAfHrXYJ+y25bcc
GurIk9ZYjTNUQ59K29FWfMaiUxh543QY3/J8VN223SbPnIdb15ZL0a4C9L8RmB6WfUWmI0hpw7qu
AYW/mtgmE6BkeIIWS7peKhNchscaTgHgC5ePFSM+SV2ztZJw6D1JhxA8/vAtnoD1QV17gUirXkYG
UdV3Zusvn8wbIM2Pf50PTw4oTQIw2C5nHoDqLuy52bLA7yXYpgerBmH2lo21mPDiCRG1FM+JaEo1
2sBriiqEEFnrIQYuCpB/HApvIpHbAE8tl3JZe1uYG75AInOoijBM4i4RXmJAZkHDxZj3zYdVsrR6
To/yRldQmr8mhpzFlrd78eb6/R/GuOIDl22z/zKOevVz4I2DFZBCtdX1pid44oOp9/IJhw516Ui4
8r5SISDRlFHmQhTfdSdbDD7S3y4OY435Ot1KZGcfzwFmCHkU8B3emUcSGzOnFY2SeSDventncbWs
tLWN0MkzxBsnEtb+moHPah2WaSWyTLEkA1rJHTRZu/PfGwc7U7ABGZn7dZRPRXEbLq8XOR9oN3y7
8pJF7ju5WpsfZPxtvzIrNDeK9yRe9v14duLjDMp1zeN1wsxACHRUkJdaaYkYS0gtZh3KzyJrGhzh
889zVWwyLQI9EaTM/AeRhuU59xTIhiVyjy8BH+eXC4eetUQlVqKho+Lh5f8i6vf0D4jRz0tya6Ix
j0R0ssJs4hh8YJmT7MM/wpE0L4iJW0SnDZ8iCgd4aI59T/hqyAZZmvSZFOYBKTmIi0W7iofNSsA7
h4jiRfWfajO3bSO+DU/6jBgcNPuD6bfY652Q7YjUEgZrzTmdjSZXFUTK/aYM5AGhaYiWt7GWpLT+
IHm1N6vC5YCoRImOLTONfsy3jaknqx3rEWnAuzyG3i9jwLGhJvjPVGk1gsJzfr0dCK2D2wLwuYM0
ds7lc0umCfGr1zfze+HXtbp2xB6QV3744fPSYTQJA0hMgyncW1FpzztPWRWFKB7a4YHCLE+7VNWv
sIYv97FdLzhrGFAkYnvCwM8fWxVQxDrj80kb+lzuPEqDWlX/tS4s56y3PEtDC/9erXUkERBOI76+
WiHMFrCf0IeusQB0X+vAaeyUFdUlGXPyUU19MNAhfDDrvMtflcyWosfm2wtxzBJQB9cAk3r1yQ45
yXxQ6h5yXNOjw6QTxUFVBsDui/eBZP1ZgIV+sA+jN0tc3trL8dKn9uwASp2YArj8i8TceX4G4JV8
1X6+Eod1zBMMKsF5pKE/OFaXqCVsf42oRGyBQVZn3phhvVtpIziZw/f2JwUuTQhG2lC0QkIHf80D
04leal6RvqhTKh+2HJJ9owUFcemblkZ/ktVwaxnN4rTC2Dd9YRRbgtpTpy9ATYyI61ZEmxCerSVM
8R3hDpmtMSR/y7kZ2to0NtTiG3G/jrAy0+wZocwNigmBPwjaUtIIVWwl0SOx5ptyL2EvZYTRejwK
y81nx5VrdiWNMl1xwjZPbkwY+RLEe0y8agbVqKsqU6ruxVfpU3iZIiiUWRxeJ/ib3nrrgOVW26+Y
U8hV2jW/7808/9B7rprK0H9t6yek+bIlv+ZCB11ghOEZ+QntLOwYXRNYM7ZChNdgRZ4s8Y8ShbBn
bvt0R/ZkvcsFZUkU3o+jxCwQqDkoICsyVRswBRFUXIoEuAe+Iq19VfdRaxuSPue2w6PXYfvzMqRZ
elgyXj6EAgnUvstFXBj1NyhHh7A0GHW3B3p13g5URSkDOKIuQfBKZRbBfKHEEfFczryPQ6QQGXbc
O+3xPxfbpgX/aLpNQYFVyBna/JWyFAIptIDuotlygH7bG4ua8NHGEeWm75Bl/WhjrSV4liLEFOpk
0iRjVKGJavCPztsFGeAgtZcUc1PjbM44AmFTvBj8DVPqKvVrnH7EfTh4AfTXrMABkRfSo40kvcf3
ZPMgQgOTQtsnuycmVTA+s1qyJHeiCDAnDb7CxNB4xOYyOYnZgM6tPbPRuVRWupMerE+pGIirKT1z
Xbm9Z/NDBvVzJK+UqxLFnKqdqcl5aPKjzV37PBBlHpZ9mfvOqFz6Wkwuu1Qzmjg3rb+DtFIGzZ++
8ZaQKPVQPCf+rp5wnW5dAD35vJdSQcWF0QhFz8ncttXRIy2QuNvSmkXnasRTRQ3V33m+TTotvaOl
SUf/W7M9wywS9GqqOhacZZp0M5sf5fGULtLhtCxMOTIXgoi/YtTA77kRDWHuopXF/W2pgggccZzz
NDYMQOclDR0xzsdeoTNot8TSaHpSR2hPua/S/HnT7L1FKQ8CBgVrHa1MhTEzUCyRGlsCGV6L4C5m
PwUO/9a0i6N26zxdKZF8zIF7r4OiJyN1+RCvImz9oM2XIjnhVFCTYmAV5QlvawW94uHq8n94SRIc
XoqWQyBtKzOE3/ECbvBmbwq/6EyxASoAPAUndPTigLzUOmMQdcIVZpDRfQON7AZ149mvxWui+jlN
zt1S3tjfKGKGyarndiaSyjR1E6vg/AqgvXvwtQbJO0awvB+mSS/5DaUVcVqaaaCJ+bdA6n/CwJIZ
6yXkFjEs/uQLghvAl00EDo/UleOW4Ya0TKGxmXSuHTPHbZ/5ARwBQ7cqgEhObOFPSHCoUsPkg7Yc
IsVXY2V+gHCP7TAuLSZ3iruBHNfQIjCafQ/IrwURgT0/+eGdPFcx/FCSOfGiAVtA8qACdSJgCgds
vCENFhchdjF6zWTyBbU0jVzdjaEa4+XeXfIQMkfoMGfdCzz7rmVwm3DIF/m/+yYPOF0vK6hMncNA
o1kRXGkkn2xFNgs3rAo0bm8T4Pj6m59WpyjXA6tSUGaUx2KGxiiK45Z+V3UQLYjghlOO5I1ZVVuO
cpdtKuSXDjex90Q2LB08Ta9hlEL6bjg3N8Ex533osuqB3O5MQZCT1xaJnS6G4lPnqWMmNav9sFyb
6fKCZ/vEmguCtpL1EUe/RfI4F4LDE6fNgS1gu8u5zr7DhlJoVgGFMrTLqJPHCfTzrFDxVmsxdTQo
k48e8swihIWSeLlbdaB/jKfHyrDBI9pnjuUaERALurD/oN3gN1mo/NbeGAYI8Vy8BagqwC7p9uCP
LZMLHVMN9zlZfcwIulB235FX0vQC7+Q5I4+zt2DoYdkscUEdo7cKPmTze/r8VY5q6W4DvpvuOXq1
VzsHZp8JkbjPRmala0AJiF8JZxWNajPrlu36lpKUU+pZZblzqubNzlaVpDzH4ax/QK0G4iwSLLkP
/AUUGwHmtWOioFbC8QT4QBhGQxdYgB/MTtLVd33yX2gCb4/SyRLwQ4fJkB38Mgn5f/B9eAFmmyxe
fJjbnnDuH8V8kGA9Y8J7gsael0Tpt/0IF5UnGWUk80o5vQUXx97ie++qMQ54bgUrE2cuZQKZeXYr
3W+8+V5JPg9fklP2cGsd/S8glYYT8CQzP4SldwUznCYKmynOcEbNab5AVN27OAKb5tUgKApu6iXV
BGrJC0wvMnN38VLEcWLMfsXM5nETGOwg0Ixg4NaHMpBnh3BMMmOvhjkc9673CrENfIFbS0BhuseW
PHYQ0hJW0qzX3dsCBwIkDGpV4EyvxWp1/XE/X2C5glXfdVRqXs5O6rsqxeh/VNfbFEx2YPncTWiR
moRsA4ZiWhCnhzHJA0kBiH9hPE5Z+4kpfef5D2KZjFW/FwTIsy0xVqihpEfFvHjPMNbUIgx6IbFv
k8BKDxjgOa+z4YoG6Ild0CdIogO4//EYl9sGNevZ/aXKRQeb8OqCB3EjusXmk7CF7gzCZCk8yYeW
NI5gKm3xTw7Z3GjeIExu+aNFpeyFdwBaEoTAvhr1KlJQJiQe9aO47/uGG6j39CgdClIvjPSxGbgf
3s1DyJy8IHdkrAkwqesPXyUO8GZgjMsTBixuGwLBzPuVyp+1ykDPMalDqS/iC2i6rO2Da0h0GRfB
RlhGUb6EOyTSMkP6rNRmXvrS3MQ7gVLPkS9kZb5walyaTgkzRiZidtp4zlGCc47qUsTC5I/h7+af
kgJ4mAyFloUTWEGyy0NuCfjKfpKLaLNU++cYSV1DnGjlQMPcnCABPyGIhfwWBw2KnhOpvocDsZBE
+7kyHRDGKlyONyZKhVJx1CZZq0LqZMW4pjcmlUEBuYp+zmMCq3QZU5lh268Q1ojWv+ksaS0JaYOD
tSYRjDZjeiIBxrVa0feaB9az1Rjl/nlKqjB/7dkxVFQHFHbDSwm0AhQ7Ioho0S6qrLEpbiROXO2T
ezLSiRHV/sgXhC7yhPeH2odBzqMWMLV+2h+Ayzn8j+NtycZlQRhYikiqNoiwfpTMgY4gti+ahMt2
Ee5X90Th4ku/Ncqyj0huI/lrhO1eeOYNVIIk9X0L4BoorjnZTxEUydNQdO6tWB9V0gR59rzWHcDN
McAm2ceA/3TirGHoiSrIFjl5BCX9nD6BXUfZmRe7ArshtOKdj0vlyGLpaz01Iwy8ERHXl6ZZm3l7
ch4LdANUcP/e2tS8LAvwcT6Mbbpzm/5qXPQgIO7hSGF/lkV4WsPfnkgrfdNodOITr+FWzfspCBfw
oiR7cZmx6BAjRAQ5NJH0tftiuEg5h5Xxqjq6BnE7pFQd1dervNrzbvdVX0fG6k0ke2Onb4ngLCR7
ZwCAeAFM6gDZFcgD1eFZHFyvZ2PpDUeEt6sn0375zzifdoBBQHmN7ODS28leAtGKMjVV0cdAmE0n
1cfkyh+OgLxBceuW2eQVkmT32wQfVMi9FJ6MxKyYF9afzsae5tLFU66F9h1FppmBVlmKDjNupSzL
CZJNe0ka48QTU/1GxbSi7D2lxCXvVReGEyggmIsHAK/F/9D2x7OxzjQoo8N/zXG1Lu92CQRjZ2rQ
+uDcaICzeTen9rUfjDj4/7ZAJInf5e8y+gTKjHJAMCVfxtIZawVwjLHNFDXSBSQCrvUohxJP/Vrc
Aih0Q0ucluYg7rTH0hELLKbMtGhcTIzkE6Wfmi6hxc9sefqpjBnk7scjfWHVcvCqOkmvcgLWrnsz
q5VDRqyEjJ+PCB1V0uVd/5Ix3ywYjV4WoC9Ce/PCTLdwh/XR33k5a3FSgnumKzkKWjqib+qAEhgK
MGmjvjHdCCqBJ6rlAwm14AoM55yvEP1tYedkVwVA3bolFby+2gW3Yq+jeleEyq/bzZatoL2uLqLp
8G54kOxto8s2iVEpwnddsllIzXTnT4h3eeDUnuct+VUHfw+lvbVTlDtMQuMeloS7wAEfuy5li/fz
e5YnG+uQ0IA3xU8Rc3PBmv1z6Y5LWA809qukKuQSOsalmQXOKpoXQ5DnGLeWY3Y9AgqQYrSBVaGF
r7qd2i8rSvF/upu3RpIzEyOC3CSua515958ynDASbg72COR9wo89QgaEfVi9+ObhBrQD1C5oLJpx
fBrshAXmS/jZSNgr8IfUiPresFhKJibP/ApNHwjI3pvYPHsp72TXC3OxxPWdi7ODSYlFj4htK7io
86vMcIk4TWS5ppmQ9FOMAFSfsF+2sbjRcr+gjgjnbc+l8QjuOzfTip9AARTn5uT9yiQ/EsK3k17x
+fbrBo8dWW6i5Ku8MFoStWPYzG3n5+gWRqhG1PcRvkNh8/iP+ytvzbRvm9GROVtE4YIjvZe6qMFY
YJWn+T45Ku4DVn0c8tBEBbOeYb1py/odrpX6KyuhmIN8P83eoS9iJewB9fnyq983nYEPkecaiOj8
vM9sTfXlgeWvrBa87uTgSz8MLQgz+DFarEaF4cKR9CzJFEAEV+iC8cXlrXTjRqQSTAVTXISF34cU
0fc6EwNndmr2PwRPlPsaOAxGsJTRe9QsN2aS0JGdWGxk04mUE4z+J1baCY+rv4Cb2XbR3GEFRULG
6YI5lIJiLs46odhTGmdbI3bXtNPBpmLpc7pcBZVt4olw15eZErgJBxpv8usP2621Ap50LhK+6GkK
Sy6zrekZLGD8hyP9iwlGTK1N8Afs5QcQJlSU4AHFsnG10I2BtavHyxgSTepOrWbHgD3IFdCS1xp/
n7e/8zIF1tzL82ppdchQsYInEf+FmOOt/YlI/eXhqTce3AHxgvn503i15jhVHazFcUr/2BMWLtKj
YmGGFMG84+yTb5dZIfjvG5hDMmTwNDYjjrpSL5ELgT9UtImJlti2spT4Lh19lbaBff7QLiqhOAml
IDydZiLGFcLTxbCm675XXfMgVdxAvjzGQijrXQPdLw/ZX4msb8PE40NdQcLAXt8FIEf9Qr4zrncR
5zs7QIbVxtJ1dBIcnfqczuqWgPfcIkRlrobMXGKsEGCPuVyteBn41LDb47kg4oDW374b0wCGaL/k
YOUv/ARClNaleVB8IJZrwXQiiC0/nCaWCiIDdk09IjcLxpPPQUIAsVZTUInkHTtF2RC2fudfIJv5
O1kWQTZKP9s2HJsAsd3OJXTSe53smYCn1Fe3ynecvE/trOXSr4EHMCF0HSJs+Rn2BKg4C+m361Md
uDSbQjuIp1l08tx9nRdZZ5xpinXDIyic9FCrGBS7VHR4lMeF6gS36aEG71o6in5Hak43Jxn09W2B
Ab1j2xl7VeAeHx65W/D3L19c1mWpwToZ245a17oCld196uRdY6bKr8IN1krcAXC5wiyUs8MUX7cV
sBHMd/IqpWs+g4EPBUUG4T8Q4EixJFhV9G4tx/MpXNbg/A14lkvf24hHklBrUm2MmSyfQM8/8mEh
bynDFRSDAgA9XqUumryKY08rSvpp3PLGismXOQaps/3iZlLCOn+4GlKsQNxfy4KXPuRry41KK2EB
rqU2oYvJZsKWlYEGryu7YE22YRy7frQ4q5bHJFwTSVfWEN+xeAHeWlyB3oDCKKteUTdns7t0ccd2
HCNbnrr10uj5GFkKizgKH8CGrExD/UrV5mSL2J1v143xw8afn3Tcfz0iLkYk3GpI3gYnxc29BHom
IFG7W78qCXnx19MSHcX1a3JEXH/J1yx384VIZkmL4MBLg7FPEUKYPj7OxJpvuP9zpaI5E88jSpI4
ASDc5bNEJwFIuCVNCngxnxmFcR9ihNyu4iVcQD4ey5SyGIJNX70vyU1P0Q4sLfXdmReo+Dyat4dh
u0ZeGomi1unnQZiPDOxL7QlQ08PZlo5j4aUd+4AkWN17bF0+sATKhtPGHvFgiSNNpLPz9sJ/GTNj
dZC2kHaT3T4Co7hRj7jegHXkCXmUZa+RGK9BYUTJ8X1jwh1C3Cv1L6KIaELCJchwQXC4lPqQm17s
Qbkk8i12O6yTlLtfyK/vSIegc4yP9/OnBWPaIvUKOD0xNrwrnFPD1TNqxfqbffADOkVjQCkeKHAv
IpYIy2nxQFIOYg/IYChj2zqx4akmU/AWJ8y+ghcnHD1FLhWoBeGssgzkpjFeWs+Y3RKrRNCnlzLr
iQEXCozexpvfz2Y5WKGhOI4/sFA0NomIw1glxsBczgmDjhnIiBHHhoEudaHs0lY78qUHUJkaq8EV
zjUp226c2EKP19CUTnKxCVSPkKcW6bfi1wLKSsfRxHGdeH0a8cH88pHGiTQVRnsJovzMKSq92Rbm
+9ShYWgkuoLxjNCVhf+d+XOm4T2e+v6JyGKySzYYqE6sVsWnQNd9QYusWH/B9B55OJ5R965OXKAa
uwsC0+zsjMPYfMDjKW15a6WvRaaYfYOsbOrGsjlnvTQV7VT9SnAe2HOuuqAOlICFDBHnlIsZHRND
WUH4z7guEqLotiivTZxfSCpojVikVnCFwTd56v4bpCUvG+sW8EaJiiI8Hqh3D4orrBEoN9wZ311J
inxmaedIoLbiGnF6VFLjDwxWxXJjzHAkm8oTYV8leng57Oyryr3KPsMtDKPuu62Gp7LVjy97Aq6K
1W0sAyg84pcD3ujs+3pdgaMMiiNaQYZFfj9Juvp53eI1cDBoHaIm2Bj9AJNp8d+vfmvwXqv196EN
kB8Cb9CJsxOxfj7Pg9JMPvAwim0vXQxJFlJFe9QlDeK6Z5cb9skFwxAkUHQ9PVBR0rwOQf3Lcdk1
xwzD5/6M4X8rutbC2vMX+dWSd2PAmV6i3UqWtehjedL22P9rvb8lnDk8Cv932sydUtUSEu0gQJgs
qLL9w4r6oNAmgs8d+Ayk4QETeY5FLRh3kqGNkMmRJWk7mqwIufMJw//Jk/aW14oLWxD/LtLENrOm
KH/R3chfNiHUbNMKDCAyWZ2eG1gW4WS+okx1DG+FO3jIlYyPhSrFdUTRPu2w6fCOA6lr6bvUb2FB
Ji9hKJBtGa4suoGOLAVR8dBm8t4XWRwSVWLxATjXr7Zz5WaGPfYzpzbIRuHWRB7o8hHPjZZnJD1I
otmpDU4dXz8gUGVQ4cAH8lbW2HcUJOLVKanew+Y22BdG+WmO/SW0v9C6rOU7VnClUagMd0yNi9Ja
WKRSALDgfpdF8Cdmkkp0qVvHunpP0AE5Zh8M0I7pOztCA30pTCD/slx4g1blQlso9EExeJzcllYS
QHFFJhBca0B6NCU2ZzI7XppNET0sDjCvzyl4oCXHVZAeBPJGTb8OSiEh0Kjv57dRgJxGKK30B1T9
hAQtYPAKVomfhZ9ky4s5BfyTFUa61kZGwJqrGDO6Ai2mkvDhyFRcTHDPz9ZmXKDzw2MChGTnTPBa
9gkUFlqmsjWkYNuKLZ479KD8NkBj2Ug8M7FUde9RX3/gAdphBPde8kI4DuJYNX63iykfgx/hnA6N
u88TQ2yiAelTpYq7zRtsmhG4S1N8DThoueR8lMQ3AtcVW+JgHar/hPGbLtQ4A22WzYMqj9YE2l3f
wdixtGeBPumaokELKpV7lJCrStDLhnVBddgEpnrF9HlCsLuLolC+mRZDImhRChf172nnFDYF824i
BZZEtXqkJmrBXey6wGxTAV4M5ZVw9945Oax4aC61tnCF/Cj6kyLtmljoPw11pOvlHKUlq/T01GlP
53KW3gyyrRtEIZ04EnhKnuKf1d46QNlPSuEU0wE68WedW9hQQAKMbg6siLq4jh5OgUQAq/O0XuBY
Q83qh4Z+CiBgl84saQJ0+foCtj+s19ZJLbyTixuTNr+pjouKA5+ib121ezacpGv1T522u4Z4oG4A
IKgGb2RB1g6hrkVc7kOX0g8w0AiDnipExldk1N1eNNQhFjeWjtVx0BP2VJq2PPNSsRENeKR7Y/kM
Kh6/cvrJzYnCdKRVSgr/iBtMK4EG1LIk0xujcqRcK0MAek1HEo+us/HYplDnpU1ZmjOfOSnkuhbw
J47D6d6ffm+zjxUzxkZbrlgns9GtutDW5mzouQ8OfoAS/8fR64Ym1jldMoUs05lrBPaoYR+HGOJc
qH5QDQnLSVOLz7fpjh0nTK7y6d/ljYBbJGFhUyudiKG7TisKbeDvmLZAjB1eAgsqZGHL3siC9/Q/
bFWQl0jHAlWT6Cyi1VhfUdGRYx1B/dPyDmka37fP6HNqkeLwYz+NC7TGWZobYEgCHB4I2ZrwQOKQ
AoT3Zb55bgei7GEwumu4q9jjssrisP1MKzzvkIbqStOH9gYtIVoWdHfOgrIkhhqtTzU6h9AAD9QL
TG3cB+dl2++R5C925nsBpXfD17x4EsONB9aABLFIoZhlf3/tYOZzvIPhgGEeY+pUeQlpbTr8HYLu
NNxOLrqvoQ4C28rDW/HVlrynMblPEohOVhzdH8QvhAB1mno7TWP/6HvIiVAexgktFWaUXnL47L1G
Wikx5kNnyBgW5MO2jPiEZyiOUIRa6j8o6zPzsDzll9mzyssKVQ/Q+IbZzboECWSnyvA2s7VcyTfz
K3+kmVq3Ck9ph/NoNtcgYNIeGW2S+a5Z2+J9KMT/40Yc0IXOaEwM0rojkT9x9OxQj+dkk202m85J
m8y8D5Pz7HIG57T67LY2/0qsWYT6THBj67+wVYa159RjqvwnB21hWhjiz80DASBAxlUdWu5HQkW1
G4KDJST2AljIZt6TZD7AKLPWRPFpEtFoKH655+xdqYo9DE8ZBgIiNfhB9ztBCiH6MZKWJY+uvlV+
vo+mEYDL5yhJJYR0aF635rCsgjkY38cXQ8vPiIk5kkIVUOZOV9Ef477oIjtZ3f2DjD68lA9vuU6Z
mEjC0FSIsWSseg+LsjpzsNRXo8XmHQ8ixLeimLymnBQhC59850xBpshyWwSX1nZ73dDjEUdawZCU
5gx/+IRR0icuC+oNIMKL5vjs3FiRQt4YiTa4+srAYQSELHGXJIhBOr25e1j1jveeAne4GJjfOuee
14BCO22FZOiUah9ToWN9ICmhU4BZ9TKuUv8eAaIWMxFlGVtBRMjzMoOJs3Iv1VjHxnQ6MaSKlsuk
8GYy6vXbe4NvIZup5CcMzquHc0ukFMQba/IeCllLxMnAH8i2axv7lEKi6VO+PxiPvaOan9ZWCJ/m
qspcTgSk815YFUiQQQGKEYHeIRu4A8ab+hN1yx9EiPH+dw+LSnxm37OrvMTYdPMRy8qxjus2pTa3
kThPpRQ4yzSy9gnA6oUAgVL99/CXRG3t6T87M655EgezjXDXvdfqeRPjJgi0p/mw4W4jIejJXFf7
g+gwl0GuEnwhHmm449U7pSTokBDubxJ5Q+ooUq/aw/lxBK66qoBqWehJHqJX+XLGrLAsGKmuf2jN
nqZk2k5VVW29ZuxJXYKjSDY3e7pO2RNlUqumi9c0nNlTQY+9kCamS8+/XTgY1wJ69Km3yQAl+YcA
kkHuA5L598bP8foGgvMmLXWN49rixhXAaGyIp60s8H4bwaAosj0tXXlOGIfc5vswV/C8HJSRynPD
i7qH4B5EAoahZJpJsiaDTBxdXs5FUCuqDMXghn6pfJkbOiYukftS+MZ9U+JYRgkLr+3/mRijYwch
+SoQvXAyfqF2+Sep+rmaZIFEiGSWWLA18RL2low/HyzW+0Lb2+M6YzvmmnMgHzJHc/npKQb0IOyI
sQ96xU71Pw4Cv9nL5sgtDbpuWvlNez0ypBAbbo2mdDZxJzQp804o5Syu1JQjmLuFzZhUFOtwhBQF
UAN3N03OVIPlSPaN/YaHZkIWFzTDXVp867WooL+k+3aGzgp9iOHJaOpJanLogkYJBrfhN96WwVNE
sAMv1p3y9GiXBrtMSIpGular7p21LT/7309vg/sqZM5iS0hxWh8icgFsm8k6cERYLyHPyzEqRW0o
Z3n7YchBEyligKaXNR5WAn/h15INk3aI+E38YcArD9feXkIA2Z0EZLBc5rQ9VGGUsuFHY9ZAtuFl
T5x8JzSCgF6FqUUjrxBPnFPiTOgihBnVFrUSRnKLWT7L47SqSRTQ23vf6iZrjH0uy2Q+WMNw5mqe
SdGv1QgpwTyua9tQn5y07SPvWzWX8sxxRmRLoYWqDd4yHLNLfQZnsjIDDgMNfrvg7al3zn2mH1xx
b5EgI8ob9oJZO0HvlkOUuiOw2FN6ODvE1sQWGw0RYIxqPic5/LEIVKMdsAN+fJhlnetdNTeFppDN
QCgLwXdJim7RLwMU/yTDOsz62Zfbo6ljIOvgpcqadFw1ycC7GE6pIPhbslaUWiuCNyA3yKC/qL9e
6G03CoyaG/4Kih9eOpz5ExKZgMnD5HflCXoi39Ml3P6ingxyrWgMlbmXuf8uvH2RQKhKJRu7+I2G
I9zDNlh8FXx5sRqQivA4XtUiNeHW3AmQJNPGX9yZsgCu4PsuWBzJ/aZtPoql0j0AYiGOY+kY7ldc
IeckgXM5wgxoIfIvygyO9Q1GjrcrpZHez/2DI5mjAgmFwA0i0JsM8aBSVvVzme5n0FewfkA6wA42
/z1L+Vf8Xr8oiuaQLgKA2mOSg0pZWU+i531cxOo8fInqssQE1mWceoywpQL9zH2OET3mWUgFtZ7N
XzUT1SO6k5C4EhvDlSiUFMuJwqkwlId4pf3ITdNq2dHaIMFuvSArkd8nz0OTOF5XIbjNiPJact0T
jmgvUxIBKOQ8v+UtVs/Yj9CZnFSqj2P0T/g62SESmp4nFGPJHMXaRbJVlWxjypsaDXdmhAp/t5bH
FbydsiZywAnGkNxkt6+ko35XH2juX9YDXvqwqjro6yRTkGJHc3q1319QN3/uE2cgyohbEtN/u+wn
uR1UVFRdoUEU0z78IJEGJej1WTOk+luRD04QPJ91Xs4EgvB/PEkfIUknD2ARcj7ge+Rqddgmv6bb
RWLVDO9qkC81xsB0M9uF9Ceb66FD5XOvKXI6xjx9b9pnVf5oleqSeoelfY/519f4Ny5JDkcyD7J0
bLNwLhVFgRN5C/tYfHhC1ANzA/QMCxHcGpsqgN0rvtWLJdOR+1lA8OATEDG4Nsxx4hpXc/i8cBBa
6exHOvf4391upLjVjceZhTa3YV456efRY9f2guioBNz+mwF/hc/RhrPhZ4JmAp8ME21NtbWyKS64
pIykiksNG64j8WY+OG7ca0imxPdzf6dh6UkU2cUZtbK4yoDDdVnSYyVDSOuo43o0JFVWxYMJ+twL
u3FmvxWaR7ssoEnKQxBxBpncMSHzkNoRzI/aSv8ig/QBRfPiqJkfFtTYoJDqTi/xsuoezXFnQ0dz
PmvbafNXHopo7gMnAWRue4KQ/rAe+JiX8cz50ZZx3yGBwl8yWD0x60d7fuFkeWoiPd9WJ2hgdcMC
pziplwe2w3E/5gW9PxERth0vMNsaHidaWprDKZndrWpdvpIVE5aDG5IQKxnMzpwU0JVU4KQvp/WJ
zZfBVKPa33RSujbirY9LpcLTk0e5NC7JvfjAxmjElwZu7di3Fw/VYP+6dpG9d44di1p/2eKH+PGf
RsvIEdAjrXGL2FZmyBQlbL2KWaHVRjWz+dcH6cJ8r4ZbW1WP1TL2XNR2xZZgNjUp4wduf5NRMFkj
ZKChGB+JpzBfDKhD2iQyZfSrgjozj61kxJgIiCtwV6kWWUqn9PPaBLk55A8dSfdBU8Scs2+3ovUe
QgWhA/MljxMEk3QZsWV6AluEEPBQZEPE+c29YFR42wbltxTake2wzK9mbMfIMrIkMekR9L0aVP/n
ydG8WeqKUnHkeSAJyCxdTxR5BDmhOjl6FFodAKXGiGKjimr6brZXSzyyq6QzONzSEesXFu+6qRsn
ZG3cSDqu+PMDAn8dt3ugJ0BX96igQS/LXIvOzERkZUNIc9a32Sq5VbNuEFiZOIT2wL3qtJQ5Rn9g
IEUV/9xZ2cqBmbwaDUbAj/JaTk5Jyy+mz3bxyQX25iMCFhCyChiXEOnwSk52y9oNx2z1ZCLhxVy9
wTtjCfxwx/W7iE6FYbwzKHdxxPDleeyDi5sie/DIsWHzyfqVSh96+/Se9NZcFxosvKw9eG0QeNP/
+UPeslbmXwbBevNU3k6kImhVU1ECNldYXrz7idKqClsZZiWdZvMcJm00wWH/r+RpxMF6LzfCBELt
2KPhvMKK9T+8DByWK+ga2ePWAM7dTqHiR0gHEmCq4qSeUfVK/FbKvbcNd5+XZbND+A9IDPvhjgDC
pvaXSi80UV+pik5xovRBOD7Mmb+6x72h7Bi/16s74PHu2rSa2LI55JCGOEqgC7oZZXjHKZW6kriM
OCBkpLcL5DyAV4J/PV304UDSro/lbMqG8G62iypWF1w5ENZdkvOQ66egWQQj1Rs1ABOjb1670lby
8w9HmNcx5mqvzuvSxRFb0ORkIHAzisplPkMovo0KAIHeH1JvwqLqJBLJTet5AQf6qARlWljXw0CD
7b7aFFoEmPxszVdpEMnc/6+wBnYKXogZzd9xP4IV/m37x31j0X0ZQqzPaqp7CMK/Pu9Wl7QX1VEW
NzX4cuO/1JKq5nzU+39TYPsIDIZfBmxX/A/otua0gzaalouYzG29XMj0XBya+HdkA8er1FjW2JuW
Q/4WsrzYo9bl/try9OKBD8Y+uBiAdJOiY8SS/RVVgBy1tUsgLKWoKlYipEkw1/TWX+SZTyXXozL7
hXR7BjdwOpChxaIFLVkokBzPInER/cMcxXd3XYp6s8VjZ3HU1vyZhBPbyLUCuQ7CxKgXOT78v6cR
aevLCAHk9LsqZwpAsI1BVibuElivs73FiuTzAIDHxaLgBt+qzAocdeAxOl24xLwh8a9aOAcBSA8/
jYRDi72CgCXiO2yGSepNccD2TwEGxuK56euIEz/TDpozS0cYCDWNMlOTZYAllvjkkHBJAlNb8xar
k8i+lF9XswI18v5LvzCZOyDViAibarFQMkf37+HonQPi7AmALiPSnPcRQBOSV6SaTdijJNGbdM84
oksZQ159L9WLCH4j8Ka5Ie9/U3H3ufaPX4rlp9Z0118kF+lohScmeriCoznH+e87RP2lJW9zZfnV
Ylqg5AXARm486qhijYMdSi5Qoc2JuFLHkYri/dYzXP5Rfb5lKbninJq5C9uXOez6PpJdEIqxgqJQ
iXOsVJhmNzItMVcRLcaelf/c9FTEooZQkooJKDX9hLUmg97JsJT7S8H4U1ajR5Rp1Pz53mrg06GV
VHE7L9BbbHdoIf+7FyN7LDM7RRWopdiNNaLEFAMrzavr6+McRqkiEVm046vAJnOgpMBxIQpPFJNA
OYvwvzeItWZaqzh3/rapm8bcIPeu7THeOlNIZbYq5yF+lR/3hE66F3GkMzwzMhYtL7JZmQkMBc79
tMk7R9/qmEqJG4XrNVcJJi2c+l/a8Bpxt0ShJSMBfmfqCNLhHs5Iq10oGmjnsLMWzgdu1uf4oTQ8
f0Fu3wr+X4MqPBrbqIXTOg4U1Pq21uIB3X1fqoAqtaDDHAxaODQ22SPg/M2eioLQACdM3d81IUGJ
9TYloi/R3GECEnIgZhnSFfpo2xddRER8TBsu29mPHkAvGRj5PYCqMeWjvHfNVuHIwl+LVGm2sVPx
l9sfsLmMJE26RMZkpEAgy70P7Z4fomsQJsbGVTxEpSqlmrJGzWBjA7VJy4BRzEr8NRq4w89untMy
+Jb2qe58Q317v3k/TqDnQ9QvkxXJjrNxSz09amtGtVS/Lt3dFNT136mPo5p2vhpMtywL1paNrxE9
4ou0NARQriPscJsCSmLXrkO5k8jvmSJOk8ahvZ6p34PKwZSAiN2HqflHEnMmOr71+AQxvxAapNST
Tp4JnBm9Ik0IfNrWwA0TJ7/A97FxgPtac4B6dLMsQT/t+XwykZitoVnY6EatvAsP12sCT0FU5uuh
kYfh42MQANqCRY56jjy9bUCY3ROvNW7/ime4J/LftZAJtiWDYeCRjXOL2NKQC+l8njERX0N1RtDk
n9Xmj+MXOlMub4y7IU+Qdc1ea5EmXYogqOfP4wHLjqjKe8B6ncI/AmXBCvbkYwk0mDj0NiW2dW2N
u9dnLuaialmV1LSd9dnCUYeibH454VwLJZ/l08NeN5VsE8NWpZR6YnhYkWtn0VcUTMsdjOkfAGzr
ogj3a7WfRvG1/VwagCc3tZToTRzKKkFQ/Wiffu9bbe8BfOh76dFPtLydeaX9+APC/JElipAenADl
Wfv+9iV3roX/WKp29DQDN0ytI/RZoPgMpqFv8NLCz7AcQqc/eDyuSsDs8nD4npDaF+n0mh3+DcD7
N7Ckd/6CvqmkbYxx6Go40b/fyBZUuAbii1X9eD49BAWxrHQFoTM2ktzS2vv7vIhQTFeOh52xuike
UhIWPKaG2PsTSNqm/K8mP+7PLO735ciRwmSdZ2Oc+ja5Yz6XWK/rtQRdb8xqOb6/cBRVob47mF0K
kYoJYZOY9x6ogFQHI1euwXVTOUll840IriBbe+K9eGJd9NA3ntAT8KuSmqdA78jmUbGSr1WXOjZG
/5FT41z6lXUI/nsE8sJ65an3qm9s8wbnS+lqGd+4nA+CezJ/OADVjSanfo2aKOT0AbBhtPlzQ3f8
x/i5Ek+YsnjXRj4ahjSxg3s8RYuCbYxQCBP/tsRQfqgksZl+WcPDvEizCJ9ta8XrmKGcYYUewTs1
ZyzRGf6TYpG6GLBOoGu2et14VtNI5USLlzhN7aUeYFACpOBH2EUzEk4NKlXBikuUTwqiPdWYINTA
gkajmE9/rPeIwMTFIRgsrbo6n9GeJCh/Z1lroyuaNLX3qfINvnlOAWUhKxQzlzFHmpBxh2BntWzz
+foxxrb1+Ni+GRZch4oahfojfZ0McpDsqbXP2A6AIA+/CqX4jmS7Fso8hjaB5hM2cyQ5xCmaXeMq
NqU7qu5c9/zMhPH+b/pMCcubs4g1DGDBvTFWScbxY9ErOnBbpTFP+zGgS35u+WMAHbzHvYPMY2+A
xA2SIvcq8U2GQUtxSHYclaSkCzl8fzvfOoIS7mLU9njcCpZYIjBpWFpXRew78RxqGZ7fffDFIGxi
fOIRGu0lTofseO1L8oLsZ7PPQBQ9KtwYsxZ1bSrLhnY5A8drJoKEfjeGZLHvaCvMZo6P5oA/mnc0
9ykwhSmvpm37oKsYRw04yGPaEbWd4XCxg88nebXaNSS6QG+5PbbZSXqxDjUTRIJckIuUH+aOZGV8
3xLF1EltMungctjKrK7KDPzkstrwFdvwZF+Hlm3EdgByhJl2RwSduqOX0MDghntyuHMneWFa8aLb
rTx4G6YRMYazf81jzq71ac6Dpd551/FRvBJVdKH3d5k4LLiVv0yhef0oKm5NUqJ6CVZzERSBel4u
oWiJUea02cOEUGay8ThAZb1dU3qk9byNJ2f2KiYv3PQMpqnpJU8lPVi8jGdXk7Tt+SW0Sd5qwizY
hnhscVHg5el0kg7oorXHtFgarGfkLz278SrHeDH5oeTRklC260NCE+XIko8auP1i9d9vCtasmYQx
U2gTeA6g7jHaM89y2af78s7kwtnRWMkD/32ACUKiPVOcqs1ZE5Yct8zvW24V42p/614qZ2cvk98v
eA0vSuF821rXsC/hU1c6t256HxVwpJVGPyR7Zq7gYJz9K05Q9P3aMPEdjCxyYZYmJECAApfIyfOn
spfAE3DagT2eOmQyDspH2MmQkru5clkR03Ou7/cvK8td4IQG2VJThYVl/MehChCboeDBMyHoLi1j
FbIMcakD1qjEsqoz85GS89qX5fipSC+LeVFJB5FYVvZM5UiUEDYaDJHDWDOh+7m/7N+JD3Udnixb
KEa8OnGkBndrCeXZlhnwsZGnfYoFnRsyC/i2tFhahFR4/ocy+y4upTK53LU3mpPIXbVdkF+Nsa9o
lkiUfXEg3z+ioMZvCE7iEINQo9f7CpZ3XEWhS4TsfiIqeLaCU1YgD5m2R727dE0rcTjG3kQONJN7
Iz/ZTAtcqLBrWeLmNXJPaLUeIzMT78vD6xZf5mYJMUnyDSaLjn7UnSlpHnXrauo62wk00t9rNXmm
7gTja2l4L/RJAAuHZrzgYBgSwTA/REHl9MDUQpTtGyJrrtKU5dOR1cvre6mLrEMRlTOMmMdncQJT
A2FZDE17d6ZynlmJy5O0d4xp9LZ597CiLRb8scxKfGaSYFeL3g5UmGMETffo1F8IXl6fIFupUTLc
NRHlOWJJJlwL3OqaszLV0SZfNxx3m3PB06+jAekZVoRXlPxE0FVfNHira1NyI/ZmU2NKFyJz0wES
8ZTBfKg94SPlP1zxdv6o2zRR3DtDlcVlXedOJI2kI9FX3ammTILMmgqM1pjtAylG8n1/Bxmeb0oF
AkRQvR9MjAuTwOMArx9iOSpU5um6jarutBOm80JmLX3lyPtbBGsbBesADmC+NWxrR4McT96nuk/7
ypQS3M8QOKo+/TiGHiLnmLhh94nPOBjujetzctcW8E2GrARedYqY3eZFtiG+mOHS5bzamlxsVeCr
VJnTvYBtLuj2W1o5RK61okIe5vHmgMjCMU/w2hp7xd0sZzyLsEKkoPeM5V5ycdoZNhIVdrrHpLXR
0skBpyUiSxBJ/oJdUi92dWlLukW3BaFwNUH0azjwOJdUrJ4TL9AD1jhdG8G7wVy1q5fBdSqmVSyq
6PoaN/jhwgflOL6FX6WnWovc39xJaVlEoCpNkXNoFhd5At6xKY5+LdCiMAkO9QvFrqQ/3OUiVMKh
SQUD+66VDWuO1fCwJIxdY1aZsKGfZfD9FITnqelE2OhV74c9W1eSjVmA4ym/KpWSFypeMC0Qt7nC
wYO4KD/NjL/YamJEUsy0R3/XlTvLJTjoE5G9s0D0tqnZTOmMKWG1xtVIn0nAGGSi75NkjofWJhbL
0JrVTfb+RKFiu4cn6E5vZRWUg8YhIYlk++/83qCMELCX+W0bOkJYTngcg/N14TKEUcFBaGXgqWVD
kFbOrnTBv0zQYUWoVhJvzcQ9vJUkVuagqja+fXy38hbDXw9I7/vC6nIisPrFAnqBj1zrbyuudbW4
ii6eg0Gp/a8U6fo5BSpEVcPG2b/anmU6E/wrjjQ/qfWpJcShvts10V25QpDwZmHeC5azZT63w6dv
BhymZVzH/wODY1Ahi+hIhYQGgbHLxfZkg8RScaUnjoDwXSTqohH7x0GnQ+dzlsi+sRiQ4uVnkM3f
zWWJWFV0Ao2vZCWpizOta98OgUs94MKb+fQRaftOOzgbgyO3zmbg5Z+ZNk6pOC2Edlw4p3qxLT9j
cE5O9WN26nSyphA5YDsSI67zIFvqm+skEB1y0ldn3pMhKf+mu8B2lrrEcVcHFeTw0wYeTiDtowg/
wWQWH8ayTLJTsOlk13FJxRfWVN8dsdHsWF4JfilBZJd5fwAT8E2ZRLuiiT0pkUW3e6gvWxxY2/nR
avxux4FJpcFOggR8nVS9J8rGKOv6iuaa/UvEI2OjjBLA58sHlzPw+QZrBaIR/8H3wBwZKOi3Low4
gjol17HNxN82VoHLvv2Cw3rcd3sizITwc8olUgGS8+TUho4+R3R0c6XDe+II5ojz2gmDDvpbOMQC
lWIQlVN8SmeEAM6AeWeYEdWrpxE+VlX6pqeGv/P5ETNhwzRi2pi5heSDEtPX7ZFATu8THwQAA5hl
l8AJsJ0iFE2re+IpjzxVFwzFVjXn/WB7UkhOjBfA/BTtmfcbQFPPtIkASixwbSLQXQDUX9LYrnFw
/QHk3SzXrhc+MlzzwGJx7IlUa9wtODPz3LiqgOYesy/TYW5s28Y71A01WlBim9hyJvVd7Td43LgA
6FhfM9HVh8r4cr7QyACAWVJw4CYo8JYb4c6SFyuFwe7nlegiuhjxgx940IBMJQ++M14L1nxJoaL9
3dPygyx4MIidi6Ld0nnKRCX6HVlgSpA7omafr0e8di0yr737VnnSR7QgevmKatGeJel2WWbX6v35
pxOlGqgHIAW5nprkjcoLEeQEWZYNINQHg1YZcvdYa93bn6bylR2M29T5rTpHi1IpR4N/65E1A2pX
cSAUcmFPmhpsmvE/gGOT6zyqUNfMR9QWE7GLfaKgC8qC2r4m/bwhEjW1yhlTswWekZflQ5z2j1AE
YCUiqDIIOTPK/6AoPcWNkEV8hfK1zCGIMXuxoxpc4RV+m2wP6VvlctNs6r1hwm75smXh9aukz6/h
DPVlytWHHAKe5p7v9mrn0vZnGVw3BtXEzTEfnUqezlp1bjMkbyhrzur5zy+MozGthDxo3388vs7m
VJoufvvG69TBTHBwTqf2vzrjkccW8pFhqMQUowYp7SO8nSLICuThW3bkVt5Mk8Q3+abKoYhCM/Km
Sao7L4pdGE8bkr9zBuZ3nc0ur8le6JDqexIVekkW6YMQEEh6/BsuUMSjEFyt277CwW8pmQoJekRT
bNvnKA0kjcGyn4vFaNCv+s+7AGg6VMwbqj7/E5+cVwAfpyjvqiNrxE9zoNhptBVeMdKiI5i/tbbi
BmUlD5STIe9NpgsvLLu6WZHMk9c35eVim+/mcfR3ezJiNz0rboqPXIQcFQIU+6JyvX0KZtzmMdAQ
alT8IegGTn0e6g+gtWJll+z8E02GInkgmpac8IBBNPncNTT4OwfpmvtzAf23fy4HPA9OyqIgIhrI
zzB8S9RGjMHbHAFJaszUWXdLODGN32x11U64US+5BbSW6CdMnB/G8xXX2jMkdJg9AAcdi/BuJZk+
UaW14EVa49Km8DspHSVhl3ZoGU6TaqvLAptlj7ehP+Uk9xpznPccvIKDnZ53z3XnGPKg4anv23oU
xrabS4JPLPk5xaTvMrWvy/E3dkWTMwFQ/1IvOOIB9xXZxeK+xVU6KeYEcshYqVpj0lgMf9VE1Eag
tJ6LmkV56GoE4K9JTX5TditLqaRSCtv+OcCuYXYs6JyWdQboGJ00w2xqUgegT7YF08gcl12XccNS
9t14SttAp524WMuuMC3LHmWS8PTh4Q18cuSlrSWNK3XwzFvto155xaIMyj8WZppzUFzXtti5duE4
waVoamJPuPVFxbC137EYGJy6RdtXhPRa1pUx03048RtsJZCQVqscduu/7F707VidHlrS79l+jGa6
l4KT1KFgQnrBQlThEVtol1U96bJPBdVLJu0VLFQ69I64Fk+7bIMpAbG1NgNmbo6JWuVajudcmW80
T2VDq2aOQyWM2gAtEJEE/gWnpKos4k10oPNKRwEKmA7tBzP0dmsO7Fv/h8CivD94xT/WZc7khdW5
IkzlfIhzsJEm8c7G/2hAI9W0B+x3VEfD4wQSb1j6tYedEr6HS9FVEbWL4bveGxoCWph/5N6k5Wi1
a3h0iMYGV+UpXI2kb0Wjj3msFoTxDFtMvEm4XFSNj3OZIjY+qbOxFPSaGLuJIyQFGMCiNV0dRIod
RdkvPObC0nXcC9ylCnberGLMr+wsTcmcDcGcsbReGeDV4EUcx18RRJ73rdaB2nvQpqeD8Muu90nL
kmFpIZu1WNSGSPQv63vvJ95i36de6d2WVh5zXJQ9uqo/J71lHvvzOodY0eEuiNSKFQlW2vrr8blI
Q61tf4+xIfigZovJkrFMx9w4L6+OBJcYgTgfE6fS2q/O70K1m/ePt2F42/Ro4zfuvoyJNng7F5x0
5Bh7gNiL21yh6oFLSzvYoOTZU1TpDSmG5YeTu/lM+iRczfXQfMUKBtjbkWTG3RY2Y48+UB8MpvmX
oNDmz4LT6PqUSGO2154AayosyX6gxKfkyPep53D0LEBSAlxdv2kNi+5a7ryWv1SIK/yXK/jrAV3P
m0zYy1sQxHUhcL7HVuDH2KC8FwgzMqy3g7RbTZhMsF2M5TkKdNjIAgJtsZNKiADeYhYI+2PgzrA+
akJQthcX/pGlApxKHffZ1GDLPGk0DTEG0naJc9mu00KG6he7KbiTfI6OtyK/lKjozzwIIa9XXACJ
lPK4DGNb+8dmhN92TsVk40g4Wcedbt15g8cx5js9E+iuYwPPsHF2UdmBzNs0H2fkCy/3Ju2qygyr
ikgsxzE5mEjCx55RpRvcaqrU968Xga8u12w8b40RAF25WqK2gC8dpApzypdeOkNz3p80Bdw4YsWc
VucQTNoJlYZUF+Wnq3QQvGA40ZOAmn1Wv3PX8FU9EOYHPFHaB5EB3qx00sABgbp+8F/UsJOXITUZ
HmadX+CYCc9jcXqCgJ5Dnv6oYKw/PSzM/gcPr1tkhg3uC0lJAlJDEjqhVZnrpR3SGFtE6vnwXenA
SnKLkUM2R4k6OctQNFNn7XGNGWCSXIfO6obmB43yIvvR3kNmWhqr7/JXkc3EckyE/l2QRQMATvUD
MIzjL2qUc9nLjhyTXCjX4w/6wKRt5hQwgBDjAO3C/hvFltAaJeR7oJUEtK8QiMuAX/U5kKiFxz40
gK9GtMwn6rq+f8zGM4aJSezXx3EG2xoTDgbwJOkX+lT2Beub8lMJcW26VPSG3r+hsR3+WqW/kw7x
0609lsZOAtk3uIHJHpI2ZxWTwvdb7jBNyP4a2sSNNKAfNlHyhuvvp42eD8LTAxcO0PjVoe0FYJaY
674+Gnk3zil0M4yAEYWc06Ln+HFswdR4V/c3bSgtiAL7I79UxRmXyzadAhwMV6NkoM0mH3TF9LxD
Q72yDnwJkqy26No5cl6OIjGh65EGy7CioIbzgYD5nQgiHOWwLhq99vpAQUPQBVPoVu0MvqEiowu9
02RKlFeXUKxJCSJ3ywYB8pMVl4XM8zwRQyka8BFHTpduKsIx7ujOpPHV4o2/vPzD3af9Zn6ptc9F
lzpLME0JdHKrZg+eZ1X50x3fJ0IKHbMH4vUuEhQboIPe7cvERfXdlIMYcG28Hkf1V7vmrQORNjcB
URKEHZWDHa3FW8kRhurG/k41OVWqErF3Ul8EirZ535kp+Haod1ID7nbZUlWfyabUSN1op51slBtp
SeODygZCapMt2HEX0BA2lF+MmPDIDkw5N9mJhc8JdH88SVadsu+9qhsZ4J+uDm7UPQeh6zJhodwj
MxBxuu/LyaM2SAfEiQcP8l+rDQxgbIVZk/06wJct9N51GS7EmSDiYS/9+3BojJTwsRV/nF2I6ndz
19nTKigQscflzbjyeTZFAz8IBf/wDP9Zsnsnhn8cZUrRlb8IRfBtr9C2+FepapPAvLi3NAyvkNM7
NtrhAscjROeAVnht5v7288Cs8rFiDTTK0YYiF9dCQ7LUlWtJveL400OPuNOK8lgml5K6pwSPKvWv
71G7JyjcyS7/YeFw0rTvY9f9ngSzEqzy9vdoSQ1jrnxlIdQ2DswYKfTR1xYrGxeiTFWBRvvyLJ9x
NiM/wX6GGahPNcpTnV7ohYnS90jS2Mkavl4GhEJN3q8xQ5ogcpA7qIRUXqRUkJCYPxj5yuLvLxkz
u3s/xRvcKrW+HH6GRQBJQz0OxMEUOWqHQvVg3QFzkP447WfNTnpXtwouTPf37KrhyLsnPovAA480
31W0jXR8JGwV02E+WElhQ58ax4owZJ1NGU4sOphVH1RPGroxJQ8rQ5RYZZF0A0X1Z8zWf1hsD9LP
EUvBGo/dDlL62IaO47E3N0FNoRvXyrOJUHYDp4LgaizVV8e4FUOSe5VwAlZKpqTArKeZvbRiFuJB
4kwZ36eHyESrvySPvz0xN7cCXnYjU/pHe/n6Mh9mUtiudkmcKF60Ulcc+0cgt6Cnu4IW/Mq3NzrW
eBwB4ze/ARZry5EFQ45hlgpkkvSd8clJEdM5xYY9kwkx9R8DaafbCAnZAyhXSTNOCSvdEa6g8Vgs
CdCs33sVYIwtHaSJLHNynvSvBNHuQHfKpRE+DaMpRlNM+Qguh3ZYnwGSd2hjE9/Bl4i6cZ1a7X/a
83RhqmpOhLP5yli/oAOlQUZVoX3EvMfZr7huDkanj81snW43EHgNGEodwr8YTArbct+79StCXzgt
IMnta53WHGvIb9xcC3aNNtJ2rdsQni+Mw11is7s/gvSXBtLxwfM0rDI+Lj1hBLR2kauV5F2tk8hb
IX3uQ94idQvaakCDH4xTW4GaRW1KETWAf+CBvcTIOrzZS3qWRZpMlfnQH7pbYaB2eD14/JJsEo5Y
gfNuCSJdVwzhUZWqoo9mZ53VNgA5C5/1tEBxYyoGYhAePwUvyO2KcUpJ7x/LTJcKeVCDkm/pr3/q
2fGCLw4nJA7bDCRSCAsugInSkV6eqYgCJB/pKKhb6BnDH0LDCl4uXTPByXcrCGree2H1ESXTUqfC
xxHJ2EOhvYYvGehde6BHlYq245h86KgUJc20/YLtPtXYqpSAFf8lA81jJzMRwc+im4QBZMDQa/CL
6kDCdmz9L2NeOTguMcIVhUkAsrreP52eo5jyrFUFFeKeVJe8WnvCYyGWOZ0OqKauY72mdxZbjEeQ
ZMG+ZxFVGuclB+Kjkboy2ekScNGj4RaDnS1hHiuWjPgy+OJDbKsGWlri4bWFJpeGbHRAszT0zz16
uqAKdONYQdt/F9uxJkv2DiRDL21ZDvG9CRyU2RJDSjG4MO2TEq5FGFTqbl83xvwcHqu52iUMlwpg
/lVyUfPCFCjrlOVNlK33GY817NX7iKNW5PKmNjNdqmEmkjrejm4TO9hUDvfo+3XvEUq0iy02J0kD
jVVud03Rl2GQimg83zKbptA3cxLs0REiDqGLKmgOeHomrMMq/HKGIGW1gUIM/PVzCqfsVGAB8x9K
HP3rdZOoa2kiKMdYn73cJS6w7+XE1dJF5CGNxLGqcxTZAVB9Y+j278JLB7h0b7wEtl3mMJflO9/v
ngw34sBnVKiSe9nJ47oHdUWzJ3vQ7Sc7ZrZwu9Zl8gitCTIw3yzAHfgxZLICRbFxu7yoSQqF69iw
ujr4QKa9x/IfBvO5Xn63/QSsfgXYKm6IihutpBZLWPi9x8rZg9ZfdbkUx/RMm9LT3PvZ5oSZrIF+
0nk8OgbAAeovBiIvZTHoJZEOg2dcgWKTGvZjaaY3M3c0sUg0Tx+LG/m2jbvrErsK22U22h6f5Zni
poKfjdpTOMDOotRL3DR+ywQuzLOabbzhNbelfztCYyim6L5PI6s4JX5Oynn7eLPVA6lCLQq8Yo+s
FlwOX23ZvuFNJWkUiS+FSihrWSerCvHdYHFIlClBlhf0d2O6FSNkVz/gKTGiG0GVcVPAzQfzrV8N
VhqAClmxHnPJF7xvXjhXPYHl1J7nuNL8ow0N31aiq9mau0nh1g1tDTFJzh/xaiEjkk43A5a4gfQO
Qw2VAWo4NeC5KC1MzpWd6nelcoYFOQT1Wa3gtWARMoPhnIPL2Mdh3iSUNc/OLKXS+TOoVP5zMVPV
y0VxA4VQWjHkNNh30NQMTQ5KkV+4cRhebvQFB8dRATiRdHyHy1NPU+rZ+1s0f0ok+k0TwQnV4P+h
+3TuJ6dpB+BF+D8FIg99PEjbGpy6LoONYBdykAT8dvJJQSLq2dcfwz5pqgKaepTFfSTh1U1AwiJL
IHebyfHl8Kir+fzQ9G+vwpE9ZrrFDusTYw18QkpWq2jL8t1gv/R7s5bbEYZt+0w6bgek8whsArDS
fRb8fk5s+5TpgiUQPWCahxZH8DAvabhPT0PrKnuPYBOhY1oOTOJdrt057+FfkmNPyaIDFU567AHA
bvFlzBeW7KsFxfaelu6wt2iWBpVtzt+BsXbhk9N8QW8VRgMxmlxWZcp9fUdATBc69MsODpms9zE1
9XbF6y3PyNYXgEEcJTF79c/VRv8tnCCOqVZq643WU7vjxMmIj0QB3rlEc9FMiLhUWbXhNCIiMRXl
Eu4jN+OFFs872QdzlfbkRs47PsFQGdxyj2fubVGuPiqMXoVO76ie3kMeQyXSvk6i+ZBBGHHXeSJz
QSmwd9Fv5Jns4myhx2m39dIOPnvjh1fBM/AbYA5GOXZwSgfHQTGbbZuoO43E75HUkXqpT1xvK/DO
j/sC6O8+QOHeE/+a2eVOhGWEioiMAUINgKWiIWJSCovthjGfrllPudm14iEZ3quw6vXEDmwvOB8r
T5FiXZBI6fcbfebg1hJtp60opezxvFkMZ9979xjuEdke71XEGdnFsWl8HzZ6S32S8KToE11HEuZK
nAd+BD8YaatUCV+oVdzq3FtB1rXHfaSB7u/P0oWOsoK6gZzhDqEcAUdwUX4N7kMsqy2IsJ+bWnSK
Dg7uozyNDa7XJugghSO2KupN9Hbn3GHu/oPdadxga46GY42QfOSFIw5SWNqF3TQ/i/9rbvy/GaXS
B3wVC8CojkneRkVQV+EQ8vNy23yxqb5surrL3kt83mm7rU7XogcqZ7E4Y7YD7V5edn81SdoBIcjp
nXPxOBNB66zmChM+84c4+++S3bvnUV+kTrpCbEMR0WoRTged1pDOZbn7BPhfegWLTAPZb3Qho89C
wVMFLHnRYh1fPRIZpXFwGRMpnzuKHr7s3SnxxiOqE8y1a2zB20tREbngBBdYI4ur6GhuoZJfhc9j
h0MqB09WddCkfwIpHkcmSICLooO3txyG4UC9rHyjdLthS8nfQVY4LDmGaTJ4dqRADI3cUubndvou
88pFrTGCA8aKaXZVN6W48EwH8X1eWSxrGH/LStGVHP89rvzvdhqXNlIgzpDcDnvbenWJvc6uWeJG
MKx6azRLSyBC9n60P+KYoIF5Xi47A31z3em51s/6R7VywWtIW8xQ8hJhIsWiX2aCVYmYT0Xg9WRD
Qz1j1SmurWLiOJgoSP97PTeKrZZddjYXVLOBlDc8RGa2I32LaY+0AgdkHZTZWSj7la5r3PNGwapY
BhJr0tY+Q1VR6U8mX384xl4pB9yhe02FCi2sY+YFMYwwbGfPqSCDFE5QEsaQ5rYRJtRHtzHjlyVv
UnmxxGVHYvnQB8HXs9tDDmQZc+pwdwkB99FScdyDGaexaJWbIxH+T6xijSXSaTBmFBOsKksxeCms
pg0Ur40CJ7PE0qOwtbWArmz263Sl6k9BBSgMVyIUK4SA5bODYzDPq+sG/MDYRwl8FLDaOB3Twe7s
aAZ2NQm7oe7f2blERZFV57tKDbwIsfyOVfJypYdFLi8yDR4Toev6CM/Gt2BHqoBKFxAV2gkXiWez
uqQFnVFFLqL6nb2EvXQviGPU9VhKrm9NEiyREur5214UTx4qtrye2FveZu6LH5IUi0x3v/9UzQcu
eHk/74J5uVHqCVp8a5VSum0D+kVCd9381Dzm9iVcQLymgiI6DspyVUGcQQ1P1gWIJXf+dldiq6Qj
Tdz+Ub0zdc0yt2wY2v+PrSbtOgC3UfUTGf1SSWX1hpWNzuDIgRxVJtGXBokH5USQRlIT+qJn16J5
dTlO+bgVMApuJK02X9Y4RrOnzaES9CFeUQ157a0B44GEg/azOL9aIZ37DkGxBvID0EYIOd43PYI5
TjfJY03dcuzjmZqeZ/ajRSpDxFiiZ5meWg9I429iVgbvMr+bflfQqecvnjBBfv/YxukMxzKbPCWB
7z4ljfQql0ViLbQxn5aGINmts+Kc1RBRBq7idM8SBY/ujWyPSQRGLvr/RhdJZ6mLWtfFPUYF7oUG
SvFBSwAl76OF2svF1bfltGlgY69cdiWO58ritg7cZQ5V76pHLpySIG9w7TsxVc/BtDCMGz8mJvaB
c/bioZphur2XyowXrRn7tXBowQlbvKCA2YsjWDqUZZRuRw6uLpudRAnMQCAZv8eoWwgcqUHg7mVv
rJSBNSU0J4NGLYrcgkEHrOEeIrw3Cz3OxiTrjoKULDq8e9H3IG39uCiCmetNIRyjQMrfYgtrXeTS
sndM6b3dH9W83MchNJZw+Xq7FtaJUhCEZJxmEMZbhT6RRZDRRIAhqdylJA0CE9SffNNWFM18k7Sk
2mOc99CH+zRssHFNGL0+k/Dv0D3Hr0DxDphxfE3innFK0Pbu4tREWC2szoM5L3XawqbGeueMDeKV
zgrl6R+giC6rdmNgjY0l9ILzK+zAGhJwNWNXRUJmMKU4nkAyKWGTts3axtuHxdfu8X865Ui9tU/O
PGx2OUvHGFTGTeGFE7SaE8c5s8Uh0qauslpN+7Wuk8a+KY48HgRc/P32viejxFN2qFcwKhXHGk0q
OvEWvceMnKEXGb1gip9UaZmfjn2sT1Tt8u5bA24v47XncDmyiBr4a5RIs0WYtxY84oGYMrtmVoGl
lYhkR1SatuQWHK87J7F9A8Hch/m81S8AVFYmJ85dPm1oavZn4j4vb09NT6u34XTKuJN7sVJM/fOs
Jl2RYFhXQ+EXfFozyPSsg+79sVSEUV8ZR5N0UANbZF0Oey5Y/gN7zGdxWZOM5Ocq1ZXiaxtVdHFF
jtUYEqHhi34NFgqPDnU1Rg2/wmwwBPR9lcY310HtRCDwjYfH+mgb2J+o0fx0LRhJUZaKXDqnx/eM
UaaJMUjF8w9iBppffb30GWpd20w68w6lNyCvf1XGFTqBL2RWkxezgPt4Lm3USB+9dv5EaWNg2iZq
wchQ9wEKEWvSuIDDPX+hwG5tD8pcSxEDPMyJ0+fuNoVFTg0RWgeQEHsVx51RTZsqiHmu25F67abJ
eoPXQB7GoRO1mAaUgkYe4UUWwqfeOShL/hUKMR8ghiCQnP7TLYKg8fCrw+vUTY4IHdgUkgvwNCpr
CKRRoipUyPqIei9hEwsGHLxINkTXEqckDNxst2FpClNGbMBO1WeJzFqYaem2bEqF7PEnetA8DTvU
skAn9c1tEizf5OqjrLfmhp5uj73HsWfTXAeFZcgqIRWAxMfg8rVkSm/gjWe1UZZOXTxdfOCDRuuK
Nsm1hlHFXttNLXr0OUDZbgt/PGfWUgLtH9eeTFvexEDxMwqNuvAr785ij5v0ANBlxfrvjKF60gF/
ea2yWsh40ExSodZSpcI4mUEfhXCAsrDc6Sk0YZq9epZlmmjUyMP1U0C/XZcrqSla5dKfj6eOdCET
8Kdm+ZkWOPpVIon8XL6LGQIed/yw1SkG6um+9HM5xgFTO/ldLXcuMZlViuxDGv8URLoYGilNmKb5
nreVWdXHkqpd0RnqO/vgQAP3gDo+UKJmEwUmn1cT4SuOQTtNMmUHdcWx5hoZPBCzt18D0rKqGg8e
gXL0BI1iq+UCTpcIETLd5oQ5Ztg5IhYEj81yzudZtyHT9KQof9MaLV6yHBlJduSPruqEf5Iks4or
IwS5YH0KmK47Flr1GIYczP9hAX1bOzUFlYnjP+lJEXKTpTrqjzA54Xo/HaO1+OdubTNjzgaM71JL
FHmJaVsorQ8/bKYEu2DkAI8Lvi66sudsE0XMIm+TsBFnGxZQsmyDU681oFtEncDLMYSuW2159t8W
PPt5ENbTonqSMV57W7cjyXU2YUCNcu8Hkt0zc+x719UGDTXbB8hkGWUGbJYD2/dzgD87Sn3QZ3LQ
HkxtFSvj9z7cD92RPTVWNKBra9k3Em//caEZUNbltwVYUbrEYDwA+U/UEQsq1VY100B9poH/TimH
CX6FLaSQsshkuZR/PyYl62gbUr7yR8JWo00bmb/uCg2QhJ5OEWSCCZ8rJ1fYk/+2b8jdLC9UZaBB
na4JZq6jNAOCuC8PZQ4we1uBV0/OXXZzy0Ki9ufh98BBmAsY3fNA3C60jBkfBCqq5id3ZfM28+TE
OHgC/H+LdhdrjgRRHnWm69WtEhjpGoA9zO6v6Doa3P3ZNUsJ4bc63Xyal3RblbsqTR9n5BzQQpA2
CcCcGCKV39IUTgCdjQncSuO7Osbwfb0Dbwo3DmA+LYJlF8jAT7wXifeuxF7V0koVdefHf93ALbN4
UshSR0YEYoMI4YYT0VQGxU5vr/PJKU/oUKFByNsTIKuFDjPjPpvI5XbOazvEIB9cVr+PYCQP5RDr
yBfKJyWVSvDnQQ07Oqx8wbUZRoG11g98tcIiWhP20d6b4thLue6RF3sszKvfa5Cx6RM1Ynv748qI
c22ONwa5X+ioM50dtVyHlPvWzUE/j2abc0y54br4YoOBf2lNiwytha6YE2fz7J9gCkdQszTT3jCK
adaO5mer1JwoDrfFFnMw8ialFIVLU2U9wK0DLyEnp7Ec1B/KT5n3n7YpxweJw9nw0Hy0jzUvLS9k
VElKgjdD94e5u+9Z5qDOPD9cs8fgdYsG4DPo1hRnMLxyI+yjyWyGK7LCg/l4rzbh/d+G65hffl8u
QEaYPugAdQvdqEJ/rbTnRDv4IAYbsvwLk7FoJsoBz4T286MTNiiOYL/aFlrv0M4w/VmMg9RoJkgq
7BZI6s/IferH4ev8m7E8nDjf+vCBmVgNITqMGtOt6zNVMlAyv0+n3y9HwH2eKvfsEI13t2zpInUe
2XPnqkSEh5H2ypE7JodhjR4ffqeSfbYRPIbH8OzFSy2bxHb4vdP2e0qwSUxAqdbwwDDUpEg95C+I
fjuI7VSLK5RVi6mGM3vZxKyeqRvXFT9pk1UfvMHACaLP8U12L7S2edU9ioakx2QA8PpEx82BFPg/
RBtXfn08L2Dh4PdcZ/soUJq6r6rIZNVQ7NtD+3+m2usnM1baCLKJEDIBOjebwXs2No8JsCjs559/
c22FXphsXdpXteEJMhhnxgeompGdTrgCKzkoyYNuraX8UFl/PFoBNQQpdE4ZLGKTc4brcGEzq540
rRVlMfv9QDDe58JJcodNL3ddROuALeiiWNBOys0KCAqZ0cSQzQUm5K3jE97YBWRwScNa4MFXT+m+
5+mfwqSykLrOXMeq5/C5/XJ0WzCU6/yQIMzoVHbDID7H/8M9nQ3pZ1aL3cUOA2pPZU/ngh+7D6x1
vRlXstwFVJivbRqr6ARi+DTO8wq3T6Dfof53/glQ5NkLBfN7Bw5mYQYIB6OpCwgPI3sHeFcy5FAQ
WfT09DYvVyrK48ttMKZ9vdTpAFPfY6ChdodDCUWyRxjJw2dxa8RRl4VupLiOUanUHbG57Wkq5NW4
Dp8GrRIl/KZW6PRvgAPcuiITYR7nsmwsSv11MZuE/kS8OSX53EcEKGJSTvpX1socv+Q6/zGz+shr
xRvmuHJc5nCwRumidQZOAQ5kvZqcP9NK1di2fdU8bk0XJZgQqULv2YleAJ4gaNqJrGPsqAAxK8ev
zFrWyPU5OM9WnV10aHZ5YqUC8nhs53euFW3/YnuO7P1ntT0UxWCUuM0ZDWzPHMHpSgxnilc8VFqv
PCG0Om4E38jXjvqoEFYHCx3lxzBLRENhTVSk6SLQi5itX1Pqam9H3X7/fqujoGHvrjaW4h/J15mh
7z5FY6DsSxmDQdTGhieXhM4u0FlYGVJ7I1CWjGHQg78fSYqKRnm+KHP5J2c88VA8xTFJwwtdMYpf
vvktMOJ1Cs3bfT8ciHdBqXSnRFQ35wkKK8NClbB6ppa8BkDFW65090Rmtsu24VmaPJt8VAPB17EU
pSLvhoaSP/FMikIiGl9oRBIWgN8Jm7Hu8ymDvl1WakObRv9H+NaTW9EeZJ8++GnwyBu9UXU2QpSp
dVy8t7J/UJtHQXT+p3VXRW5ijzF0tu7/1amYFe1deO6LOwCEwghiEnrKWlbFBDbFGKQDUcuTqJC/
aITwcnaPwhIFm4MVnXiU/WEv2XEbKdBK9ld26+9N9k6ocBCHoGSELFeHNiPFvIuxIqvFsDkQNGz2
5V1xk0RyVJokf7+uP/LMN3tTTf9YJ/Zaqn3a6PDqA+jBF7d5w3j5fESZ2UXr041RLVqoMJlyB09M
bD3k5voI2RURMptzGlge6MVhp4Fw/f8+zyloGzRe83elIA17S3rF/OEuGY5/kEXx3RjHUH8/niH+
hG6cAc7PnMXCKdtevk9XLAr+Dl251KPL/FhV6ZL79e84VdcK2xQD50dnMLx0lDhNXSiRtbdn4NS9
p/+io/5yTNnbXmtmVjEa8WS1uy5plG4biGNLRP1VmgHaeBFzhdYBscHDGQbKvBuSHNWuTDscHd09
AoEUJtQVUCF/BjCkdMOwLg6QXFq2GxOda71h6dD2sngvRUsr5JKXvyEp5p2v/oxvN50jQ2DzLTJ3
6AUJx6rsC8pEAL4oXD+JsZitVqwlaTuC8++F3T2rpZqkXGVZvtFmN62PmIGkN7dhg2oAy8cQ3IZs
YMZAc5Jp271G7/haZFNgIIeI8pq+WX2IwBajLfWcn8c8aboLIi18QgqJf7tyIig02QoqnsRXAPfG
CRvDGwasa+nWyVhXVKxPvVKBQQma9FvBaRyTUaGxgWLoG34Xc2RcWetTzm+vC6RxGUR9szoxMczY
6gk0L8ktx7R4WvonN004qWDOOS/QOszy+MBXaFcjVL5Uytp0IbAz6sFQkuCnvDIzQ5M7hLYjlKX/
SGNf0iA2/cAF87HSqnbeEBGfSE8rZqOGOrzjh+hKmLc3VvKmjX5SXv01HGQTAdBWB2Qf+v2itvhf
dEGoSjTFXlscApIq7GFVV3zibNlzxPcZ1qeJGUHRWvELcu3r0dx5iZJYgqZdvAL3ZxlMU+m6lATQ
p1/dCsL/kV4bprhzA8n9au8kbh+ZydoW9kINUPpLdlHunKtE4eoGbiDeigN2rYBVDkr0N53YQnKU
dB+X3lAWWUhdimGkDwgpfBF9TD8L7yyNuBZhP1ALBw+RlRg7vR6f1vJqRdHA0sU0zah7HWZFkhPA
6qP3tFVZNNSOLKV7m3yj4ZslaXgkZ5EwBG0UINDO8vUw+ftZVm774tVmvC8o6hQMItdnnfBKgsEI
/KK8WS/iATEwwuyDhKTKwEXTGkWknBtnqtAtgcEOVLzqTI5f0T3t5WRESB535TrP0P6dK1d8YkBr
h5+mOzJfPC2512bdeUyuTr95MDjGGtLG5J9SGgEdX0gOGkSRODhoa9j3hpaAjQY6nsZJvBKHJRmB
lg9piBB2VbDnrWWs0xBs/yH/VXhGtA9gEW39rfWdeKBxyhzK1iwNPWjt7uYl39NY/qD648ye2JhC
b20tQCOoZ/T/H15k0z2d11fd6ZDN+CNFhg6vgsBIGsh9pmgPuOzc5HQJxs1XZwa2TTn2i4G0CgU+
SPbgDH7OrQ93Qjky2bvSImFiKKfNfx0U8K9UEyOGR1bEeBA146OkkSE7n4DiInqU1wd0pMjw/9mG
B6mF9lEy4+cYPfCkP8kSpDnbqY9TuzociLs9ni0QQ2uf9+slo5c8YO/KBvMMAOgC+wuNOkkhU2xj
mtY4dCrBaMo72SWJBw7C2RqVdlhZ6QWobr7QrKixoUyWDSFo1i3UggHEF/WlP9apf4DZlBe4dna8
nia07nVQIn5NqfH0lTiCfjZ3Gq03V9dFwe38tMvVSBPJHLuRWA2lxFaMLTCJFQLMQJQv4gyTs4tj
CjGFWKX77BMXM9+TATjbythHs89EHspXjH8QZsqp+XI2fMLDoA/oDoWzk+IA9uBe6KbyLxYYZP5g
H/gDXxtae2D6bPRl0PDUGvxG94XTTea27qoBrjIl1zUrIR988EjGrGfysX4bL1FY6dPFJDgN5/UD
DTysFSFqgjVHb76+9riT6uBKGhHtr701hFK0SpPnHsDxWV5DZruFdXCGkP9oyfXhCtkovaJ9nhli
HMUr7aMBtdWfVsHPc/foOkI90SDOIHX4YFQeYUdY2wj+DxT4xbfoMTizGSy08EHJ/ZcaX8r3CSLk
xE/1i3pVSna2hz+UmzLjUASA7TrhsWQEI7HkkCEgBFFpHFGLDOEG1dd5+q8zyHYe0j5xph7os9tv
fA8uc6UuBwrMpEnTyseTFfncQOBSiFmK2IIirf+DV16LPYUa+cTRSqGseUHkT5Xzza1u59Bi3hDH
pZVc+UN8+w217DVaqVUwE/5eQSQoR7cQeVe282s1yOu6tLqawFgUlEzIF1XED7H52/IYhY/KC2uc
GmdeG/1NgTGCqzlp+//yBQia6hwJQPiZwDxMoJCBGF+df9DLT3wqdms0Gf0hgEKv4NHlGO2vJYIW
J/43apK+EFlQWpD6msuVUhhk3tpZc3IDXd+f8vKgwku7FcAz1bSqWIe3En+WY+IAzM1znVac2XCe
0xq/XNfKATuJqIgFsP5PaWUc0JTX2CX0HaCUGMeOU5fOPFXe4JDfDL8dve97IwiARlMMqTObferY
0932s/n5wAVw5R1rKtCUVKRZmJiwIc/tJpAqyPBE6XbEnoKTIsW/D7xKw3L8Ku6SkZkTOnOsM3K2
u3xI2XGCV9SrHm/DSKbA5i6AIQ/yEKhiNW0EyV9PQ3+c5+5l0d3o8HjqV95P393VzXLHH2hU7GOQ
25SnjSsjkVIn41bQzWTVhrPH7Pl9FQ14wwFQwE5DVOAfe8QkbwdumY++Bsz8zfA4BTXqdBVTclhi
7oWyfCsmxW5dta1e4uWoMzWI9NTrZQo/mHQUQASZzJEy/mEKnjuNPzotp1DfUKEqIBTPl1nKZvhi
RewouY+9Xy5n8QKYLpQcHbTf3KPCtl52RC8xJXax0Q4OgmG1B2tC6Envx/Lzu6+D+XQ5kEjwHmtX
PZ8eR5e/qmMRc/v9T5MFQH1vbY370oRm+1XyLhLixRIDfNSbO31I+0RnFJGistYygKjP70Et6jGY
aj5qn8bjKVmD3aMFsr1FwHbS7BVmUsD96VlsWS6h1J6BtAOE+9lQimoAtj+qeWGvF52yvKpBLxIJ
Ex4Y1MEOHpcWLAjxsUmVRrHb2bEqUBVDqYU3qYniaP2oyMtUuESfh6NTu9usy9MNBeI96oa7gl0i
rHHFi9lKmuwMgN09Xq0jW8S+umwilg+5lWKZPqsQjET6b+eotUv4BwYPMOXEOA1dXiha4GWPeQn1
RKBsvoMZ3QZd6oTCywug9b8n8k93Pn/nuM6IWBBiVNyyIFzgpya/8RW68b+aIX44v5JSqk3uoIDv
OVn1FBE1fBLPNaeOIxB/wLzhE6h2LBQDEcweb0ijZptP60uUJyz4Mzqq4D6GrvWv+PkwV3v/5hZc
QornanD+UIbHp+w9kuDaxnXKqvlP3gnKbywpJoBWZjosWtG+znKF7zELKiXNyx5v0VpLlhcUH0K2
TpkJZgiTjpwv8zhqbqyk2Jqn3nImeCIUpPpWvyQhJoApT5si3l1+SOFty6iJ8R1qQKH3+JYDQYA5
QkkbUrY9p7yNnUSeGTD1nPEW0Y9BFdaWLVtuy+70yOjw+0E1OMML9Q6X+sDhsv401jJj5OvJn8vd
5oYZMxGyZfCtH5NJy4oUb0Yzc+CadZ+46YMLFlIO468HWjk0PKB1TLKO0rQJ4wGMFtzfwJauGjbp
xMMAmQ2bKQ3ot9TKt+oDHSvUfAbcjp2SikUn8CkSZtQ4WOYs1n4jAjR5dvUG/cjj5nHhdAu1j6TY
9RGgd+qvWlSUom9GodL104gwrasvkFJLonOvGV8EsQ6bjT4MRFGpm+h2Xu/fbh7pfcxviQnCkT3t
fHmn1qEqbvh7lw0+T81ZM0gwY6R2y9c22Sq8iQYWnC54lC+6U0WWja3tI9NzT2nBfrbMKotjEgQE
u44V728I2rsBe8g1T+oRhtcjw5t4Rg1MlX6YRf3H02X8G/oytEqaSWieaRndt1vt5/PX8KdkUuHI
pdtY+MSmRTiGuIY7PAwuFVsEG6KM43iXyD3WlN/pI8p9D9HlLXAw076UiAhk3Byv2bWo0TGx/xPI
KLfnY9706DEFbBtJRINELVeFjjBGx0k72Is8Bm0NUFiF8wLn6mti6cl9Cgo8G8vMfkEPM7VhCart
LDQI1YOolrwgKWJiDkO7tH36edneeJNgCCGmLtN5z8shhEkYyjGbOLDEBDD1xbB7RpdCHvNIZi45
xJCM68KNYE56iRXLkWASryQhdDwZaBV7A8uII3dRRN8wJhrH54e8zUm7+pwGqGWe0MblzUBfWxoz
FNNdMhoJHW/Xz/M/M/O8+nsKAL9g1oPLTINwHulzJHBLIZtO7plcUShg6pA05euCtIZehPMEWFvg
Y/lvN5hFHcIWRcH3f/DpZTMDdNS0o5BeMjzlaAcUxWvF0FJpSufHdnl6AFRRhvmY+MJxZtsWwXK9
OMqq/XYvBR3+E8L07gGG859YWwkKm5FJZAZ+/qDkZDVpsL6+gS6qflxOrqHGYz1XE1TJC67NWiNI
myboDvUE/Q8QRqtfCHmInRPfFc3DiAUub56NfA2holy8hVjCP++cScPEq04BgcXqipiElhXohwnT
tPUsxCkZcnUlxE4XFxdhHBVl7noVwW1XdO9y9m0B1e3GalLwAZkJvLIpiAbPhHJlsYWLB05a7Z+l
vEdkBWIViGchorqTwJ1vvXwp3Mw0G1kPcOCquBgGFBigfQHuG2IWnFWu1yY3xogZc2Pz7j1HpJKK
Xk8+iX+qMo6zHZYAk4Uqweuh82yM1tdLXLS3/9YEaObiwdUTNY3oy+hqK7eInk43dE/+c7bv1uOO
yfTltK+A7bojuoFZ83q3eVj7XhMxssOcwI39DOGJ7vpKHFAYUZbi+uLnkVKKZI4CWJ4UfPFTYqUi
JGTuCMtsjFk9GyePOrLrG6wKan+ywoZDWoFRTJ+tQilQ7LL/H8Cm4PyIKJ4IgANP+YwJGAOs0Fb1
LHtPvNLNoNp01vKMOa6X+zVB7uGo3MoqxTO8lhrPSXB2998TadH+kpUOFdCn7KG0k3DyOVhdfaCK
nwcWzhU5uE+EGLDBcLNoqIYP9ou3ezDAy2OpQUcqzTx6dhbuIUiDGAu8SA5+8V38Gh9PmvhCiDC6
8lKYRCM6Ia1hyB90VawaJoO/9PZotGpvTIo9yVeaAxK0UMdUJeV95yckHd4nEb2KoQ4KUWQAAbQF
DBqTOCCXctXXjGcE+rmjcMtv1cq7oVcUzFj5tPMs2H525DUq/CKcBT8hHfjDHuebaotf/TRRVR25
aR1KTtcnJDtWyHmazTSG3huddlAZ+WZPAk8ES9HhWU6/Rh5KKq5WQj8TMMS1VGG2Nhsbp6LJMdBm
MMIUmwrQhmKF8Lkq8xWnY1glahoTaU4sxyrO1+RzQb/owFOj0r5LL64lDWPmw333zJC8JxI0z5TM
JoKUc6EwtjBbQ9JwPx3TCF4J426mP0htQaT+nBgqhGzXw/94igAJxZOJhSA/8xiBelEcPxwL8cp9
VIquiOxqAjtUcwFzSjAc9aYZ9KO0h3JSbFyqKB6Y93Jb6dzzw4HNrRTmRlm4amGq4FV75SerqhZN
mOiTZY/RhF0XMAM6gAc9/SfAwsQ6vWkfosdw1SEUr0qenYuSrsm9v3u3eV08mHv09ucuEXgdhCbF
O78/vUv6Zf3dokwDQMzFPLfowla6Sddjb61PkHCnv5zc1bQdEdgpfdOrP4ATVaIwZF3HNCduB6KR
F4BR4eF9jiJ8KO08gXHBiRr2NRmORaNpmZHifTwVuRVTVt5YoY5vGqP+32JRJx/YziPsNyg82mSU
MuHp32vhIczR78E/7TFEWPsdoAS0DjPhfG5MAyZz+2vdqz1eydmp5D4UF7MBmajd/3Q2sleqDQuA
7a5VxAGHMlGoPLY1sKJLOiBGqKX03hwxkTnpjsGnbXi1N/BdngYpinnv3MNCsbX0P3ITboukSENG
ZhyXnYQXAvmYyff0iP82c8MfcUfKEW9Fhr0+8LWap8AoNU+hNhsruFb6xOCNx8cApdOvuPU0NvC6
N5B/qlsoQHCODcLC9D6Eef8v7VF+tmjCjyWjMbF8y2+puezy7CEz4lJqUj1s3TOdkM7SQwvvAq+m
20DvoxQDobXLoB1DTQ0D2D11KlltZt1Inn4x/l5QLmkyCJRN6sBjSX6N5EtwLmjuRKiaVr1zz/Nz
FhI7WYPOTDZjdkZe1YLrz3r465iTfOUAyy8OTHlDGbgRJ8gms1nZ7MhaRVhMcQjD1XrYS814D3Wu
8V+YsXRdne7m2k8Rlb5ameYhn2oyVi7df5oL4MzQJgoptrHuS962Occ0LuU18dEKbJvGWk7S5DS3
XFy4DLUoVaqPKpj7goVV8ChLDvly0zlaAovuQey6fIs2D3eVabrTDkMBHeFUkBCXkfH0eXpSShA2
fuB6hxttLusk/etr/FseGwmD/REoySz2pz4XpsU3Na5sJbBjKHeFL9kUH2omUSen1VdKLxOlgWVO
9aHb0ersQqi/QMiN4rP/IpO5dRuJ/bBayobalv90ITRYolTCGYfvX7imK0LzmdtdxogGN0soh78y
LSKH53W2jGLD/Z+txkxekjwuxq6c7cg6MJvVAWsuCgjAt9fC1Mbyv+MeZGEc2MsLvTuwAQHJlSxL
NmtLFCse9J3ebIyErQ6Vd4kNx2GBT6Rk+GS4wwJq8D5ogVGB205uPySjh7hHC3zygS5wpEyJK81Z
+bUS4sxLVrdk5nu7Oo6ylZnbqTYbcxIJwrD6eWciVmu9M2JRA4GufGZ45BnRNnVXk1JjL+2Gfo9A
nG//Jh7+A5QOdfUIUkXxt5xTHpTRBuOCvMbyxNBozKuVhu1BwoUg+kkA2YCv5mW/VQYMd64sRPsi
O/TjG49ZFMN3HqdbFNM4rBe2iyFhzmWHu7fxCKiQbtmldDElWdAqGEiK3kG2jl/Q3yyN8aTHAwhX
+2tu0ZWDS3GejFK+ixF2appTBzia86A8w8q4T1W7jAj53I8PRzRz/4rWFFUJ3cmdqjPo+NKbwAYk
HLSWReQjY0WgFU35p8FoFuIH72HBBuDSaavLXkZIGKwhJ5HcTKxWbXg9mFshgazKCBmjgKFv89xb
enk0WiRE9TDjXM60ZI+SQznR4Z8H18iLG1K0zABYNMlQvSzRb4FnS5vffswOszB0DdJvu7cy9Fwb
K5Bmu3Y0975d3/6+FG3+Ppx+bvLZgS69A8Md6RlC5KypfqYgfIpUwKXP4rL+tYkxiolFLbqD3zpR
7xAvPQFdrp6o6Mks/TvpRhbznXTyRW/uekgBg7McvRLLsICId6vcSOxyRO4pmhUlEKW8Ginku0IJ
wwLcAgSOX9dtU1R7262vzxihTg2NAgqKSxILbFcbqFrUDJ0yB26Ty4V+nSsJGrFXCU/aT0dGwlcw
iiKAV/0EvnswdmAJyDHFOPM7I5eNPhZHwE3uVD4M31vmR8HOlfiiQIv88oz8IwnWEMHP0Th1+To+
oawiGsOoBgW7y6LPecxNSUo6WieroTo7/tpg+gEN6zJKOAs9v1fFGRz5WuDhn4sBCVVeztCjX0xk
6b8a7N9iafIsPdd/9a6RXSKqrQKT0h/81ip19NVFZM6qMaipbcav7eYGtpoZ/KoT/dqjxGkJx3zL
Ea1FGCcnUnCMa4h513v6jFCXVYuIgPNWmy/TLsUU36b+feqJMwnAeEr0d5a5iMtXvktW2ZUmmX+E
Czl3VHSMLdjV5hIsJRFFiZtu1cjy9VWINLoANTiv9x+vqyipwHcVoX0fGUN7fueEdPicGx0vieqn
yZtNVnJneyrdCpBJOLu5Rp9oxcP0adT0tIJ9tkyIye3OoENrhOhTpG6whXFzOwGJ2zvB5yEvXd/U
Wsy+jrNWubr/vJY5++BIVtI5mpDaxSIaEudrWjd71eM8720k0a5MFX5JLOnOwaiqPEuwNk7H1Q3E
ppze8DKu5vvJEg62zHAfvRk/Bsiht8VB9d7YYzT+R6tMSuJlCBbKwPf5ErldBkIuxepymZDHmisW
+gzl3OeFqf2bPXZIuuFUhTFE3shA8RltAMY5YF4vQ3+03Mk0aIpFbWpFgrZJTptemhOZ7c7yV4aE
A/2wkeW/hf3drH6+eVBxyrnX1UgMLktG85BGnQ6jl59ysfyy98MlDDxefRNju0R9jniKPcpLzbh3
SbT+qdw34CE1ORvZ0hnhk4aDcMXkCITnR21WLTTm4/RMIBYN7KqPoeGBUU0dzUakfOwjE81NmGSX
IOaRVhtHkaMVOBJYUvjkPjSsHqPF9EcKimGGzCBROdIFThNqKXbF2Cb978wQ5zlb9MT5a5e6W4+T
5+hmUscXac88CBnZ+0LaBIlle7baPXChXxwiDIJMyl84c26aBoae/XCjvcJjx7NDBpWwsq0tKWk5
CnzQqxGO2ZOyf70D0J5qFC4BRr8w99BbYBT9KQ13aCGqsFdHyUPTA9Mi2HCT34cZqBBxxLb8vIGQ
k68rwjQXt8ro3PCwS0+XSWTXCNAp9pLrPRVTfcT48AT54SB+/R61rcAYx77HI5yarqBHqdZUmdyV
4gREwHTTfIN0nXNNfVrtIzhEBLGbwue76kWFCQxtwtCoCBxcMDrySAXmVi1+zcpyb5zxov5Tq6EK
AGxzSAD2alewU2YVjQQx78c8qMlKmQZ0SK5H9TKS2bQTTrKjcFswMTpniG7CfanBLXG3arhha/zr
HVDEu/ZKXvNuqwlShBb7czP3PdD+e/R53hWyxNON1eCak8n7CxhTouaVhK5q6S+cBGDq39DPfKU6
b52t8bwYwwW2PeHA5SrWClsL4hHj8U3GBP8EVTek7y6uRSrpIv6At8QvxbyBDQGmc7RjBASiKD6o
pChM9SLa4ID6M8+RE9Mg53wgUtSCnQRxX6bw3EfkHC/Pxnd7QnLFXICS76RYGRW1ConeTnXH2vgY
aFY5mkAbUYLXXfYruJUohDv3lmgGMlfbLukknC9B+HlwFca89N9duDY2lTc7ZTCCrUnQLFy/APYC
i6qCEJ+vtORIc6M1roUwGbLrP1i2WTsc9cU/xDStHHKiBaPhFIKnPQjEuCt54Nq+eN7gwUQiSqiQ
Zs28UM8vihJykXKLg8GtQPhK4tKGOBwOsSRaUqFxqutnHnbzenavIOAfxN2q/GJH2lmiOwQfF7R+
SKe34TVG2565fsbppmyWG5VVfRrRbzujm9wPzXmkPBseyHBF+/xwh2BUrMOymyz0HNi3CGJgdOs8
0du0dHs1EJvmOFGAym94N/FG5txNmDPLwu5dX58cJ8kAIsF1f4VFWxwMmc2wIkp17ek5qNyDhHFm
OPaVA5FgEC020gvbjLcTYWEI0JIQnYXqtTx/Rd8mSJFW6w7nTaBCvuQ4PfuYXfe/SqzB/FMOTbMc
1FbNmkehUoNjrZSub21fyKbb2RfIZVWdFdPksM80picmNtx5YUFJVWYN92blaKHo6ogryv5POTWk
/ganhVZJ9NzU9jn5DbYyJpdEsXCsfLjzLOFk+54QPcOuyrPoOBbvwExRwJYWNx5bq9M/sFgq6mZp
bqtaJO5RzqqxCrg5Nyhe8ESQHDp0rzGHtxPyznvbXFBmo/NGQBeJlslfD+oBuPBIqPPpafXLu/jY
XkLWEOsucoIN5b4FgwwBpcDH69YgNHJO2jtk6+dJs3A0RYqSl5yqa88BkPrwaCrcaeC6krw8XCD1
LupQwEcRF8JLnqCZTirlSoMSTc/32yRwxzj9Fp6Y7jLJkqH2F+i7wgVnYop1DEv7ymu3Rvhhty8u
HeQuTSfrGcaeAPXlEUVAP7yleWuvPm8E7UhGikwdxxPrvtcfy0PKhlO1+PBTgoLCRjbXHFTvX5Bc
xJZVCA2g1eQG+4ZNSYlegG6jjeW/QoO0vZIUCmF+/ZtHTXC5YN+icMD4OAqJnKWPnkTfVobbIlvB
zdTlJqz39/bdHvTyBse5NTmfvT1d1rjdQwQfbuSbxIHCMYP8gz+I45UytnVSnmm9vyEFIgdcp4E+
GNpAgSa+iu5ll4PJ5fjZz5+bVfUiEadsEZzosy5v8UB+4i5oTxrI729T9Va9GNSoWwYI62zQDHy0
1ijLS7BRo/CbAccLZQ45C6VLZ1RFJhi4XG+guuw8DCUReVHoazjIlR/Z0KUQkB/LMfr9KGQjBxV4
0huGNL6UtG8MqKRQS9MJ/PljitamfHvA8JzoS+qEeMR8i+G0ceynDovH92SdwqDgiDG58hnysh5E
HAkppif/pDbXbfuOlekRrGIKFXVbUd7k7D/gxPI0YOhwxhXakBfb9J+OmqsXY5LyRACXvh3A/foX
9sOI/nNm0/JKbJmZ1/RstNuCKrLiZ581lk/LDEnJEt/WscEVS91fC1SXbe1ewM1zHDmUamL7F/xj
fYojPc5vqOH455LvaZFoZv/2v/iXZ/tGTGsvpVaWTRHgUu1Of7jFTxHxgC2X74nQadLGCN80NsMP
z8DXy1FXZfop4I0EOkKzRSy2t0ytUGpjpT+zOPdVCiLxqIQ2skQ+ZNFspYLqmVF1g8UDB4OE2dEz
+DVy9gHDhWPQjjf5Whtm6xbgqATKAJU6wa/DUZzJ9Z8YqmDALhVevLI9yLE+hjhCC2tQv5bJ26Wz
8tKXJPvtok8oDAxmntMlK7rn1OZdtvtKw6zrxho6OJS9I3mYReNuwmaTM7XONWSeheHnGBOO5cFY
OiXdeQcwyZnAk619etWs+uOO7596ZXAp0L3lAwWAYw6OdEeNUqvHF4buTJcBpCSQwAtWOkfpA995
NRwZDG/z0k7HpV/ECd8WAK8gErQi1tUlOgmpgw1lRRk59Y6AoQLa/9jBpkoSbjjCrxwjejQMjfAS
h7PGAXt+QQC/4oV5mv1BSrSnIlqGf0+hF83EJ6whmbBQ90xRN4ynY9e4nH4VAdLW0AItYJ8m5orQ
T4M0X8qea25XceC8OG+Y81/lPmF258E3GU2V6AkiJzlzfB+nGI1R53nsqrX9REv5YBbN6WLlC9jA
DGND98ps3aadc2lx6e5CyEVlF+gtY2EUF2RO0ZnscWlTSshHqYGC1uIrDaG6NvmYPgbc48FLna7a
vnwqT3l6m8xWhA/N4+wcHVa73rsV8Q4szctVQOUtRcpm0VlkLpC+09TJY+q9JWLR2a8T5s2SNWvh
/Q0gwmoWJ4M2Oh0xDy4zcsXxMfrIDxSSjkLQln1hZhzbG3bmGBQALnKc/nEqd/04AuqUK2W5VRFj
PY8aRjxrAT6q66dcV00zTxzejN0zxGe1TJD1KrzET+dWtDl3VindKzCMEgAw/lipN29tSf/7mQkM
73sQD3jHlyF89lXD7/Mrwihe96JK+cA2g9hT707P5ruPIAOf7T+b9GzM58Y88Rga8ugBwX3P6kTz
MBsld12cTlVNaaFE0tbb+gOIXFs+JbDxxefPRr2+LDNo+0Avn5EswEjKO/igm1UgUMNiJHn6wU0Y
LUYDLZfU7ttAK/uywfOP8+sIBCoJA6Zz1yF3vN7UkKYCRtRBrWuIBNCip+Vxv4iAsnqon+cczFha
lQlWZKolC4Yte9KMjLNM+4MNA+DEVidZ5iK3W0u6YTQ0UAnXJV6NWAPhnE0qPCHSBTFxNcSR+Dj8
Hx8C4oKkStY3pUlmf1rOxd9Qdm/T0Ix/iITI1qcdlvGvqHhqQioxDo1IloMQzO0qW/ypb2bISiB6
U1YPfBnTgZceuliNsA+3eNU7q3lcsoz+dWoV3gEj51ufW8feTKHH9kQQugFDKvw573zGs8uD9yUQ
pxi8YXMqkkEDVgY5qzRuD8oE0B2L/rUn5Wkz0Eq0rxSk5cFKkqsOxxDIalO1RWjPrPWIhREjMTaH
y4IKuNi5UaxXSrfnKsm62fA7I+Rv29YDo0bjftianlA3EJ/m5F4N6FU4KhEf7aK7lw2w3qqADvm6
HKvApksN63hgMtliw/slrGe0HskdVijwCkjwhM7ptSTAq3vuqifv95YZ3R+N0rp+RU2OzZBx7LjU
USD9MUBDG15YaaBz+QPGmOHndzfDgiNuk9750YNBcJctSnG9gNZ4xc2ejfBpqa1p4kYl9BYoDFys
FMrUprj82Kv2zE+Z09khWmwaaE55cYBRgy1d3UdQrYuSkfxVCrx9Nj6uRVfp3xuLTeOB4KtQYecv
/jKCQi/87Atc78Q2nyg75WWPc5ghVpIpSHe5Ikjfk/KgIcu1+2qO4UNKTi08jW8bc2JVtSWMtxVh
iUyrztRrN8ByhfsmPtYa0bD055Qgq/KRi/ne+hdZ4axSX/AUkSx/4Kt1C5l/FW7EZvLC8gmMn4V8
YiOUrRAZZu4CfXK4I801dgIIf430OrO6ibQyu1stL9zIl1AaeD2ykRwZvMFjnnr1QmMs2cLxPS/X
ctsBgm1M2sizPG0zr019rBiOqQvS4bs5WlZBhBsCXEWSBMNWxUfhKhFYKuPy6uPqyCZVSY9OgNGC
DYC/IUi/em9gjFSDLCkgGA+1kLGTDEiqHVa5XZQCIPq/gljiuBXAw9MvBNT84bitO8VfQv/56fUC
506FVbh/RzXulb4SJD4KtTrbH5O0ukKJjPTIjhf2YztpYCMl3pvvJD5cubaN3KTQcCZswBvcc0ER
0CSQM2TlrnU0yhmh716tx6c8Nzyl3CTJDB/OY3vsvXWvy6WsZmHPtf0WfwKz9gZ30njIUuJXjiqt
1tsQSEOZlreu6865MuIlhkkiZAc0XTOidXPvzjGpsh3KE/lA32TP8+ReDtX/F17NRnutCOhl2kbV
HY0qCPVOfKSD1Fj+EPyfP5hu+/0JQbjxmyU0AW/10JAM0kkrMI1Kdxz4TGCU4mF0+tp8LUuAwSvJ
c5CQPmZnPxwhgbyGLOEbBtWYue+rWzYfn5CNOJbw2ihrrCerYONisxetyPac31Mdd3rFxFT71gYU
/8Z2pwruBvBL4kNxCU9Yw7XUpavvCzVSHsxXcgUq2D3bjNyyE25W3CDc9lkJRgfyuMmpzsSGvrKu
1qPOHptlgktq+ko9cGbtofRSeqpwWXpS8g1GmW2iH1u0biBW9VvMKCNu+u5FsmqzCEyWnYlhG7as
IFwgXnj+ZyeFbaAUWCAN8jh4xiAGU1+S1AesMkIFRgAD6HGkDpbf7Bd3TeSB7GGQLqHtGCKf8j8D
y1PW75r6kHJP/8BUUFc28ebTuU4SS2GiHyVZ7TQCYBjvFOM7bxxrGarEoHS/S47ulgLt9eipw5IP
7f2RUQJAljxQFA5G+HQQH7Y+5+ibf5dSwatVA7O5Hd0zu/H/Qh33g+Q0vOISBKOBWhP9ZIE1ch47
LsbnavFo/G3gv1Fi8ZELMxlduZ4LgHLwzgMDhwxcj1Eh2fzV7NTdJ8R9zgOUx7R4PehI9+aDu1TI
XLIMocOqcsUCvP8UepFKEmJ9yXdTFLOUS8PkIy476tS5Gn8iJ/+UFm+fUDTGwURu9EORoMh+g1yC
NW39zpt9+zAEe/avdbXt5LJx5k8UIAVFYpLtg8BjUQJK5MoaM8cniuH3HezNX/GSfgETXdW6+aSx
Dz86Jg9hg4Onvtvu8rjT4yaAL1soSpf6yiRwc+HfmeJ/0mGNSbQl1U7EZrrX8C0K3CyI7vfRbVyh
32Er0RKsg1fmj8lFGLSQrMU37kq3UhNMm9zvyvyCnj+Sff4l/S0QpPxmPOgVWt2hptPB1v3PjGge
z7tihZrB4zWvirdClnmrobmkrtnTykfLzxilBoSyygBkSqjd3vTNdkPphkN0qvLwxSFdaCYY0Wdy
XLHVmu2tkaaNPK3K70vcNBzp/Lz7+yeDuxMm247wM75m4H/5LSQczeHshV/Gh+7kT4fTIYtcfF2D
jQLa5LalBuKjj5NVZScCp+mvaILhSY+xxjBOcmiV8sL9uOzWif7LIaBCGUxqFuodtazQNZok5sjt
HUuMxFwUlhURzYFmSLeBVXmZIAuakk9Oyc1sXvmsfXN4xn3hGeDgncrRasyt32lu7KbKWcJ6RUm9
2pfGBHxH6VYkPi3an3JtAOTRhzny54eq1fMZ5wgJq0uTEEqEJqTJjA8Gb1iVCuQIfY3H0ZA7mdmq
koCNRgyER2F6vQkw2BpnyiJlL9EfnaNDCglb81aSXEMTn5dvPBEp/S/tUIbbCwadrgcBPs4HYDn+
j+htus3+vbp/yNIrjnJSyEHFApuQNqtrRBpKPLMHVhswJxfcBigtns42857AL6zsGpW8leqEmquc
DtEapUiAItT8F7VnNvqqT0w163O9h3pt+ZXwQ4Cpe8WSnDQTC1N4ObMomY88a6YqOCiC6RT+mUpS
9h1nCL8DZyI699Y+luUrhT20L9Fgr9VSuMUpjfQi+MJ5pAXgP9iz6PfCA1WB86xeG8p9NWG03HCf
OgC8HgqIvcf9+IJHFuii5f9Qm4bOZMP9SKlOWiMC50ggE3SH1zI4OLzQZml9UzUiv1xrgN1X8bch
po2vAmcSrdaOO4POpeWLSL4Mp+J5qFUszgGpwz2Qg2hOqgtQ3paqmCHPV/m3n6gbWFFjP2jCrDoK
O7+sarP4T38R0yjKk6D7iKu8udW2owj5U7rasGmrsrc3RD3ac9VIdG7NUs03CbZ3kxjEzj9QrmUe
pVkB7fFuoRFT1vUoa0A8rpP18ehg3FjMj7q7F80gAc0fFpZUVMd97VarvnDhJyplHUDZ4lbWZkpW
w7Y+eoxd2UhgDrFDx9HoDrz9/4xUXAyl7LCZQOpdqkWu/tpLRcbSOE9oL9pcFo4+LIxKSOQuGtGZ
+Ns63otxyoVLhiOQO68+4pGZeQL2oYhESTGfE0jWTV+ZH25aPuJrdNrrGPpCtGhS3Nj9Clfi18+b
euAOZb/ZYc6p3BdHuKFqxY2psntqu/G+ypx9qmJkpiIGWfaAylNEMobN9SJ5p8Xp4+TwTWtnPcmR
IxC0UTiKSgitl2jWYosrljF9Z/YbNQE5KYNlqR7UZl7MJyanoaLgO0S1dXGr+muQlkkNMvyUP8Iv
Qqem6f35SMJNbHmFDHsDCFdgAZRzUAkXCZXzqxhSO/G82n3AVadMbA+HuD8odTk5pu9u137cdXiH
HnGwwoFcItLs/vQLbYhSloqSo7AxbqAka22Nf+jsxLeQtRNzSNNo4N5bPGvSz66jgO/Xxw8vikMO
vZ60c3XkzX63dziAMxVcJvfIDOtnoWODZKtXELZzRnRj3xYO33/mB3ZWiidA+JydL3yLg1KrlFN2
LhIIxHjlduQFeVqbhjy4wRkanp9kb6e/HKqjk37+5IIHwVZ+zybpADH5GloV/P7n8hx3/X9jTChl
oAOhX6BGJD+x05B36yDELCaNg916d+j9f+kAn4AVlbrseGEYdhDQ27T82J938bTmxbzp+QDUYXM/
TvYpsxEHU6bLUvpimrTH36jwWdibMUBUiejh2xhvSNnoBlO2b/SM+1HJ1omn5Ld6EJLBuS4w9vIa
zKNTF91q81ri5IgFT9uRGEnL0u+00qq2nMeQ7tVWcujmy2gX1kpxqmQJgOKMTiqYKGRmRl8wqTOc
Q4GkSZE4xolR3v1FFpA+ewORfgF1et1VqooFn4f9BJlC6maPh1gXgWmS5skBQjZMznjiEyjlYs70
OWe3oQgpOagnzNhy7PBZ9l16C9FQklwZjcR1cSJbqzid5XeDfdOGrSeFoaVcaQowZnX1iOKhJZEt
pSXl724+0o3EDhQDpRcMFvSnjxACwkGsCiSnkbduSXVFe8gRSohyGHssL8APa0yaP4vuDv14vsBR
v+MTbX010yVml/6votIl4m+214z1IIzMhy5YG3QtzmdQI1fSE8Wop5y0lAbC9VvRJrXGW93cIHZ/
KGljJco4lx5gBNusaBwgqlSFlKeI1UImMp1HLmd4Rud9QtgFIvR9ZhhmKAPwAEQBmXZDWC+2Bb8M
Kss5EgXzTTig0O+k+i73WIkrlbCQmSiOKOZYdrarhyYby/zVmihkKR/zGtqEtyBJHivGpdvNUXVV
iUbqmBGck4DEY62q72HMgCTf8pMEg7oHt58yT3+NCULrR5tRx13rRtPDKdlJwarO41HK9DkUDCYA
i6F1FfZlZz709eVcDnat7cgkBfAJbwY/9N8L7F2MdJvKYm8h+Q+rkzzqaGJSJnAkAzqU7Iy8dE0Q
S+GpBv9OeaPgut/gwAc3Wa4RAkpbnFK7HnUqQEmgROoy56dUPdOVfC13jrJ9VGm+0URdEHrjsa/6
YAhyXaLzik+eVLP7zSmfxc7R+H4+e7ONZkfG9McIdZ4zyRYe1U5yb4q8tKgmuMFWrwBUsAMjvuio
9yKqSJsznQ6+ncIkumTPTamN1zdt0hM155PCVqjZejg7KzADXtd+nrzinU8wFQMDKyXQX1tbllPb
Bb6oiC7U2WAEwi0uxl1pKsm6UW6wbZklrpOf7vYzivHhB7t+Ynybk7t2ug3lv2vAYLDi0AXBXLUK
PWeu0PEgc6PpTtOYoB8AwqZi3O3J8IovL6uDwbBIaDFeEP3j8jea+Ijm2YArZEohlcPiyYqaI1S6
9aCljEzf01V6V9gwtVF8hZwK+T0PiMxsj6MMF9KjKV4iaM6RLbf5gVswJJ+ajgLgr+V/MrKRVMHD
62RYmRu4de5lY0q4K6tYw9ho/BapiEijqOY55Png0FKF5fp5BycBKfzxhpCJDv6dfP83ZfEPIEtI
cfTSna+doD8Qjhvn7u4LDwimidy9jaht0T/VAFormc0ipXDAEomOwgcHJ4R9nSOdomxXHEdQB2Od
j5QdnkgobqGc9tohvNhbXA4sJfhUBrPcuLPo8tZqp5I4zhSWFoGwcTjexSVqfefGVdR4FWV5KUra
SbkK77XWokVbd543pgGQZFpQkHte+3f9zUeuM1Hp18uYJ+6aU+9D3Hxf1ojeGHZQZKAaN/76+1q0
7WPTYGzm7y9/fYa/v1F+yTWTIndfFv809t1dfsnEJ8/UWdk6dw0CA9/ozpvwI8zXXF9rx6p6nfsW
eaQejYlIhbCwYFL0KutUmzBSJ7NkliOeFr1obEm1ZebIh7Hk6YPMIBZ7Yv/WePS6r8XSt4jtc8D7
uFP9UVMW3IPYoq+cB4TCIyFr4Y2Cxw1hHVP62Z+jQfggpoZQ2THKg1J03wYs40jRAphJC8DXJRLm
V3yHOC/SomfriYI6P25B4LF71h2zmufYm9VhwLrsDHSk33yu2MYnE6zGN2zy/xqfZxgp/vQj5wQN
7/0tTfiKfBMGjLOzXBVF4SNm4Rl7qiJVH7ic9hwDDw61eevginhgihLsHayyPWjNODglPoBJ0pn6
XbMKE4v7I1FtqpGqlw8Cq0YPyQMhvwkkoxaE3/VMCphU6Tqckj6MWWRWhfjYhlMyU7X4uh+JS4An
zvZyRBZ5uthQzFW8YCgx17CW0PnRNa+8fmJHlSHiNkLq6ynlsbKrbUcs/KrfFHL2uZhpxPzG0aQK
mBizNhcne326lSnuSd1EY2U2zhEmQvGKQJC/bxmvDgeBKpWEnbjwcQIqXgbMxc7vGgBDbOPLfYVz
V0JfqiXgLyfvrJ1Zvz87lwcvqWnblFh19m2Vzd4S22EUYLNLq+NLDHf4SBSAmKDiE37GrlE9soh0
qAaFp0D2EZgPqhrUd4nRxdsl6x91XfZUEvVgRaZpXc73kGhpZXPG7cw+SRP/K4QCoYw8B7Oa+0SK
qTmv/bcjhuLv6OCsDO8Mvr3LZcAY9kFMWVg/B0lVDLR3sO5pyGCsvea0b1yg0qhG8C0XrIyCw8/a
JKA3+1b6iWJDXrInGci/+oI1Ng0WVaa1jNC5GGd/TUKOLRtI9sNCtIQI0gGo9UWXC+eDmb5VVi5z
DS1nekwNrEbfCFO5pODPZioKQseUYS0r/8NHeehAo+wJPSRd5sc04gSoxIslNLSo2JJWjoKygxKe
FTLxMBX3OMgBkCt/eZkNacZVH4p2NhAVh9IDXsmV5Yyf/0dyguuk5RaWvxeztF4JKTtLuu2nDhtS
CTMBwdoQI97IuSDCFhXriD3XAGyYM3yvmb3c2egX3eKOMtNas+YVwsA2U8pMq62T4lSyM7VvuV4b
9V7LNWdR/7E2Ge7r4//HEQNbqXfAdv2eBuRa801SD4LNBfmEvN1YToIFAu03cl2SaIgE9Mhiqxc+
apHh2xNHKH3HWtC0BQynyzv6o/yuTcEfU8vrSTBRHnVBvqRnchpuDPNEVUcRInQVuREuWxwidVxG
9uLk5K/g1yjq2WMfxq9JfyCyqsvqCBYNppwgkp9MJk4k+pxs+8JuzSm56qc0lFGsz81yDF1Acayi
y28JgVyDrl63VhQfEJ5C6+yaUlwGibIwu/zzY5BneluEUKrV/BR9NWIkfDcNSYgSxPy/crzTZRku
bGKO33vdhYW2TQDhxBE9w7qVruGw62xgiZswxUC+DAsXvI/L5QCrhE6fSTY/miga+CKx8APk/oxz
eDA7x5EjIG+WcBFMS2RnW8ngoerhybQrwb0VewwyFna+gLm3lu/6SndqMh3bRl3WoEiemYHCRZsj
YFt4nJD04diS9PKxCDqDJvZIcBQ3+yly/GzNzaxoS/8XqoEMUov98SplvVEBUq+Bds8h/5YQsdJh
aZapfw91nt9W5TKBl2dTvPB72LxrrXIvkD5XCORVKAUQx1Kg8kfjVBaQeO9hrJQmSTn6jsFjon2c
jvkCEbaedoJaCfKDbsAa3I6eFXt3W5V+Xopo5LEY8Yr1ivwiWqBlwu0hQJiTtFlV8uTk8gTSFLLH
ZVeThlcCXh92N5OqihtbjD4kEybEtEouiVCgOsZvShd4962RC51NnkFS8PEiAUuVSyPP7rTfmPEE
O7utQuUJ/SfmNygSRfSIZ6gbjlh1Q30OtvcCSMbYnMP0bNA1jwpFP6SwZ1VEURnNzjG4knwcBBqJ
7oelXOsXWz+GWeW+JtrHjLnTULDsLJexHGgHen6+7crY/tutf5AyTb3kfTTaY/ANy1k4eoSHVorf
KIcrvE8d3BCurnFPP1JqDUUTbIni3EyHgqESFyhEQQx9rkWyEKwOKkRxsUTKd0azuM8SO/kZDlBZ
RShPWVKxUCs1LOa5Lao12NYK2QtgkyxJJUZgPh5TSd7YfnNPkx/HGJ+EB35+bIEfdJBDfvWdHxCs
sZtkcirp7pFbUdLjlNDm8vxZKQKi/3Sij3Nrc+kysnkqscTzcCZeuJaKIHNCgN6jydamxIwis5/B
0lliGiFaUkidAcr6hkZEnf0VjBD9BOPfWpERGlUDY6xKlJGa41Bl5gwFZWL9CP5UjOILVC/f/Vbe
j0CFomEutIIZ3YWhz3vTW3jUL71OMit+CpYEUUd5UeDcLtr2WZDUeaiuGOalgcELPMJGzZ0z50wi
NXH1jJci4E0xykzVugrz+zCHyQ9A0IJpQ5u8TLsccDPc0C6c2QJ+SPHgC8eWmYmzL3NXI2KZU7xK
VjvbqDIISTx1xDAdYEJwrDb2nflJDnJmXZKa7yd9vVZT29u8MOKRUnCNe/DFbYOfHb9L8XTzt3uA
kMl2q9KcYmEzLv4Vf4GoOl3VSjosRXdFxH7wBmcRd9GIpA4wf8+YlbHLOC2A4KcWR+pCfkc9jpdm
KLIBrGBSJGz931zicMxvb0x9MJclXv8fzCuwld66xmAoVr9hR6oJ+Pm1P7Nr3wolR2O5qQmCcRmf
QbUm+3HTaw2CIj5c00dwU7LYunkNNkbYLDvvNMr61Vd8/nNFhr0DqDcJpsl06YN1/Y+ewmcPQldg
IGTr3gFHbL/riSGqCyD9+8ZnWG3Ua9+AFKtLn/HXVwEgffcKc5rL0iYo+GngqyXIJcpcI7a/v1/r
Ft63ymCyfXycofZHv30Je3nUb3fpdOWiCYgDDInadLShJEatRkbv818t+QTQEgxIQoGBliH4xxdQ
L0UQkotHmFbqtWB5zPozv0plGnfvP3CSEnkOO1QPgScCiY3xaB3y7rbmAmiD/YS3kPb+VN+SqbNG
K193Fzzk6p4znKCYrJd1JQ1lOArrDW6HvMQDt/AFZdzYaOQTylgyDemcQ2IYuA/qkKeESTyXmjFe
HDhK3BkFkv0NS13355TkWzHAL42u4oLk4bIfaiotV4ZNOm6KBS2H3GKys7nkPhaBpRT4XX/+5mDR
nOsuW5GpEOdw6QRLMU8fY6w768Egrd+XGg9uLo3PI/d7JHyPwX98sSZK5Ky5nQfi68Dh/Pf/1V+O
rQnqZBKqQnhjKTSD5d3uCK74XFSGFsMNRj7yEFkL5SAJS6+7RPeyxM7bNgwICA9acDtPVeRvQJKH
rRsgh3JCg8og7Cnv9MwfI9X/A42C8eiEuIKW6K9N4DmZli6H2y2lu7pMNtH/iJsHFK1AGIyxajwQ
vdufs0Et3BOt+ZAZ4aY5RSf7i+TuBkRs7MixbYl7xMEqbC9T/aR96zi8vS58i0cUm1GlnWaXL6K7
fEU2iQlawjnX9yHPU9GB0BiXxvieUt+wGW+a+qxvbSAhwpQ9egzZy/yeq4v2xBbhlYX7fBcuB7bo
XSpdO820GqU6oORRW3Yhg8hRT+rh1OibrrYnZWD6YWXrlfforAQRSZbNEzKh4ymu97eq31LO0ANU
b/1qNu9FJu9fmBuvdGQiPnwSwIHQPDBMw1HVYM2P8UI7i9f/rgB3BrJHfFlfpkb/ZJ2RC/CdAPO1
m5rAgoLKkMZndbkBpjcamYEemlI0r9X2nG/aFM8ACybIVMj5b8rhmI7KQs9cFbrCkMeq0G/xO6MA
HAha4fJSElVJY59Kstpf4vUDsvB4qkEu0aEprrssYEG5ab34AFXivDUfsZjwvSDOjUbFwThmlKwz
CBLaKJzZR04mEHeeeh1xCURFmw6JMplLab6jEDu0dxm3cl7YmyIB85gm2IDb7ydi7jx/7xQuyEFO
GrUHNZhy7s1rbaBj/rqConk7t6dEGI8jbIORFdMefui3VDxtFuHsm+BoE9Om463GNHd/6pq2S8oL
UN7fCLRxFyzVne1i0/gSTpPDA1TgJydwJe3dEhw4lD8h4jcSNrIfjT2NsEyag3oXyfpx7rz21xMW
6Cne/jZiX+RFjrwWGLnDIKbEAy0xfZEPkPCvuF8lUX79dDHKbflRut2hCVuNwg08+c5RbqDmBe4e
xVHKBhxO1RMYNJft2wcmgKmoKZtVY8xn44FIL8mpgy3lSTGRA8IyAQc/0fkdzrbiPo6e+fuwli+6
B5TalbGluzAHKeTJLH0q1VEeQZyCvq0OcVxqImefa7FGiNx1arKvK2h83GYdmdW8qZPqg4WuEfcq
Mchx8l0TO6G/kW85x2JX28ax5KO+kTUpM+75BeAQE0DUN97U/qrXh60mpywrEYN5uACDAhkNBV17
9+fh6RzyWUgOLMEXuuCZvnmqRAw3jETPG9ZhvqF8Z/JQQLLhODZMj6p5yxLXhvel7vb+3/MWCRLa
BsTRJtWdjb/J8bO/s+IABkcLaTolIuIVXcdQh05Mq6b508bayNNlQ2JA3ATojH02TWqFyp62h0Hm
y1COO5oD/OLJOrTK47ZyS5eP8uRZgaxqzMYg8UOl8b0GlTFUTgdgEEK+jY5CB0ANgXlQD1iwv38l
zEfbzAu+Ct6tQQbGzElgSVFMf8X8wX3H67DLpK3W3yz72c0rUTNJmPgm4iSLjkaagguJObTr6w07
9WL4uqxqe4UwWHZqVcWqG9eVJcg/GHzig0t48naqAc0wvhAapEpsudbJ+F93HoxWvVPwQTvp789c
zIfQkzqAHMi5QhUFqwg3528e8ebJf52+24kWFkaxncN80JFWrjXh1n7FkUGzJtxfEChf+C6eFk54
gygEcDdpZjbpNyR5nqsSzBHL30w9OFWBVDKlVc8PtvNydFxHBLb4R6oixEPy27KEC3S9UY6q1YLB
lL/Qdyb2fuvf5SMwUQ92GCYRSEUPWjVP0rgzaVFKYKyarXtRNvWpQZ9nd+NDLqzoJmGdGdVOIY9M
0sCGleDESN3C4Svcx27WRwMtcRTACXxiGVh0sXWtgIrA3bcFBkrvc1yhfNVDAF16y7QvnUsAEVb9
bbxPopo27/ECA71qU6gXEbjUHLL7yectyXpRGj5oD/wFDUZzar9gchGNanquoTcGx8FNFpQZ0VzY
GrAWHvXYHwQGTKdyLiqiHdOMSu2Zyidv5FEQdVBQia7x+WAKvcaFKsUu9iedksSPO8C9LQi+WoQL
w6HdtsgNr/oxmDbAY8u3V27P7DBNWp1rPeSR5XvX3L1SIfCyXVJok8zMQTA4tp1nEGhnRluHJ6Hu
ZWTwVm83bmYDi09vbO8PNzi4JHLmAMCpL1VBwO2vnsbYQhukLL9Cwup8ze/tpi+LaGPc2Z0V1fYu
pYXlieLQRIh06X4jzgPk6B8Uvy3PPdaBQpg5oNG+uc2537rfv/b86fAlQ9vqPLnNhlL7TrRCV9O3
Vy/7ngtvxzM8s6hxPDinXPN/d2rhgbwxXUR6Xfa9UW0yXh6RKI1KbGYhKmfPwExTKWT6SablKc6J
Sle89///F1ZQrJNYBT8tHfJbsbPEAL4luEejSaGSGJFt0o2ZCjdQebnkPqiNlIHO+6eIpDGmextD
I/bXyoaigLiSFNCr6qruW1Q+RvLtJ0fVktpB2kuOVmb+0KMupeRbydDjjb0n75YJn96zWsxocX+S
kRCPUnm+9RAod6Xc6QTwFXBfzajQhOVgGvbn5Lj31TczUxqxmqpLjtbQS9NloorARYqxlYtKx6iZ
70WKKIkDgmdZ6U5i+5yDrmfhC0jnaoVKaw1eHUbVLkx11TenkyDzSneHpgtVvaTXoOebReH2LGmJ
dkIy/rcODuYv7j3yGTc9PxGrPIlA+403qL1Z7uFCHyKKZnVVDHHGKdRhVBpm+prVpQAICHSd9vyl
k8z8Kn/TuO4kC4EYsdublRhX/AXYzQ0D9eeIGH3s62SJOLeqxxaxgecZQlb0tGnaUUoBaxYrj5Jk
Sc3S+S8aGtwLkSmy1xdjtJsbHJ30ZgGPCDwct5nt9LECj1wZLvKypnTtVi6JI7vJcdxn0E3QUWGh
Nc9dbugZtT2MT5lEVCxDNd5PnhkabJ3T1oBRoMo6xu5l7Y7rm5LZLhLJYGYCG0enWB6CHgiZHq/I
j3otAupI1MY0QHu2mcCX2ecyKRE+MiD7ZZmbp31CHmiMq4fA0v24Afm2+jr5YXY4ZYhY9w0ziBI4
vsCZYf3e8LCCdaBFuFS4RCkYaBMbenrA5ma25+iRrjmP/NQlEeT2zYB9K3Bdca4MZ5HAY6+jKRhD
D/ti8xHj1g9YMhOpiB5OnfEG9v03Iztc6a7MuQs1UJOXZUL+/kwUfOor/QiK1ZVNr8N8iOXrSGyr
wtDVjEg6aDVekLCO4EJWkpyIGxpjjCusec1t8E0Lz0wD2S2NJCMa9L9Qet2BYsThesgtRqxdw2QC
KN73QcTF+x0GJksemP55KNr2t2VGI5fIu+MMQ8R9otkQykGMA93CFPFWYk3wFOO+gahkJoXy7smZ
dyAToGGU8yvfNMlw0VZ5yBXZaJqlhyFNJYf4lrjOV4fOFTuH1YVpQPq64ynjdFJ86oFTrv+W8c/k
OnN9xUGCK4d/yAUQ7w7YIBnGPii42IjdOvIMC5G7/3ZH6bEM7m7ud460UpAXTKBPaw2O3ehsJ9Ek
dY7CGcguX93ErIJ6G72CejMRl3Cz6jb9UaNEetDCtWHU4iitg4cJ5Qc8jVzhGPaATFR5HsYqpJsc
Ujpgkd7eKw/8jEa+RMvQyCQf+cWXIxEJdmvn6kfjpDWqql8ukGQw5e5mkCOQX/4TCQF93wtGrdxL
vMlpigqMZeDpW4gtqAYG8dP8M5aQ3ZaMbeALtPzTSstY2nPRmNYC1kK+TRcPcmJu8s6TkkXILolC
S5No56w/WmcXvrQy16z9i/LrZnyGQ99DGG1VQ0QM3GXUntSJTa9yAgx4MEclAL6HZAlJ33qqxA5t
qoxMG6P8y6F36yx2zbOQUSjpEfaDRC59b80ibAP7DBs+WHjieC1B2wfBO8+3ubwHPfus9+1QH5pn
RtwP3G/qXf13kpx8CE80BY2/71cGfEoMv0+9F5gxs7LirLeyN+SUMR4ZGKtywL87AvgunSYAaVeC
d+dwRDJ9rRCw9DrrPeugaBD68uT3fzcM/YUXCeNCX+0eV4HTYWw5OyVd46YF3onjWxohscLDA1mD
IvqBspfpRgjScRorxkxnfT1uc4HjbQIHi9dIXjfmyREzLzJqdYMK4d+0DWCIbFn9EQr7DFxX7PzU
ePpik92eyv2lgih1Sn5fv6HQvlbCvsja0MyHjicfMm57NMJ/2UrxmNb1VrkbuYLMdTbZFRHao3VO
nHJTVLPjxnEx3LGfPJAvklP3NEiyEW5L7LxsqYK95emwfrX1A3DDBWLMBjBCz1IwqGoGQq4n3c85
Vu/T2NF+uBp5qQ+k/kGA8spnzFT54JHGuBaIgxT6AXpJiIQl/ruWY2A31xajudqEiOxN46Y5fk4V
Aix8LuIaxRvbmwpInPxjSve467jGp4xG4lVlACt/zH2hoDBFA+faRB1Wozma2Ize3IpJoiQTUhX0
x8ZPLYzQJNj1/Fqa0qgua+eMF9s2vNvufYm2rEDFbGU0H8I9x5qnMiBWA6ewDrNw7bzUNWmbwO1M
h64/JMr1DMnI8tZ8q2tEMqr1wslT4cqmOAxd69xvj6kdoL+P6jl5orQppIznExfjkBgNGCJF2KUw
xLc1vqskabyQtXy+EP5VQCQur2HAwrE8FqBXZGll6Cx2dk0LTUzsu/JcM+wuHGvHMrEL6+zJNfRi
zBQ9VjfD2u6Qw490WwTspyax5Y1ov92rniHvhs3M5vzlCpExu4NE2DhTmzD3oav9axg2JWdXfw91
uRUw/wczxN5mHMQNlpBgyzwbROHyyvMSYoBCIeRc4tnK4j6GOLfdGV2hhdOn1HmCWONCINmQbpCJ
TvCN3S2nBPXfVSl42sUYXs9+Z1WKBgsAwY3ZeQ5aELvSQ+ilWEptYoytU2dYsxoAyvWmFrnQ1IsO
yDBnGgJhDp5tpMk8gwHyCWzNxI6THpYADj38PL1hzL9qJcuT4uAdl/plTp3cI1zwo9eGajyHvQ0U
V7qX9BxaPgBpqm2l3OslMXbbAGiDVV0fnav/Xdbh+Pfy641qs9x45PmPyCjNo7E/oO3TSFxc9IC3
OKJjaZzKbjBGhRoMcBbBLme1eFawcu7Oc6hso2nZfc+Du5sP6CwezyaYYWnxRE2QHL3G8t26mB89
HMh3Lvxzi7Grb952M5xQfl2q1fH2ch6A2S08ysa24WaWDidLfKEdmwkfZgg/HG++eLdzIjqnjeU7
slMaRql4WtvyYjG35hEvoDfheW7aeJe+dXgEa1V/0WV6xxpqhW51RErYbOM8WtZOB1XH3bM72FLD
Wd6dOlZznIe81n1/w+nBhpH/Aw6oENU1npf40kV0k8bB5Ttueh7346ttG8X9Bq6BGb6Mxbh6dmWb
7hopNdfETcDK9v02qLjj5ME2kzebvJZJM4LA5t5F5FFjeTHnf/DY6Yrmu1GrQPpo/l/bKQEFGiXo
sa7Ez8s1JmeibVOJCpH4Cjvk7Ogq6DAbQqUj8U+6OSMooLmmD/RhcU5JAZowWuEvLVxYCk8g7DM/
AcwuSWGZUUubJRYaPHoFEh6DKZSBlcmWTE2dk5l4caC91g4FX1RdBpHRpORIkan/NEK+JNyOXsec
mJ6RrYTVEEjnGAg07oVKRIKdJo0GEYa0mIdzctDMgBL3O89NGcZ0sj5u4dvZy/0Gqj/oDaiEc/kQ
iOfA5o5rKI7vT6NwQn07x7Uix4T00vY4ODmkOrH72tbACP1CRjkwy1iIIugH6KPQsF68h/CXbCjU
TBExeRde4Ay8bZ1lfHBncrExQiI1H+bl8hcmUoPZ1oH35DWVt5d2sRnx0/U+x8IRGhzYX9ith1pu
ytTxaLByPw1Jg092rJsHxnyF4Ap0O4P8K4AUj52KKMz+OJc4u5yc7S3zDDLqndCf/mDaZ9EzICkR
1dsisN2glGVauchKQu4vXHJyGhvYX18CS22ugNAtmRmV9tn7wX3IlteITSXV7MEZl4yGkKcowLd0
5sT0uDjDl1QQMkHWWJIUDkflWNIfhJsPQimYCaV9cNCG3xDA/vXP8xSqmdMVTj5EPZ3deN45L4JA
wQQFKEb3iTSXnj8+F7k7WVyzvXVLPjc8ABBntvFphRTNHteW/LCtffex7JoRnXrRVcojguZuFzdV
wQ2vuIDqpWy/msz5/LPSbXFglVOQ083YTuIyPJLubYD9MmHKPnsHDXQxqh0CZDQTAmvpZA0jE6ew
vctQQBcf71etRPE5iG/UMNMc3XaFg4q17+qYH611IbzWZAl4HauLqCFb80UtUtLaElfl3LRhWd/o
La1I/7vJrA60Sk8AJUsCoRCayPK+Y5jfGLzOqUJ6unmCwJIZbGvt2yOTsZd8Oy/2BvcFdt2JiHFj
LVZoyxY17BjK5Ot0h5Uq4xzZGKi39kv10cRdv5FgzuA5y81xDBInL7iDFv7FxEciawY3NjlSj3+Q
+AVKo3Dod8zMSPoXJZx7OAxhK5NI48zpxWJ/r0sYawCKOfm7djJJjycfiF86yCV7yEPbzThFoAX0
4BS5HUO9Ieh+DgFE6p9TMEwZ5jYTZlw2DgVHUU5H3CPOq1XaGUpG5qAwLZXlXm/eNLNbTNkGel0e
TyfDFYc//tH4Wg2O+x95yFLXkm9U6UuFI2YC1TU+kp2aLIeLJxYtXbw4KsouvS5LjFPwlYMPywcQ
MQ+iZjd/3lP2m0QTOE1XQHQwVi77jV/0mq0/FF+yvWnTQUEX6pRyZ059cZ/t8d472Ct71Nti7w8r
ZTzte9MX/M8WE5w5lLce7oNHFyg62uPq83iD1d4Sz/uhhxfTdNOhNo4Z9/kDPiCTTFi1bzyCHhZd
qiwCi8AXlZFt17QRkd6bkdFjOzaWEHW+5dVmmGz5Lhj9QVc6NMZqrMn5TXVUHh2ScermBMRz9vHU
6Rxac5R3M8UBZGAlhcwvOgQYGKTB01I5YwCjLIIHLFFNWrDeXlWOhjjQN0Mb6WHs7DLWMT8F9/Kd
nT32a+F+ceZgXOAHZUWaszdzIArCzDaQU6Zv/OF0x+J2sS76THWs0KzRZhqazf6+tJJFBftP6C24
z1YymiNKe/DhkTyJQl8ivcYsvOhPNLy+xqCp8sAtGtmMcKPZLHtOHEampIjQLvfHzzRvDJ1fjS1g
mN2kdWgWuK0uf9tG7NVLqrbT1WSSQwF4lDtBfdeyV1Is+rI9Ee22Z+JGCBJIo0vbs+vpX8P1ifXt
Vp/pdsFJJJxVp23OPDoN3NYoVkkXiYnyu4SQOlTpq6OC1cT/Hg58u9W6SYEY4Vz1t3MZQByoDIBl
lQQgQcPftwp0N4ouw8MM1CHI+vyMqMeoOJK4k59YSXYhK7tjxM44Hr9oAIpDZNarOiubGHcOAFks
/Pm2e/XhW1qsF/tO2p6f360A7CJqJ/t1GEIpj1Ev2y0LHsPOVtOfCP3YhWB/nd9/X9fswomqJqi7
NqyyeoIl+433dcJX8P5rblyJhpvi110f2l0GnA6/zRXPXPX9kPjHzXtnkSfoQ2atbGE7maq2qr77
PCDu/VC/Sj/jawBWUObAIig56uKntUV08cuWSsFJe+Q8FX6NmGX8ImKHgf1pf832ivQhRH6MxUWT
lq6Mxt6Uma1dxO0jgMXuiTs8n+eo33XItTEy17CXUFhxn7DKzyoYqXUS4+dY9HYOkhIZgMUk5okF
B9FrV2Z6uGmCwkNky+d16AZSyEVILY0tBbePbAZzLz+iGMCOWOoTqxqwZmCNayG4EzKx1A9+Mdlt
S6lzFxW6/onV7ti4uApEcKlQXV7d7zg6Vj4SzpFe0HxNLjHm5sOyCcSGzYeOsntL1H5pRvzAVDZP
XNkxj/ydhE+eILxA9mkTaAQqKjFcZsJFCh6yz9nDCrHxQgaZxpNsv3DpSQdpmXHfQBdaKURoZy+A
HDkYQRAnnozcO4I6c10RpDlYqckTv51n/ovvLhyBBVwBMpz/rBx5CAApGClBikvV7A75Mpq5P+gi
y11LKw872TTe59aCkv3k/grGfAet//w0+PuRxivUFky+iDwL/NteSZ+ih075xoowHBOFlrOot253
GUSAhHh+lOAhJtCIY9rA4Swk/oMr+KcRoRKKJDebZycblNFP84r+AMG6KreMny7lxapG4k5ifLn6
YYHQA6Gpx9Li5pBPGPPXkl3BVQCCzMpdHfbtvgcEZacNQ6gnSzgyMiU2HRWXEo5XWCi3Wl4FBeVA
NoUdBBBSxWU5WL//7bqvanX9sKqaZaRvqFpACMJDHJpY/+KWUQ1I9gDHtd2eUf+VaX9KaxgEf1sE
/EkpcQhybUq6M+v66BnoXmzYrlOq9aPh+gj7R4Acwtj12Zj9yBFZ3/IWwBC8Rad2pHkhfC2nij/I
IIQYxhGHVbQpajG/KsRVvTmYRoZnR/ytnXrF5jMMi6vXlZWfq3BAUYpCGmKDPxWumgM2r/QhzNyh
Y/1DRIRQY7KIsASDz2nbA5j+HxYpv1I64FQtvD9xpLWRCpHBDO49j5ySRkN6IWg+royBZMN4Weu3
5ElrCv+3YIsi7CdZ9AJ9tooskOcoOzPMaWotqRd0BkkEhEVkUvQk1QxQ1toChzN8NkCin08jqEsp
vX6rOA7ljTm5Wv0nKs9EDU2QgChIG5k1PaOsCUUqHCTyZ9IHkLSaSyAXCNIwejafhn1CpcgckxSq
VTTTdNiX44bcuk0422mHFJi1AoeCB/GVbNS8Jbfl+VQdI5iQC3H9W8FMoLbpvRRlU7xS9P45aFFm
5p9k8OQH0JB8gwxOyimS4aHWZuYNsIbuz5gwzWJfxrOgnmOTiWtJwrBG/P+Y7XhVR7D0Fazvn3YA
+LyIywcSdLE7jho4T2gjuEQAdbw6v9N8UHCUq0Lbd4IM7EHiCuKvn9HFcy2mRza4srTqQz16F71F
ca8XNlqn1UN/ys1UaxpNwB3Rm4LgExvO9/vX7glMWQYJNn9ZfLj40N+uqta9KKKgHbdoqjudknCz
KJ3oT+2MCKbXoEhM6w7e6O7RszXfBGJsCzFjrAPnRPuSQBFn2E//Y9Rq2uoy4iHeWNza+qSTavQ7
wQn8a+5UPcJdo2nEbY3rKHnFO13ccqDNo4+x2fcTDDKHOC4rn+WPCoObQSvZlo9x7FwrVON97V6p
C3s6gg86IiWmvk6MRxRk5wxkE+TIgQE5+Swx6iVSTjx/WjO5vDT2lnHab4Lq6z3PlVbZVFAoWIms
zZ+UcKJX/HJotZm725Tf2/lulpfOZcJfO55/V8XluDs3HUReE9cXz7MYZ5qT22vG2O7qDpxia3TO
KWAd8xLdjp4jjpnIDVA0EhEBfeuKXWVgKLoIjj/G54rvwB+bmJTrm9pNdnrffR18WiXIEEGCq3Pq
y8x6BkAktp9c23qenfolJSPXD9VBo2v/jDlMdUl8kpRl5y97orunzLdjDm8lBIhSHd5BYpA0m+V1
IAEdRQQY3iFAe2QHLHRrYs4mSsNR9TTx1tvC3G9u5dU1tyh/c0AuOEFjB+rss4fI6o6aE+dWmeA+
KvKaFlSxybBIH8hX+fi4ytdK71B2vCvEU4FgvjP/JdA1dheAjue7ea4nh7F5gmHhVBagCh118pUG
r0TzIZRYZBQt5Sfou3hQoElbYQrCkldkoL93ERU/GC4MdU8wuDyk8dIZZCSin7TN3IQHufxMb7pS
3zEpAyZQ/+1DdK4Dw5XhIOf3c2pNDA4dzSSZNr2clPlLU3QXZbsmH59zq2lLt6dtXjooJ8WvAvls
tPST6IKEvyNNDp0m9OWbr1MBsyhQe7/bUKhp1A7eUxCmFnFDx6wO3NFObFy0Ebsy36oBD4d9ga9X
YZ43xVq+GRn9Zz1dcltmEoWesDvbkHWWR3x6BqO9015QNGUwYH303JoPbILs74lQp5FTi70oTd9E
dQhX7958QRS4s2bW0mH6bUVQx8imT+/BQ7adZN2jdI3MYf6Atl7InP7aheffCLNz/GxYTn5I0Xy7
QjB+4PSs5B4yVsMMyjhNKlzPRbl/nuK26CnTfUHANKTJeI8v9DAvJZjNHsoV5YF/Pd06a7W1L8T+
Qam5c6JW3SNbQZceo9DnvZswoVKUR+xhOxT8Z+sOfTZf2l8P6zPM12iIQhOADGKVGxBLgaKqRigg
qrcuetsIddsLzILXGHI/wuqTuEAqN9igJWRBCvmK+KcSxM7u0RJTGGBiR/z2U0F5vmraiMst3N+f
9YKC4tyEi6zvE5Thc+TDU2uW1dge3afyNhBLTGpy6PU0uQ+IWX99Bt8UaIu2Qy1Q+XtxCSXiYELY
qmJPo4xznr5Mgikr3SIEJjRv3YqTy0vN8gSRQHFCQv9qC7ZW+02VelWd+PUb+q9L2mv314yocf0V
vYmdsvRf7UY1jEKHoNfaRyKsRYL54OwlCyVfuVrxzhtx4gVu4/h040L6/geXIRUvhSoTRokZI439
SQE1rO3Tr4FV75yPyAddSc+JritEDRKOIjo1vAv/T7lWlSEGjGw44W8XUqYBC5wvbzPWMAj8lBch
242p9INuZtUNTlNYIC7jeAP/oEV/NF5PSxqeyy4dQaV708vN7z0ZawWmrDlGgDZldGTjzpyye69D
XZoi+vRv/uao1zZlojOfo7IpBSCVV1HdLtDCRXBl8UDmwZr9/cjCKooimWmqFkO4e4ivKaSYsanc
VZQOOy+OxUhHgkMDckDZ7cS0UdXxJL1BQRIvwC1jO6VZt6StH2ZRMHKS+kPy+F4SYubzAn7dB60w
iz1Gqr8fwX13yXSQmWlWbh53dY+CcAjryq86y4tM7s/EBSoCTrs8Luf7qQ3pDHdk/VWsnPQPD3Wy
HP6NJqSFtZrhDz3rr/Ti3qVxnTKjKHZ6Q7FuhyK8WMUrCXwdSKSJt3/KlcrajOlFWJRVanrp92Lx
zCs6+ACVia91L2Fox9Oe0xCiFiAryLZQzchcmZX38AEYIH5Hsllx6WsqjpJBNSK3mXPwnNhJHFU8
sInlNwyVLJF8GgXF0hEOBnL+pQbzC7AWW9QFsToeV9fAaPzXX3tfXcWwFqty95CbrzN57nGaLWF0
Z3jWpQsk1T/yft0BlDp99GU9lU0CsOI+tGoDW2JSjekW4A6HybrMQph+JIn6QpEFsoIZe6aMCp2z
pt4fsr2MMWYFCWsa34lA8CItdnG6/shtiouzTR7jbvkrdkVK5PxMVUVBpOk0mFfSVEGak1F5qPUC
iF6RUVwz81empVrK2spS5KH95KllSEqiIgYI9CxjpVZYxYh8UsleKJ5iAsbZlj/+HHXDauWE82iL
PbioYGwEj5UbWhBBb9ro+TUX2Znz/ncH+rW4T6ZdmCqMp+XFOxOofIe4TdavJXr3r9AJOu2HvBBH
U2f2bTCA7weN2FVS+FMuNs5U7IU6Q+WJ78k+2TPEhlAbJnv9gP1n2ZmnN0NQt+CUEhU0M8bbe8Db
RwAl8PqfGwmkjt03O0sZK/T3JEZkGJa6RIbzHQUqBej/VaB8K0fchWrG2nx2GapceA7/zwqhA13g
+J8bv1EJWEfY/jlRLytA9YBYptVGX0kirBBpha78qpYhn9D7yFOrglhC+z9jTV6BFX6v71rsUgq9
jLzjLeVdpa5fIbnFKy9CjbXp04EZPT1ESO2qROAFTGx/K75g9X2lmqz/EWRB7vuHOp9Mg4ufQ/7s
tX6tshrHis/KVDrUS0zJ+arNTvd77PsBLBU9+dNsFxyfh2q5DTB6aGN6EdaAMHA6T32Hp9mRVQei
Foo6iDEspT34bbFCLFbcOSqSbjB5FcCynhLm4EosHYt0eOiTqUH/87LCTsQfUJO+IhzbAnLFWFSq
iYXsgBNjd+UbZi/hEtO2f7tpFB1lnzLKgEW+jDkHa5n6DETOWnlE8vyuHahoYzWF29NKcj67oJaV
YeJgG8I4iyDIe80NbZjH7D3gMp1B2y8WjzskQTqMRQcaEh/FXbf9JQwdGlHev67fdx0tTlSsyEeC
114VupCXQgr94alWQeCayMA59mq0FTSgLVF4VG5AFx1LJ5j+roS2plmIwsompQotJJAep6Iaau83
Z5JPZrOSIE6rXqVIfaiLFtbMWRwzlBpq5WWPRTBveYEOy1oQZyygHfrJ/qX8jiKIIIekaf5M7jz7
HzjZoANMOFg2KaLEHV85ZDPm9tLXq4spcN0W7wj5qVYVwtMsMHmkTKY7WkRXMMlLRfClEyhJSA1r
oe/ZS06ztnHpglj1M1ZAAhTVIE5waN5xQ/yR3G98AS62gRSz4c5pUbt/SrUMdH/KqHMG84HrOn0F
4/lyRiphI9G7FqDar+0UdfXnD5etDnsp0DsCBNPSQ1glki0Zu7tp1gZs1lgqhOUkfKjJqG0kEESl
UkAZK/yg3HohBCtodrjgADYqqPXt1DmNIVEqjeYOUeBixqxiWNclVdxEbc82berSJwJy+ToC5rnE
oq5sOVcZzXVCSFExI76Jgs4M6z34mvvFuTPM4MHOJCQYukw3jYFtwEVa77iH+7z3iSdXgcPtOUGz
GwNFXWyl22prlyu/UopIO8YWFik1+F3zpjX2PFkaJSbwh01sP3nLFBvPVhOuAbXh3rg6za9dL/u7
p2tz+2pkUlPlFROqDKHb+QbS01h+3Jd2tnqcQ9qMhYn2AcWc+nvnNt6YW4s4pQmuFm26/CLXssjK
YJQJ2n5DesDXfqMv6Dp2iFi/VYv6G+sY6dkM5da5Nj1F1F1gv4+KRrCEJNlYgn3HNzEogwlWdaO3
TanQzERciG6UiWSqLK3ptr+mYU/95GZM7QqAsxfmE3vn21T6KYw/7rtabiEUsVPROUxUlMvI3eWy
pWCKDSIkcaZ0RtsGOxqE/91DUC+nAZNTkoYxyI5GfE5MfDWcBqSF4hLcxA/MdyfovAqHk45Oas2g
JHrvMXDMm/unrC6LdFGGUClViLoqHeaEDwJvNzafWicvFluFbOTMpwbcDMfAN8iBgF7irP3TDuqo
649vvPp5FaMoMgaUFb/soReSXwZa2tMVXH1zd3sUi1I7b0/lyk0noFCFlrw6Y2KmZvlppgNxZH7X
L4k+8fw2Rq3l1olSnqFNy7bqrtBXuunRbShduqJR7jWbMd7ClzLUuxFOjH4RDXdTegKtuR/OhNvn
IGA9MpPVdDFu9T8kzkyTfrnASA1vDeEk7DgJEKIsSUx9Fd4MZelpcH6lQ8tv2RsyUmJKP1dWgh5F
cqc/27zQBBa+cQ+KX3OXFZ69D9M+ddJ3gm+RyroJPLmUKaZ2KN2AdACLQLvQhcHdlzTDoebby8Qp
7mdLNwfWyP/UJkvkov/L+EcAYZ6FxACfCn835T9rHKaNPpbM1i8vDaedbMXHw3Vv94Z+Spu8gUAL
2z/Vt1e5Ns9yGEJv2M/0DYeT5xDrPddAznKAO/JvRsJ/8Ua5s8dyO9txpQs+tQSghEhntZ19Imz5
fOXDYeJes9US35wrnRc0MMx2gxIdxOH6oqUt8N1KEEciasVqnTomvPKnesdbPLqwdrjwIxLhdEf2
YPFTqTUBxVZmkAPlVceiU1Ew17ajPDDMo7eyXn/NmPvx4YXg4dbq4FFIEQPsfogWnbBI2yisxU4W
7sXbgz7Hl1Jp9qEMBWkTIrP/C45rA11fzVfB2+CQvHlXWM9IvMVfrFHpazneBl8DDk4oEu2lr1HY
CXFOs9zlMsN04Wb8jCGyVQTyGPsF48KLeGGyncMTxH+kvr1VH9Z/sjd1hMbGnoBE4rJJLtK3o5+U
AF9BvIIg7w7qGFPxkMSsRrjg3ZAA5KScat66WYxo8t8082Y1Kpp4oCc2VgXb8T3Zc1rOejRytg+p
bIoQYH9IKuNurIrSyi5RWSP0GlotuMwi3R+kOtNn7BG/J8YOxkDL2JAbsNNUdDalRYJYiCcaCxpJ
YWaQs+LRS1YvgUALgpyY94qV+mOSgpWzol9TPO020LjaRhP+WJ0Znj3Qfhmfpp/UcSRUOij8KE9V
MbLaNncR6ZMT2dJCUZLHRAopP6yyYsVIyfm+KNgG6OH4+7jhXWzj9y/UHcdmaxueJo8+yfXp/kqb
dxsOq3UhMEJFYrSkkF6bHuewgpCH+vNRWPsgBLwquzphM2Cl92wkNyxLubUr9SL4ApN7onps1f8H
q5O3s840ehmHSl2AN2IAU0ldu5RWL+L7gdOBWyK5a7Wrnj8MXl7rsJjTqvE7YrcFzd2zEkNjsWtp
WOIUYfgfWRaVDO9GfqKxoBivt9aRPhtxkirlgFSPQwebNFJ7WM0lQ5fNV5BMdQ4L5haU0lmXYdXh
03AmKyEFlqNUEEsC3HJT+icwBmyiVJY8AhbAk3g798Y1aX0LcjfohY58tVnAUUVO4KNvS2tCIKc2
myyhzITPJvKLLpFfQWOlrB6DRpxc003e1iMFn6PyUn+6VQ6T6MOg+VXvnAuOGXG/PVqqBc4z9aRn
w4msDy3r7+CzTOfSkYXplIqBJ848CgEymZZd0hrWdh5mb+p9ORTeqOxK9q41gNbGDwJZm+aoUNqx
/wOIuD1KLkNEJxIEyGJ/GN1ERVAKD274C0xt9uCDwdNqBOKwn7Ot9PkjERv9Lypgvu+irdxdWyln
ay5izH3+U7J0W2HFLUu/trd0ujfwbLP2wjolycIdt/Stq5KYsN6JG3fzp4hw9Rq18BIbA0kg3vMn
FV6c7rRN78vv7ZCR8R3I6iT/OsOoyaM9nvrLgvatnXMUWxmVGxOjc1PIfcdQTIbJiOVwPXe4kx4D
yoenqlXFsMQpTQkXk9Imj7onVDgBKgGe2pH+j90T3F0ylSyWbmz3YQbgsETY7Z/HuCHLoHqOvh2i
hxxy5xf7b3SfQ7rTBsPh8loVWO/89FcdD954QgtZCurctSRYWnEstTV1ERNSvPoUZHkjl8gnkCuV
7yRsTa6l/AixC4HE7dyFIGQ2OZNVNuSR7UVFCOyvQtqOamjzteLLIvIyl+5Sgtqb7AgBvFlYwXHz
GXUjK08aNEAPipfaVib7YEn4CvNby8GZgnm0gyQ0gxYSUw5rJd0AuCmYGtuCEy5eIPDsFkWt2qSO
UC7PipGlNI+N0TROfm34tGndG9QcLyBgdWsuzUoYpNjoOSCGKIz3o226JIDSBD8GZZdJtMS7faV/
4aCVS4x8WDbFTdTsPJFHotX/HuVQSYvLPQYf9HxY+PJQmUmH85CiyoeYN9Ru1HhR2ZGx1A7Rw5z1
qsRpPySRhpusMWEREGts7LU5FNLDgquUXtrUq6QxjYxDUolbS3U4vh98eGcXm5Hy8V/SJ3d/Zf5U
sQM8sKJLgC++tTcMIDjKowaxMOXgi+0jw1VzBveLjtpceoOtnvrcBbYPW2EC+n6MhQ373FptR+zk
eYxf4/cQPV+IOswquNCuDtZY/8kB2qxdtImsjQUOpB9YlV4sq7BDH0LatGsPlH91BxPNYIw15+90
PK4EtcyYtUXuJqsCYOg7syPIweqBv99H+n3DCwPNxOcpjWtp2SQ92mwsTucd3GhrGVvkpTj7uu7y
YsCg4C2zudpCYRS4uTpTBYvrIoY+MCm2DhctonGEtfkW/xOrYBwqwgDprlMBGZzdOnJ4BFaqMxQs
P9Tkog8BKQtjgbfcod83e/Nn8pqTftix9cJdp1wpE0MTzR4nYca8pbpZluZwgVqNRJf1pjNeBPt+
j3uj1S7igTaPReUyqI4RmB/SCKBZjpkx5y+W5LN5ZJILHKtrMTN1gqiB7j3KWxej+2G5cVWPBqHl
xKP6QhtmHbUsTHygTeJ0ci2sPBUfswX5afq541CSZ3VFx+lxRqqZlzH0EXzObsfWx55X8MQpI9xU
eW3kCLDDMfjqRslYmxLD5X7zZ+wIprQZGMTzuMSIfQTK7hYTpGi08FNdnVxjoZ3Y0cm/5wtW/CPh
3EFFio3Rcb1X4311HY0ZfD1wnVnp2Zl5ZbLYRYBUO7kvuRfYSuknwIQ1g+VmcoZk7lFyeRb+qz89
s+Jz3W3Q+bdapiczxkawAQzHMWzqRwHe1HNCDgFyKRQ0oO0SYDZgGxG1m+D5GB2r+6BigMkUwcJi
5WS7k7BteUTycrNZzvGf4+YGXLDsHZzg9/Oefdub/7E5KRmEc/ds+aVpXSgmPdiG2XxwhT/RaGsT
4PZK7axqMC3ZgyMxsXBHnYHOCspD+azscp3WH+nO4jta3xAuqnpeJKn39EGxd9jsaBHoHirCQSyc
5zeVOm4F18B4DrL9AFFXhYMcH7cB8JwkGAQf59gAY3u5Kk9nRMaYBMkYigU6bJGXxmHmi+X1hAF3
3WmvNufNIyKuDhfINRGNHZd28gjrtaWALlP+JYZa75B6k3oMJ4pYAAT8bm1XgM9fx5lesMltw/yl
99dUDRlBl4sFT77pdJ/jB808VkVAaLPVStWcSz7GUylb03jrsDeF4lzc/n7I/VfHW7jeDA//fQOq
jLJo8p4fqaSMNHKxJETFxe3EgiboKdSeaXc/7Q+JjgznEvimz9jaj7Wg5FbITptYbgDhNCkXeI47
rBvV8C6N5FCfxjZBQoEe9J2zvo+IcYhNI55riDO3bnez6u2vi00TBAR57wEie9Lv8AwUrTyWikQ7
1lBnmiZYX8Xx9Cwbs0j5BeWcRqOU1gZRAtK6AUjdieX2aQk0ladSrYZx3VXr0ssVswfgNHQ4nxRA
DrOXZrKk2LSAIUwXacLEJyeSHI9t0CltbQDjNExu8kt03qiZBaButNQRqYwRg0iVGf4w7Qi0gMzK
pH7J596BqufvBcgoWno47dBIh1zSRN27iSQSnAYiaz/MwF20aCMmO/pt4QxiePyMiUT3SzxaklAm
IQvxXIGxAQiYjVO59ROd586l5EldjiY5kt+AFhmcUVw0Rh8jTeeU0Yr/uyCfbheIuCnn2/zfATNs
Wf2Qg6L0JojamFCsVNjRmydFxDKMJouu+/j5YePuHPJjbZtW3/gMKMJ+0oo1bSnFJJYW6aMJP64t
nHIx+XnDo+JqWnLG5Looox1IFW/5MWWU67jsIjZERHYFRikkMQTeFlEAaLsa7nUAx+5d5JSS56WA
7zn/EEaumPJdfnL9fau4HRyoas4rihfLGoCgoXrf/wVGuPpsKtyfWgbZ9EGM4SVmlgEsz3ba+PLE
0TEx7D7hmpuPmMFzLqYDGWcGKXbKrkasZSppNi//3UkHrjxHpt/Tl/m+nboSysF9kXqPXD5IFfvL
A6BRZR+m1Kk3ooHBdGKDldi65HgcRMOvhNydA8NS8Rw1VYd9qocQS7Gy9McEQ0ohjOko29E5R8bk
8nP9NC3PtXDgEI5XYIYyCsBImzHAKFNXLl7G1m1kswkGTgBlzS8SCYROCCWasN3uh04dIJNlBtYU
DX5XSajdcRuLKgYV+KmAgyiUxMNsID8OHGBUV40U2MJunjg2bkd5lzXv2oBg5FaZtdiRF3Zo/kBJ
jxfXVNoJCbbtjR9Jmqys06WJIXbg7Ioo7HMhiumuDQU2AxEGlp/uP8kemPXi2nIWRGlRXzR1VqOl
EfusZg2QUT7CxvhT2+1A9BFmnp1vxtDUnoTovJ9LpbMAUOSTyVMDQEi+rZ0GY2T8WqYJGJ5xtpKi
j88/paA78CIjxMVVEE/eVLQPe9EDaX3o4Fp07vX1Ut7JDUR9nOu2UPCYuFIw83LIxsuObXiQQCZw
U8Xo0WPDHlsgz0gEfEYlIu21hh82EkgB8rwttwEzhDWqWxUtjQZwEVJt0ZEEQBIwuu1M5H2DZMJb
mOZc/PJ0XnnwiZI5NkYzF92sd/FFYlstdkjfpVFFE/G/IwiH6JO6vSvlB5NIaeDYP1XZJWRxqGRG
Kr+LiZB+6eFZrBCFHCRTIud+2kqWdLDir+m569t8gnPzZt/YIXi3C3CMBAa+vLzZGzoPrrXQQ1iR
JzCmc5q0Nm+Worcpidn2l+QOF/ZHXuvQ4XuY9hbM/AMy+8JKuLwu0glJg9fwWXY5JxwC57sW4H2z
2YIYTFf4+ud8TjcQoehqdRmQtRhrtWW+fXuHnWmAiYFpXVkCbrmQvM/66jnUnBuDen54YoJLyFVg
ZMiFxZpWjJB82wNIJnGqvnXtA+44hYf2ZZUgAedd+hkVVc4C04k0yYpMTQjefnfsa26xgmoSqzgG
JDZGC6eGf2WB49Tq3bGkeBR52DPtMZn9ugf02XFZ7Xec8nJN/sjeN7FY5qWjhl7jTAUvChQv38xk
ci9ZBrpOhUZQf9RGED6t0IKzYiOhueJbLknLsRoQ7W3DhulDKEYC3+x0MooO1osjgnGW9tIGv/AA
+fx2v3oGpOzY4TkyKaQZ/Tn2tQmTtGAO3zgWBrn95mkooms/uQoxt5YougeHHR9BIImuXpeFQb+X
xLNc5ZbDfjz3z4w1S6l3yP5DWiikEFfuYEc0Qm/Nmw3neprYiWFy89Gejr8zItGl2sW8ps+UGPoh
OlJlte0QLKMGCaJVYKyJxJ5wv/igJ6NSdU3mat1zUw+Rh6Ug/2tznco/dyjOrMS5ucR591MNYe9K
yit6Vjwa8b8S5vR9s9wKAuVwwYp6c47kovZrOHpLbzqPSDlXX1DOSsGPb0t1KazIp6T1txmofqzR
zS8WJ8WYxa0YhWWxEwej73xtI6tF3rXJrpEFnUAHFFP8/tYppQMM2o6TkxknZ8jyQshhNTL+0D41
R9qN6aUiAQXBObQiKKkha7OO1UPqmp7SZcUkBTr3u0tRxKqFZeUf67FsMuivwVg3Qr9IrAdnt+Nn
jtH7QFuic8cbflfxjhnRhxbQpkVD17PBIEoUPpKbPz/8PyfChe8FVrxzXxYxjg6YfwpoxxnMzuqu
+0rbvHSzNMGf7cXtIEpGsaBmQViDPHMLUD7t1MCWMbINCrPbmVV7GKSBHt5+v7NMSCGq0OJfl122
L0hIFGlcvKrTdUU0iMEk9ORZALKTYu1/46Re7mnUQd0K/LsdIPYad1hA0tSg4PGYappaswmvfAXg
ovS99/pY8+iaI9bO03hdT0H8c2kRgpSn2iAOrJDfZ1kr8kzRvU8t1aXOUscZL8FpKMlmcv1CqsC4
q83NF7n2UkIKxu9x8vnvSwpQU69wXT0yvW/32buzdHAoLwSZyCDbFTn0+m4Q0a2n1F2Z/kTRHllK
cwBiKCYD+JfaK58BYilFklZzhUlnmZK9KhwplxkYUeCKJwTa18sf3DuyATEKztA9RcGSZ4dQP17s
Xry3YG8TyK00Pe58rIAw+e9QorYFxvjsYPbh1yv64PS5t2uqLr5jEnlpiTf/mw/4onNrFTzOWEZp
d+7ScUZq/0Vea4HPwCkcw44V58nZZM5Gsjeno1DH/6TQBXNnd+Qya6Y/B6jBSQFnyj6/z2e1WaDe
k9kKEAMqTNk4SxJVpytwteupuCnZr/6caH5YmHrM09Z468XaNb0A8ZNeyJ7UgkPAjGMsgJI05BiY
vLUJmbTOgRPDK5FinwEDeuPrv3LdD9g50FOxI0zBln6E2Q9C0JqKOL50752YeinEfSoJA8nydJon
KzCxu3fQeHxdlfYwB2T11WEE4DHOQffN8M85GWMsarj8lRuJWDw+qE30Na7IVWh93rtnqj9uw/8o
xAXcvMA5j2np6YuO+jJYLIY47ILyHFmU3Edsj2UAV6FkxoS3XjMvfwq105lMJQ0Gklbigb8UIy/e
0uSxNIC3uE2OA4qLwy9SemD9HeT1lVbZgzhpp2P8DRX9WL/iNhFFYj32rYTczuca2yhZVDUJcB1I
hHwN4eYqoOU6i5Dhy4ESc7K12yGRv0gVrBNf/W4OXYjmtQ5IALtrpFUGWDiieCe0BnkYZLYnUsuU
FNcUL+7yxB2jPP7rzMBHi/D/pl1zjZalzqGH8hl9vd+MsINUrDkhY2SHXwSYw1mKsx/rpGQ2Gmje
jG3ku3a0QKJZS+9kXIuqvFuMlGz5dOWfDHJWGWG++eqz6eWI+d08NwslBBg1vYxClxgWy56261hn
jRTj1YNxAXm/NciiEhvFMb/+EAG/pj90EfmrL2WMXEcK11P34E8UJsV5T9puROgRldImi2IbnP1T
YyUnlsLj8ERXebPzIJYuovKwKvJaSUqclw7l9LuUdSbIEcSyl/WZkEDoJguzU6sUUfT0+HoPYnJN
AecbDyePf05bebldnYqwfmL/NHaXDpl8IzohHn5LeoDv5l/lwwSQfohYR1zyUgoZF9FxFBLkQguP
Qq+IO11bMoDAxLfWoEWanHzLUQvWuh4uz0r34O0lExHVAQZWzDM/LuKGjGXeurRz1hfUfWCFx2oX
52aagB+PZSlk4nGW3NMJFVynNRgHRgKzmSn3wCQvZFref2WStAYM1eZM41TxE9O0gO1DoD/XtJCk
47JTtA02q9X++uAIjv7dJTL2mR0PJAyqg5HSHfS28cRrLILgtJ8i0DJ7ac+yBwY345PtHuM5vzBg
e7vIUyKb3xPa5ju7o11PFQXbz8fdRrfsgxZi7NAn/vaCCf6P8qByVr8tqn/w3m6XKb+681ypOOSG
zwb3VPVDCJWyngdOg9okOXWNWr5PVtK4VuwM+GdlhnM/JvOf+2c0C6fScm3FzJ/BsVBK9bmtzMwq
V3w8EVmhvQLlwCjpcV7KsB4VtxrJ5LhgZMuYWTIhn7/iW9dyr92AmEgQD+4vXNCsvn97BzX7zmbq
SLUCie+gjcf+jw29yXWH7tv1XQ5ee8wEcIVfBAYWtHghvFkrmE9y1HwqDnXcZK9ux5vxYLABMfXb
WAwUJMWxo8YGpqdmXa8iVWLL0vZNTMujfT2P4rCuAGcVF9YF9lkhCbwgIvn8JgtelPmWBlk9xYL0
SjA65d8vAxkD0vSi80EQExtj5OcMxO1hR2B4JvRTDR/4m3JHEBtM42uqH1fQMXPiJR0qyZvSE8Hs
TJfqpiQ8f5W80YGuKnqGsfukv9pZw4VkSpz0d+vvU46LpSfUN6rGLUGGlQjT2jZAig5JAJsUI3Ia
9kyM4+ebWlUKiiySOUNoo7+//MnFKF1SmgeeeRG4DNR0dZUbbfxe9jlOe3N5K3QYkcpy+sczCjUL
jWoD3PWfnvEbv+OJoKsgCUhH+MvPjqnK7W7YveOAwByCZtgfrxIIkgAqwuf6YK01JXmJBvWL0dRw
qUaXX6/s9m6iErlvyBx/RcQBn3bMCxZAteKF8pULasPd4F8b/o1c3u35yxGI0mASGktqyJ9/715e
dCrmifaioYy9krFxg5cb7TQoCq4JHr+5lf2Nqjxbpy6Hv+SCV4kQNuW8RtpyaT31rGeh5mRoXtZR
XKiEAJAa1WnJC5iDeIeMFJs+bQpJQ+4QhmiHvEvFmNk2KaE/irlpBaiPjFJqvAtHaS8BVvFAGQe0
IZXtJ27CMmBaHgkBWKg8EvRC+YmdRYYN8xXqGo4PWI6aztwzlTKzmcEoq2BFvDchgKYAYbrcICv3
ruCyX6EF7xKXuIzkU/sePpL0Q0Zz1wIsdUawInx9TFQhtOs/3HwB7E8gf20OVUwMpuWXudOS0a8w
tWR8UT4DJ6J+D1rzrv6xXN+HmfIIseHSc1wrvjkuQdrUVfA/U8OcBDlHr9qjLZCQcjws20+6KKd/
FLxAD5Pq+FAgS4RGkRGDpwBJAH3jC7NxzYdIxNeDibi0SE8F06RzYTsLXlV/tvVg4qsnuK8cfjRX
SiAQK+iGosYBqp6Ah8MXmn/5R1nvAWQ7qGUpVSw1gc/eRUfq6Z8fxL5Y/+OxoACa2tY7zZiYl3CB
aWCOG5o6N5CYVJ7uf+Wddwaj+jHoDbIVyQc4hXFEGa0MMyG9o4LetjgD0Fa5vfa4zwomwIuLWmb7
wdjcM94lppBs276PCbK6MB9AMquO6brC9E8tPF44sCRaXyezlGpmkcz0YhuoJcHlBXc8vJps5sHj
tKCAL88A53euUvc4148+zPcKYwYug7luPTleG1BmbiQLRf5s65djPUfb4yCtKbrS6sKXQNmaEI0Q
yqPE3y15XFFLH7ubQ0y+5agTWP1eO7huScDo9BH+yzjWiT62lD2gUTc+RcU7hdkSLgDyUL4pTytx
8ay1DQpXH3VrpsU4WoHetfQU5lVr7QcHiOKW4/wmtkIulJUUX9j7HOtHZEYAZZiVhx+kke8cbaWI
dDXZlllAB588N2WpGm10TnnScMevO+MwQ+taSFNXbSgCZwYJ0d0318jl3+QPRDTEQRRw/fJ6ynWK
SiCQb+NuwoDv+NPnHHg8/qRsoFzee2j4AMGITCvMG2OdQxwVrfttbPyp3duefXaYX9LKrblDmesQ
36C2l/JstxFnbvVPCtl5fFTigefKjwrUy98CggQRshUjlEIzsMBpEo0jmxZrbhNJrWyLeBj/QJR4
IVYftf7N8Qi19omBFH4lyrnbqj+wycq2uYyYymatBpcEjdkJ8g3AN7Iu+XEiGbgO4ewnwak5wk8N
yuOP3K9xr09UsgkPJyDO5p5cy3GUxzSx5/Rv4j7fOVQymt+rbUxSV7FbpG2+l2TAqCALbRuqegkv
RRf5oz3rDHvFhjRT7o6aU9VyQm+DCEZmGhxz4qNRZv4L/8q2vc8m2HKlfD3DQgXEuHFRJlUFttrp
DSvMjZdgXdkaqgewCKz1nvV5LcO9E9FlpJRYdG7q57CWEloHpDvUmurYy23exPaA3VChtL/aezgA
EWL+EFznu0U4cgahScXkN3gKJ0wNCx6uj8hFH5C2D+FqwAiyy7K1nVPzrZzXR9B+NF7B77pChVzf
Zocs7MpEblmKXsvtYXZPzH/Dcmpi69vvZZUX6OY2/zrGxkFbCN2yX6cle2YS3djmymOFxIVSL7V8
+qeX+tYy9z7E9eb+g2uxSRpKI3i8MsURV95N59RbJaDLbM5GVJigupYb8fgXxG8w7Gn6amaK/mgD
Rzt4eAdDsDAytzTTO/Ygh58taGzSu68KpPh1BqN3hrzNHY0c+mmw/L20kcBvhPHjLvQ55aFguEOv
nrQaMGCNzVAH1ZBVz0QprMkCWhSYxd/fFkpJ5b/COhEf1mt482yCmKYflYG5439WdAXFqSvO5v19
VWGVGAsfgayDzGbZs3ZrzbxEULR7+eQ7F9Y+jd6T98eh/PtbAsz6GQb/eTEFAsmVK7ZvwWPdYfdX
i/yXS4dwpPsVcSOFEoYqU3nKHeyMmx8/El5GxAAxXTjvhz5mYolGJ/s/WSwa4RD5liT22ljSUN1J
oo39l6tyIa+TOsAGmBCa/Xn1z6TnaFg/hxVeg7lps6XGd/jjvXTCL34VZz5xTv+qixI31ADBu/15
mEPzzJTVlVM+lCOrTuAAvaFffqEu0x1YonNyz0mnQIW3HGmvf+ff+D55CWbdSuccKdBxbMFtxKrX
jnbKL0pIPsyK+Y7p94akQDpIjBcFNVm0SFAOHKCj9W8IyCkG+R/2bkV9aTE+ShJhjinDFShAQbiD
SprnRWc5lsUDk5f39CTKWLHb5bqaHNFA+5bC06tkyOqTqexqHq3kNfp+NSkAbyqkRCyd5avZ/77C
+7ai7txb8w+H5JJ/IWCFGRwQu+G/K2Odbg4EpBHh0TlTdLe3BnsKslfetXClCd0zi+znxnaB/5Ok
HxzdVDwz7bcx9OHbCyotgfiaoYEozhafiM/7vAg6klWJeCmIwprmoXwO7UMPPXppNUYE5BL0xDwU
qCrF7XvOx3Z5IfHFqld4w9Ng2S75IWj8zLDUXftNp3CdFOzVilgiZh9JkbLMkO+fo8fqEUKTtlKw
5iWP0v24uIao7gKsqP06AbQ8/CRDggt7HySfpbJo8H+TLdNbSSQdlqMwXzZssmSZ0IhfzcOI4T3s
EwJhkv4fotHeu1dYV7lmiXDZYfeZnrW6w8F/K4rRiIfpZYS/g+SfjJdZHnra/oIHSTmxKTvl+62F
r6tV8rsKY8pYP1VhdEp9fQgtt2PEsHJQdx9YeD3YeAH1XQdC0HNcFnUpdP1Sm7Gcd5toc9KUzKES
hfxSBshigf1lAauik1HWYXU0EXRNZSebPpolbOxR8p95KpYjc77xlkbwvLkBZLPkDB6yiDgvUtMx
5+e1N+NxbodrHsa/2OXU0TKe+LiQOB1kH9/IVbr1n9E75e3xqcBFte2fcgrHZMiAhnaDG0xoXsDn
CUZGI79wCs3tk/Uus7FvCt6MFbDlFQxeF9f1Zv3w6dpz5+ioAwm2Ayq/7nBx+lHMcmMGJG5XXIvr
C2vjcTasvoeJC8yv4osKXs9AKqllE7E/n2y8YDZVP1DQpNnMN4q3EAP3ZM8in2D9oqUo2K+Z7vCc
mH7EWB8mARE8LcyGGVfTSlhcX0gm5bfMFGVOBTc9eTbzlJ3lW+NN2+EZK6j9lDF9f+8lnTRrMCCw
7vMTJelI5DUST++aY6XKO5s35yvwV11i50Y694U1hiX38yDv5p7e+UsY6rTK5pWL3Kby4sI2z8JI
yaWQHsl8Bf+uHWOoRK5Kwii67fjsxnqNuP5TCCL/G8nkxDOXbII9Dpocz+v4HhhZndGbMXoMxxXU
Nd9XILgb9aYvh5tUde/G2JFnZ0b+8KhpJTh+SGTfcHKNe05AgrFRtqsxKAxncQfAF+v1LjsHxPcB
RuVwxlbdK0zoAU7KfUFf4Guhb1hfu6TuFyQB8WEo+v/aYjZ+XQuck9i5P+A4fORspYo1Prug25yC
ZqsltKWqPNN0O4IFPKc0xygEos6bRIDDsm9rp6S8Myz7djfcaHTtTT8VCOzjrgfZxCg9edOlWUE9
HYw1LlM8l/rHwA3O53Zgc7mLH8tPZ+xpzWJa9oX98CFDF4bxRZyxA7HbQipUfOIyuh8+gxPQGzvk
uhWsmEI6+BYKXk+x4enU2fXaYASpIgMorureU9gNmSg1Tw3lGT+anZjSAlHwOHZh/VYs2YAmsEsT
+F3bQSEnevgA2TykvtXX2ik1sdL2EVW1j5T1LiknUEMfK+THi34i11HXV3ZgRuAn0AqCPIm+HAAz
MDy7ycP/7Vo36ZgeORsqjQrdwF+OqFP2EDqNE310d8Xtzuob7CrdgSzLJC+IeM63XGrOaK69AAn1
f7UPgK+Jyq/CMTKpWjgr57SLTUOYUseeiRrAw0zX9ds6t83eGM24F2HRXrt9dNMUzD6ocMvuWxZb
4LCaYXLHEMHtjSsSnceUg/YhXriJWnPAbiX1ru+k0PHB9a9f3Ns+Cay46OLUyniXzNAeGUKZ8Eer
VQERih0DT1qwDOD9qezmeMisbM0H5+QyCq4MNEgnSxzrG6MeZ+dVp0hpFJPek0Z/x79RBJi0mEiR
R3A4RCEw5+byiMO6Pta8st9gs5T+MWdC7mQPWZ4RgGHV+Bcibf4sXhbCdKMIp6XGken7kPIp3iTn
OBNkvgnJE0hlJ17jaoneHr658R0un34EZbicj8NNu+JMSYrTXiPVocnTdytjJw0ipEdLqqu75IFy
Z+SEigRiujnpzl4F3cBeWrpQMXEwO12otgK8ieWB/w4LNKn5AJUtjH90ilgG8PegYRgtl7CwKLS5
Nl7ugfVrt7fvspyO53vO+Ofy/x8cKlZd/ayWCVKRZe4eG+RCxAzd86vs2LylbtJAFs92nZYIuDrn
rqyfzBALMso936e72ty031bCQ/zT7ZRmDIxt1qcxhiWKMK8GapesgtSUTeu4VgpDqda9ZD8aPt+t
98qFV4sYIQFgkHuzjOt07JCUdB5CVQpEOfNAuF5dbWeOla1quU6seJoLY9fmH6F3R/wB3OzOYqsF
Zd06BY2P9bm5m2iMFzsO+lQkHg4yfF71qGKymvp/lB/ZUqwU/bVgN12+HbnK62+slsahPWfuxadg
yOnPPjN340awnV28Nv3niweU90khtiYROGfSIAUcFrE8ob1Rsj1s0U49hLKQpVx6RQOTGpLqiP/4
iPD3Y1d1hHqX4osX1tokP7WsXD5NBCpvjxTNPCLOLTPWeqMaSAydLtiFexIVFXS0TOfKz+lBsiWk
Ci5ZfurbEQS4ItZsp+pmlLA19I2P1oKMomc5wIM2T4LblWzsq/e8w90J4ZtR8u/NYOHebJ3OwXep
pFOu9vfcJuJSwWNxeOEhJB4rEBG2zGNcrot4xtlfRDFFDpXjk6KJfX2kwWFhaDuZuN4jIyon6CHV
F3+7zF3HxJHnKOgWwHGWRo6VE7XBzV8NVG/FdCC9ea4nEQhcTcI/33DB+F99rhC/duhEEutrgkfg
/BRcG2/XXVYdWCWWNaf6GF7gdIuYHkEiSs4hAYRRypv+lgcWfiy32VhjsTxCgKVZZZmTDcwSABik
ViL6pHS6UvFZFRCRoGJDIN8dihyqsBLe2BSArlSM4u8G0V+9taI+eQWWhYoda1hS6Nld5V1EtFvN
wedRgQ5P66b6FThxHdAKktFDRDPVO0JFkEU10R9GckwgnDDtZqJ8kcBeDd4tpMbO9B/eDM5gVmaN
x7zgySazwgi1JQlKh1lxJ04YoshCDIRk+0YV2wpSxkPiwPltrniuQz4NK2CL3NU+4+6nUEsr6wW+
Z7reg38dnHqYpcE+d26Vsp3qn4lmg+oHBLsxRjwv+gxskMpKHp2dNCuLOf7OsRz+iv7VB8cUXTe5
kZ156d+dj+IJQpbpdtXmsmHpHM/cCZiDf4dZrUftks25UahdZYwDIY8llOwU6nv3KbYEUi6BNUtT
kxJGppZ/wBkKmRYJZDrMvlBsopRJRPCS1SiaItObZiyvz6twN2AgoMV5Y2SQ7GwV2DpkCqZYHykx
LxvdlEoczWPjThrFUolTcj31CW4JqKIuKAMdzud1UVlJdQdahncaRFQAov3Ydoo9iEyU62InvZpS
3w3HQAxrgWJPBfz+1TUGZjCH42zrQ1TWwkpVI+8yu3jaovgeVcLHzgP4HVxKraNkF51mzQNIMIBs
NBDMfZYis0pIwd7PxgLhtrTtNA+oyPdTX5rBMo2JazPnkonbZ+U18I/y/g3lwqNCPYzRyCWjoHaG
CdMG5BjR202/GxyLxwrp6qPTIRyv/wWxNu+tnLvcp2me5f3G5EYg2YcigaZ53WTX1brwEVsi6rcD
MfT83shzcqi5osfguKYB/Ybxz5oqkVkqu9z4J3Q6Y1WzRUSKT+znOigg/lSkzap8FNpCKu8ZSHPZ
wM/nMaElnGi7vPbLlv5yQrrxi5BThNYkzi6UnO7d8M26gCOfJdYbQmLB2W0VhJpCdPJ9dzLNSxDD
aeOBwrmgKu/I7kGQKLjnLM5rD7T2D4yRR3PRyBt47GwQt2GcpRFV27vU/wvWLXQUYV2wkBdwD4Fe
9aRmjiqzp1tbM8SuhlNJn79unSCpGcerpHQcFRYWEpNEq3jv8qKImfmsO606dLWMFUNU2ulhTmxR
RH3d+TDwOgtHCpSIwUz+MvjaZ0FF0vCi3DbA3zhkrktcsBV31WG8o1s6rEUh8a5pjXxNuZq0iHEm
8WNmU+jhyl9d5MyNHs8enkxW9IGowu+fHSpVFq+tjlHsCnmCLdiIG7l9kesiIOpbk8mggKhOV38X
QiejAq28/1+zZTrkhugQZBSWLqxqjdwGl2VOEf4K2NDdxGSKmgckAQV50RHCmcR4kuiDOouRv+2T
zy8txSnr62/sw90Rmirjh1DEpe6/f6qGfW5m0KWZ/uTWVqd6TDKWIIAr+VnWMf0jXf6EjSdxKhlK
TMXVHxoelJirNNqDLXPxYgubrZmrJbewO5ikfMfIJsJQJ6PeXyt3cGwtkv7obQYWP8jrGP2PedWZ
04zlq58uXLKSU9evNM/ZCu9VH38zVkiLgKSJ6X9KodudtJDcagpg0EoGRKMkZmkGvdGEf9YFGCG5
3+xBKnOzfA+TQlbu4Z/1mGXPK7ssyLLyA4xSjFP2hxZ7UDelkRuZl7x5K/qjcmw3KyMi4b5ty04I
qUfwNyce8aWHwIO8q9GIHIJsD2OYp3UQdk/OsDac416eF8GJtpKaxOCpS8L2KJMwQEBALxVDYVxH
6V1UceEFYOgjAat8WOGkgH3tEu9D53C1uXrnULN3uky9FsnGZ2olsrBYxf7uL7fH+RusVzeeppNO
x/vcQ/j1IoYIV7QUMbr1umjRyNGf3raMU5tQ6d4VPPzCdSlGH+K7yNIcPqKGlYdo0gKKvLUFeovv
Hnxqe8qJdlbHVU6GJsROBRGTeXomgtxZrlkQxF85m9aYrNnqsF3TdUpONPui0J3eH8eV3enFfvnt
yIFaWNOrbQ47IeCQ5XTuAOzYeckcKjbVx+u/QrPfNbXODlr55PHVbp7thFsmqMCec5+gku7KzcHh
Vsu5jqPR8yCt1Vpln72yyTZVvv5uNDCyl2IyfdZ7gIOrIPtof3P8OiwrDyUtP+lRoHePvTo1Aazn
R4uv/5eC1KAOCG6euXeod5xi5rdjCSD6C9Cunh6+8Y02pdrO4GpI5rJUnYF0jUcHqbstFQnt3btS
UrOCMdaWmxZbhWd9Pac289da03omHRtKBr10cXweeIL2rnGtwYzHQofShAkBEWgMPw2AbGTstmL/
qL9Q1lNq/GufBGSPtoyQUHpk73BbBp7pxntXd8QFa+EvWuOK3noI6hN2Xjjx5vBPa6iSPRnWQE1W
WDyAZxJauXMj1MJkHTHLv1ulP1w9IX4uNEeBL7DKLVHIW4iX74nzHamY49gg1EyPZT9jZ4aL+ll8
cjdon3VlvL9QNNWFXjd5wyRv8IvQc7IPSrPMAigG+MvteW0xPhFQIafXHLiZ5n740SZdywHAa0gs
ul3IluRuf5UsS0q6bPO8U+ygzPQHpMk/O68yG1UgiDCbR9MVWG50zMwXz11bG3YE3Jw3M3vKGwUU
DZNImecMjWnwBim9eZi2Nc6I1tVZPZseOqYTV5KMVSLvFapJuVVzQZX9oq4N0g4fL0AqfmczY8Hw
2WBZpm9HFFW9S2o2f5CyKJg276sU9ASXvH77d4Bzh2Ths7wCrZ5Vje6fMnlZW/b7kgmuMVXET6to
sEzU/cuuNHazkFizDkOUwKsuTzrkgmFJVrJ+wt2rYPMbxYghkuPWeCsIDsFbECG3JV4MCWxODxwX
UTwWOArgLhHNED4nQRO/i/iIbGOXaOiqso+4vd0s7mBrGDlskfa13fLea5uHerWFgEBPW8kxpscu
l8M8bYaGIyR+ZhOLlrOLhxYyLyji7ONtKdrYa+WeLUjlatfROMN+p+fXVRlf13MZmy9KjOFPWaQ8
3fPk4et56nyFPTHUi+D5JrM+ceEcMuu2ru2onKs3SLBfzBPYOUgD/eMbjMofNoPOgwMQBYpINwfr
35pTSZl+ZfkfpTinQipnmVkqy5m7CDNePbDVhZX66MQUWvUrsu47so8Cm1/glNdMsiSkT0DQs0JM
naNPo84JK38t41wveVHzH5LmC8LgxpUIem8Q7sO+MzckK/q5XY55z5KHZ+gOaOiLBJL2NBz4j5kv
+fe1QVKNOmvfseU7iwi6yPLew7LluwJ964eKOxIfVTyGybfstPWpgMOrWSQmNQsSTCd3k5K1LQ3v
PWAN+vlecwjmPG7vfS5PyTaGHsV2FTF53CKFqXA0qsn5/2PP8CEet9JgcQWifGR9az7rgLBMEHUI
d2v0COo9R59U4aojsPURhmKofmz+EacIlP9vClNWxnOO/3c01I2ASHmur53XDrYQF919iXvaSg2g
Cnl0BtB12T49EmMpyD1T3LCvf5ogfmMsTDIfSzhXNe8N6SZypvNLlYKmL7SQQvYZ6CBz5m76V82+
vISM0mJTPWXc/skqskPCfIcJCgfRFEgJ/l9LXA5eKS39I7AdvBSmVdi/oQE0qH53fZ1chJNawgiB
IJNf/1T2HyIiP18wCp6rPtR0JCenpRVke+5T7WGCH16fV6ALvaYiJOhi+9anvw1w9Oujzs+AdYHh
J3gerp9lUSGH9qpE3ItEncsWCgUjiuejM56Cw93ZuIIe7xnfWQQmoQCv081uvlnOe5ZW5cKD/wBr
Y6+fOzL/7EisAIf8wJ8vS518x62yG8h42C8FYLbnVlFNskWZzlB3h3RgKMaPbxB+WY150dE4f7AF
i7JO3n2r6vMmOdGQsMeBbaUiq31BkBQdDWPpePZzogSxhOUa06aM+2/aX2ulig+Ry6rF3TUUIH2B
evPlVCj2pInVDKqIQ48MjYwU+ZNsI4W29q/Ks4hC4HuzTXq2Wdsbu6CdriwPWrpwDuHkzGzH3uPk
QdIIhiOCkdWvPrIEhYU4EmuNC6bcYBcVDUjmDskQ6mMZL9eDFaejSvUsl6JHv+4hf9kMuKf0rskl
EpEIO+x2AG465ub9x5aIMtDExYAfqsrQjRlKEkmk6rsmYTpsvwmWSagIX6dzaRnbMrc36K1HTieM
nc3rJz51qNySwMCTaR3BPZZaQmRjUqcWXnRwM32rQvLKVb5k3Qhk9mUM4gRs2Vp41m4tSFwakxMz
Q1fenM3nm+IxDK+gY6qTUksZX/x9ID/eZMu/ods/rjh+/qzRgSAv45HBsO/sSPKw7qcbW3qY3+yX
/CfI2VRIl6To4yvvq7juD9/5BEMY1fAwvk18ATlFvRv4KS0CVOchyiRJUjdfE/FbfQFjl5NNLcXJ
L/KNggm5LRV0/3S4IcqJVdr0Y0MSwjtQezpo2srTg3N2uZShQ0W3rg4uoCnIDAfQlJnEWNSk5aOF
/BEA5nVj+KhJBYF5q844Gpl80C7wsSnyKTwv03tPF84ursL6b9a4yGOPU365J+rlCM0R8AvdCS6c
w4QHviZQVWhtDt4O4d1xONV+FUnMdU6/lIUmVmTFmhjbxnYVmmz8Xpm0gfXf8XrfKSmta6oC4vy/
zzNB90xZ4c706HuV4DQ02Th0V6AUmljQau0so2mxZ/ocTqzxhOjpfRW1UWMtzkZ+nvgasftMjf+k
0C8CXSXsdYyX355Yctjf1RPRMv1eGXNEcn61bVNd6ioBkFuk03cHZbWqVbpFljnCTjuZkUsMvheM
xHPHP7NfW4AwhjhrdcqviGoCwIQemFhJ4pAxBtonesMxtx55cxBgPeFdAGKCMvDDqLjOGnIHZNgR
ZrZh8m8xPJABGLXmjcjwL/1tCE76yL9d3CsaWYR4Q3f4HavgibsxX+3qLDxMImTAICXE+lqtKuae
mj421GSk5DGxRSJubQVF7+N7D6h1QjxXnm1dp7nLK/wapPIggEeRJt3sBvuF1h1OpqoI14z5QfXL
Ol/2RKxtVgEusVLp8gm92XDnMuBJ4Zw5hhMxzBU24RJ7RZ3+JUIyIY7qbFby9zBsIUwEVLwZyS3P
vLi9l8jjbN8f0EgI15Al2aEj6u9uwsCc0fTU9zRpNwvw4sJNkeg07NKcfOwlBABMzrMWBxyd7YYt
3v5zmXuhboSe8F442+QKeKdu7rvk+D7WVnKpSy59vxZxmkXgVhoujlIrIkTYxxkLEMtlNKujhB7M
ZweAgOJtuzaHS/oqAonbWXcn90FFwe7LrEjMVyJqiWqIDwchwtHc4kgpnCwiu5MonTDT90wyQ3z5
+XnEUbA4Ag6MCVvYgk8QZ0/IzTHIZkOQVN9DAzB7+suSTTOYerZotwWc4baBC/5bLD++a31jtBpO
/KKn0f6JpsO00nM1ywKkTH2DbBG06dzY7aluNgnAlTHr523Me7Gyhc2KcTYjs75JjvRX8VjOpsDn
CPaU91lWOGbVDbenx2W0LTpTlkrQgSYNESGavZ8/nrVb6D/Rtkf0AhQaAcaS23WFXMRw3KCQGlIJ
WX7vfv27uY8+79/zWOMO3Jt9wKYFQJ0EKrtwjN8rZ8a6kXRhLiJnkU8lvIrDccCU7AKbkbhSK5yt
aMBoEfdH+ldswJy3tLFL+JYWrF2biO4GzSkeH+o0p6g2xfQKULlO8/n1DusyG4QecHz4/ce6Pcky
yv3Yu1qCvjvap26zVStUvvkIQIYlICmYNjMsDeeOZKsBXIohqLr2wT0peFzQ4jOfGmhLhZXPG7Dn
pXj6wXzcSIJKIqDgylbTy2ng2Kgt7DeC0fQWd1KqBGXga3BTsHGmp5gXD6VRGHGpX1OWyX4z6pEO
PZA9x05zcdIPMAP1uSZ/m8x4B4xy35zynvQ50sn4/x4Eo2EqewojtVHP1hEWw3YX1GkZzmODoD0t
1jbxsHbZsMmoUNf6b9dsiM6h4owAolXq6kpBaIRgvGyPeOx9ql4KpZqo9kZRSlmqC2qRA16IFQNn
A8B8fnknj9mx39qJepksz2rAOfxriC/f+EWqFRgte6LZB2YVdq9sxBkSN6aJf0Nsw6ZeRX1v9ZRH
nbQlY+4MJI/PGvNfSD2xx0lCqyikBRLeI7Yso6xd5Ot6JNbXPYQrSoO936Rh1WcmK8KbFWmhyZqa
Scx1k7W1L/+/Ap5UxVqpgJN3Hmzp2E19D+hLZaQ/joVAx/VwJMSEkDr2I6WF7zTabq2XRiE9Ap5O
8BcNG/ngqtyN7UZq2W6rLL2GH/NPvClPtAJgN/gkc+R8V+x/VPnAWk0s2A5hWV9h7GLY3riG9wen
fYsNbBWE/12Q6mqdO5RSFLW5lcg1IcKuxuZlcB9uctv67ou4ePlH1zI+iFMg1LxZnG33ZEtXkGFr
P5I2wxhSHKNxsusgKc/pi+5+oYzrFX5fGwhaQi7JV8DHmXX2DMyGQp1lY7aVRPVG6660xhUsztmf
FFYpKqWDrpgxJaS/vBNGDq7cYqb6KUk5mGANcAFp7xFAvf47ysGaP4IARdAn+Tx77oxSJ2jvut8M
WTZL4lA8xR+Npb+YShvmRCICy0aw9kvbwoh5GHPCZMBhisz4sHYPP4KTUFiVjMhqL2uTDvLaFfns
WEO9fUPm6ACAKEdiSigopNMAuYzwjgEyCl/R6T+DEVqARyl863yzowile/BeVbSVeUE5ey6wU2zU
H4LmG8/z1r2SCts1wmbgFD65GAZlkupUwMOmELnbWwatWvGgNYC1LgdjPpMOeR0/qds8rCa2cXOx
3i1mNidGnzbmgXiag5qoHoPakPQ0KLjKHA5ND7W1vU8ROc6ZTyr3T70MOxUqRNOlPykjhpjAJCRS
Kj577fA4Sk6G+IQ0XTOC1/uCVfrL7ubR+WUOTUeicYIzcazjFC93soeUPCFWPt88SoWYwtO+S42O
gf1k0k8nZbR9sskIxkP0qKloRwVbXL2h6lxhpAV6aZcoCuAJJb/kny/bpQEVDSwI34Z0s8S+LCyB
63bVE2o/hD+p6Au/UQ+uluAOplyNAJmS1pN1rGYhqraIxQVoIe+8jbojYez+ZWIqjTjm6FrKnH7A
5ucrc5piFWkryGMsQkr+OPQ5ksUJSgEB0Dgoc9MhDA55ETsUWE93mYNUopOv59ethsnfcjhoqGAP
45i10SWy/c3iFCvQQ3G3f8Zh91s9Mkp57JXA/Z87PX8ReIRweR4pT1Dg0raqKsfVntkErahBWKvG
gvEjS/N7s+fDKzfWH4wT+PYdhmXRCFcvT8ppuJSTPuksE3kRLve/cI72GgTm9gBXoGvFiseZg+Co
jMWxKR7s7Ej9OO/yG1OHyYedOXWVG2cgGlZnPxG8YIWh5EZB8Jhf3JOZC2S5uYjmD5DYNaxEsHkA
nRag6JtL/nXp15FcJGMyU1pYvH3kkOg5R0pV2kXemtlSfF+IIqEf1UffCbsBsK0LivPhndHq1Gul
inBWbmo/PBYhVDNO0R1/wtYCsC9Cz+F7eIANbdMq2HSXBWFNWqimNJbkAlDF5j/kQTCj2R4dFNmH
Ecoiv9y+wT0O+9++Kp4tmo70c105O7sD1tq9ZQsotKfnfKcISTKGg8pHcTFszqtifV/Al9q0lDbg
MDQvAr2wrA2tJuvBbS65B5LweVCqMwcQvyOCevhJKOSrDmjFDYhO6lAhf3Dly1+ke357kQzr34OK
hdqs1q+UlXCamD2Kv4qDBbgI1fetkW/YGFc+G2EbOwThJH448pScSfMjU88xNPCfvTIysJ0srSgI
W5ea5Md5Dvta1RT2WqgD+VeiefisOA4mTqEgf8S29OK4Q90WYzT/sy7XfFndtbamQ1DnPOD+LxSV
dp3VOhrRfnaFdNLyz79jxPAB1hCsApDEVvzsJOtRSsEVhW5+w2+Aj2dj373neEQvcq+j17C8Q4kQ
y23/3/+/a+dErb7orwcARrKtiAvU8QZxKuP3iO0OOFLX6PYOL9MUO6QwqmjcldnEI529tPisHwZA
7PUO50oSH+NaBvNoyBUgrF2opiBCMX2JzowkjRclokZ3ubqHlz74i8Zhi+HP5N6/V4HjgHcg9JLx
cXB90qduoh2qgb4hHrCFhbgQjwJ5UXe/7upk9xMMB9EgTas1e9CY+d1IJkZ37EsyFnxRQGrCSeuI
aTuWdiUGZshOTeC/YTz/t5PbtdvO1LOlUBg9I7SUyJM5atWMIGiWG2egO8kVR/Lr6eEt1RdgoUPQ
KiXEJ92FIwYSk4GjDmlCWHogEoHTkZa6I15awjl+g7s+mZRbuRuWf0OCgH0qsK1Z1yGGxnVs9Bqa
kU38zemMmeWqq2jvpmMV5c6JCDWBgNShDxyhWshpADM5S6N5U0V2+njYEczZJo8T5jtB5X7gS4NF
G1YnTOASWyEycH64oEHmy2OeC6N4BaUp2OVzHmK0eknZ3igzMpGESkaj6VShfA9jB2QYgkjnzYmr
D6CpoGjpAcllavy1XWL5TK0lBROInJtig/AGU2GCYnVKWRisVzPWKGcMLCp+YmFT1ZFqY9B5zmH6
WRuLHuGEAjybkzRjm85RJyfarNOmasu9vLuzbJA6vwNSi9VyrUBxL7ix1BaDw1bK0+IHOk6fbkKA
KYehzwD22/f07c3zp6jcK5iMFcur7XgfSlsVCCHCexOQrQfv6zGi4I2rkf0zycZlGiRid9MIQsPu
K9a3qUFKeQ59u8YvAMCAOOyP9ky1iqHcv1wmZQYm0iSiUE3lunX5/JGRBX2EiJs9Vi5kxEVj0L2f
r/Z+J1xTI7Jku7r+IJ/bL0pK9VOKoe8nPMS6uqIH+hXpBwxqgF8FtiRutRyhv5FVt/7N+W6+Jf4w
ASeQGOaKNI/c0zB5GFCyYFVvdjuRgfNo/Gpm8G9XvYKJxdkIy1VP8uuoLakyizDqzQ4HPJwnDtKB
vSANBNsp2PQT1DyvUpNOI8L1IhQkRIBzILYcMM/46ug+2tRTTD1iqhv1KME1FJ4R4QRggNDqHvKv
3vT7MM9dQtAVL9hxm2JI+v3nEiIH38AYSagrKms+zBNHa/86t9TaCdjy8FJfdOzzrcJ4g6Bf8iby
z92aavL2TYkeLmJhK+tHHP6Na6yAAhW36JGGHYhuxs2GIAhDsiKQKoUkni1NO0DCDv2kPTkBdKfN
CUiYEAF1zF1OneKZChMJ9L/f2N8swY7dEBWYMTbgoZ4X7X/TwsD+rvyNfrqCtPAxdeOvLTYNfeLA
K2bN66TKvsHwKaOcFx+6JqySS02xC1LQl1PK0JflDXTVQIKfI+UKOLGbPoFYfUzfJwIm02o+kYMf
rlg/eIOPDIl51iAxr0Ijh6hvghwc2ItAjDL7Ly2ouyco6pzmVcYtW1hNGrw6yyI7/FhThhCgXFyn
f87Qwjc/MyLLQg+3y9Dac7v+ohACkeMYB8UyAquQMmxdAkb/iET3BDxPQsX0A669ox6hj8qk4FpT
e41NQN82pqKHaE5F078pDBR/GtI4cR3Xoh55hnHvhiLZFzt3jRc9dCJvQjV8zGxujTJ3k9+3ucSz
v9bePI7uAR1MNQBYGYPvPoqWmildR5iXszjrEC0gjfbCvfKuEM74tsNMI5JOC7Mbu4X/drf2wY2e
EG9eAMaGwD/aBCJMbzljP+YwxS4B9eTXcU6OduKE7ogbUDs/2E78hTKrfWr7gLS/hMbXnE4wldjT
hVkOwZUXd5/sPb3Pa5u+HAtQevON+VFzHX+bVCWYR6QaqnJg+US7uLi2O8ZPpXuxhlT9IMpWGT80
2T4AqrvvGO15903bBy4mOS7kbJogpvVVAIdcwbs1bb4KQs8u38ZpAmH2OL+LSu3m6lWywHWlmTag
rGXdkcYtUAtCJU8XNahsiTQ+kEPtjd1UvhFFGiUqrufNGbcZcDUL5gcVUPOOc8xbN0a5OtnH/aQj
koBcUTHF0LJt6HlMHl59HuUcCU3XgaDub+85qq+PuIIZgyZPn3fJkWRC666K/zzHXtpOvOL2cLom
3V8MFKU3IPM5Z68avRoKrJiH2x7uASxlB7rksBglxjUM7Li6f5pU1H3Ukxb7mKKTcyowVw2ii0gk
24U1Nl0vjvaz/MtHBM9tBPkbF46wGjZg7k4kOBHiDuzAvYhqcqGarXESzOFrokGsrOUZnLMkcd7j
v+9fND/DiLWqYswizpZdWci+qDFvUwwf2Rr4jpJ8SV1D7Pxc8CtuveOuwCk0NABt+wNzHKVSiqO8
0KUAth0Gx8a1oMQP1SJnjt456HCkUEx3+cg1gukIdPqvs6IqODovi7Jouaar3xckwXbUMmeetj5q
TRVgbxOlkRep/YlHRg6ivL5FGhcnZt7jJjm47ACt+ljmZOTO/khvwB0ggGVOSLG6roiiSql8j2lr
LygZINZFmTPcYFTaETEE6jbUMRYVZBjp22w/0XEnws07oPOnR4OAKbwxAVhC/Uft9k8Vf9lV9ptS
5PPLMRfAzJsdKJaK8aEuW7qR6xQYhFQ+Zn2FKcB9X7cUU4I3auwvgD5CK+ontg/avzqrjXajju2z
37hBSaReK015GRRF+2q0zYwPNaKCqNF6vCfb50vwXwkvayKEx+eJTQyhZPmXGPvwCgNRuQLqBRq8
aHx1LLT5ErVNbU7puqyVNO6pUPr4bALWaPLglbkGa1SqlUPKuLDOPzY7G8JbA5tcwEJnNe81hXFT
WPUCsKju0gotUAUTY/RwoiifO7KmuDFpXh8dnhxlUTieENVHBgA5mrFqSp7tXdQYdeGIBTjPBEgZ
CyrAEJbgOQtSxIXNGnsqBCaBn5toRnarqv8cLg+Zp0DW/kZsGa6nXE7Wr5HL1nHhBKqfTOl523iD
z7lwUEEAGvDhdbSjvSrMEc7054EEaZ/eRFIIJ5bQRyCHzzMVYmuzEtOxMW4n1DTkd4aY8aiD6D1U
o7BdEVS1kPgIP5cxTHCbPmedg1qvKAjJ7qEHw7jtravkuCZw06VJ6+eAA+zXAypQwZBIOX617bar
UFhEasV3LiNfAziYX1kL20VyaNnlQ8tqTHOdk+Q0C9gCglIQM+cM53zX1GEdgcovtxAt2o9shTi3
KOQvqr07IFIuHylpOmziNJ1c+KbFDhSg4zcMxMVT5FA+gdM2LMdIGU7bZT+fd715qjJP3V5JN+iP
I1iVWbikCBCqxwG2o+xh9tPENA8q9W6xQlDS4OFZHaClgqE4B+la690Bt1xzyNL0GiAVlVsOfJzk
Ut1/ia9tWDu35HkHdZc7Nxz0eWaN0z0QjKfCsD1DQFjkoSNLa1Dd9r2yqhpH7SelpEC64DGOn2da
EzlFeG/xUuculskYUNCOiUXuxv6SmZMLws2UCDnO09rvFbqNyQLbPm4mcjIHqIEz/fEqfixFB2Hf
0toSJ1Y7nON6gHKO92EE1YNjTuKkIPB+s98fe8xHQXNQPQbY02fHGzXWJmYprPO90EAUX2C3wGND
nOuSMaHFSUJpqh+CHTv2HDNgt1z9MLKB+QcxLKzX/+6izCWgfHE5sPsB8NCDPHdWtgDA1S+9FZeF
kHlZ2vjfX1fC6XpDLEFlsqnZhZMrvquiD64kVgP95N7pKjMad7/dppOrXeSzwJdn//nQ1VZmkTKW
3Jm38/ML7DxpklTsxU+PiKDM4+wXpSnNJALtj8Lk4Ca3RWfJTyX1JNBKWpy9wQDAmWwoys9CSjFK
ocHfWZga3smq/OUOYNnO6akpEylnCV5xK5XFl7cGfjxGQmW1UZK7M7PlfmEbun250/y0r437z0SE
l96w+SBnPdX06fPtwNIK9Mx+xqZTjkHNSiLgRACnxOAcpQI4aFS0FyPOt6/YbEtMuoyR7cNXMt5D
+6UZ12V33kg/Bu0RfYfhOkCRlFA5TP1K2FnGSNumn0/6QCrskSDcqgKTcldGb/qgvvs+RPd3Q/cy
sg42WIV/xdzNFt94xJaikCWDkJRKfoVSg0SawglNuJaTPnEqfjjevO8i3mFwwaDoGR6wC7cPZdjF
sAHyQxKLa7QYPzKdX1JybZ3W+qr6GGb5s+AS43ta4ezEUWXC8gmED2h9g5QpklCf4OhYqhvAMuYl
FnpZJdYC5pQjffQLWYQGBOovQdEUSsdUJdUhokK7hIfKNCSQ4EG5/7YTJ/pYlWhFL04OSYtMIxGx
40WxSEaXufJX+c2ae7W+bgFHWdoc74DDG/n9u4sV+N7C23EalKXqIC8Pf0bCxxTK9DdQC2IBHJq4
+nXG+71z6Qt5xJC87re3kYN24jaLlb8dGOwpoVpZcXE5ucYdTYrl4ex7B1KTg6Niu/6HhWGWI3hI
RmB2FQc7YVkXgEGIM82+IvjENFvK8EZ1troEmOhU3+vEE5KTCcsREn4YEzE4Sv4oh1f6tRwRZcEZ
ZzRLNcSHDUD51mTz2h97oJc6uTfVLMwwgQ5eT7gZG9GCzKu+ypnxqj/uaxb9CAOAQAFpUy/KmFfg
ynoXSfvLjvubbQhtI7TuCCw12g+M3ir1IitN51ZED7Rp7Rte6o80AV6ia2wJtlGFQuf6OWTjXMGF
5fkIlypg98EwnB3Zk3ui50ZNIsUQbOYPc2vC/aYVG8rH/JbWRRvVPXfPaaa2Bzo/7MWZbVvClUe7
WcbGiTkdt+NeXy6x8/xLUp7hVSDYUWx38N2yukMI/RTNXvwSX4Z/ZWPm7FT4bizg79XqyBg4ydO5
reRZsddLVPimgVKVD1MAa7jM9r0cnz3o3Dwt+vdVZqVAMZDse5KDWFvJMsl403LUmuHe1kXFNHON
zsv76VIxZvKmsWAuGWGrOBv8xgBTgHx4Y94MubPPIznGI61DGhXcG6NN/dSwEgGRH0vujSCuZkNV
z8z/+NpHM4Ci0R0SnSep0/IB8YnoUUsTLh5U1kHv2FQc6oHNTRpM6tINfsJgrdQebrVvT8Du4QgS
PIBWDNKYhYNLTNFDv0Txs8GbkEJm4JpzadH6pl8RTM0PP1W/KQSyqPqMcE6zn92DtLPOY7LPe2WR
Z2+D4maxJlOvVzzQPW+WjD1qhQrMU4uCkPjoD/DF3jEYIc2c1H1TMl+kPCBTqj4Ljrw+/cP4RHyf
4L4L1bVJhHOLl5jp2TQ5UKMNL83d6z0IsrJSpQQ8GPmHIdjmjxpczv6PnoGBxhKdqpYAaRqjBPvQ
CM9MJ+I9Ges6y3BUOMtiggRxBGbGcVfRcsdF/BbHjjv5FV7u0o+AhHa60qF2sVC9NcBHK96DfIRV
Tk1dYR5jWGJRKSqkZm9BMVDFkpOpoMRcaU7lyww2RwYf1F5FrKa5qRYgKRg49pT9IuRwxp08M8ws
SgPOSXrqXVW1bMPpzbNLVGIac1kzK2ELde/ne0wjjMXgEc0YtM7GfHizQpufcTBWPUKUr6vwC55f
mf0lvleLdcA6W3OkZ+3C3D0x6x5nPyjQposPrOTX9NgQt3FCn3D29Yv+oyjmGSOejmk38zhe+/5a
0St0hUnSG2puT3T3rStl9xvL+yT0lFkb6UZUnWBeX7tUPg4/PsYr5w9nidwv3pVyNnJ66XJe/xNe
2NVW34rytPowZr5u9J3NRGxKJxDPLvimVD+1GzsdOdkAWVOrhYJp3JjmR+GlggErjqWm/P2GSi7C
36SNGylNEy/9gVsDaL8tr1sIZAG/sDF4Izv20nzW0UNVAgjNbv6I+g18/gOWRXe2KCk/t+1/O7Va
VcV/jjGK07UhbCSZF7a8Oh5SFwHsAX3eAP7dTO4upOJzUc/DQaOOm1hqcA4R5wL9Udx61eqGGysl
sELub3qIuB6nSuVIzRfrTvA7Lk2Zyt3O5qK/6rPCjELB2shmKbaYGElcX/iogICrZsCDYL9MTYa6
MPlPdm/JoaEuBtnoVFEufaG0BdQw/aTn42bunyvQwYXuuN0aZhBSOz73iVhPU7lzuafPn74Y9bRW
RGNSrVIOdgEmUNyeDdw3Qy9d/6mMSG4kT1bX8Oz1lXZbxf5YYO3DY+PW/TKbiRmcW8ZCkAzqCFrM
dR8SZAPgGpqdz0H+mFJDAJ7C3a3VHAuhR0Ry6ABtPkNpjVDkRAqDHts4yQJdFTmllxQT7jGeA6yB
eIF5p3m1x7sjKMhDtZ9oBHRyDlsupz1POyS6Se3hOwMN3iS3Fyeh3xx6G+SLxua149klIZpUMOn9
btxLn2pGwwezPgVL/smhSSgnV2shHpjQEZMfrfWK+4DxBhqyWXB0ifPtrXClnjnv6idkXd70F4bI
wQmusDVrSUZ5AlxJo0dxAIjV6HkwNkQpRbgQp6e74eJx8G+OzgMxByVrHOyWr8VDaHxnbgUBlys1
rOqtj3geuvhqMFsoSM2p22VYsZZHKH6aGR503k/n5whie7LK8SL3ee5/6D1tBotBEnIkiqKU/pCc
NhnnMapXTHG7aGcfFJtWAdCsMIjMin/8YJz/bCPHKd717Br5OW45HrxUimWZRB8sq+CyWOmEVIIq
QyM8laP+RIsLjCPsmXs05PYb8LmrqudmA0TaPG2SNkai4F2aWepzoiYYINVSxtZXFGvqZDbV2f47
zZ+6nmVOkQbaxZhPxRXJPxK/l5H4SPflLROJGxXzf/cfcWc+ABSz1HZLdQpgmcblgEaxKCm7a5wv
kUbns5a0tzXqICiT6oOIzhVjw8NfGwgM96d/IZPBZWjI3Mzm3JeZ0MIklP65WNMqA8+cRSro6JI/
qB3sZNRpPCqcGa23HHB6K/SRm9zjGB6wpjKlVhSbqvZEki7AS+oMkiXdXjDqj35COwhyYO9TW1Ku
/YTCHRmi9fFvsrX+YyNGKFK6jSUsp+MtHmMy7bpbF6RMIE+41Xgl8qIVWnUMY852my8iYy0Nvm21
Xx2++I3cl9w2qMFg6OupCKqoVPkV3+N5xcEnypUIXuH+WEprsk+Kk8miF1DsImiRyBFNK5aNYaGv
QVMTmCpStxG9i/J2v1AvvHd76I+8cSZRSIFeZZNdizFdrzj9Ljwf0SdfiP3tdQIE3fXEOtiiDiqw
4WxnbgI2VT3ZAhCoCOjtQblpDOnL3Wwj72+JilRNscPt6V/V544P3EmDgDkrHDsqqTTvlbRwsWUC
6HvY2IS7f4/1VAbxdus1yj5Zp5OWFDJPpWuvisQEqbTf8GjUBi5fvCnA79rox6Row5TZrWJh/yto
+tNcKJyPdIOVnF/vXQ6G34bgqbkWa4FTBsYBbJpKVc18Vsm9XciX0520u0yGWgZi1Q0rvtflidE9
UlbGX0CqVV/EbBsAIkgJ6MOrh4EnRUzXvzpqdzKcaOOdWSAtikCxiFrxchI8IXPF2Fm5o4qUYDG2
Lv7Y36WV4g0ZYAkC1gbkKxBASFbFmKnZXKzhBgqeL8UVYx6wP7LsjhIF5bGLX1le4yZDb8SfjYSQ
6l5Xw+YK8EDipfekrXJosLnTaN91T9CAIrop7C0E4Na9pytPlS5AGqmZeByKVaNiYMmEtwdbB5Mb
/hLeIogmByWFOD0pmorHVLpxi12JCbI43eqhg8UdaEvhGkbrP9UmsvwWdm1u9S94aWO02voVvqj6
TqIkfRdmtOypHoBKm5fzv9NMk08x2GkRZVRqH+AHbhXjeMmq/X8fvfV5R6hI0mscy0CbHM/l6xeC
PXS6upp+F5rtW8dKPPq8kUWdV3SuCOWXY5ZVMSEcNwqvlLwlv2UE2f8ElRJRBHdXUROptkKbCdZ+
OJICzSH8u3X1CKSjevgLA5nbeZOxpU25phVG5qcbgRGVHEQUGf/nCjrf0LisAXsyB3iTvxzrKiko
+aoQn1Wc1bY+24Z0fqFoCgwUX6paC+kUaBBIcctE35EuIJykaxabJZgo0au0FX84EiBrEaehCWn1
V8Bm7My7OD4gZPGgOmI5ygFq1yHwiZruGWkEzAPbn1n8iS/7EakyhdsgWwBs2RQisBbCxolfTLBH
PftoVYJx48LtYQmp0ieHf0CtUMTGEYFll3gElw4IHYRCbRQCi5cqGPmtOSPMpPLEQ6JX+24RykGN
RX04EnOPSkJkvEnUlu4xVW87/N2nN9af6pAR44XCLpBHpxNrEgzIzMI8MYk3i5R2NTsOQQawshYA
/8zMfokNwtLJIpXHDPmUrRCgFgIX4wxp36ZGP0g1acV4mj07gHnAVD7NkygaoMVnRgUSlWrDhfm/
MtlqoDsifkrSUV6ZCWxadt2FTlya9aVMYrwW7IEuKyKxCxrFLkhYXsWl2omxCAWFbxYy6QDQvFbt
Loz4lllV7ODFQy4Btkk7BzDZt5UVVnNcT/5Ny5VHq62y27b1pRbnUEfGriOzFGYF/oSCOtH4t28y
Bs//1VocTMlyg77hCMLxagWHuks7P91EzSiI6hnIlqPVQuFNQo4lz3iCZLcMPUr3TqC3+1w6Ft4h
K2TPnkhPVVeFwTQ3GGrHokO0JMhhYixbjdKFpWF9O2HT0xYjzdzYX1hQeG66/A94tkwWOPkOPrvP
xIaTEay7NJgyGQsjEcNJwmqmonwCHhijqcqL33yKwhlF0UwOvERDnDmuQpLbeliywYRIOIKU9NKb
dBvHQMrW5w9bNYOv2382kHSX0AvgSNcpdY0gT2OKleuWyN3PzrBm/ZpVt4GkmjwjMXfTVN3h75Lj
f7tfPJvGcqYUsFHniHC4+rXUSsOcjLGck+DcN+9ytntXsV6ca/Z9itlYyBgFBi5lcgwu94Phveq0
YLoMo842em+wivHPL71JZH0SomRjnQRjZP+aIkJY83cr/Lkrw8gbwPWDX/kRVC6CvxfzEFauzzYQ
xPVXxJqGz4FU4CO31azuf0o42Zan29TfRo7fDGRBdKg0v1r21X+k2gDNe+t046gkGTwbNU0DyEXk
zfYIcvjNBNvU8tl9iTWCrTF82t50MXfEqFx1B/4OYkykTb5NJwTnAF4nZpuM2i4wbKT6fKjazUs0
cphLgnnLoDBOWXGE2+chhYq0eb1ouG4aOMh2VojP8L7ikjohaitcqVsfRThKnYUj43+zjsrL1uI4
8Jg8+gYvE8gTLvBgJqCCjerq7s6ORD2ViGVS6qvg33ZCqDldKG9hP9XUndusQ+IhzghSvWkkwke7
C3+FgoX00cP9hC6Sm5insRNda1/x3dXVN26Ys2dQxvP8WOcC6OlwhGmm7R0GQ+cVVUmawbdsOVWp
hxnK+1DWsdi/JSry+FpU6jirT3wzA0qzoOpxlp2zrTGM4dy+OAZ5mG7O6h2aipivv/GQI6NlHRTN
/vULv5WjrGTdq5x8HaK2J67FNXvPhe556tXFLGuFbpTiOoqWWuArP7f1pibNbGcC/xBwFANxiSVf
j1p7GUPK5eeiwWCO8SyO2ZFFB2+PYhoeMrV6su3rBPoVfTV7fYF572elzxXuUPxHbIqIramj8+zK
tK2mon8KIIaGVlpgcfoBZsERaD9G8GUxWa36ucFlNpHiL+Nbmas1D3Lo4mBzCxzjTpYdoKNfYskB
TSoWwxH4j3l/vVFsn2iMiKF+FT/nARZeQlJ2Xuk4o5wt1ZwjW56L9Ljv0swDQJ7roI+LEVwGhORz
mRmuFbxw3q7104tUn2Yz22QYbR8Ranz8TTbZaJ+0eivoV9Rwnr4n9QDObVkE7ytO2aceJDwkGg6B
f8l8i3u8K6xiamol/QnRpSGsJkHCAfDQ+VaTP03d6NjILqMui0TbGWUex1wA/UkU5TyBAXAb2CMD
EcN+1xJPih0o0F6j+DMoPretemosJRv8PI+Ybq+C/l2u0228dYhyZItXusvbKHkA+V62uU1F4Mle
jyuxqkpCrBbnYMqjRlkMw1CnwUyM6OKWcgIl094lVIGaeD9ufldYPX7AnW2brka09WjXyG5XosnK
7DqCSYaTileJIbN/DpyDW70jrnp1V1DB1Ob0W4MAGxLDosRiDlyY7EaWCONLxrbIYOtt4w/1+8pc
PeU/gBJvuyTuwsoh8aIHRkic4hFgDHZrTKSR2b/RmhT01u1kXvlkiXG0PhgxvLL+kA97Ncbu+Ri4
zli6eFT3PwA09kOe5PJrt5I1Qa6hZruOz786W+9LIuX4bW1226Qw2b3HFU5Md6M9y5Q7qR7NEyz/
PdFN1JJno5a38Qv/26JpqX3qgKnWWwzLpK+v/eU67CzChJpSZfJGnMRnVvyfILfTpKEBsZqs2SWg
uOS1DO0MYD2ReS7ZPIHOGjjIDuDIPtaEtHsPEZREJr6zYxUiKkKtoS18SIUea6I4Xs/KfIWa4w9y
FR4R28bxco/NgEk06W+zbVW9jDMdsCz9cPtX3bMhFV+6FrBP4lVVts0VSsEuneoL5iJ58G8Ln3ef
YTNxiuPXCklFx1LlP08nIRP29J0Hr7EPB9CX8+aoqFc6SqCg10Q2RpypV/3JJKfU/0xIVPNT7ccX
HTD5QNLB2bj8B87Lz4oHBIuLmc5N7GBxwZxEJcAZHnUrqFnhtxOZvbz+9G+Cc3U4aIZDmi1zqCdV
PUtsnwG1ctXgVSc9cnaISGu/8BcUt1//+2WhinRylUuDDW7uQb7armkBP9ryrKOhA2oq4/D3cegG
7MuqW7mtcH2sj5I/K/vh8NZRoL6OGHvlwbAKdts8k37RB/6nUmkM+LvwtCe88zM9oeFm9D9ePq/w
yUm0r0235NOLllFd/DfXJ7WJlg09B/e2VRx5OPUYvpNTWbijg+E9H0cW0WTNuMEylMnff7he9fYn
rsZ2KGHv3WX8vi3HpAq6vCObZAKb8PVzv0H01arQfAfermj6IU8tTl+h+DEg6CZkmNtdQHkrEvof
wpRWipWYUBLSUstjWbu7wMtJ9P2nMCn98kW/TfbN/O6euie6H/bCT/tM/0wbHyiPB94ZBuXdSQta
3WbbU52OySocZ0nUwPEnZjfQQ4QweADmcjrNAog4v1J0s2q4FrbJmqhzT3+xNZF9rH5Cm51L1T4O
XOhV/5+oDwK/Of/C3iu/rCHC8/E5wgAkb3aA7VEzRwr3fGOH17hn4f1ZtCNpDTraq1BYVrDf8prz
/EYgBG0LWdzyi3/TLDR4nFwJlBDcPLRk3He2EuWNrsds4m8znis7tsz41kYm71dIzUY1DiUYYwIs
kY+SYkFXks4IFKPudyj8uO3Riar3PdbK9WUGBzFyDkecjLA0g8EwmoW8tisy6L4mw+1CSOZicZxx
jBg/4WcTGGlyA2ITVV+weTlXT80FXRqwyRJI5C4CUuax/Ty68qUIdaR3sbf7e0widV1Wr4nn8KeO
3qOFxdhLD/XA/JS/ofAs5Nw7ZHDphiD7pXKqvBANiK95Ohtb7uXXiR7eRVdPM3Ps8tXADvTBNXv5
J7SDdQ/EMM3d7mgZTZPpIoIb4GMxCoS3nlz/rpBSM3NZKSkIaDC0k3/ctIyQtEMGTUfmn3U52mOF
T0oTkYpKnLkv/kj5OmO7f4gWRuOX9k+suI3tFMfncCDpp9neWmUsmo0TWzqHe+y5bCpT+RGHxjsh
Kk9M/EiafYwjQoV+6DcqDioWnxy1XqGzDIrdgPUp0j0N5AM829jIgCIeJzaQ/s+CpWr2pHGeS2c5
n2gk9u+W0N9oT29aDG2ArQGyiED2K+0r7nD3XqUOA5d5HgynKNinH194Qwf4sg91DR0VCMG8qMvx
lj0hE5WDEbABrz9NSGrZpHwti0X+En5hgP8A0GUb9xCddGEUjm5FNDkZj0ifBmvbalovtitvYHrb
WrW5kWOsD3GxN3aKK52lf0F3jdmGtxhDT7+aqT0u3lXs77syI+u7hIADsG2RUphVNbGY7bwWJotV
7AEcJKyU/tce24YyWO48aHLC/jJzbVqM9QgY3Tw5ilZzNvJuGeno+vlNl5qNrw3ypJ6TtJqOnSpK
e/d1XfNRUba4eiXCjeRJ6oBE0h55RGm+BHwEqm2jNtiiWivQR0UDhvKwnrL/83r032/RDwRdv2Vc
yCvFWysbGR36+0cw3gBvLx8VnjPtVemMONVdZ6NCfCpOVlV1iKNhwye4oRUPtGXTxs5iNF3aovb4
qyC0R4XbOAZ1CAjEgBDbpnCDKDNX3Yf7UhbBIQTOXQEtJxM2RWXp1lZg0tRn3jM4o1s3R56h/FzI
1EKv39Jh+b1G5d8eshegUoEHd30l56MEVvQXxk4yCEA6PNHkILXL5uG3xFzf+WkiNRZpthaZtHIT
ye7U9MG55ONGhMy8Twq7WSxaUfepx2BN8c9k9gEyX7b+/h1aWljSPICW+gB03eNK3+Ws78xUpe7D
CuZ2GIN1IR+SKCX2nFwlzyvEujinNTpWWxCyM8ajBnojq//Z4bKFpzTNuxeRgQGWjaWz0AWB6fvh
tHQDAFXLMi5QmreDWoOme2vxO2o6jg5oLV/a42ki7AwhjEDrSrLdiols7mhLTrC73gY3eocvDXeZ
jZW3pKDDKHNZ8ICaTtTtxXUrecpRRKC2/stir0m+gv+UIGL6Ig4SXt9OeQdKNc0ETqaaZKeK3jlR
jlbowV117kP8pl7WFqzi3IEDnydClIeg37fXG3RfITkEr4wCvR0Vs4FOdyYAU/TdDxZpGkT5v2H5
XHp0HXSUSFjoQv+XVnE49QjrCsT8tbn8RpmgZnVrD2EXykwWs52B0WMkW9Xd8QSX5GehhwfqfoTe
qSK3bjL+389cz03tptNCYvZzc7UD85tv9kwlP+5CjyDchErFj1SD9z5HvVmJpABgy0nINDPqjFrU
2OF1Urcvds7drATFDTjPEFrOloCOJX0UeWQRJ/vbXYYjZ4zeMhC4XcwRjDYOgij9f7msduohN6CQ
GXBeQ8l8Sq8jpBlUT+ZTLt9YM4XzrtLG3KPLkYljS99kFxoz5f4cBo+UDfIar3d+ngOIuGSOk/tB
uhpUudiKyNEgxIbROGI0XnhipOWzl//RRTLOX1j8pZ0y25abXqW4BhNahfSBtRgm+4ZgF7TBUy7p
Zi3H6gXJV66kCqCA/9JvcqPu8ncaxx3CI7Eb68cVNNWaPCDXryFW+Y8COUWz9oC/LSkYoC+VT9FW
OFWaG0vw7njng/qeRsZxnzTPe+5OVdsp7RoUs8KfOtayhRdJiiPBDl3Whyjt4dW82Peb7RIU0Kv3
GHi5ttO2jTM4d24vG/XXrqpI16v+zpH6T7QjxjweCVGa1vLJT/v/2LLtzTVThVCvboEiVYlFtIz9
hT61s1HY72QfcOUO77A3nwk2YRZe/is6Ckg8z3tqTH5KsEOsIDqeCtaVoLTzWNR7b3eDY4ec1SRg
pjYWaTWHEO1bqlbrZ7a5nghyo03N7JRPXK/3HhJNkJFN1sk896sF8BX/FsT5rg5qljeVjkWDWQzj
vkRhLxftz9zyBCmVHh/FCGQw2am30tREjZdWtfPzLkNOohRIq9p3zvZWjNfCSyETyPkn1xq0x8ST
A2Ar4sJFA6AwCoQWzQYfOhYoIqPwVemuxQ9HkHa91G3ShLA/FRazjZ4mGFj7VZxwteC4jVY8SSGN
a95ceAxHGk8aHaBjRAuT/eoaaWDHg6++LF4sXefHb0ZSN2iISUBOn3B8uDmIuktiFM6xMo6u5GFX
+DRO3FaXpQReLkqW/1cDMUJHoIXOpDqY4E1A46XgvspZ8jCO6mQMBiIoVmpldKXx5TXWsfN1e80A
e2e5Dw9O82cn8u/I39ORn+dbu2B+R4Uvd/prDTR6MPLs5ZgUMhdG9LxCo6lK4OW5Hbu7hY5bjut1
C0xtreu0aASGkzNVnkVgLoZ8mAMrdqVoZBZXQU4i2ZG22cwYZKPwcwMsWullVnm7kTF5W/QNy/5L
Mtmy6nRpO7J+vsgXvpY009lOutt11Vek1w10K2csdhFGosabFmtubBSZJaGskNQozxQxZmja5MpP
+h7O3iEhueaIrUG8vt8hrBIVE+3B1xWlxJNnaztCcC9lSDf3S8wi/fXmxpfHpsx3P0z41TphYyAQ
lTbxCdcEbNqB9GpOjDpEQdMQYhIzGn8vYSGOltlX4jYPUKehGnRLTxFbvhfeiZxB6ByptEaePzbF
FTho3N0Zj7fzKcDMtuvQusOY+yQZlTNv9nzt/ZlQ8tF9OtUBySuuYaWxX75RarSVSosAwWBScNYq
432+5GAxHqRtyul9uN8pGogHHhmm+JQiyIO8ElsV2tAZ5GcuEAbuaeV+NG30kjLl2Rcko/4Xx4sX
BaEzwmkJ/rSbP/8Znobzq+5nICOQpCGQF945w2TxX8ToqWQqjPCXGI6Hl/3a1Q6GtqmVu2lieh41
knl9Cnkb7xrXJjnzQWhX+AYgd8qWrtQKHvWiGEFVoTs/+T4EXrQcokQ0lkDpB/BV6dx9pJZJ1LLQ
0t7mVdMpnaTK1+nnK2eJ1FTeIegvvUSfexYp3JEN/p8th4Kznf+CYFXd6FuvVdc8K4e9jMrLdN2s
TAvFmGV385JpTRml4eMFsnsCLS90Av8NqHzAoEiXQTsPn3BhC4B35Bk2fR+bDs08h5TZuxVhDQd1
uCLOhyFh2TdhfnoBpV6GRLyvZNL23nsrjDA06ki3kb4jfnVqMrZC+yFLb6T/SjmTt8uMzeQP1ukI
RqdSUU8i7X3MW7KdSb/Doh5EqNP4NmLhWD5eLs/o32FNrhckQfGHIJMRLd5dhV8lVLxELm1gTtHQ
ofUC4E/SGES66Hmm5z5G1kxN8AoJT5fW9vl+2MjIZttvzlTmtscEr/GIQYa4AxsUYHa99t9nop8e
lLaKYIOOyST6L90hW+DY+jqBSagDsM5JGBlvhMVHwgefEJK/aBGbSJqXOqmtLLIXu9g9Avde7jCD
9aFA2aFOKtZGxgE0LcVzJy/LjALIMTHH6El6BIGQ4djehDbLJne5PnquSCJ3XOEyxiT7hXhUlYbM
sHhqc6PjRXjT3O7AJKm5LTOV/STKynDX8oEBi02thXFTuDkIJORfWvPmuI93yRHBKLzbaKie1Gc4
IYsLmDPcCpPdmG67K9JQlQ6zWKkDJ+GKFyiZh66gvPafzaBz1+dJhIvKjZnjdc2sz2622s36K8KY
Jxy7gAUJjWH9cClGWKR17f3rKtdYWqNPT7Vm+0Zx9gop8RyCW96vD44wZXycAm9nMdEW//IaOz61
WtErGdTY6aowp2IThcZX4z5HOmjWf4HI890eF+1oeA3TJLM2eD13UAetrRLkViz9cf5lqhEvWLmq
aMGoKE7KNqwHAcerl6/VMsxb4cAJ90ebwMl8PGiOa4mWbAQwf+kkEOGduJFIgbmIhJWWeowd9suq
HVQUsYZrAJ5iGK0aahhWfSwW33ro7ycmcJYNFSxBHRwL7EuCyk/uXvsPKgL27+7LQpWZLC4MfBQ5
9dgODBYCILrXVTHObDWZ2d9BcNzuP6+Odv2f7SrPe1KZXLH1sVN7GCdlPDTxAjdm4OSmSEHWYVNv
h1Z3U95oX3U1C7Y5mnhx7uVIk6BOKz7QRdTIR9XbqVRMW3JGryUEo/MHKeVGJop4FzNGPImw2Asr
acCca/cuzwwMjEtG9eVm5XHjHZmmy4TsxpEbem4h79j6t/nmTfZvz8h7LGtSF7nxstHrQxfNN/X0
vkXRbVId4d/WTSpvGqqH2m2dTp7T7b+Yu5N1tM9rgBPr6xojG91wQdZCzsr/bMaa77iVWEZ+12l2
iNQ5I75rUqLQxUXOWzbqYtzyeQwCkp+JIfsr9KvreFvlu8wW2nyEF/EiRB9cShgjcA283MSaJ4jv
n69LCGxA3CKfS7oGVXaouFERGFm7bjMFhmLo9Y2OR9mLFBnJGxQyfBaUzBHTouXsri9PDzMXSyXH
EPhQ7qQ+1pH+ez5UipynwAaEfuZTG5KKl8lVzfAn9H2sZXuxGb1fZdkunfGtG8EYd2eIYTuxH+Cl
UIW1sTYkD6euv3FUlmJsEENbuhW9pHtmq08xyJcR0TGDytN9HNxxTDNQgZHK23vfFBiNwuEvnQZF
ePX5wUB8JxT5S3ztWw/aeIYJlHQffP36YYmj1PIQsvo2KMFrhOyqiuqYwBmcCirHcklrQ6ZTfXwf
sUBwW0Ll/mfsAsS8zm6xnzS/N+mx+ZrMOzy7worIeitw1JWMMJroP4wJ6nkH5V/ZRLM6ISv4CTGp
xTQNY6Sh2q8OhUTuOp/aqyGYpfPNbxoNyYwnlNOYIQOcYAvc0mwGYrwL3VB1QXK1IzyblDFs1U+B
uvquQRLZD18xEa8SxRTzlt+9l9GUt+DyOOXxKDCNZ5ftDcUil12n2jqDCFZ5dlvyB1Tx/DryDjpz
5L0ykFj3A0m+qrUj9mMoMf4G4dif2j2mDTR0sHSEGEDpp15FM0mOwRgp8vtTSWM/u9DMk4AKTove
49p4vk1ZG3p9Kb06P/Co38m+K75OEPaIFmGk2iFenRZS8gCf4wAcuf+qp8wz59MiAbOtzhXkaK+W
JXjrUamlQ4JjrySev4PpKrd0BY4Pb0qbcvAax1SvEWYyQFVe8ol3hb6CXtksJ42EblXa5nrClUXz
UfaTKJDQ3iknXXXFRRq9mY2/QpTw2nUfZKoTKQkRFq0kjrEiGSCH6j/3kiwmEOsMluBngnmwk5yp
XDj5jyQzGLF0E7MHgIAJrUfIDCfcbdT0wei6/8jmLG9Fig8po3rfNNq8Mo6Of/5v4KZOW/xgLlD5
i4HdH0lWRl9fkjmjrO/53xg62PgeV6xiFvcMtjWX17o0XCM3s7WEmQTytjacA4Ph+7aXll/Sdaa/
UjxFMbzpgL8SXpfDWyQpQFzmJeGs5nRpE0f7wzWJ6UWF+U4n9oLifVazer3Pe/z30GyK5Xo4KaU/
ht9SSzGYtViPFDOZtYqoEy8kC/yhWOZ733VY8xCWtgKt/acCGsbGwjlUwAKv7XBRI5eGOXfL+Det
Y6ZXc+7NvsYdW93IGtXKD6uv5YRF6QXbaCShpkeUB5hrw9f8ryYTUEB7jOTBUWZjBTm+zFo581gy
z0PmWuxqZxlKGXohDZzBuQysdqLKrhz7TxTpSBkRd5kRXF0dG9qqOGmG0H/rAs3LZ4U+3bXVZpyD
5ChdNs/q4G2yzynMJfrENq0dBBoSfMX/SQHakUg4Fl+LfEkwiePa8wLedxZATSf2fCH6H9K3xSMC
R8lL+Qji4GESooKAQ+hfSMTVcAhuQF4rpKWY9orSuQCUvZrsHN5YKFvhF1bUrRg8rBmLdevhhDVo
Ky0n4922MdzveuHrtdULlGE2KV/cTau4bmmf5RsCnHS30tvdiL0BqkbpSzxtZO5hHklpCZDCl4et
3tBOHZ86Maqb9gjMZ/b6dpaD101M+HvMDuFWf7Na4It6D84VbQOzfme6qdmE8AXxtBhIfuOQTFuD
q++DAdYtCd6fhr4jND5aGkxzSC0sezkJZhQ7rD7Ihd46bJm50lwqRhidS6waY1mhWsFQ4W2PdCUh
v9rHHpLleH+tXmtRdU6gmTg2C4LepMEoqT4UdQ1w2fnThBzuJzXlC5QB0HxkJB1BZwJBihrYG5UB
4NqVtWSzvjrjDrl/tY3WQmR/x86Kzma5rILud5z/3u9MB5qYZkie8csWMm9yzWcNwDUBgp3zlj2c
vDBg5eqwpey+CfDov9KI6BWpLTBoMIjYc3qNAk1wSr3qu3Q2JyR2vZnT5tMQ6lpwj9d0AC9JSIGS
NjIIwzbAAsNR6Z95DKJItqI7iwYPsQgAys+NEbt/Vhfp6GpsNe91v3uoW1d0UTRAwIrKNdoXzttc
8vNQjF/fRIvFi58s1mifPW8l1LgDXOiWVLOyxqJ+RiXQo1g71CLsnuPbnevBnAJeXf50xacMihgh
YTo3GgNqOWjEFdY+XZkMmqwNhmyzAr3LexOmfu9MZFDGVEfwYe+0654HtRTviOICS8MpDgyelepw
VeIYXg0wrZVrilaawQETK/EujYvD1mGg3dgCIeBjuc37mRmOkE+c4CI8KfOXZV4SI7PjiduMnczd
oX1514XcRw2KPDpV5fg61vHKVUQjCseYRuqXvXQ4nf5V0BGNDLC0gJ6AJ6oHAF9KMKDw11eWgGTF
q8HdLrHKFXP65HV6fOQvKo7OJGyW/LtLNOnCAijWlvA8Z4zoCz6D0/2vsGqKZEJAkRzaQQgyyIeM
JVeYcC8df8DkWLvvPe/9ENjR1yqZ0VXQX5BlgMPkEToayz/ldAc5awHWlmoOYOsfViCjFxxiSBZ3
+Gees2djTu6w1Q1GwsuY5iAgNSqH8fkCobkeuYiJ+1Q4Xc/RTwq0tHtWxFbtoTY87e4jIbh39gL9
Pkh4xq6xXHce6xia4fjWC49IAkfD5zWv3n2Hn8Be2VYLILaWydP+KNIM5BoED8mVySE3IIZOXnaW
imRv93X2fdGlLDXxGy8AHxxC/7FNXEItfQZwgPu6BsifV02ni07W4MouRQnlOBAsN7G7qPOjxknZ
r0Pw11BaEuYEFD+vs770YYwlrUNGy4pG2D3BLftUongzGGGs5kcTWrI2+BZiPaaAfIqcIb0XZzb1
SesOl/Yq83sSxO3xUWvbTmAACEJJkpErL8+ZkqhgFXiE5xyK7OkfK1uWWH3LITQZiy3EsGX70IUi
MoW8w0/JxH++YcmXXsO7/4TlZvqteNs/9Dl93q0o8R/EBpka7DcDwC6j/C96vzIensYqaqfIL60u
8ddrhmW0Re7YaZ5avDyObBGhXrKGEgKJPj2pJe2PnpscPhXZ+sZIUGixdF6ekijcv7e1M2be1pAn
FOAjmDTtxusFK84NKcKYXZKkAV0DQqh5MZ7c2sPbzGDoK+JLlnuNAsQDGfDhYPuatbHxCnBuXapJ
4BolBcCiOsojFfyKd5Y5AqTFqVthznfR531HWiFJnryafzR2fOzTQRLi8T45iHOMsnAxyvWpaP25
PmXWK3tLwL8CzeUVbILb2XDN32gnndwzuPCECEMI682lv6Iffwphio3+Et66KqveFtDla9TPPgGb
KtM2+PyHZi08xwPhAigF4v+/4N9xjz3x7/fi52XVPnJB1QtN+Npa3c5eORj+N0YhIbldJORTSxOG
9sojlvhHJxK4uaxHjVgEJ2QshIkWRlQ1V/DpmILXc6+0j2XPjwZA3IZSG1Zw7DSalND2Is+DvBix
LGb599BXGcRFTsPzZ6L9Xs3R9ZfknpIQ+pwbrxPWpFr9QAbRnvlMat+YhdKAP3FzVsy89xNzfH/O
6kBkKDLeOg0b4YJ/6r8A5j48bcM6dpQl6GFRN25YhW8qboEQcKnNq+7lc8MTQXc1+M5xpydB1bJ0
VS7oqEC8SdnjRsr7Zu6u6bAVH1v9nSdJD1JGuXZTXx5O7dxSdv4yT6PrZel6r5UPlbehrUa+R9qo
Wak2Q5i8PFpl88Rhu6QSujCY2mH5JOxLPHL2LKGAw20SnkPKP8LK8vwDpeOG255vj1e5OY3P/6RO
4HEOtvYFPTeBJUlEaaMSwYLDCEZG+VAGECh/w+c9X4My4LOD++n0S1zqemapt2gTqUzVzUxkV+he
PZZ19pTlca2ZTglB7cKW2YttoRM4B/Ql9LvjLfZRFlEaeTmPafeLAT6vatK2/whqkL/qsHm4r7Ql
rT+Ksen0brtN6e4cDi7hPPRTVxygzTn+zfjH28dR7mvRUw1lkuo4oA/kKb75SMsKg88TcMXk6HDK
/BYCXeRKQPN/IZNiso2Vjv6BHsHRNngHus69MfZ3a85gKLOabnpOLZyOU9CVDF3JzaIk6YXfpM8W
J3M+dCOt6cVkjg6QB6Ggc8DCZAMkDfHO0Ly3MTMQQTooIW7hZsteaRa5kLAj5jvbgap24OZfhZ/C
58fz3gECt1AACoXW/iLKmi2zAKtLTiTRDBUHlZw7QWOQFtssOWMDz8xvCB7mX+KbNnYqXQ8g16vW
O37LR2f3ncyr88+ETKWgdncAiIsEu7VVOiWMQwc+wg57INh8iaN+o5R5hZ4NloW90RC97BvK4vWU
DIs193PayIZrvDVFsp7C2x0P4KuFPlffrMql5GbLjjuEhF8+7c0+IaFF9ErrMyybRkCUMQn03aQL
fhc9yBxm5eAom3AwE2KlPmmyChlzw0X3OGtwTLxRNoSmAs98iE2Mp+B2YboMry5YOraAZPcCexu+
+8hHcix5zELCxCIWmFyNn9weOp1ipWl8PpifAzy6/MGyhQxBgJO+F3ALCro6gkkcK+tdi5lr0/QD
oW1kydfZJwkpIwKBK/3Lj3wYcWrgVpuxFLeH6lJm5WXNYZMBDaXy+8hRPL0gX+SCHSuSbT6DU3O+
l3t3A6F3spIlPqoBMrFpRj8DGJRBSddKhmPT2YyAscQg4E4aoI+mD6FVaWFOl3ysrWTKiJSf4F3R
jaGb6HhCxs6ZtvK6F7Wg/lcGhF3b1rZIrneem15F39Ay3dDJyYiwelpA5MazexsIoP76ejTtsITC
VFjwlKleRA08fmskoa8ml06xEW3e+bCtNwzvPtSbJeJg8QPCwwlrhXUdrDDMIpvTZ88E20PD02Ls
Tp0fgkUU4bXlaWF8i9VpXlhT38tmefdOEU8a0mUfNXpvGZWsTdeqE339UquXCFq/kWuU5rAMgX9X
/y2yErbOAHsuJ7RG8INgtoy/0iJkQgXYBpntafbBqSk861fld+GKdt4lNbw3K1FEiXK9CofBawH8
7foZ8Ihp7nrw4TMSXow6EDTmUmI0oiUMT/6SbGYZ++rYOwMED6ucwluTyzgeQ+csuiIajnDCa+Ky
92EbTb8K4ePXferqt9o5oKpnPjdv26TWOsR/vzd40/sRoJPpcgqNS6eyTji2jrADrwDI2dpxZZOh
auvJz63TmO18m+YPl0TZT952QhST4vKXmiEtDN/tCIDcBDpncdl/9gHFHAx2E6at/odwMs4IMIc+
yrgPfnrO7pCB3sz0Ot6JAQ75AGQRGX3cEaH2SXfmq0km+Aep3YwndbogknxepGXu+ZftNplDjs/L
qV/m1BRGZOFa3CV6qjdyYA7q9hzS8Zol2LORDUQU3xZZkwbGJ2S/cIY1WGGNLB5JOVK5NZmExjWe
pKdzFhx255oS89VSJOM0/RD2zJUUWugq/EHcORw82EklOm8FTwUBp1Lo2ObDvUZ3/f/Vwp5jzaTB
qDqnJRN0ETBicWondCZT9g31Tf633embb049K1cwhwOhKHHyQ9ZZGf4tWhT1mmUOE8shzexUuqsQ
cdImigPp/QZLwureGNMRfBzb0P6qrhaVUv7nYzLARc80b9hzvOscKXSSM3PhX+SQRUaJG0unCP4Y
LlkBdAQqu1zPWriC0Cp1Bk8pAou/9oZJDB+tgohFsYoleel0lzY0F6ZP3k39OF/8so8maQFWVikA
kpOHxsKlMyvYRHiJjaFDpYPtFJYium+DtE4SQTkShdmrjrPvRevzhyJW7L6mRBNgBN9vTnVN5z2a
p8vZ0adRqGEaBuLtVLtP+1YTY37GOc/sxni9ztELMdzkZcWYtrZDvCSIth5YVwAXNHMlTjUJAOjK
9DTiM97KRhLikFQcN0v42gCKvl3gvo7Ah9gudxhdKxFBtU94hWAmfrbfyza9yFOA/9gZHCC4+wAe
DV6uC+ofUhhzQghYD6vz7w5KnetpGNVDp8FvKoDCeS/uQucLxVtvefq7wPK9c5izvzLZ+vJWJt9D
b9vVkE5+DplgYgN5IHSoAXoi61SxEDaQT4AWjFyCz3IPqwUvrbrTo3u4+ibP01Oo76zRTif4C5v0
DzmlizglIN4oQB/oJ4g/sZ5xsd7Pi9C8e5x3UpCKCAvyRVosR2tbx6HEQiIvuBIFt9EBffBYwtdB
vUCPZaEWKFhuJ3oMyGQ3mdVchQGSv2y/c6OSXj+RhRuNEapv37/CBqi6D1chEsKxeA/J0lc95sp/
y82uf9kSoMVtdTwHzGhLibaSlUMw/luUf55Dekz1/PWdIJd9pJSVO+RIs5FG/UZp3BlO9txfbmD4
ewa44cuyLovaow7vOAGspMLmiCIahD+2GB7zH2ay4HsLeVevCqbOAq1mfHfmX9MrE3nDXmETC7Bk
JByk40Rj4ZvyArn77d+v1bjsTtZByfdSdHxn21Jks8t0GXPRNi1EtuJRkth/hZ/iR2Quc6ERMhUe
zFcD1QGIn3vBZ6AJns+OqQQAJJk4n1TjYkj7DURnN3bnf18QlrOHLIHwWb1DYcZweUEKml8NNSD/
ISPTnXMNH9PCbRXQNc/avW51oE0i5DJtM27E6OkBy0FQ27OhVAQ/RqyLqptNC5RMPSe5jAlhZrnq
Zx/ZkIoYFkozUnec8XAeNiCLe3qApv41HdwSH4RlJDPXX7XFBFXFiCFpDlLTXhe4ewYWZOm74cir
NBxo0N8EMh7TItMBQLM5NX3lhFak2mTKpJAj/UwXUkMGZJLrmuRoMgx4J10lEF4XNmGQ/DmRGDvb
OJWzudlZhmdjHU0KjrbkyEZ6iTqCD1XIxichyREFfNxNXWPSFHb0e9D+4hjmUXhZUtpT0s3Ivwb/
SKlmWbHsKh+8iQl/+feWlgCZntGN3JLP5N8euUFACr9OKHg1VJc0pji57UbuAWCp1hyYUOXWztiN
GNeGf9pHNl0mUotuPUvhdXmdpwWSc3fY1ee1glQ4ms/ilSfxYrYi+zdCTT5SQS1Qb8+FYiNWXvyX
ORuukGkZmOXmYR9+dk+0kSmX+x4aS5aVJKrULQpLvlPQDx298/FKUGbIRfale0y1cxHunQhboRw/
6XjuXT2Nhuy0FI4+iiOhA6oFf4y4jYi+lI3m5HPMY88YS3OiHFJt9XIJjCdcg7OftOxtx/MpSjLs
XsPYzDVf3DPGMcq2nBVaN1acXpw0zCc6YlQ1o+aIDSn1zN3ddZaX/9IbhEXaItTPRKWhIUhuKUzO
4zgkTA3AwK8MDdiV0s/FO4vV+Nf0L5aabViWC79VyrWI/cVY9ICGKN7mNYYM/Gn8Ago2iDz6oSK+
YcCbzddJuzooI6B6ZgjtEMrUpfj8ey81kYAd04TNDcndVS5Io7hmyMTIzzxBd6iAaeBkI3arYn4L
/MVJtCekNn3xAy3bCrIYsRQgx8G9fT4PTGdRGWGZGH95r9V9c2ivgG2ehajfNVUeJgidRuQFB2Ow
wTkYh7hyrPbzE/NjhuXvCgs4Dauh8R7Cr80rcimPwlOfbKAS/+fREvrvQHPowxp1rvN7same/k16
4pzhZVOMgsdGkLthhFCpsRSM1wk5HcHNpDx1rzPh/mgecwSpiK+jcqXLa4BELuyNowhDmTizTvEL
bxYy9m6bm0POPzuNNbMYCo91YhybWNPT73+L7vBRzSD4rB1YTeYgHfM4bZTpuCcfQ4a8G6Jhmf8e
5z73DUvQ0PKgxBke1M23gLTpB3U0AS7fFZHsJ9gybFXO4gkxeGIuUKXDZgJULEtAuXoECGo2MWVK
JNEXhsD6XoZzEyYAQi56/12ateOey1XWxOHdWL6OqshYBnRc7vQwnnr0+E9nxOD+LstVbDqmmF4G
/kF+rCRMF5p1JayoNGM/3CiTdPt4YgRBZ2vBOUMuzhND6NKAOZlxJLaniNPWXUzNJLAtsiMvIoU2
qYkhHuMhNoB8tUFncBb/HU6Ytngs0f30txTLs2pcDvGaqPlHTTHayNZdUmgIaIaJI2KlZR4jWdN5
axIJH4QCYOJJ9/RNplIi9LjhC2Bl1CtGZvAf7hrQGViUAl+X2t20rdAa6UMrXMsQN3vczGDXBrQX
Ocos4t04koVvH2Wju6PdmiQJZwJiMan8FT71ibU8KHMBcKYqu2jI0YkcJnJGFZ8ZqRR4cgR0tIm6
NO0R/vdg5hgL/WQI1CMpweknrsPyuWkYHa2uual5FqLGP70nm3U/4WW1BYJXbe7c073Re98eJtpd
W151DCFatPH7TEfY5vGd9fhLhBO2a6ZFEqTz4bfD6ITqKzsptc/1QWvhY/5+J4oCx4F3ypjC7xp7
T/eaDPQa1kFAB22cgcxqOYMZMd/c8Dza47q158OhIscs67y5VOQAv4PW496+QNiP3ytwQYFsFCQa
CO3D9VaSRMwTij6GjC4PEDrZuAm3sEuj5NgPWpqsEDXCyoxwziCKfnzHzEHv3SCbXdKOg85mUMnD
M6+nyNggrKuUWrldsgEp9kotBjxq8xusfglZyiKV3zoVrx8jzyl2NX5COKfd2ZfGE5ngF7Iqmb+E
Mwmk2+tlrA3XtpAZL5Vsz3NF0+sYuekjN16Q+64YFpAGRJe+lEXO8y5egnQ5coaZkvIbwCt2nCxj
mbuGRkceir5WL91e2GOPjqi8OUiUE6E4rOPi8uybfBTA2bHAaCUenw3ywn8djG14nX0M54jLLRfZ
3i/U8O65zzUdm5lxP5znmRfCQlP0W8quIswovpwSTKEa1bWa1zi3EgWKIjFPjn0DFnpjbE+oqai2
YaqwIzxHWWDSt+0HiWHwkDYVLEpyN574kiIn6yEV4SrZczVGhju4eRoOkMXBgKp+AFAgDatDYEeQ
OSe0+pbkwjhHAv6UyBB5JK/CyigCHp2nTtKTZK81ZPuDuckuahIK5c6F+muJu+CbJ5SwXZZaym1a
0vhr9MIIVcpGY0TtjetpYkPNjPrkJ80jnU5S5f1IwQsNKn46WGsf4++o48aYZCnShxgDNWIEMCv4
Pe6v41Dihs4nii+xDwI6fVov2gHNm/voW3T6IfE6ZN3+gF7JIv+j9Jzl16JOuWh4xNGrnJKQ4+f3
wa9t/0rCmfBXsbWJaaG1CyciiFCAgwM+HWSPtaL8zsHxCvuoB4PPhgq0KC0V4hTt6ziA10yr4Vi9
N36TBJ9JxAsN8u6MvseIBH7GduJwrHSsvsa2b9WZBhVviJSFBYNLHtxP4FjaD9m7kWeDngINuO7t
BxkqKwKSSJg64tTssSj0TXUW+iHJvF1f2TqpRdjWlOlimL7Rtcamf3jUbmaIfsjWd9ms2Rzbjhds
dJ4+Xxds1maUDpxYFMxIz36ljSiEzaCBv3O8Xe/vDSPmqiiV3qYZ4G++RpTWDikafvQSw73mk0zd
ysGXqmYuM9STZX+TCiwYFcnU2YmiO5scf10SzRcaVefhYFLcWplUXQy2S8LQlv1rm88Gr9QBN+Sg
aqAKDJ99qiUZvG1jEWJL5DAkNkeec6iXKinzO7NLQ847Yucia8UbzW0jBSX+U5aR7/vvDCdau7rJ
jOjG/47VFt+a2ICaWkVP0AA6QnS/lnFAXvojYpmkvJfq9ri3WXaQGXhssRdijeoAAxGCAKGRU0JF
AiEx4J4T3odmOTM/4Q0wxLOTsaDoNHlWGpUqeCOdA917Z5aovFyn9040D7iJNCmcn1Iye9Cv4jux
rmWwrRP8WOKzII10HRBumBghpenCa8vR1HD+FkL2cVSMxWMs5MAbZHliK8vsm94UvKq4YMZL6UeA
UCPOdE5BjNudArtaK9/5gj1k4cJgwxL9Ec/bKyCrHWGI1RDKmTbTmzCOmFL5d50X9vPHMCdsEgQN
xVBdhrWKBQcZR9yAQ4EtrEIu0acKZ5i2Bja8inpg4FUAE9zfo8BzDTrcQ8T02YlNsxmyGMzXWn8d
IPEoBA8XAIYjVvMAtaLNFYLsEIZoXem2KpF1RnA2N4dUjAoVqoBkF6pgVOjliOlJGJXgYpjoBqoD
QOGhixEAzmnXb4vrcLGbQtUcLNkyBLLCvXatN8Bw1yuqR99KnasOGQa1j9SQjUphc6dMMmoXchVa
KFeMdvXgDjM7dgHbFK8HKZtA138AJjOnhm4eom3aTC8qNpgUXucvUUkKeMN4ZEivQmHNZB4fQDUU
u0XaFuMk5vDMdXum28FlksFo3SeuLG6XFgUXguogJzddqCcB3DhXJNe0PNnOuw9hCcy9OI+Nmd2E
XLf1mnYxc9e/wPEwkktBFaafQRB+JR3JixChmLDgCnLCucbpPY7uG911JUSAJYQMGbdK3PPIJut7
CFBUl/SbB//RsCRmRsJV/c+YLRdxxTq/OFbYSkgHo7rJNrHd95b8bl4Le2NFQui33ncsQHcj4POL
m69QfBZ1leiTHUaKYHOR+Os35UmMBytAR9lwxS/sB+OAkcokk/3TLhojt5tfb6KkTbl4/uVC2y02
1m/qQ8JGC6pZwAFk+gBPf7O3NUDSmZIVHFzKwdo8RoU7uKs8Q3tas6qfwQ6jW9naCYVRshzfwMXv
oGp2PPgAOM0ZZ5C+h2ioGHkeLFwyI1O5H2R7Pz9yDORixyIv93pl8zCmWpu0Dd9OYXuW1BixLQg0
tudN3R29APR8X3riDZdC2/E5pzWb6hMhhCfrY6i6ev0zqK6ZDJI22iNisoGPANTPgHHpbOc/JGZJ
44WiceaEoZyVo7lm9iNTJm6dEiTPnc3yMcNea07YoO/swUieSq8MgnGa/9TetABVchVcN275/AOf
/N2RL9YK08kBWl2lIU1A3EhwPASYAlSoMbdUY4eRihjGW7SeX/PD63bSYPRfICFz9i2FI5piFceg
n0KOm9Cu56r+6V5g5PvpI4USpSAskFI+ThAF4JgNWGQ0X3/QdgVzLz9ikc93xbAlbbiKqorc9Mie
rA8cCk9jXuRqBa0wBOXDsxMQRHA7SwTBES1B4GvZq2YF70okjFZlCE4celKKg+CIHlwRxdCYT0Eh
VmOw+AYFXAJrAjOz+A6PT22OEZDtlhha19NfuShw7zR5q93FflMegE04J89jF6mbOckIPU/FpbAn
jzfL/DnOgMqnVNi6wOBkC1gnTYxsY8dnhuK2QCSNAxdLlaB7DE2lgIFfF37n+SmMUkAIaAXM6Vot
eWCTvkhpQTUCUHmAWzkQgbwHlhATF408Ap7jQPeKSb5BVQxAmGrKmI8oz5zwIN/WzPJcYn3Z9yhr
056l3X3hkVgdvGEuSODfDA5l+nqne0gb5ZEliP0T19lDg9CKOuEW+xWNdKyHLalbh9fYRAdiuEj3
fYalwVnxnOBCfSxgImU3Abii16GHQfFQdjnxMheD+xSHOUMSNmhghTgXBX5yBqzxpUtLFhrxpOaS
s3Pyd8zpbP0R+8y3MGWulWqlffjvCQ7x9h8Q2dEY5R70LF9eXJ1O7+0ov9t8JFsTRpays0W8CK5x
8OI31pnHGGOzo1j3Yo/M/VIftT+jJVp8/h0DVn4B8GCjO7TXwSTgT7w9J/xPmyK/SU099oYoZmDK
KxcrfsSHHJzmUG98b53tBbiTye4TUHigy+NcMZQyEmj02khYCnRJZ7NeYJmmvIwzyGI1HyTZSXhl
vrCVo8Vz86YHmD0PT0XrieYoj6kH2d6/WQHMMlNLPKEyC+IvXZ0n8Hd76Hxh2+ZhLcd87yXrHirt
ZAgDE8fnbPLxmKAOAjs52pSypHRQPK0NAFv24x8tmjuaEysLwQQSlOt/UzO62ab1smj4c45NWqh3
Q83orXZyzJx/eUHgeGKSHeXLYyrK7vDvEbWR14OAuqUYlnccW8BqxYx5i5o4CGlchESDGmoXiId/
DG1s6xfry1NRGfipCIUZBwWIMm/9lONnH9ZYQ5pXZfCgYOedzP/GDbLARIZyrgOximnFc5AeBPbD
CLznxjzfC+OY2NOLTaLPRQmhvRE92IswbgKGz88D21esincE/9zVgR0shJ4q0fSZAaZzQQ+p0DzQ
j1ARFUD9fdUQW/CYIPFShIXbBul3BIJk8GDaxY+LsTdIhk60sIvfRR+6iYwau+qHS3wO2xI/i90n
+SuUdRKGY9YWuTBaRnr1WXtJe2vk+tDGzD/gTtxi+jXpUwxqeBR/YOpaLduVtCIT6oWdZ5Q6LYHb
qtA40raifL7K/QMjNmyNtZkkGDSWxKXVu+xVV3o4x4ad7s/xMzEZ+mngeyFxs0TQzUiKrFu6rO8I
gTETNAwlwLqZKbD+ONyGXcOL7OpH8zWQsFk9wvtx2qk/Ki2GvsjAoYAnEx3O0lNrVFU8pAyA9Hoq
wZKN0D0GbGPo+yGo265TqyqenvqGyHZqJ8a9PuGH1qf8QaFbn1p6pr8Dovotz8JamMf5yl8GW3A+
wDaBKf8UW8yS0bYz/n2NviBVZi6z9d6qCTZ8HA+DiDsCK7vP+DygpT4atgQh6/CFMyR9Psop6T7b
sg/CXGVXLfGZ6hX+OfllhaSiWgS+ydreRF5uFvlqG7X70Xo68EKZkFsPepFj22rhhfhCxzNliACz
sw/UIU/20b5q/LyjQ7LdMBoV94j6AI3I+Ptx/4TvAZMI9f1vQ3u5OuevWFcKzwoahOG6YrgEKXMF
47jHSMTzzV0FjTuVAPaTGUG+NOuZXx3B6gZYjJ/vDaci9LDRTlCNrVEHI99yTCWlZ6CpKdSZkA6e
4zNyQk6fUfOZPYEskESgOXylmcKPQ+1T5dewCs6P3rPNLpDfC1wZAV/3yiNGCQkQiRPX889ywu3l
NLcTMC4wKfqNQOzIbBcclbtcdPZbsMWOQLgoMnsnIL/L+Pw7phS6zcGnFyNWWFfMlCDCjUnDqIXQ
VgXgtmJ1wY+B/09hXaVvPxddUD92DeZIiz2lAfYM0W5tPeMIbc6bszAfx6StRIgF3HU1Mk82Jvyc
lYakeOtoh1WddNsIpLKH/lGX3ICGH8PcULD2Ld+OJMelvUzbVr1Mj6tjRHxT/Tv52OGJogzlpwGe
Lp8J0x9Tzzd9fJDZB6TtRTjoUBHtLAruESvvirkClwUCtYywxlu8wHtGsjd+77KncT2SYbU5oeYJ
NwoFVD4tNKvIOuko/FPcBIPfj3ErVrcWesGEWX929QSL68PNK9OwUg/4QmMFQrLwdYM1TbpLIa52
d6xgSj2y/A58TsfaAIXrqw7JPR3Fs9CuZNfkOx+B2PhuW8PuCNy5zs/p18yhUbhTzE5bAgfONg0z
c/E9qR7yg7EJ9LT1JRNTCA6IvJP3dw+IgRPVcLNskZMO6XyVNDYbQDcdSAzyx4z//Ua7nbdormor
KsSRXeOmJzepsaYgcf7pGDVtf/ES/6LA2O9kLT45UBAO6S1S/In6mMg6VXz/enQ4l8K1hRdBDmzw
Fo8FQPDwwHrbRwVN7BHR3CA4QiWH82YTftffHqSNxGDk+4L0+TWnlKmC0euxzSOK2Pnl2+eozcbR
PF2X5nM2ABd6TQ7G4oo5qZNWG96N5kx17aL2EdXZXpdkHJpxKTPB2xvh44J7WgswmkNmGeAt6f7A
L2SzIw5fiyAWmHpiDz07EupV1f7ZBGEl6fa5Pu4p+it14XNMU07hr7cwvfB6rEyDMzYMnGlCwWHz
oDUULnOghhgMNolOe3FjCDbq7kkNSPg8Zn0R/IwlMmhJQb9qNKrtWhrLP8uGhSCOdteoy9QvN4pe
vSthP4hDYdiGKkIsHlHaQC5dLMP6PDqxhAINuSawSWOdNrfzwXSx6ctapTn9KB5C7xE51jmHQ2X7
RyRlge6Y6Utv+hy9Pwbrnk19qm82sUbv/H0stDvgV6QFG1su0bmDfejjYQN+N940/f438TjsKB7G
U/eH1h5qOSf7oRVJcKOI8vyGXIhVhfRFQ7m/rrD5c04E2bsbudOUGHls5G+x4d8YnZ033IcJjlyi
nfNlRF15BoY+kN2BKs1sYikfnf0lk/+wnzX8PLm94V0m4WJW29bOM02HjRdjYSDXX6TkS9wXfA5l
1NEFSp7s+AtN47NP3nhWqfkZG+K6vXx9qf87/PLO2dUOJND82TKu0Nn6q7AjCpt4dU2fwVw1WqLN
fbGqh0gNqRsY4i44SkBEUnaY6bWdPXvEchwGpXCBcEXAXMqjXNdp8VPb+j/NnrckcTiUSxATaW04
MbfQ2SfurnO4tl1GwPr5gtngFoBM+PTE/YmEd2dvJi+F6IYx2RpavoriGqqHnj7j3glpKZ22bDUf
roRQdBF48fXj3hUiYPCPgjvSvVBqSwvXh9irqx6g8WTvaaQ5sVbex68zNxgnF3SPFqRGo8/Hw73l
HupnE80YFP82AB9LwP+f4AWEU9jrNl0AEerbVT78csiY0jkRyWfQXFmxaGQzd8l/ak7SiyEGbOMk
7tJg56p29RcmsEpOsOVyp0txP9FBzVOeG/TzEBYIC1i+d6kEHsc9iwNBsaVrYB7YAIsSNwDeSVSs
aXwZV/426iOCz51ggqzpTep35qR/4xryG6Q4iHRqKaSutdFgIALz0vRbnxAhH3jiVhJ8rvy/n5+o
IC6Y/cVSMlYLQkY1a9R5Qbak8ealbtDxVK/yNAR34SPcffkF0AZuWfhEG0QsolwFkiT9Z79Nuhlt
4YwLYGsOmiSIMchE8G+EKH9iSU5ZdR9HbU3Y3iiaYNKM4wXeb7A3v091VWNF/Qq6jpvJp5lBICMs
KnYmxxvGc79T64ujWYZ4a9m5++u3M04lMIZ9m5mYLnchrH48EuvVOCkD71XJpEHA/9Jr45PoyZBs
O1no2xZt93Vj8WwZuGaeIS4ScrmqMxV5TCsLWr0uSsQrl7zrskOEgZ5Hnc5nSQ5vUzjg4YHA8kPY
WBiXWjawPrNm2CL5Rc3D5Gd8pIv876iFxQkN8bTF39e67oM5ilDtWHDfU4HJ2xtSfxzPqUKSwkKJ
i/X83vmUhR54xdzsSnMzNpIjAdXm76koUAKALZDfNehTrcIfB8wwee1UfWzB+4xTM10H7dHIbhQV
Fgd+QrBj9KSAP8QB7aXsV5t+Ld1l+8439JHU2DjfrkRbjXyZNdDcHeHu49QovNe0uwrG0bl3nbaf
yEJq2Hm0DeE4B65me8tWbqY71eIKSy7IzOifYeoMU47jMj74+mCnvaR+fvzKSNc6jYg6UDFjcOc7
biUUXfdFR4UpDUzExwXg7qxI5o+WdjoaZW+P2iCvQmciRWHs81ZOwgOFgcQO3fZ+MLUUvPLkZA7V
sjxthaGi7fTBicDZ6aoE5nUf+f/hkciQrDHljUH4el7cpkBjPqumv/TrxJkr+zkP+3QLU7L3nW35
d3C8MPKEZ81irbG6hvWj+xeOOcTk/HcYtEhxmjko8SfkLU7MGIsUCpHQgrkZkO6zOtMVzxpKayUb
XguYimJbX6o+B30E+rwyTRsvbPlPn5ogFX1H0sVBJIONOB3KEdy6bXqcbFH/UUk7eiQ1SvY3zUK4
VfVMNqb8J6osN3RIF/mgYcWj+YOVUhfqWrqi2YzROCI96Xz0VYWOWXhcS/x9hK4ZckwH1oTd1yfU
SsbViM+SnLC1ZEedc9Fgy0MPHspr4sWrtf7zctZOwYMh/7yIVsz+cvrZ+0pEt43R1KGnZs4qvQJY
naYuuAU7XxJy03NN/iAhArURcyi0o3XXfofoGA7zP8iDNsw3V7C3l8KElb5JyqP7jtpyIZDOj9rP
/LfsEdm5m+fK3dHpN6b3wYFJa716qkQ6LhV/MJ5rCqKGVYygiNYtB48yCAh/hVv5pdcyZv0CVmlA
D9UyHnbKBSxDuj6sc95QAboHipFhS26KNakVpRvO2PJyPPHhMs4lmuaMXY7Y3f66b9lI6vAk2V3Q
RhUXlLDU71yWvO8Vtbzw5gYKShxpruNXl4mmYjwRb7e4bpxJSkc0E7xB9IfZTnVkPyaHtPb9HjQs
pQtD6TvSPPwyf2G8viCzAv12CLix1dVzaU5xlylRD40TkZXoh9RYPjhPHEhgmfJCnxoNtonSMav9
KFaDEiExdSzKPVipNd3jyydwMR3CBK80qMEWll6b0pFCg3CmRSmLVCwA80jOuV80+f+i/6oGSeGK
ldm2wT7wy7bI16PjmVoPXDgCgvczxS7UXvNPWr2VORHWfCjpTFGAHgGcs8MEafA7WVGMdyU2bq4S
jwyGSQdG63OmyBT4ndSzLW+7yRmqtE3FpWwEnyUmrq7sjsL7zjiPn3KFpXU5/3hKcNgEQES5W647
3u0fPPgvHpdhXY+35ZUCyp6plGsTSe5Sui64D8bJyN6JGAdv3ToCtdkC9UoIF+zf9YY6OaSwy4MM
3s2Rnxa5ANrG3SNR/lT/Ci9eGnCIuIk1LSDczHW3g6sr4jdiNJgOrYFqeSDxd5KXr7aILa79L4YU
XBSsZi37DCwVuOA3jHv6NElOhMyxcksHgxpHR+VmX0qAWqIdkhNyme43ibh3U6HElOzChif/8/dn
Vjm8tvRLjQUOF/p3J5PXhDT2AZuTUfPpNfa5Ia44D6DakQxv3tExPupFC6dcWzVEJP1UAWdp3dAO
kfYIYjDgI3UjfVJNp9dAQJ1oHPsCZMfhmepy5EQSLJvLDBDQ23acMDQcRioYUeguEHYbsZMUOk6n
Sag+6mnett6caU58dwMUwd28opydor0Yx1Z0TWXZEPNSeFKAKMNu6+azvVozr8+oo4QZ+G+yOrb1
yjeRfIWX5ymbXOuyOVi6nTV/UKRoEgP3aypMDT6bZLp9Qg6U5zpFdQgFGj6sw2a7LvGMp0G8ta1H
Sdrjpsj3ga9OXbytz1vYcLBpSJN2WsfxVjFuG5S8KZYff3Kw/1Qzsy/wI27uE5L+4e2pDLYh7A3X
lzZUcIE3eKs+WEIWKRbdcHuedNt6aPw5GBcEKSn5uMivA0G8dSTNG0lsfL0SSSaYZyRqReXsZJ3m
tkJMWG4RqzR0N3+m6AxiIqtyR+l2vpu+fk9rRgXGSLWT5xgJeG6ce9VuNqBwWyUbT/PSlziI7vnT
Ur2LMaLIhwHxPQqGv+XwmioBepiLGW3uZ9VUUqbvWGBiTJ3/TYFdECuEq3HAl8DFasTvksbtgQrX
UleX26u8PnD8sIK0OE0KI7T4CYYxBpFV9nDSxcSD2bxRctUUl7Ocza6uHUV2QWD4/MTE1bjc0ec5
shFKosgWnMI93ulFNcf6YptdRYEvdQjoPjwwr6DP5zHUGUQJMy5ljXR7Q4lHIgHCzvj4RKuJOChn
OVumXwUV6obJEyZhKS6g1N25k1MRPKtdF59Cigr520us/CwkXzr5WO3b1UXmRdbhptafmhJcY+pI
1RI8rYXJIoIS9Q1S7lec2FV9DjG4g9z4q99zCZaYHVRVtUNqSyimmUVRwMAuyEwqgtoKi368i/Jx
hEqQgONtxqMPBt/iS+hZ/b8kRT6t+DbAUUJUOMGOgXl987eYM3r+oFTUuRVWi+VGJll3I0VNOVcs
DJpDPoZaJYWL9c8OkRMN4qEtbG7NZUTOjHbPhD4u+RUNVO31Xd/wWM3D21C84jTkjBrFGY5wUZv3
AlsdFVmtOYPG439CMNFJ3d5ulnMsFThvY+5XLmNu/uExZG/UBlKknxbEQJ2WzcyBB8vpZ1rHDd8w
03i+9Y534y4oJbiv3qfn9Wx2888DhxFMZQLg/PjATlyLQ8K6FeDxDsnRv3uxrnqvbbPjHX8y/EeT
ZZ7WceDs/Eru8R0VOxWnU3Ixd6qYVinlW55IfUlvheU8QfIaGNq0UqPztta3rah4TCW1HNXHfiS8
YGPn2eRyiY9ux2o3QIeQ1/kNi2g27uE9AV1Dw9YbMU0PLoL9P0dW4KSBAKWujUwHRB4P7CobHipL
7ItL3vrnBWbA5ulKABlXDWy70n8jzqCs88RKwa2c5PgfhZjV84xWZQcVlyEhIHWNqNFskOTsf/nh
Y1XdwkwdJrP9lzfkg+SMOB1ycZFhNOe1MYpMSU7mJo8c8xXMZ2EHfBy3IgE1wY7m8OazWxkyEFo7
YjdkNSojSitKFEH348VjF0mzFoQTbaNKZFB6oFa5iBLjSWJmixrpD/75MhGEvAYq3lVfHvFobOMK
qbvSuz2kVHRXfdAdapne2gH6d+CDSFm2pKW00S603ctfGGhG2tiOBLayVcWVRrWg6suEfIHHHAqO
jrUjI0/VlZDG/Mfxe3wo9pmK3a4uSwM+pdTFGVWgfhzJBDp0L+GNduXZrtWe9hnHtClcnc1RWSDu
GYVh/kmPgYzNo0kElGXDfkhKbd+OpSsqH+PKoTLHrbCFdlknIxlwpQNBrLJwk6UKQyAKzWm8USKR
mQwez2/WIgvKlC63FzK5lcBERFMGVx0KhzV8tkvUMaCkFpVzwZATyS/8XiObnQpABwKlygILy0Pw
Yfcc6TzzQDVAVuixIF6rc5zSBxQzNuQUNnaFqpZkThV2+4lqHBH3fFqFvl7D37bVGeNUSmbbPQAN
jK0If9FBH/rLIri+6uxEW6IOGDFtrQ34znXeZ4Jsptkj+xyKli7iyQPjmlIqOP7kPFBHa0LVWWY0
1qnkE8FlkWCyNwGDZSqknszILe+LtcKtOgC5sxoh8Uu8xrX5XSFgdt9nMCVkOzV5C/r7cRHEkolx
VjbIZkX8xww0NsrAsdnMT+JwRJPCWnlgBMeo7qpmaozdk+qWJ0LHVFddczfswmCGZzWsAS0oMGdr
+JAdBRdnWvBmJ9A3uwYZ8luj7jrpRYYT/0Ek3LNpK/pFQ7QK4mlH8falQ8FI0Tes3XkTbX7H3cNG
GxhWkho4AUqgcxtQElK5qytp8DMIrDyQ1WIyHIegot+3L8OLNDo/P5g+dQMD0OLhIjWNStvBptY7
H5pzlILJqBCkhxhfgyT4+VbrKnXWc9WCSxfBsp0eGtsN8TavSxhoJZkJf/2toAJxDNuR5BHVsjIt
UfIuCTO/8MQDTMJ/KgP0jtImKsXipoI1H6YOQPSAzITWTSY0esGtmI3+BxFxunPcL2oaXDN6eDp5
V7f+6NqRIBjBda7DJYfDsJYMEqa6+NARyKL2TehHtTWrgtfU3dIQ3fdjFUntJ82fuRK2BsipRVqH
/FWYcT7A8U2txBzdQNrlDjQ8ERJwNHIVfN4vEnEh0lsBGtqHjIgMpTSoUB/6uEzyTK1ukvmS6IIz
HIzKK6Wx+O8h8ab3GT9vPbXDc2uxrBxOee3Av+rP+JMxC3TWnxjjMLZqqIXmshGp764nZs57IGme
wndKQxJk9Q47KvOfuWwbVda76dhKnO8dImuV41g8Ob3JGzwzscADDrF2ZRonVg72qASefO1u12xx
Qf+ikMJkcH/yQ//YgaGhDrTJMdyEm+hzMqgWGsxL9YbiZo3Pl0XiXFRDcjoNtUy5vtQXVp+wXnms
9CkakmwrTpArUCbVp+zwmSHsJHb7hOFkS2d2Qptr6cwJUWhJYqoFY2V7VgR3Zwq5sUDhVGhEecXy
x7nP6Ar/qWQyxopQwMwzpWFccki2MAPhxr0YSX+V9qXNDy/Oglfv+2F3oiTQ/9IdiPVzyJcS8Zvq
nECXDdyO68A1k3/AIMXxzIzKc8cGFzY/wiK/jUic0A8ZUXO+58Bz/BHDP8VBcykGUpGghkHYXzwd
rYkhY4B1AzuHlKm7CovImm26Jtfk9c7IjHd9MtVUIy+wIZ/T88IgJIABvPEB/whDCHYtPxrlvAJj
7nc4vv3UVDY+JE6SgojOvE6ju6KQnFNfeOcz6UyhcSlriYLWYwg10+XvogqgmlYhqLZVzhW7iFwK
OkV5bD18P/zClmSWvYDpHalI/gLlKbil65+GDbmGp85lZDEKnu2sD+pwecQjp8RFe5L7ILDL+CE9
l97/PI+q6/DiNEk1bBt0D0dngKuJgrp3SVEbtyogfJ7JFlyfpwh7A5eznXy2cWucsoRm4wdCxQ0i
2ZA20Dy6BAXseWJ5SC5S4JhHjTVyc5rGdMYIcHYXVU6AoBd6yVYCjtb5k336ULI4juTbBPTzCf4t
40Cjwe1arNS8olbnCtpFSWxyFj7IMius99pT+nIyMbQr8DH7l2jgEqonpQntcF5bH8BiZ2k8UDq6
F8GpBDbVmSmqQLRNDhRnMH70UTes48W568fQ4/Bo+VF/6KXk7NyrznSNmsir9gxP7dxx6lzb8A0W
TuSz2CGVbydHbWYVFenN5VRw+LmWtik5sic065q6s7wNLAh/M3efPzhmQ1HNlhFp6RWV0feexsmm
UE0OjJoSXTpCSPBpXRV9KNb1RI2qXHk7B48Nc5kZSs8jNE46Dh0kK1yxJ+f5IvCfIpfLmC3vVaHO
Lv5ofo8cWe6w/jOFvG7Z6kiOKvn6HAR9QlrKRG/ZDvVi7F7V4Bp4vFtDrrC3CPK7VX5/Zpnwkl3W
qFIsw6T+yfA1bV1udLGxMAOFBhDD4xkJP20pBxPahgMZoJ+JPlin5bRjOQr57f6hUJTM/6sDp0BM
cdLe7fsWXWby+yihEFIl+oBMFHrUdH+yO7+8QiOFgzyxluEuP5qsnUbWpRqK1v7NpuRP5CBmtgHY
HO+p5dlshXc40XNOqkDyGQ5p7kExHVPUXjuKW4rIYPoUd0aE7GDaCVQo4pzyEyXgtTbggsqgbzMj
mvCPfvxj1XVNf4QU455hUDGiW2vxVS9gSqp690Z49XMftqh3tFDiJg2XDQ6f5aPnKDaqWMgj3VrU
bGkiTYh+RySJdMVzYFdXsbOdqmGt7bNVH+bb4zvNQD4JtOO1auhNnf7SkSHd4W7C6lv5CxyG1Qms
R+XJKYtfo7XDzJCx4Bv3Oq01D9xYPfAtt5kr3Z+mCtdQgMLfsfDO9QOY2nKIjYj9WNqR6CYBAA0n
YGteb1Vr6qfJiWWJH/jwWgjGs1GXtbO5AWgaySrDztYOPRrUGCKe44hRVhJjZSt5n9muHWH5FklU
92vg9wL3KNUSWWNgl3rgk1X0ySEc73hD9NTJgmcjOUdc6gU99OgjbiuYWg5Qt21WDXBaH4mruQRG
Yj1ymDpoInPUbmHz+08WrJh8ExmoMhmfokq4YttfwpjnUzapMI7V3aZROmS6L4ybqOxf07B9FgeB
TP/2K4O4X3AaWJx9f6sQPJMp7/z5o/WoFJt+L/Ol8FOoEkqMB4T+xy2pj83iI222HrSJnXBkZtnj
mYIBGgrRZ/qvG+uYliaLxHVoFWgsa2YH42hnUQ4KnAUa4SUoxM/fvbDE6L1+Ah6onU/4y9M3lKF0
S140Go4zXI/gJJ+4RUFvs36v5PpXTqEjGdbStttgZqL+dGVzdNvpTaGbYOCKJ67+dv4QA2vlzAnO
jFNcJo+BlZ1rQKG1bxO2aTBtzp8abpXBjYt1ESBEmOBgqRHMNFaGP5GCFo2Jn4sc3p8AAQwBr0Le
WnuLXoTohfnZh2wLf4iObfGiNU3eiKU1RE9NIMb8W8XW0YEACVi9rbFMLlcxdVzMlbOgu5IDsHK0
NrE/35cVc38OZFKupVxy5+K3cTyY6WOEpZ1TvRjpdUmCBfGz4L13V2+IVm/IPPqZSDbbZtLfLy1J
YJoOBMbL6f7rc1GnHxT3m7l4/3vA6cNe8EO4z/kl9PoqRY1ZJ3Z2B4ysgSY7ZhpyPROR4Q6zqOFV
lITx/aMPR5Yabd0ksCgm88mJBxsgs1DOn0+UD+KvnPBwgSgAYXiy8rawapvrMh3XpEhB1Wptbg+Q
lXOky/5x57HYHjIe9RVBuEwEqzALbACgE5n75XmFMUbfV4Tclu6oOzG82vUvzqQxv7xnLunAWa76
pINwJYOca+hDLrnnmAdYim+cy3oFJsPI0JScX9Vf+BJBcvCw3l+fbsRo8UHdL7D7V6bUrgc8prsM
8Zfyr+dc6CpzGp7uCVjqlk6O5SifA/Vk/IqYrUHlLtpPYgxqskmOUgH1XQbPWVDH3HD0hI+op1GQ
SvWmdNJfAPI0q5d/akGj8YS+2m+v/DE0w8edkecqIcD/p3VayG20yI6FJv7dfT/F2gGEDrRd22an
1lywxaGLAs+wPeYvgCKbt5yFqtzzhglj3tU67Lc8diuJUVHmLrf5UikaDiola4JCVCnrtyoEFdnu
OnWUdX8OKQHlLjYPP4ZXSlumtq5qZqqZgROo1+4TCFwjO+Che1FkHOhILIRmqHPbmbTAAtxAEo8E
w/QznP8qRlOdEAWQYlGl14eqgBQRYMQ/1gDJ+wgTYAedO9Ubvpi1x7jd7QapB5c74vBGZkSWNlGp
FMi5mfLnFL2sYZoLyRHKSsRLlg/dx2bJX7qnPhHEnAsmGrPCpmF398pQI4tCb5bShhldEL6gLUKY
u5i8tBM8LH2yMycDpoyR2O4nU9OmtAwm1HJaHZn3bPX46rGoAB/5mm30LesIGN2FRwZZ/Io6T1Bb
dqORgNk1dKSpgvp8gCdYRHyea7z9Znn4u/Q7YO86yvpJZN9753a83MVIB0tTiJT6JMQWB+h5u5GW
bJ5zMIpFJLDVGHFq6bpkEI+cpFX/QYIASzys57FDOf1+jts723BPw3nklgPzEYafNdft+3RoP4GE
fUOKVK5MryzXY+alXad2Baj5xA+cAz+78fes4TN0ZAhAZ5cvpQj/VOmoPT4gYrZL+kMCBzWhY+0r
4m0aQrMTaMsEwWm5utZaLdUXx7YSEI3LCFJuxvILiQViHMl3IvX2vzX52ZNK9YRoqeqP8Gk1twv2
D9AmFTmBJW4DHRSi/d1BG0gyC319rK3GUehVyqv7NY4vSHEErudWXNkbFsgSCTuqb2cXpCCc+PNx
t+g0IsWh533R9hhHacJCLwk/O+2SXJ0Z2+7vM9H+xHtpd7X2l1PPEAHYeVBnyavSWuu4r+17nqRD
A3sQKdSPIQqq+HxL/HE21ZQvbkkfLmmCVHGZ9Pfv4CJzDkFlrHJKOoEyeUzUnx+coA+MJciI4mc1
+tez4yNEvxS9tP6jlRqqIUKyVnTlzdKpfOaJvhJrpLg50T29ugQpBXJf0355j+QF/V762l/HU4OJ
rU5bJYx0qQHhr/ElgCoD+r6OIbjLxJPYfqrEvJyDjaCo/446r3h18XOUnAT77MSgpEn39sn6x/kv
J2BjcyhK+AGfBgfQpAd9yHbQoP2lT2Drnzv3bFliuUnvojNNdVz5vSSD++5h3TERy8qZQyISCqmq
y5l0O/95YSKwdq5M8BJIcndCkmS+o9Y1NKo14XTywLbSnLINsFAdhs+KuyBTzJSXIkARi0GSvskn
/ywqSCwYhESTqIRUN9k7XUSudrvLC9eA5An+iJkjWpRh/my2NbMW5cTkq2ZYkFfrbqS6h33B0BeF
l8x+8xYxkVANq20XeKXtOKnLJN513oVq8XAIHuhwPxXL+RgeqSDmmp0a2rgMm7vg+U7izfYCTQat
hFY9l0jwPgCjNF9/rSKovQRKojaLLW9MY5N5irYAih/l1WlMAMC5yGjFBVQkrRmRaHSdpZ8rYQjE
idQAIJOF1uiDKCkDc4xWN0oafhPtaXLNtNK7s//azpOSnYDfFyxTifTQEOAZqnlS1Hnx23ja3hrI
G1sJSU/72o20rQRhR9aCVXTFGDrfbvDODm9HJdNBMPTOlsl5XLeoL5DIDkeYTDcYggVKaAsvvTus
YeH43PUecpJ1RLy4XBmgR8l87RaHACt++PTPmWXl6EOVwLa9yVMg3gvQ9VQccxPSraP2mkr2el9M
84OfOXZ/Bh8vxk6DZGtVx55UzN5RAyaRiZW9gsoi1ghVLhMJGq69f1cvX5OBT4oWNYAvNGurY278
FtvZb9Tub52yOc5iBA/i1BXuV9qHtgaxi6QrHX0X6EG8IBoh3QSBt1w73a8jmQTifNNdqU+HSS36
iYSxwKYdx9hyT2h+DxhnwMuFo1KLPY4YaWM8js/VloYeXsJX+SJQnPXH5T8RN+di/jP5+ZAp70g6
bbe5rv45i4xEmdgq/6+U8U6Zg5OQThaencrqJthjI5DoBPzHj2BYc1cu2R4rBanRugy1mGzF7Ffd
HIGvyJ58jK6mOWqtkj+rSofsaDGCP3/bLk69aQP0RbRuoVHQCayHE3vsnzV+gd5geHhOSjsn8q/F
MAHUCgdQuSe1BIpyIUkHpg0NZMSmhrlym3OJiV9XdbFDREBOkTNBNLDEo3lbbcTx7MSmYFWSFZaW
bbQBfBBYfEKJVjeBaFMxUbNJKdIUrMq2KKCFmMq//o5ofdjHE0IBDdj1Wh/i7pAXNJxKhBFrtHf1
wnnGl8yYjMdYkMzwXYZ2rsmrG17JZVu4XtMrGGLrlg4PT3FZtAtVAii2cVEHvOg3X7ly6WVsvpPG
ZMtSdzbL/dH5ILAaf+tC7INIRVK/pGRAuv/JxicdbIHanIBfN593lAIuS0WeOrwGhfE0yrJn7hvU
be3MrvQ3mnAVNOm3rS9nbeZskb5IfqVBtv3tC+2vXIv+FIfVxG0+nljoOLKvgmHJppqcHg6WhHdT
EhVnka7Gj7cmcAy0o49fm2ThNgiNd59zlXl2xz+kWmsqg3DCJM9Fxo5if8ii+jkhJUIuBv7tGGJa
XaWLLbSjmTKE58WQxy4Mc2aTa/rFUsigtfp7V6pdY4am6UicPKNFnGBfrJr4orv5waPCa7oNueWc
ic4GBsLsc9BQ+xxJ8tl8parrLeFgmo+oUkzz3/Ha9Q+CHfv5iGvwnHMO3jJcEm3sGgv5QvYlJ+2c
8PrLhe56oacq5sOlMonn/8z9HN/Ckcw8jOgSF7aJ0Mn5DrVvAQghYJUUbMFacFmnaOOVyJZLtEW+
s/ZykqjTZp0B0Zn9bvAJ/eZUWUjRRwSWZ6DknRxVZqpfm21c1iqOQCTbp/mxlYSncq7ijppvkcEn
TWEle6KJJTld66rUHFTJCWlUxkRcn/c7LAdChR1Yim3TGIxufjTm3OdgGdX2nqI2YixPUd5ZIcxa
dXjxdfy6FehdM/mRZcZHezWVxYL/44B4pEMlESem7w+ImnzS6eHTCQEB7AW6cP2oXcrRNAl39nXM
Lx4WnU1YqGOccYEKOotbYBDb7IpsZwfttu4w5yz5j8/u56OaxIeXHTJB30Tr3HfOTwTBMgCW1uR6
BH1PMMk35x8rT+pSuM547pq+9NIMBrpBnrUOLZjQukKEYiqcePNKeU8lIR9DFqkkpgAurjrF+/y1
d7fzDw+NdLrfNOmrvUpYS4QxNdokDuKZQP+OuGDgdfhbGI/EBtwDBezyf3fXsmrjlNPiO6fX4o3y
EBF1MDXAtc5bnUEAlIOkdUjRtLZwRCQQ1ncb+gQVmpftgxD7m1OmDVgWhWDopcqiYBDMHlNHEVb7
VsSCt21gr0pWugl4ma7H501SUG6okRVMQU1Rn46FzeP+mll5+U3GtrjVqPiDFXEWWcJKIT8ZA+6I
Svt3eVMo19QUIgaoCXWQYeyjjTFNuWU3Lhqg83ngVNeVaZxgt83d03JJe5zcNACl/u4Q14sgjwXq
2NsELsI2HACbRU7wPmtjk20rEOzNtky3c6rKMLlNcbSAUuLds01mxvIVr3VPG6jAZKiBYZmJwo7N
gs6Oum9p7IRUunioieW9SeT4eCp74GZaEGw9QBn1D6cazx0DHJMMht9hdkz2vcTxJcNGcsbb6JvW
dl9iEv/0QXgFJH6qNecrqcCHCXWG4Y2n9wUz5MG/nvobFxgKmQXHnMATF9BpqfZDfVhxQU+1nYs/
Z0mHLpSxWd6mx8HhJzbCB15DLXdNqoDw/vcWVnF73nreYp+eM/mcrh6ikMRvwhthtYFL5d9rSRe2
OmoiEFx7IBUWYc3lzUkhET/fKv0N7f/S5mXrOIM0OuP/NivZuSSwfQm9xNNw5aQgeL/6c9M6yqjS
MEcwEjZwywRRUBA1HYwJ+haYjXO5ZLe8+q49X3Kj7/Pb/hQWc9RSzxTQrgKxvV7AtRHi8ZFVZf06
P6kXwzo+ZkjjNxw2Lh7r9tA7zUmDLzhdsWH/LCdmIjiVWF/LMbwkIWr632Bf2zmXPCSjkOLxvvoi
ZHpYYIbdzpArG1Am3GcZ/Bhi/0oecr4oJPM+hbaiUyDOWNu5UaNvSx5Lj6X3YtSADSanubwmY0+R
z99RiwrGtJ1bf8+Z8cQwQUsuZZtwuKvJdiZuhEalUh5LuePmmht93ZZukVQxErgds6LmixlqTl5W
YWPHhv8IPJPw3GUf/RI875fhYnmPUSAo4S7I8vqgDd/u64ywtSadXhhhpJ26py05U8vXrvKwL0LV
sCxoa/o7EiOctWS+vnwf0S39gHuMXiLKmprLQbWlYaitFh81BM123cfJTHdmuIUHAnIDj8HRXSIX
CApfDAnWRalyo9yE1sLx96cKW1YerG6vONFVlRpZgLK7BsyI3MeRtECyiDCn0wC3RuBaZm35TFUD
oF8u50Ceea4Xxhq+CWS6NTyuNO9BGxvDWvvqNUVmxL0yhqTMy+P04xc2tdHai7zqGn702IR8okEC
iZDzSHsc/Zlx680zV8SVs0ZXtpjR5h5XWHMlJBMg9T5FtXTQWn2rF2j/SXW5pKy4GwP4FaRUvAVt
hQvGwJn6mcUIjdV8iDicWa5YpiL3vcUMkNGw8XxDbq1K5MxNS4RnoMnwmYXkAncyFQOGx9809eIQ
T83NAfv1ZQnM8q5WgMrycYS4v3LbcQbAG264U6B2OfKPqCwahiIjpFC2iUYr5uTcuxC38wc/y8y5
bwdDBS5I978pMX1HFlZjk+asZSGXpfTEExGZckVIrxMp37S6g8VhnEBTh32zf9UPe+qBXe3YOeYg
TZ/fyvQhndhwgZ9Ev8yNgJagg0wn9KBtosUEQO4DNtzgWEoDafwvh1L+pk8Qe78W+LuUTD2s+b4w
3SCZeEAn932CxSpp0rytu95AGEtLBLN5raJbMT7HS6TuTXFiFtds11675TOuPHVV1yjZyhyUbeTo
sF8DfmpYSN0CJ2kTba5bpWhtVSDKnJHtDKFlxHdq1pV2v1aasdYJIU84i6RFStrKhqOW1VNACH8S
xYmA5r3005+I0pqq3c6N6l7pB+MrVQ8FEG+63Sl3/U7RgYZNrk913orB+yzscleCMM/J/ybwkPYG
Ti0bXpzuTE2QEmN5JbaB7SYjmzax/3MFCmLVAyc12KsQhGVgcmMaY7MAazG5dlgH7O7zZ1LoinOP
a0qa7IBCpv9j1IqXe54VKMIon06jXD93LjGMQ6ytPvz7xAjTasdLq5zxX8suJ9LweF5CGxCsF2FG
+E9N8WxbEIzhem2ejojG/Ct3MI6b9s13mgl2nYSDv4kYporKCcAuqbvthw1p4cyGIOngTlwd89B1
deRyBl63wZDtxWIEJL6BAZnY8IUagevQVlfXaKZUoSa6nkrM2O4X65lEQjPlvGNdBCs9QIXE6gpx
dSG1FyHexDgXHxfdZp636MoVOrg4vh9AbAUVmrHHmkhy3CA+pqEHx0E+n6l++n5yQt1EDB6ZeTBF
8BhR2Jy7BQOfuKmQRw45Ja52pCV3slYURDfeRnBNWZUa2hccPl5hqdh2u/mXs/N93yPAXdP8hUXX
GXbBmcVPUYqhuq8WcJ6X0u3BtqxSiyqGuc8f8KLz0qUB+tmd2n5QPM+i9JEQpuXnJovmfdHI8nLW
YJrDNGvUT6mxs3wjMW3U2n2vGxywodaNVD/MqmeCUfdIYpw/OI5CLBU2NWBZILvLEO86OuQ4gGJO
+K6iGDeJ+uPpJEHPANBUmoALm/H6l0HB24q4U6q0WsIJhjr7ZYvwrQHOZxJNtccD+UkFT+FiAu8v
PexkLfrl2RCWbq9A3LgeTNGd0zFc94MvgwNI4kSa3uZpPX+bMss/izlCqX2GXoZedq0mgljx4ZAx
3d4YL1klQSLUMfC6b80w5RPYGzyHGwCynJmUWcRmLjeR9tvRqBwa0bqNnPVLxEnp+uFo4BgnfnLI
8Bo0WRwkV14P5WXLdx2L3fuarzcTAUVom5E4t7LxXpZgoT8OVf0jDIELdoTd+GEj4zhFJhvyPDkc
/kEhjZf/r6snS5ZwokrLMakLMt0be3ra7qKHY9Ey4KOyTL0cGZcHuzbGvBjb90m+3v4LbHHFFVya
muQO33VwFV1ngtD0W1ooUL7sf4QuXLX/6yl1pZLUj+QrYGjMMd+k3+WsOUvWsPEafIwQV4jQ+Snr
qHVCP+BtEW0w0HrZZtnGxdmh1gg33LAn2Pii5+E1GWU4+TqP7o0kekwZWL4iY7pllPNIzhrhSBGr
bqukHIg4cBvzedswtUZWbBug2N+rrnySkNjgdak9Pgj6XzW8XvvMvJZuvjp6XdijNkIgiZl+oufg
4mAa8tA4nfnCTNK/NtDUXTNd+sE1Bshqam970qX/XBIc1vhG5xQk2yaBHHv9nPvYqaT41ZYOqTmL
AI0Re9ZT9+/6dmiZgRttYKwdvlc4BUXPJbEgxZMDpl07YdlK6ety6GVxZblZlkGOXb/uY0/5RdiK
TaivbEiJ9uqeA9C0dY5YM7y8gXVu1EOMCw3P4wql/gitopwVxR+cRozK9cH+l0XTOluH962ckJCa
n+N+AwZL0uubbm3FuxTB14k8CTR7u87PHrxs/+vXdeQeJs/AhRlsproN2iuJ7iNqvTcOSSMizRz7
nPVNvMlJGaKOBdJMicOq6h3GnpxgmBmePoLEx8QjZ9TDFlbrbj1KvmAhJVtijJWr3K62I/ucZ9Im
+EhezxQp2cF8NO/C7KjxwKJDeyTfMuZg01Mw6vszEr6WL70iw6j6uoDcvf8eT4ESYurZc6M5KpcV
EbByl5I12VXO5LVavkZg++XeSzQTX5QTWJ1aXcGcvcaW8WyUFPi64x+Xs2ad1sZQ2hz/wdIywwpT
tlhrpAer1m+oNyvbH8an4EzLkgo9OqJwfrAnOv530QoHvdDcky1vw0CFFu7nbToofwwA7/j8D1vl
cIortZ1xQ3xZp3i+hJ/BIyzA1DQinCl9RY8AiiRfIa6SH7QRhKt7V2G0pGaCBoT2ypmL1l3rBHK4
ZXPQDvuBhK93eOcy2E+9aqCjSk08KEg3WkuUhq9MTXzVkV0nl7TrrbwaQPoyrEeGFVoMdrx3eDWq
mTlWvMGp/LSnBN4sMqtQiR9auTxp3H2yA2TLCljv65QzfLHYJJvYVm2/c0qkjT6gkLFtx20B99HW
61TU2dcBj+Vshr1RpvUw8AvPR18LpTU9ppjLcz0EpzXukdO8FBtF7e9FJ15Nxex11/2ER3b3jYn2
yK+HnBkZOi9OLQSFNMlk06EHojV9I6b0Q0cu0Q7pPQQBGkroSJBLPPrbOAQktvRRZ6209F9tIzoi
o/PjdgN81K06eAEhCv8fNcLXNY3PMgylfKB6QftwWtsj5+KqnCHrZ0rh1CRbPRDsYbiuZYEs3Pp0
M4UFQJxgZshD6Z/ofbGtUmnTY6NdFFqP+9cq+m3sOiVH11G58e7/O/v/5nloQuNihph3/5cBgIJK
sKUC+vrJoKbc88l3XbgXz9V/PSlJIpZIiuK7Nhxx71iJtHruClZbnSNBxdStsVCpSzPPovmXQBe7
FZ+Duu/BoDT1mr+pnPzf4hdIy/XNek8DJaHkLJXPOfMwvVOIKoUGAFPnGoPRyprK1TngWj6dy0LA
d6I5QwTi6prja0UDZPWV2EMomQ6rdT3BvieRl0t88a8k8HaoMUfkYupVVN/ZZFPJk1ZYot0t9Rdx
rvLj3i0Uorgkm6c6ONinET47RqGPSvHk1EZ1A2HKzQV0Jsp9EJ6iLxKLGmbzIWye0f11jHXQtfwu
G86kIzFpks1ESRt0s/Jk1hBPhHoUXnNQI9UcbTZvVtrmSYEUbkAS2YhEWiC010o3AsHu5wQ06cmG
xOgYBHIMiKOwFS6CscgMDpE13HrfHsr4aYTm24XlR3WNA62G1C+CPhFxeNwTrpfd9BOT+GCnS0oW
zJhrVMk2Ey+AvSrKtaHNDRMEu8JuBBWG+ervy59aDRUMTQ2J8YZeuHVxqsrZJMuksP4QzwU/91Ye
GT8cGtYiRvvaf5evs8DJvcS9Vt7QYr2ceMce56xXVyFzt/dyvQKoL5+iZfWPMdA2H5B0EtCZWX5V
JHGqIBiwCakwzHbePBHWHLKW5yvQvQunfGbhjZ2DGf2R/MPT/UrIXDIyjLWCHavbv90iKpXQfOKL
mqvaI5B1vCkFMVcMGWnQSdyIvOySPVut4WqzZGWsMwvaLoZK0yHR9+36rdpmxoHTj9JRbdHcWy+w
qJ/nJHphR9boA6pU4QURqNQIxImcAJEh1PiE81s1SBK0HHH0cWYH2Hd42SKkcLu6Pl+wF67k2hOO
PDytPPsG7hU4zCJTp+9remFOrKSahHDdAi9u4aMbCHPhEjxeAqKM6hzWHlzAoD+pfJfBMYi7JcNM
TuwqWoYqMrnNsMc3PLC8DtCZXkRnMIEly0MbfuQ+kdO94Eb4F3ckhZTKaYQ0k47hUOe5HzCnpNoE
kRoQrljHd3Eq5pNUD0qVLocVVLGgxynmA224F4MrOlL5k7rVGcZmWH3d0Dwh/iRyx5PG/2dZ3p3o
oEfBXT8Z83fswa1vIA7yFi0gDSJIvFRrb17NR7dcs1duZtL6r9gKb0NPehL4w3kFz5zIs9UWA84t
+ZwVtRypjludx4QQgRxE8lvVygQQP37xtrcr6xFKa1zrlUb4godG1hUm+10dWsmvBBuc1j97FOiY
yt2uFSt3+kQGBJKQhzEhzdSJUphIuyUyAUCQW+raBAaPxVUTJLNQ21GG2RAP5rNNpYpac4FwGA8D
n9FoV5NDduF4+IkN7u5Lk4uidPkQlDPrEw2VJZQTcL09YjVWFLPgBVqF2dqU/eY30gl+o8ySmEqo
Nx+UbelIm1ykeVmIao4DEetIBv1bAc0FxzrW7ZaFw9NpDMCv+LpMQu2u0H0+e2a63+9GmQBOsSwL
YjPKKbtk2hGIVTCRMsatfOdbBKUqeqPzbM8sG1nWa77OL5MdX9QyHcxuOy6YCm8yZJBb8stDOw4X
f7YKonAGSh2PIN1C4Ro+QAVW8d6LfydVAIqihmk0xWW2vlOscbOepHJAXwU4y1dIpwwOf6Vcx2KJ
dM5I4RMBqRc42v5xxBCKqvtE3jZkjJLrtVtjC2dEuvseIGiiHNLBnnmoihItx/cPQoNhcsp9H1uz
zU3Za9TnoPJANQcys5dI+FUZ231uukqbh+DtdOq3drBe2RPY+rG/LUoRGX00nVoI+vuxTAY5hhO4
Ar1Fps2qu5hMDelpKeSszyHCL2HySeXLutUS6/77y4V4PTUM7DFt3jvi7vI9MgVZeqUxqBByO//j
liII6+vCjpTGXTkaKvTYKiZf69docFVVENaUaGoDSL7fg9TBraXuuANzoEcv999X/6124uUuO3Ve
bfQ9eyEzDd8fQgJUVe5ZyKY8qx++CmILPQ/08J2fPf6v+E0p33wsNAp1env8EUzbQTfAJvwn0aG/
mRrgsdx6yo8tGdo809cjDF17IV3ZOIeJIh147uVngYMG7T8AEYCGC1f1UCLgORhdSLUYjv31gvOg
Wx7OEzzacZ3AxfciFm76+1z+AjvKKjnNqfckHnp+y8xr3p14JMe5MA9wR9MXu5vr1nKjbRQgjqxK
ywMNRymji4PW4HRwQcNwxHRJ6oMR3/9ymBvjxpvsGcsHmVaXQUAWrKhcKcaoe1R8CXQMIUn/ynPX
zaYkHnwZLfZInKktYvARjDqZhsrixszVh6h6n3jTElx2/nEQze59GfNym1PuPBbQjatqyoVKBU6k
3ugkzp5YBfHJvDThAlKNdzrNoPYvz820g4Alfz71+40riTLmP8YUvUheeQEW5Ec5JtLpbNKWe4l3
fYwZPrrSw72Q7UozDtbrJyMaQ4vQyteko6Xk9Ye4t/pWPdJuyDYsvx528buExvsU+n4g3YrJLUfy
2zRDC0QQ47ZWS8z7hSsPdTVabP1oCZUEvERY0rGJxVnf3tLQ6/HAuVuACHYDfM6L0GitHbnFZcMl
Fnv8j6/qQyahG14E2toZPWLw9shnZyO0CDU/87mTr2VTJeAoZ2uYSsAU7uWS0a/XJxShdv2eeq4A
5RTk3j0BuDN1Joy/UT8DIyOlvL1LYF5tNpOnVEE+rg43c/qPxA6/RGs5fiCZP27D77D8puKX3fsC
Wkoi2T6ujXVEZstJzCZw9eVIGWlpxan5i0uOE1p2AtwiplN7WJrw+FpZ2yBSP+i7vxn8rpAeXWVV
3v+92RlZSpRmsFTqyCUdL7U6Ly5zDnIpZFAHSap6LD4V1DoV9WtekLtVTmPtekdL2DeiijR6O/gu
JMKd4k5hNcp3L0Q5TjfI4J1Ou/bG2P4KBSL6DuMQcXg4omcZ+Q2vTO4GGdROx2ZJ0f+u8Y2szvbt
+8Sg5NQq9Lt0QxgOal1y649iZg1/5SjpfJc628vkZ50hGPoMmOGwduqyDzaPsKHA443EDGaVLgO/
6f9xu09CABa+M9oxkg/zycbrvOgDXQAi3HfdvnsQRXOIerwHrTFxTDknfuWn8Q9uAtYZOpfgGTAS
u0+c9q0SHgEbm8HAi5rbSazCNWa7z2rzvvSbOb7aHKsXCbDOHlJb+nRfqa/3uUytBzpKXq6LXMsJ
5NB201qVIEvu38hXJOuj44LWAZo+rPptmrIiCfL5T0G9Kw9FgwLJgQO/40yB3yMFsP+uRf+bB+Zl
mYsPkvwRoMarKxwuaXmC/0bEMkY5Q2AJJC6CEc+3CthTW20pjDpLcj3mt8cZRoe1COd0cWqVQvcs
q/ekWyoem80JDhh5FZmvqBXp2Pv9TVv271KmsNpVE2YESUklsA+UlFLKTrX73LMAmG/CCtOLIeOt
K3R6wbd2wi4fqD8hLqXJnlOV618MMiOvPJ7VOwIJHieOoRZS8OuaGgkv+dRj2fHEzbvWK3nlWzWO
pdh4b/Uw8R0ebpOpNAGNzTe/GiE++909sOC873h4V8+679WTBvi9rzjM0juHk0Lt85iHurwjD52s
Op9S3NMn42Ou58KvNc/ir+jwD/B+FCRC2xP0bx5+vfnu9xq1A16DqNCGd88QvH8yEpY5zvycmO2G
Vj84jWfcMipipLhF2GusTi/GPhqZZKDMsxbPYSpcWymyeTCPD1IQPsqJhZAznhq+CS58fW5tvnvm
TXI94L1/rfwa9XwQtE38jnCwn0Zqmydw2HIWtV0yh+jYZM/7Eze1PZVWMTGaspNQHc7F8vhnBgYr
k6tsjShI3kIyl3N4GPRj62LssnVzgGjFfIm7rJ2Gc7REZ4W7Xd/2f1Wd78qwXDcYOB2qUzvTs9co
yjBuu5/vIMAFjx/rpIVZfbo/Ig0MOa49GeRmtQJSJdswmcr2YM/S4RCXn8VHNy4wXqCnsLbRfX5z
/47IoKcX/saJIAgrIVTNT2uxKTjt6gRdn1Z9RqC6SgBlr083aMKeV7AobulZUwNDiAd1FC/W38j9
lNaH12VRt7/V/jondxKlBspjPtIaGjT3ej79yE9vgzm5B+1w38543tl9WQvO8l//5kAMf7pY35h5
Ek5ylh6tsFks4zqMoxnV9ZOOTj/j17/+XQ+w5grCv/n98m/RhCFm6eIwnufT0n5ydt4JLXZplY+G
snG2Rnt8eu4u6AYXwU09Iv90DFEiFYI2A40sFMkpl5uOU1W+Bmid/TKfTVhXNpbsXktv5pFUVr+c
W3xXCp2qfSH7LGMtICUEVc2WTSpnvubaThlCrqRAvDrcL8DaqkqlxoqODkEReaRsVXXUepraJBEv
ZimXldOUDDtTty9/7y22B1T34cNmw4JO1b+dqwszT/bkFWfrkouDPTf4jPv74jRC1QTRn0bR57sD
4RvuU/LQt3Dvykdtge46hnwgGNtcfEktE6GE/x1jYGZAo9evUPqNW+l8gapCE3wXDzk1tdYFJ4eg
UMFhCaIdWmK9vc9OMgSsl/gm0uvLJ0RBPydjS9R7PV387KdXyKEss/PIshcMBNg37+0zb74LKAC4
W6C61/dWEq7CTRgX2XoTL2DoRNjvWJdbNhndtmkqgvJ6ZH23VoHa+tOnCty/WhBOdylwPGtTXKEO
UFhUQfn3XQziZjuJEtgQI1Qn6vTAx1IJ4aFBz/dNoiI8f5D5BB1bIoyIuhaZBYWDHY4bTmVvBOWv
n+R66wIjP3mKmh/Ngg8BUsz9IOaK3rF53caDteSRXhSkktQux7J1t2tXjSRkJIRVmHxY74fnABAs
gcVGkGQexWuaB0VCdO7YDibuqAe30TmvLPA0nZBEo3JlB7aOKI8PlH6KJEJjqFVPzVeTdvdLaKFE
j4XrOyWv7cYTn3QRgdMqDuJXryGzaCby0Cx579emgsBTO5BdALQ28wgl5Cz+H82HvJRY4fo2aQI4
KiVOjrpLUP3ojQcIsTy+q+bo29Xw1/9iJgpfD7VaEENvywXRUMjlhnYly12oDJt6dtRkv82oF+xX
UMJngyI3FwiYt8uOz44b6DUtjH/sIUEElAerG2cOR7q3+lzWXH2/mjZAPY+oZ6adRo7Q/2a3BAbO
yMiA9IrWT3EEEEjY9X1C8rbROM0IEpmJ/WupsZNg8lQKjgY2c+8wQI1uRS9lfGZbXsfRDjgbQp4V
W+NP3+Dc/CPXAHJGh8TZ2D7Qvpiculak27RNaHP3zUVShpkUQFKYlpA5UAckd8we/sZ17DwIt1GB
IQNNyKv4ZZhEwZGVOiFC1v9sHT1gNfzH5ur02TQhBKu6hl0aGMBL7CT8YRDg6XpcDqpLHN9JJ/AM
dIWOhDN3j+Ut+biNkQnRBOx+v9kDNT/PMtbM8rjc/2HrrYb2XlFfArLtIEBrlMIpdGm8dVqrHgps
zVxN2Pj6QpcRG0SugLKzlecalUj1j3Wi2OynIz3dTlfU1bHCmnHFhSKMCHUYDuxHknrWkDW7KLj7
HjaWqC03zFJfpmJ8yNhtuNGathKdwGoXm/vJ0HhndzzVvMj3seKTBEC2V+/mjTWk0RnTYxGOzH/5
9wRRjFpfGaMh5+jJ5DHqlmZ0cIOJ/YeVEwHCMcwPBNcvi1sCtxRnj2Lhtjt4VahEpGoMchjN07qP
t2ZHGNlFYMaN6aHbaM+eJmF5zcBNlcLxXUXGrM+4018YH+hhp/kAvNlhGEHwLqmqtWCHXrAiQOLw
kq6zoPDNK3o/KfhZrHqnESDXACgGWo3iUJnjL7mwqMXyHjZ+hVMxrLgTKUpo30j8vqId6HBfVyz1
vSyDIX3Pp9qFAs0hEYm6hvWrN9gC/KC7w1rqRgr+aLro7DKgxqM0UzuCsqnB6LoD3tqUvVEtChDi
db660pm+ZBv212hQfcGabJ0kge4wXlpGzMl93gn2BehXQipRJrg88aFZ9u8opEuX3jIMsSk4Caim
02LVaMH6hb8+Fv6f4YVYpx6xdsJasc0eHVXNk55ZISiib3+tu22ZcpGQDvaEXSAfHRXz2dTC4OBn
vRt6C2BnbgBzAcZrcA/BX8L4RzMARhQ9fK9MXxq1TiIwogaYKyMWBoYH881Vt7s/TnRujxaYkwd2
5Ygk39ZtANwGPCRUqZXfm1uB302kad7vQfYyb2Rg6xYoT1i1VR2TWe0sNdgkDtHfvQJ3pFdGL4+I
9N4RZKIH+fu1yOoA3ssGENwLMZKWNIIgDfj4Z4XwANa4VGAFT4U/OEjRYYXZIt8i1wnts1pA89ZU
COpRPmJIssE5Zc8dP5nPZ+4GH2sFKht3vMTHzPdCxjaVBq888ltZOIK6dgLd0XxUqOOXPIzCjoCb
4zBTYuTlBpq4ninTWHILbIlK0ogDmN0/uafYx5/pXuHp46izUWWn3CGiSloH36MByg6QglxEOmsO
wUoj+i5kUuJHti5LBI6VJoi34f8utF2CmfjPwzFin0b+OzzsKgtb1L08m/IoZo2wV6iwDKwmGY3l
bVVyDuOYUY5oNCw0G/9QUvWS33vGgKLmagrPnOWhd3v9yPXK3h+JHCloCcujDSfMcw3XakZQEkI7
0x/XwDJy8/KaWWnHHwHVfwlupCqr6/5T9Fn6XPruW5sVuZg9d9oMUA6VukOCG53bfPDvjL1D9DFl
0WOdqqu7JmD+K1vMImocZ6btze00ZVvuoCoeXVRBHqZXCelcaVAxH3Mv/P5akfod7XsoWfdSUC30
VxaVW+eiUTyppYGV5PbXfP0glrvD9Sqg+3kgh3Zr88+zN4nzZegCmw3zrn6OvPxmP9JrTgrlkkx1
8Ctjmlhxu+D5PaRuL4y5Cofh9KCAqru56DiulOfzPQ9b4GIa+krzxbvZzKF2BAqH1YrciwKomgcP
bGPbceIAL1+QxYFSibSH4avbV6pXk+7zZU53Mds7pyfGIVb+TXodGGTYuQdPEpsL2GSW10ZA7ru+
gE4OLFJpuHm5/qzsxWUeWEjqwvuW4MfjuN/z0RdEUYr/LGTkUMkC23XZ5EHJs6o0YJy0dxVSEWts
5KFh+AfqgxHR06w7hdrQ8CHQjJp5fa04Kf6qWHVogd9aiXjuTHLeMudHjMWxooRIR2bCigLLhgkl
JaB5Yl7bYnTYoVuMnyi6ZdO1t69M1Q5cMKrhncn6i98WjqF8rl3bmEfDURtwIUV39i/ZWpH+Ttam
250n5HwK1Mhfk2QQi1McoNCN6cgjv6xy15Ovj6lX5R219MAiyRayDLdgVGkbjesYHEPGVFaYPMaU
JfnO+fGSxXaOwGurAuPdArYnpI7hwu+o8YnJxrlEU4OFEZ8YOwYwir4+6OusxOtQGEip1uy+N3fd
PcevGwBVvNz1oVZ6pvKsaqyO8/V/gJNyuEGkn4KeVpEOJ0nnb97oM9gJ0svBMlNcPrfdlXo5RJwR
hTpyHqkmHv/xpsWcV4xdKS1EGbu0ylifxyNeAGAhzY8ctfNX2x8QgwfE3CDhSoYxAqP9A75lLSG4
aPO6Ec9E96jmgbohexK7Y4TPBwY4TBVtHcLqkY+XeN/MQ7sdeVYUUsf2I5M5daNysr7HlpzfSD3P
5JhF8WTDKHGiXFpmy+Bl1jqKxK5hQdJcHGJGZqXE2OIL/1jCOIX8/4yia/SFtlwvQ9CmQU0zMhhW
V1yaWRGYXdSFw632HwUxVvUmXLy9dRFeV1cFdRnwfiS4R/weBXj8mweaKyeHeKAmIt+YcNUXecV0
Vweb4tY53A4Xa56dUmYYHfBPq3qyaUTAJzZ53W6ix8I3BDyB+znghDy48tfFwnTGkOM3EP8rLi6f
xucMF6Y9CARW6aD586cFwRnrIkuui6b65nTkS/Bm93zlBRLl8x7QdDWkgmEPhLPOLOCFefhuRHWt
xyqQmEm3fg/zXaRlmjAQd0D9aNicoqd6KeNmh2cxMxPZi4MkHAecJxcmGVFw4pqbCL14PIrW6XmH
+4h8AAxWPPXhyhGTSBmJslJB3bcck2VyEvGECGIC1dmLnLERn+4xieruhECin7vApkzFlyTvJ+//
wJJ98Ui9Bo5Gdf4YJ3yHcBSj/iHrL67EfsgRO+I5urMLKYLWS6yatTw1VdSkCc06Fb3gzy4gIdcl
N1GVXseDl6k0fwt4YccPv0t6BK5XWRcnKNGZ+7KKYdrmSFldM2xxmTnSL2A+r4TU1u9eKoxdSnXo
nU/mBbKEdkFffjMO8okVgITdud5ZpwnS/iXjIPaaoWJKDEHSUV/LaozsLn2U+w1UAaZsS4x9J6eW
Qqt+R48Iq5+8TJFpimHNVIifFGQAHrG32ZtsTlmiooFTZSToHtn0ujUVMMtGFc80fXdKIn4L1j2+
vUhRV1QufHcA65baxJWOFvBP3b57V6yH7hS8cH8RqiMUyE4FTHta2pVUhKWv6g0yvl2UbKMfohmo
j4Os8OMpeQBI3dXa9JVuEHG91OA/pZJoMQ6tRiZ9+AjTX9oQ4bjW5Yz5CNBAeVK6sQ3LAcK9qf4B
7GIYezpJN7x8pYdKv1BoGwYb01hkLAp52b8HI+AO9E3SPB9CYlp3zTLqdgZjofac/vs8GjXJaDgp
45zBRNg1nvNilINprAWprg/F1ysXiuAKCxtMKOvcxHLx5JAa5DGOxK3M94kIn8cgiYrvzG9rM8LK
iN7awZfDHyySGBjNQv4/Vm6P00h36P5fdGxesgq492OT5M3jSy4ssMq0qZmqeq55fKqjcc60qKWU
Zjwpvm8CsBT/mJ+8YnXPIfnMzdOmAMVFyZkGkimO5p3IKPqtfEar/iAAK7kZx8isv95WCuIsYeHQ
oEca/wVkUVI+b3aBde+kEPNTlva8zR7BGIb6vo6nv6gnakNimAEBVmQafxnllK4u0opMXwqfS7G1
dJ29f//DnoeJ3ZxY41Z1h+TdrDRbEGsgHQBaWjkmD/h6Yox7lCc0VA6L38FD/GyBME15Gki11VnI
u2qmktQhSajqvq2LiNfMs3YJvDBdBIDKFL7hBhs9N9p2Gkp13kz0WrPEnlhAIS+fPUIATLu7cYKv
sF6qGRQDfzMjoDeyBJk5xN5X6HDn7yv43ivMtS+ign/Q8C3DyRLf3yJGf5MTuWelYbXPdmZgWzBR
qwbj7LvuOnTzOJBAL3RnnpJohp3/DePe1VlxBmajXCY9wN0DWbv2ugZaV97XMYzn7xrRYsMQTuHM
EFskr95OcNYQWo37Pxch3y2rc3LDYZ04fRy+89ml5EDfu4SstwrrIHQJ4Z5eYDZEMkNx+OFUC2Gk
8BQvKawJPCh2uNwAcCWlrKj2cseQdCb910X/0z3THZ6Cu2EX/LAIaTOr10SM4JfxftP/mafK0G0t
FljEe79rtgVIXpTFJIxEsfs1/GttoRsVHhkzaBBKKl3q8Kg//5vUkSkzTv166hIAO8dh4wN/kCr7
GL/5XMmLJ0Dz+JoEEsXm0Y8lFDx/gUfF4KA9GNzI3I0W2eAv5GUh2sgUntBXyNtflaoVHRDIKGEd
+/ipNp58Kb4sz4LOmBc7FFYMre4q4hFgpfIjt6njDlLAOD2UeaLlwSo9bothKXlhL04w6C0Kj3U0
hX5+/1D8SyqaYOLG8DiP/hQezkoxUrhZOFCk2R90J3GIst8ualwEpi0KYENvGD1AgrhT6AX7AYtv
kZNgSCP68ziqWcRTOu8KvukNnEfPO7pYkSDXnnlgwTgDhX+KltIr8D1WaH33GQaEyjBgJbN4q9vJ
QE75MVK5roOEtTJaBArwjGGMkTOkamBWeogObJ2DAo8p+y09yc1Rw50PkMjVUpTBK/KBcp+H/8AX
av1oHNDi61QDH2nHVz475OdnJAUdDaZAzmptTDWoM9+jxWSuUKLTBIiFEbs9+3vEEMzJ7CdsjrVF
lrjzaipuD0+j0UzDUEnYhGBKK4sT5+I1tzEfXV3jZbGFUQLKxsYKxkHUgEjuHBUzXfvByZBcM3W+
IjK/DUXtat7pcSsSq0Eoxld+86eAhuLtivmwnwtLy63FRkvZZ9UiJyJ92Gupxugnis70GB0gQcwk
fkSzN9HdaeK4FPiRKoo7m0WUdeUplEZeqaRwWDyzQNsvZhHXvlMjjmnhtF2EScByClQXiz6nhryC
ukQ5+MlOHzZVQRZkIxl9OMHNbiTei0y6g/NJ+3GcbHwGRlFQ4JZEM10mfu2BjNm6EOHx5TqSg3nx
q3fMW3B7h2IVViLKHOF9KftoR8ETcxbqG/IPFmdlXBn8WLqb0GsB+Puu1t8N6GT/xork8qGEOrXE
hNDUb0r+LLlIN94HN6/VoVnOw3FkJEIGNHNKobeXTu85qOumgV8NV29t1EVcakILrSBn8uDAYVKY
unlAy+RmRXt5nPGOLMCzoZoY0EtfXb69s34vQvWNqkHfsGH4RzQOvpXDlmRyQryIXDfI1PRB1zVG
6NQ8KnPx5e2vD/1sNHABItfnicuA5/VYP8PYj4ivdYcMdbRBZJjI5TbwNiurW2Y9xjS3KXAfGa6m
3Detm/sl7d04uo5gi9yVV7rdP6guVXsKUSgAXjOY9HSTo4zrhWJ5ZaV9YMSp8S5CBTr0UEs3kZd/
KV7CzhzxOlAr4gs4BI7ty8A1kTRelB4LZVtFfa1BFToGE0zjcXgn1z1N9mJ/1BtJ5zu5Xn4VrYMv
0mJE/IqpOuDsX5cG3XZddaZupK5uoi0w/4DnU9TmQKTm1yx8m+rajrOjWe3dBj138TY9wS2h7u/5
yxIJrYwiD4w9O+esUCtsiImuY8NNMjAd32jbOVqjyS6ljzQVSxw6ErZ76J6w9Ex/Hc0CkLJMJ6lB
1N3PyvUUUEfwQBL7ud4qWjd9yoCBhRKl8q9PLbYSFIUPHtMRbMhpG54tK3KbHChwEXctU13hAf4g
GaI4G+7Ici6Vazlijcg02LuVBYFPyhoKCbRDVU/+a4yy6mpD5yYP5q1xSM+JhByKjkWnASz6wQax
UAatNORfb7MXUj+72baGIrQDsl+KwCQEqk1+6RRFZG5fYKAn2XMOFISN+8rTXpgfTNlHsfHigfUU
3bltt4xm9oqo90gDbCqkyqhurAITfEgE6eL2HJpR2lD5I6a9R1u9nUZRTmlW4j4yCrgDOF7KopUM
KxfTLVaE1pN2XuRJDscSHgshmuNmI9KUP4PZANLRloDNJUovaWYPT4bmbBZ9bRiNNSNeIEgkZgzc
5t5Q7qUkVSAFXKUR0WASwYzuc5rRzyrG4mCI/WptHpzq63Sg9dEfTgWS2tcdKCnxvlxfk3oJDESi
vly7vzEjIlUnOhn0CaeSn9TfTaomWkMrezuzyD8yDBqGGRoY7Qs/+yYjaM2hMzP5XRVYMVFGpI7F
IwKAK7rQMGj0CdknNUARB0VuxXeELpnwBEjssIu5ftNFOJ9TZUxp/dTDuhotb7M9MB75ObT0P5GO
5V0ajWQFqg0mU2PFU5B7yCaKInxFTbJ60uv/sPlZ4FLDbbX4bhvio4LzgCgF4ekWmn9hLDhtbF/J
npdE8JTM5jwVcaj7SIvKPq4Y4d6/Qlgk2ghyROeg3kmcK4gKRj4KXqv7ROJnJyiN4ujBI5yNJ2in
h1CYyouTdhQTZ1kSebcf49fRchJU3oMRS/kPHzDfJulUPXerlX/lD/xXEpm8c4/mD4QqTUUfiess
/9A+nxQjbpJae+ccFAIAk3qPAkFV0aZL3NYfCtzH2QhQae/6zeHri1LCd4+JwCokw2nStwmmqYqQ
hqVIB1Z16lorCSzN8xUFBuVhQ+WVZLNRujDYmqIbzy6Gyk3BkDitul5f1BMn6MQOyBZAqJxf9tUQ
XJAOTYXop38J+s5EwVganaMgjITXL145iEVOmxufq5i+ZTUWwSP5xzGvyvFKQuI1kXWiEjPGvGJj
BbSzwZkK2AZBXLfqB0Pe0IHOo9vgHmHRyVE2vJpAUwLwxSH0rtr3sdHq82kxrSC4yFsCfu0ch6NK
unDf3ENvgXXzokSjCsf3ek+4/CExfv0OQGtN5ZREI+9daTWHDIHLKr9MNTtRq2byelGptRkV5TdL
fTyazmtsGZC9QCGVRnuF7/wc4ZtIBIimEO99bWyPCgwFf1gIciLYSIlhGv7aaTIDDkAX5xpAsFZM
STFRV7jIsZEIKzxacF7R75U2dnWlTm9KzzUBjBBgWftp773bGT+nEhmCQYtZ21DP8fnimG6fLVoh
P1Otu2my9wqrgaxc6UITdn6WQcobnRNanlmrjT9VKwp0eqq9Tti/iS1ZYmK/FAr1DsJJZYBwY1C1
pKv4h+1HG/C+9RT8uRUFbo92I0HXkhpXr9tK89p3YQtVdSyxs2CVeKlOrsU9ejuOJiLopLYzoMut
yQtTCi5gXv+6Ks90rNg9YfjelyOnW69HX/PH5ice49VoFIy/HoJnmVlWC+fOtC3uNPzCrYRSXt8+
6fodXd4976aOOKuBTIr8VUHx2PRzul1AYLm33wsfkSfZWTzXJrHbuWYk2xR/ccBEZTJxxtlYltPB
Q1CtS/BQhdKWH8n6A52cIYmTsRJC/BCWDKWAL9MsqbHbiq3YidEJAEuKsL3ChzyouylaUZmLZiMf
mlEKuoM9WdXV4zVUlJ3ZPb7F3Y2kokA2q1wFWXCgRmbOusK2Nk3eWDBF6gMoX6UlZcPD/EOZqtOS
t+6jTIAAdEgVmTk1lETyJho8yckgoS2oVBoRRwtv7W1iCVQb4OoWg5W91KOZceYfJBEoTmbNaklt
u/YGV6aCA1/gJ7L15TCeakRMPwi6NQkVg/OHze3+udL3aIMI3efoBcbIaFINrAlGeAU8XI4mj4RZ
66kaP9fW46T2NyZlOkRl2OSCHixm5gxD96sCggCzHK051H1NRH3FQ6pYMFZaEiaRWEK3VhB5n1t0
A55lXWvzYAuEBfvSBBN/UDwyS7yU8yYLSKSu5pEuhF7Ey9hY7lea905nYNqN+nvvwF+Bf5k3Qqus
a5alSIE5qbuake07RQr5ryYps5Qgf6dxuVEVIz8eC9nMtG66dmnmYK7pyYhQUvyUI5D4qcNcr5hf
O/r9B6Ar/HSziq4Locmna8araA4cJWtazSx7O/RfmYPy3k6eS4tXYrFYFcMkSoO/OXqWs1LlyvI9
HrmtEX9k/oNYDgfNLdSbTFyxi435M3Xi+3zDopiBazcMSeWQDxKnPPj5s6U4/OeGcUSJwq6XWj35
ZrYqyKRTwKG/uYCjWmJHJRDh6NQSq+LiUCe1lCyUC8d67N0zr9JvfZ9rdmCsxc3XOifSIKnpv8S9
hWe3AFqjZIM/95pO5fsIU/fQ3AJ1Qh3x0TjzwdWdZ1VLRNvw8eYSgns/mBbKogTEpxe9SEejlalG
42AmQzLyub/wE8F/8ere5dLjh3Rt/+mR8jY+ZrdEIcZmW+H5h9kubywWqUXKQzYIad+tyojv1eGw
xjtj+qK/btWUpQft7Uit7r/VH3PoeRmK/5+FGTlE1o/mZziCAPqDxS3tjrqpAayH78rmn8TUsu0o
hB2X+alGMKGnii9M0PR1kFQIH2OVkJL9vhqaQ5G4PkPMgLEsIAkVZhRybJxLw4x1cNJe5IQrCwaD
CMflHKtM7mmVdpM75LSYUvLiaRDuWDrE0sGZuXTBPp7ttMHVhMq6eR20Bm8ih5v/K+a2PRhmltOB
6q6CGmDLRQpXwWAYvj0lGQsPFgLgorvHjwUYvPQPavmzPht33WWklTCrfUWx8ey2Kcr8LsVSpEHZ
2MS0jqtZSiK8nWdViYQAJuTqlt6M3Gzg2VaW93InH6oD2t9SxlR1BimOXpng+3hnzt/CAuZPVLc2
eGJX1shgXVWFQ86SzAcsyh8DrjIclOyzxwjlOF5s6ydSjXP0G1z/DIfwH1VhsR1MY9M4fj+b6pPe
MpVPWNfOJ1Iyo8Msmj++7uuNhbIcyyo0hzYhmPSYo/d+7zNnlPZogZVrALsBMlNWJCw2/Ch7tK16
uO1odP5dRiL5+u8PNlp2Juwwg3Oc/OZS+4mpzcvH49S3lELgObGNnscsCjm6ACvEsW+XAZKXK8tn
89iEkOLHkWAb6r9nsjDOxrBl8dnRV3dZMzm9931iq7n/v7TFSycsOEs8iV2YRvHPL4JIujaGwnIi
DBauATXddSqFJgG4LBbOppoA0m3ov48JSYE9K9KE1l132yWO4foEDuAJNiY1l+SXnpc/K9SVB+VS
Dn+2SUcee4jUfsS99OjqhlL36zBW/QWhUSt7vDr7vcR2YqMQplVDHisqSws6sgeAnvUa5G/k23nF
pTp/UsVxv2JCfT/RvSpEyCwR5MXDm7BAwvrdm8h9hjC1yKRSdNZNwTYlItZy4kqlM2UGNbfduauO
9jmodsoPLRYt1llDfSbh5vwhxX8AMH+3k5Kxhb0mXA7ayJg3SLFoCFxizrUW509bMOonlwy/jRKj
x/uCf+7fFYOZxlAHKZ9AAZy+8uG3iFmlRAWPo2BDsCbMjsG+3K6/F2r+ytGFFkDXmcQIzi0bip2o
WELJgYoUw30iXgwhZxTWpe/ISZ0d/jFIq7Yjec0wXPzcU104XXXCRlZ9r6JgIxRBLD50DdlescXc
5oZuwVKxpRlEztE1H3Pn6DseFn2uaTg6m6+dZb3uUObrulAPR2HbKJOGhh4iTP0s7d6eYrZPiZGJ
9Iy41dpXgdSy/WLC5LDc/7uVUqfY987bYDHP2yltTg+uNXBrqoKnaXqHKStFIaAI9ZbpXIuV3E92
016QMCtsoCtHpvnhZ/7+X8dbEVStSwdm1mu3kVKXRTB7/GFMuQ13D3HAzQLVlYcWZqe66bXKCNJn
TP0u+LmBIP6y3Atw6T81W/PeiEVqtYyi1KWkx5gujZ/RJE41912kYOr5XT89XLZ3/8A1TW43cRe5
fM5sMWO966CNOpLH24L2nZqO6i1HtNjbiIc8z47NkABjX/6F0XTUWT9octU5Oi5AdDJa5up4cQe5
pZTU/wXVXQxM91bF7PAoqn17fgCzOKCF1j7xwoDvtFBLEA1Q+X4H+e0o7ptaqhxgpYaVMswl6aW6
ubHyjEFOn1G9THKvoWA3NqTkTIaasudCl3Chy3VJBxEwk/RSl0y2xSKyRgSmHIaMmIX9ML9tS7Xn
6PLYBR6oMju+4hiNml7LH7ywODrFa5+ZfuJ6gRhhlo4y6h77rQdXmyE4mhbYlpo8IymFXopdHiVv
d6teWGv34erP23ZD1QHqzb7LWI5ku9/yNVvX7Uc1RTEArJVHceYUPZucZdCrD4VvO9t3Lj9SUgbV
dXDwIMdhI0PZNsy3qRff2W+pZr1S0c/hodkRQWiaYTR/WPpc3vFH/PKeT+BLxuL2fTpCLvGaYvzF
a/xttgS4X12r6TuNz17NZ/sBBNu45KxyBu899A3zgRoZ4Z6JRWkjHw10+ZzTT+4AfA/m8zZdO2RY
FZI56vb3WlVFS+SzGLCRWqFFg4sAYGKbJdE9g1YJFvPh+4dXbc/3fJtA0RdczCTpXe698h3Fv6+b
6ehV3xjuT5Nvcrn/qe330X/zkxGL8Fn7uZfQ+MEZ78AcB3AwwxxoaFzTFS86xChChEMK0gtDcBR2
8AGAjj62gqU1eDDee0nNrXkYnnwidcQD75anlyP774lhHH3EFVgp7f7B/AAtIUipnErYXDdK6pFR
2ssLxDngqRhH39hkK3jMzZF7X6ouyzP6sXERnFblOji1IqM7sVgkkJML/2SCjtB0HZ5NbgEEkRTq
4c6yx3iE6xXtQYGQHkysNesdM1YoKaVfvMHeXgKNrLk4Ms0AmcUjcZgkSgTeW6sN3an9YZlxwg8o
BjpyJ/k2errEF8znbvca1hZxScgL3TA/ts97KiuknVs2at/fKR2YOWpBxaKfYKlT9bNUUycotaSH
3nBxWU+JzG79rfviqH+FVaw0PfOlcZA/P2wZqyjuQE/ea8fTD49z/OJQWp3nj12JoU4pcGE1vwC9
fqIqJUJ/SVJCgpUIdxE8pUyeBIzvRYo/GN+g3CmAsGukhsSsOuOoJmjPi4t+NnxfTUPn4yCgiI2r
JtKpe5xqYSvi0UnVpRXy1PZsihnErpZIhugRVNc5/J4uj2caJ04xiXM8smaXnkgxIXQlD7hnXY8R
hJiV+BrUMPvk6EXRC+dt1d0UOVqa6Uxn5cryI76xKBlJOg0jWFQ6VqT5HlqtDmBypW8lFnKViPhh
oIlzsP1n9v9COp/jHQAAvpxGboKFZwqjmsGTgnR/HppDES/9ypGZKnlIXmu1D9BiJykTS52xDtF4
q7GkpPQ/nsk7za4NsvKtw9WsiHU0OHcfumHMFe1/9/UN6V9klknPJ9Tt+KOUZWcCDDLxGThxY6VD
gOYNhozVkbhsTRoon/JSN69zApL5CISHqyAYWy3vwuOscCShQnIpImsI3xGM8N2im8AYWnXHXU4z
Qxu05ddTHL6wtOW/f2zRQmBbQWGKd0VLgBkkZaOTIKY+arot/5AaKFUhnN3GL8ws5Ure9x+QS6q1
/7l6JGiTR+7F+F264zn+xbyFruwEpLKKuGOiZ2iV/koJUGILB3L3Jk3l9k05tx50X0q8xpFRQzc9
xQz37a1Yoqhold5EVEbujaajvlcYJSjqPUdo2kwBYcYCgXCKWMBdBETVovP8tRgXIc9yhG6O1bMj
vvZASezXBYtAlAU1uV7KVfZZEGqHZtEMophEkt633ZdzYOwaoCrnGZfr/CwROyIpmI/ZMUX7sc9H
mSZ4rI4YYQGuVzsXvF3bgSF/AGCW0GM7ZCK9b8bU56CdPPeELnNdGU7Y4n+gdCmRr73pEeyMOZb+
VDFs2J3o08GE+Ok9atK1aK57GhiY8BrLhw68SG0Eol3hbzdp6t4nyI4/IneLRlw3XlAdCHG9mVEP
JRO7q1U/TdmXs6kJQ4tvahCXQnOeULboHTQgffwjp0uOV8czeiqLoMHtzPbukiC2vXnHuTPy3HSA
qIXdFgQGcwU1xJ25yF1Wjm5yq8iLmd+saPlXpu8OkyNsiGdRgAsKag9S2xRHF+PXYF0iUJPmuKL4
N1sdCV4iy/hG7eGIpR5YOjxQ3zJFMj/84JNqFNFVRFOpNzoimy17k+wWGcYzuLUaHzxqHij5Z/wy
Yir+dWXD0MZZCw+Ex/YrG842YOzVlDVSBgf4OkXK2R1YZ9YkNp83/cHJZVWQcwu18qECH6umA0Ha
VP7rOK1xQcCyWy2TtRBf7bTSM6Lhn1UIzmiIAYqswzW+vOVcjkScIMGJWZoIcxllwu65y+payMtD
Fu28WiiObEDlDf3wqoCxDypFGPZUEsW1DUBWvDjMDp+6+B5ir4xPqJQIHLnPepShKVUC7MJvWHjF
AVYhJF6CRIPXVu6m3oYmgAUJYcsOZRKqkOj4aDmccPJLQ4Z7Lc4lz2+4pOrshsatgZXaoI0Eub17
b2XCckgGzcl/uk66J152HA+1a66QN1ohNium6GFKA0rSanKnV0nDuM9DccHklT79Z2FH1RKRVh7N
BeDUMqa48uLqNAb/iRAdUC4iEGQE0f3cZR6P3Gn0p11+k8ZsjGcqAaVTkO0yomaMhDP1RJZ8DcnL
s6SyxBwL6ej8CcLbeExor6iNRffI6okdCFwJTqElIxZsTqoiIzaldHV6tTVaovVsi6RRUYTGZPqg
geye4FC2Oc9cUMmcbRoautprPTsqBFT/YB8Guwb/qSSPyyGjMZ7lddAEL5MiPCnXf+ZOGSlKsMfD
F9iek0omBJlYkd3pl1i6j0y+0XutQ6EzyXLOoHYIdMslVAG3yZ/HkbAHGh6l8mIa3CONEtFl6FTB
OkNAgQOdHHnxDV/sIRUvRJ9UWpWlhgkPQNcuw23buKi/6exfh+5rczrmxjIi8NcZRpOgfWX9TcZJ
0tj/Vta4i5WHFSZX9laDfPTNrHvwVASl30LreGlpOh4fc2VClwVB9G5bX2a2Vd8QXJ3rWei9BlNi
+xCkvCJK4Nb8jnARLVFT5iKn/kpXCdkMmpBsFXSATxAlZiM+3HOTij2Y57POHQqwVfozf3Yr+xua
1swnxcDXcnHr4QpKVeenbRnbD6kacKktScKOKx/eLI4Qk4oEe70BMh/gAlP3moMhbZR767UWHnTn
hQFfXA/Hbk7hSDOnuJhhe43QBwZsLDNm70fEytSkcY02jQZmiCVpolGFgo9qSgUhc995hDA77L+P
pTU9VZTOKa242vjrQf36+/YQjQL6GqdUder/DQrAtNVTLcdeoXdDD6QteHAAognvGtwEYGHO3R7h
cwD4b1kyxeBAdKGAvyJh2OirVFpNczHtydR0iMinNQ9VWAUfejs6Qj6BlDZuzp42Bf7cAndNE7io
F3fhU2bKTomIzKMB50+F5gyIykuE8e9TpHBOi/Dvp8DoIeInCj4psIrlObdYRhm2whiUJt8OF7zg
NQXAtrLbkYiwkcKwvz2NjCF7xzFCiS4RtgqHnX7f7QnlUdNkG56gttTEqo1FeVyBxSvIJu/x+gjA
JQ0LOIDlDDc+QK7F5JKRjJJvxkQ82frqeGyD0qS3ZPdE3ZsW3smOc1gAGXEHKEPwUSRsg1Z4VanE
fo7OTml7hGu6WLpKVbq6Ouq09MWfITiO1+EfoH3z0XmLrs7nwhD4nPbpxZEPqTyF91+Nc/Lw8ri5
Eto6rDblZ4WuWzs0ScuEG+pNfYvK7EbSSvXzbWk2SZkIUrnXQsCbwVz+uO4cvGDMgG3NR1SWrFh3
wP4on9ySMrF2Ae+qM8E2Ah5qo8plnLoTISEUV8Mm50NFFU4fIOBqtlrO+wKdt5X9+YkQd0j0IrfL
H/54UqWKcJwsnoDxR/n9BQ7Ucl7B4lPXRNLKAnb69p3SnpoQzfJboyiR396bV5FPmmbidVJv+0Cn
g6cKDoQnCBvpJr0t5bnUdSQmF707VgPuKuP5+gWqOuwwUXvAlDrTqVFReDtMaXgmIyQyj7NzHE7z
TKh4IwJEXaKpNOycNWVjYWG0RatiY7jwUc6exWEUCdaWBHdDOZsADceMZAZLbsM8ByWym8jcfjy8
DQQrkUhSdJ9T+jcNEpNj1kUnvI0BHbx+LBPAYGle38ytgiPA+3MW4DIV81xqznLG61RwhtDGMFhk
kYaWvhb/K+mQU88Cji28J4qcaV8HZph1zYTjHwebOl6XEKi9McP9oqVcVVs+Aam3SizSP5vFcIMx
ZbAfrpoiJF41J/FNOi+O2+wgy805ceIYSxKuDtDcnPw1grqUUPqK7EysvHXt2tcC+ig/a1hrGehP
ufsuBcpvuEwD+jF/IIh+DxaWO3hJPShi1kJ5PMRhUx4TtYjL11heFvIpv+BRYhFAJiRVSWdy4p1J
B6Wmoeps1gx4EkH3y8Z4fWQjw0E1iQ5l6V2CeUIdtp86+BuRAT3tY/hAd/Skle9BBlwjA4G7i/wo
QsvLvrjxmcNe2nDHpK98gBOTa8vqmUaD3Do71+jl0jWrOuUx9E0n9ZOnhna+Gk6wgNJ1SPkI4YIw
tE95M2yDNj9IHa/clk8MMnD2RO01DNlbFbKNgpNN9wlFzmMoTiHxei5tDO4QEKEQAnRIAwez5e6C
HIaKZSfmqADOttnSalEvDGziWv+yzP5aTYDuNL3PUnaPNalPp0Oej53lqVVLE/dT0q/QGT3AmGnb
QNsqKFJUXHSxpWpBstuzWC3j098CLoqzSPOY/rVjzDnyPK9ZME/H1jX5gPFNq57WN8VSGioB0cEY
DiU8yDbpsWgki85SECenYFzluYfxoavZegw2+BO0bOfJZIsxTnE67PvMlwmk1K4AIHuxE6Ypt6/v
qxzjL4zxHIfQaLOrPkt19ci/iNW7t3cj3AbFehI1cktkKJpjRobHcEsx31Rn+haUxnmN/yiWlZ8h
3wF0od+iCNqa4M7OT/0l22n1UlZsa4ntsGcLbBKiFmQDsaym23tMXbiFCk0yitbY3/VojQCLvCnz
weuN46RO3qF2bZLBKXrJbGEqUQv4iwR8t+a0m2KTthAGCC1aNimZiv2QDEB4h1rPbRi06vRkoQC5
3NJva+x3D5d1PCmLWtSayDTqQXL52+7XYJnHC85RfMZrgo8Hf4SyRsXLitEQIlZAhyq2Oy8WQ9iT
lIHblcYya4yMcdod4PSBOGut9I1ruavDzS+BUfqN1R03nm6PDRJ0vim1qWLoK7OwKnubsUYCruSR
0yEnCu9JgBF1+OU6AiQVDZGDQvyH8s5UJe4FBMOq5jS3SiNtgQiOh65j8dZkq8a2SNuVwaTC3kuv
yzZBbBwMgDnFvNB2yuSRB1sDVRdtcF/r9fUZtExwFxv6V8b4hwkFIUyV8kxVjLisMm2oNONtlEHL
oUGmcOlrwq2ak+fHTLHAqS7+6bpvz0POYmWeXH9IoEOn5LGsrXY36oRKtsUO8W5XzlmbTuHjyGwm
htLLdf1f1KIBcS5YkGqa+isnRMl/zWpY3VdCzjYcNfz8M7pPk7UL1gEfjUQdBBL6HGUlqgg1nX63
Z2YKTVLX7KGVXfYmKV/LBr6lMEQKoJCjm8+qHcr/2UCVhroo9dzGytjDAdpaMfE2F0ykEDlMBMUx
i1XWE7RfHDMCmJGx74FxIR6FSkmy+48VL1hzbXmvpKzPIA3IhBORU5j9ekmwM04sm7L4szIy0eW+
0UYgAqc2lmDT9A9fUkNu/rI7v+434kl+kOhNoFwZBweawZjhhbY05nxQOudshZlAqEMZqRMXTzj2
HqW+SgBI46GKIzo5u8qbGJZj4//wuqG+FqLZ8mJJrNom8Uw/l6PZ1WlAAKjOA2ptCfKkgkpm6jy2
fj1akh/x0WZX+vRiuJfzEkUBHwi1HyjxQ0F0dfbCpFNQQ+8RiiiOhL8msMhDAyFmLIo4LzSgkzRg
freMmqMw+wXqLhspY2eK6/IE2PiYjeS3XzXWi29Ggw3IqSLv691Cz2wfBCCrleI4jBp8kIEKoFda
an8Fif6kjZKTRytPpECQmyJ9FHQoG7uEV2CuXs6AdpZ8gJXalqk9K/UfD15ZhzqyVwr3FgxwnQPv
Y+u/OVO2Semw0vIWK4rkL7HA351qmkFOS+MV23oz3xQvolAT6Lyl4FE+XEW0U42056Fhh/yOZFmI
hbkAlP4EQKFptJAHhQnX+xJvYTvKm0FVXOy5L8E9qkwN+bQlrXZe7EE8TEOeVgC+TbYsY+3itTnB
ZkEqKPcLNVsxtFw0sWqUDVM+ODmV9bh5fmTlg5baj9Sw/o/DvrOAxXjolxNcbFk1wX8jaz1HnAOl
idjqEcTbOGS/lL6L1uDRASYEuAjAj4OUK21xfYSmf3lGXNjur/So2Lwig/oluoJkrTQMUvejFXKf
mgI3mUTWIcdQ8j3PQf92BB/hbdUHyWWCvUmjKHuIdKL+rLjFwm26RFErcGRWPppPxf3K8QCZZKaP
39Yo6SXbFbqaVUhuQ9g13UbUFt9GWcxyg3hEn62g1Ugp+RaLgXquHuaeBfAswX4E1KTPfLsYydBR
HmMjaZ3ocN+Yj2zu1VutZyjN6oMviCufouIz/tlW81j9A6EHiTpQnHZXrihW0DH6dvhBdlyIko8C
FYhHnPBSwwpATA2hK0zazcEqkjyC5QKlLbmgkhZ8pKpBmTpmVHGFzey3s5niiniNQs/lXsl/dToS
S4EWeEKCgUcU6IGiTby+FQznPSfnN6ngbV4e180AWnG51TR9aE48tMIkldUYar4mrqpt1KArOG7C
pENsAxNLvG0iJ/9uQyg8fCKsxYsYGzyIlKYQuzIs23RRquoxonQGhBIfbu9iJUgLi44WutAD87Ua
3ZWrKeOy/zGlfz2iB7ngPOsfYMUCknD/UEpUK8qoJBdgAWbX1mnjG2S4jDsi2G4Vq+IV8obciR7c
Pzd9wZ07r97k3vaC+Hou/4qEbFy+PD7HWs/lsZEeMlY2iyxxWBzh8eKU3h6j1dTsGABpTEKesizY
DFoSdc7wbjDyzAet8q7pywQr141q3Z/J+6EUG7jFoSIb8eltnxim/BkwlrBAf67D+ge5dUnT6+30
nzwpaJH19/K4B/35DQV20WremXyTj1hHLu2RZmcqB/VnMX9himnmLMOEDEQi9tQZMNBDSkRjSK+Q
bzNbLN8pkmjFkMnV+2W6RsAKeguj6T1VINms8NyjjeGf1Nq6e0Cb3oNl6aK/qRQV1vQlkEDdzQKU
+E03+0wNS/U3Kk1p8xYdQg3cXycXBRFc+CE72QTTC/xstbYrTIt7hjj1nLUa0kh2M/n7T1VE8Up5
91weMdfHsuxHjcvcPwgfecbTakqd/sIPXeoQyjxOTu0sdMOTMxnKl48m+1MhPR4GrpXhgfuqT+e2
IxOphfWj0Cd4w8UZPaEBW9DPeDj4Fp9O0YT4DttdQICwTW3nBo5XQQUEdG2aK98HIKfZJX/+jxzc
Hf3JfdYGizEXKT2iNw6oqtfnPU5fSVFOnR85myEvTiJTHxDaTQUsgtPt3WSO69RR6SAAji2yw1jw
aVr6SBVRBSP+fnTB+24xO83d83bGU9YsxX6PJjwBLLKf8jupvQQxIord6A/turrSWpPELkdN6jQU
K16XHXRpbHq/EQJlQGguwvzPb9VHdFc0eoGnT5nxmNEEMF2QjNgF7M/2oTWN4xd3oUuPSoQTqXiU
agx0gY8wbyGmONfKf4x4FqUG3DHp6kEbdmVDw6AnoBMJI0lUUWeWJUL2BNsI/dQRNn1CkiwyiViM
Wv1ESzenVOJQyoS0ZgGQSKg8iBTWfNpJmquQyU2qVhcKPl+6txQhxwSWY35f8/lR7PsQx16WsNTK
uZvtisENoUzADfi2WFdpUazLeDTSPCiyxOafkAkXU8HWY2abj4bn24wWCa53OLzeYilq2Kq77SId
shp3jpOQ0t533xCjuqwuObwvmXCHuLj7LDZ5DKtnWV/F+gEL7WP5oFPLFeVId065BmfdWQaIBHTD
pzmKcG5xEpT+Hz8djJn9KyPm73dxu2bZK8u8rlJ1urJTuPZ7hs/cqBQYzxkaqsAWGB3Ck0oS8Mtf
2bQjN+GseXCo8OT5klav/6CcTU08lZrxliiWeekRmHND65oQosvDN9REbJ4uHF/6eXU+ka1nNLVJ
noDXRcV5/ewMhRIxWdzBhDL+HfE2Z3P+JJY2A6DHS5gfCNNxTdfaQSJmt0MSADojCFd+6/5lXJrT
NfPe/EpGcKnrKFBFGeo5/wbNVWAHxiHlqqz1QceOMQnxr1/xAj+4oGkYofA/LPee/ZLK4h98mSs1
QaiN1BWKmElhXqS7Ciy7YI21Kdn2fiZoezbC2p6ba22Kbrnp94n4qKXHsa89GLz/f8nwTtdFSoQz
EISWWLUGg7Ky/Jy6/QGBOZBP40bUBXoIb0rMUWcEvJ3BwRAyOqJG3dMl53UxxiXZ7M/dh2OoVJtE
ugno2B5v6i+1C8Esx/Auh/6v20lt1E/4pW6xW6VP4oAPErXzS4qhbQsTVhx/j/mLL0Ed1Q7TzrM/
2WlRRdv+Uaj+MiAnQSHJ9orVKxhaKybrWYgTdDZZFT1m2LyZeTQKzDUmcYHgWYSJ6uvBnSz13HPO
ouQ8XpRKrcGpa01+wtcoOTQP86AiWUteWuDbBU51at3msGqAhMa+hDIY9TyprYaYQ+jqpzLf+sa7
DtDkSTxGLY18pK3Idybo3T1ZSSiXgdQGl9gKMEP/UatjpPkqmqOxSfGZhXXIjU6feAOPWiprNuQe
dcaURL6RPwzok33gfdx6DGV4uckcnRnLMFAjdTgRmFUNh7uAey/5w6JcjjjEkFa9h8vhA2urfSAB
defVWTLUjlpBGr3UmVdQNiQXfR+NACpq3EOO2/HovEyMNu5A7yOsXgS174zETPP7ZIE46QINjNCh
LcQRy05nJ0IndK2VG7LcnP1ZAvX+8I4/dl6IFFec+GzJ1jZdm6J+N9vxqdtLb9oddYFdG380FRYQ
cODhEWozCYPhiJD+2W4qHchk1aRhRZa/kCc64BvRnyudKusfQL2HCdu81qxr1PTcEvW+EZrOiTA8
mnhQY7ztWG+1s64dinG4xNHe15tOztkXRMXmJ8f4iW3osVX5OxBbMYy10Yzs8vIO1NK4SWa9xvD5
MhSi6x97pFhOSpERc6SbkEaXRj3u/ttjWZW087MO3EvQ/wnnIuaBRZ0HXh+Raocu0b5C6t6lqRa8
EGlY8EjSi16AKB77nAwOwiJnL5533tsE78KqN1iE6Bw29Eeqb8NeKB0jICZkUlHzjHv4SUUfVw7h
3ErinqHdJNwvAkniyt4q60bh1c25ApYxHvND9trPYAodxGJ5SFmsSixVEekZoFij4BljRqqeufD4
YBM1t05/skRFtwzZlgiv8yusdrsweEB0gmPlpt4pwSSBvthxJu1zjSIVpXttwfD05haV99zRfoBF
3VVfvsM4cjdaAupzGOxtgZnzMeU9Q2ft6IntspYtFaCSSlhjhOC2GFFhrGLt90SrRzXpNj1EP0L0
7uantOZviriHp46YgcPKLZtEz5xfiTPxO9kWvY1qgYlLBkEglBGliXVjvUB0YB6+SZN81TGHGmI0
oeU0oIwXag1MDj8GuWaPV/vpIq3jTW27VeCJ6NBNliQ+PUGRH0EyRUirfRmqdMDoIJ+7bItWXm2x
GYY/FKyE44/GIfcW/WQhWkTTH6Ijvs9Jdh6OUwpEbBAclJ5xHIPyY3RV5lLjsRNE6H52ivrvfdxC
3wH70jibLoUMCsNNXRp6sLDz0JLDUpggAA3qexZiXsXrp4HiinmgVJ6qyhhkOGNhNz5xZPTKvRvb
/gpqu3sYfD654WBOk7d9hN1/9BK/0Xw9yaG/Razi6hOSVYq6mv9VmYZ0P7XB55VFGoAxCeCAKJ5r
cifksH9qm6Ej2jlzGj2GBQGtPVT0hwSdrU9nbw/iyydFow/i83zakjb8MGxIvaHVGA85y8BywE0V
eDCw5dmLjrx8L9FWvE5oSt6oV0MStRp2MQfjBkKlCVahMxPphzI3i4PyV6GX1mfuwjpls5LnKbCO
SB58urlc+mD/wVB6RAq1f/3I4Wi2++qaQLH5QKkiwkh1Mc200SHTWZqr0WNTZJBJRxqA0qsQbChw
oqLJNVB3KcrgSalTImFrXyXxwIEDc2gxGWmVQzIKtJAakDvjcThhdhH1yxpyqvGz+5TYrFqWMLIf
ca8RlRoRuiYjJiLhV2Uih6kJA+u6WJ5LA0QqZrC9amqtBrwfAKHyMR/CN/U/Dn+mq9mTsKz+8VJq
VHjaIRMyzhWuz3SL2vEjET66QlKtnNm/zhMeRFltI+ehi1VsgOxtlKM3e+GiVvmmRAr9nOM1TCPW
DxJxeXpdJ/uR6Cw8PoS7SVuxG4jUf/DPxahjOScl1g7vth71a/4XyF1ZSARTlT23U9NLPrMCHAr+
aHv7Q8JFcSnpWxNL2eARk4+GIooyd/GWC1EFo9PC+ZmlYghXyaSi4qeeADzBBbdrRuZ2jNxRhdWy
kiYuoltJhkqIb3aJ5/a5VBdfzOQqtyqHcKga+0DvZi4d4e5kjWLqCiWClqWx4rxoiq5m32kdszAe
lMrjsFyIO2yFhWxAkMi5hHbR/88ZALnbbY0hpZ6eHXuGpoqX3m9eGIbQorzTB4KzMzRgDgks1/KO
i/G0qMTUytQKTIpADQ06wdOSGEvlp+5UdIG1U2e1Z3s2MHUJCcDAaaXMsn/EJZzGZlI+wcv+1BMO
rYYeWlRf5It1z2XpKA2+csgTMvo/4ZRHk1PIHVR8Yo9Ucge8VM126tqlk/l/EvrJxzPeqbyMEPL1
Y2lLCAxuGA21k/9JKV5HfWn98fPc7e8QJUrJSNBhITPx8b98r/k4cYzuD8k3cgyU6rHnkAvl9Qbu
ACilUCQfThSNPMpn69N1HQtS1+pWZ7jCre9eYuLdODwSE2d6KRkUIWq55jP4DiYOPtB7FiZqSyHY
5DDYNJgJugUgP6LhC/1SpNVsiC8owfdwIcLHzVpjRdQOAWVshifVENBiqQcn8PLGEJTG79U0VaSP
iqO0HGnPQPg6bSRRCZEttAGv9vVP4HebE8gG3yfUqp/EdlDtu6wvNDsBta6GA0Z+SbGWgxf+ZmCX
rPWH4mpkIUz8V4uL+xgWZ2yG9cavM8JrP8iyXqQqPqGSI74un4ojJs7xjy9ypE8qO4okVH9ZliqM
Jwy5z7s71aTLytThRXSdyL6lw+VLDwea/okNjibvD0LSMe50tqavGnDkBaLVd8RgQi/HDDDZfzYO
nBm6UA67HaDb8FDEGOHXjyV1y0nd8K6z11LDI2GBUdnRE+iOdQf6uK702DBboPkdtxRGHf40Okk6
CsEviWYJbBGjlF9Wm7SJ3anUkp3H7Bae3yvtkpybNd9m5VZczt0PFs/Pu4nWGS1c2M8p5oZ547ZR
iX77zXIQUnhTVc78PNeWwbc3fSlo+T87Yuf0rqT+8IwF/FHogJUfbMYSfRhuy7dqKK6sIvVPVk49
5oWLcHqvAdzPFCqxy0jQwUDUMPKcZmr6njhdjeDhy5lUrKbjWDXYXCsQolMuRlNxuEsOSV4vNUZi
Q6Rt9Mf6UNAzjcNTJbE1vU9ptjmkzExUvKyVVzCY2NCcQlTllmRmyMfRilS12nZcDQErHqGzPcZw
BdC9GFr3Z7fiU97ef+HjDdqAQ4RoyM6Ge9g6dJCFxzEsDLxZaPDgtqxP0QYAnaltp5Xm2ub7zgnL
8xt8yc0yWawODn/ITNCWbhpcI1F5u3SvXzZoKXV5lg6Tls/yHlnxGtESv+kGFAWjgKqfqKeXkd2j
Hh46VX3pjstJb/eISYvjdTAE3mbDoKc3E3wOCdr8ksFWWg68BymSeMYVY3So7BchgF3g1EWezIpx
Ad7fuThxAmb1JoK//rXie+KprkHQW5owJuqzBQokqzgVhTPJfoMD2Jo6wZlo4zogYjdmEbY0+iu8
KpQy2ZYn18t44M0vrm5ao6cbE0Rrrcx3yz+r//zx5CMGFsxbM4Iv0gvNwrw7MKkMrEsk+Xwcg5F5
5R/lDy9r6NU0yGLqRYggujDyVm6USGci8q00GqOTrgTAFA7aqTIAbL5ZClWV8F93bBfAfQyo4WQf
v3uLJSlWo1ppc/ncacyyT3z3UGFEq6uaewWKdrVkDKoVRIbEHGVQ5aLUSZaUXTKml61vDEenAeFV
ZLAYBFqbCif6jqTh47xaZ1ZCVNSIj/zgIo8HeiHFyUE34WPHaZT7tM128FZ5pT9bThKegpnqrwCX
0dd01CZFuG22qPOuFFTqy5F4IJvDB24wgP+TIGRnTmXzzIP6wP+OdwpQBpLOwFZrhkOkkMJdP8VB
+RX0++Q+F6Uv4jtbHlJPP/l0Ua+rEybIcgFFkTp9EeWflxfDNtq5W+cXRxOWxHRWpSMABnINZuet
LNrIGN/639T6TGd3MqScruybS3c5Xj2AmAuu/T/ix/wCGmPIIuQXa90fCUOW/WOlIiET5Do3q5hM
PuS46M4KzapiQ1C6T70ZSqCUsYP65Xer8CFi7aoRhu/mymhJvhfg3O3tIPELFEyJPjlb70lW32Lv
68TzV57Q1V0H5mMz0rAxCcnLJ79j8lw9510WvHo6BVodHPtl4YJKWlfnw0zCG2zEZG/m0s/eDF41
vSCnnoFK00BR4Wmt550p2mTkMkghDdP5stJrwQPdtEOak/DwoaRhoc0BBkk1N7FZQ5NJ+soELH1M
mqVDc3bL2B9RCd1F7wNSu0wrc63BwKo3VcHQYJF11R9FDbUyZG/Fltjs9nvWu9X9q47z17POP+sl
R10DTwImFXxJqzMxN7f6rcUTuZIjYhf/A7+rApUdR2EfFLoox+0YR9zLjH/GJJoT5e2vqYkwen7M
QCQUqFY6ySyY81MRmdmqR/TidwxPGfyPI27fhXlNUemd5Icacx62AsvfabQS4d1wd4X2ze4aNxge
/rPhXH9ey2cm771xTcrunCjPcGL+i16lnyop5UtOxA9LZtqZDT0oDNjmhWsiFK3gzC1zGIONhxA/
X/1Wy4Xyj5z2yUdkelrrSTTp3yBmM3qHEMtM154aN6CYWDEIZjDzI7xwy0hDgzSP4P5jt/d6FyX2
blW5RNmfEllJRz4buUeQETOJUdpV3dTPbALF7dIbB43bdhu2ZFuivlWpFmLwvVAMspk5KHzs4pt5
8MGmLYuJ9tssLZ0GrgQtnoTveXSUFigkDDwUV454/xCZdPXrX1Y4pB/gElI9qsfZZmpIfFjJkajT
yw1a4o7cqM400UeluYV5zIPctNQNuLwan6+YOJsHTgaTU2zPBuQqNRF+P1El/9lrCMZXPjU7krrF
93P6lcKlKDDo0VhA8+9uqvIcSBrMWsQT9eXttCuR3VwMAgU65Qs1Xb34P91LLFE8KxDfYgjP7yWh
EtcEaFLTz2RDVjcnpgrSBUU1lEM+jhI+RPYHKWSyqMUYdmNg+k0puE3Jkds1FKjY20s3qRZyKlBt
60K5kzc5FI6h697jZ4/dgqN20fHwQBDK+XocPR9OsQaATiLhMnmnn+ectMAmUZuAPabQrAsQ92jq
IbIIqLkZIsGYfcKP6Xul6DP9wMm8epcDJt//V9ONV3dZzBCsFJQ5WzSqVT31TX6YuKFfyx3wyxL8
hPhFKD4wSCPa+5NaXIatF9EoDVq/vQBr5QtPdNCLSfjhk5KeDORnYw1/MKLVv4NabQRS+8PJqtRb
YzFhIZDXs887AdZVNI09aXXqUpAJbaS2nCDmm6Q6aGfsoY1PnEbg3L2IkqSbkGLg/kdmeuPdlp1g
a2VP3gxJmPJY4j9LwjJooiyi0Vz/CK8d2FVz/ogfhmfIVmzAqsXiUvGX7jlqnmPvnqk3JfBm1hKT
WosM+z01ElzM8LxBZWNLRsjnibB3foKA6UoWPQzMST1U/kjWNFaQ3UdZ5V7MZX/+FVRyQWB63B3E
YppAgPqtYaBlSaImMavp3z+MW6oAqan+6C4u9uaTvmD0YPG/rHiAx10OLGlnQfQkFzaE836IULkP
ZjXsbwuWSdiqf2AFi0PRXQnueaoL1yFUn//iYrXIATqHHGu5fncHH6T9lfTqo6HKPEHLbW55Fscm
jiPYWj10Men1NsCktsgV3O6DNeN1V2nTaOOqfqyOBc+0bj2mKRqQeol+1w8fDEdjsplWPkbsf7qQ
3caAZ7WP8CypzciIX+HpBzkUNlJ4CQWHCkn0s2fsO+wla/Q6rjBapsdv3y2RcHdWBmrwTNVW9Axd
PMuJyq2vBRNePLgBhEJmgJhUrJ8OMm8atbv8b3+/zFiqOvHdt8Zoch87Dp1SjRMnA7Iq/TYYNB5h
rKiR4zgtvlij7x9OR6eDMyf1w3swG8+YYWlsqlkisoWCf2gGnm/QSIXqclU7UsWWSy6rNQjTsyX2
jYRq3h5eHx1uKK/L+pndavsKOohgWt8PG9cRbzO7t8ZUah9kWBL7kvbPVemwkqv/ubBA0mL7+JQu
DqSpW3e4gRGLS4ouAj2/8Tomw9Pi2uUeb3nDZi+jayCU5PIQ14KY5BhmwPgikAI5rWmDiAQ/BZw3
qdChoch/emhBQFwMvSlKBU+Y97aPtLOByfPb1qzwhMVzPLzNoe42QhBoZ5dyMgP67CgKWmypgYfH
ajDIcV34h0W0ecaJptJHAGB7Hp3DLdMbPhxFHUhJEjfd1xh/vjRubmVbwzOtoAGFcsqIJ1tEmsyY
FRx7m7x7rmrnGxBzHS7EgAy8elGiUhAdYDn21kdIyH+WctsjI7wNiRUbQy8xpxjBNWgY3mHcTjem
aP7hpEloNoTz2msB9N+CO2WntsC0F1piwgAglIuTx90fZSjMcq/jhczXu3jCyag9N8O5nsXHuYqX
yhxaOg4dMVPGsMbm7b2w+jCE5heXzMtBUE92wC9HblioLgp7lq+igbcKzNwc8/Mb/6SCb84Q7cDn
G/d+Kxxx3gJFnJCT4SnAp3jqmsLDTj/o3O7F7LwKdS68sZ/MXx5iNhSvWESRu+3KaKzLEBUNfOgp
kG9yhf0sDemnk75+euF4D4HcxDKapaqro8Z7N/PzzK8lGVO1H2wTC6o8v3USb7DIsdKvLTpB1w20
tLNMfQCTGAw1dA+E/yqDTD3XH+MHZTiJ9mz3yMLyYn8IgX3ussRzoVhXZthH8435fjK1np5llLEl
/MGMRcSwQs5LkDCATbDLnVXHuO5fHhTZo7TMPoy3FpyKSLJcR2saXaTJGAtMWyBl+ad1odHSTfjN
9xNMeKIYhkk7uMBLq03lmLFS9B1USS4+f6vLoYYaCiPaesqgyVUIXzzFB5mU5NcbBINLac44ZakM
CowpJ5i5UT/HC4Hk9tqpxZSq1+gYkTPx4+JXVvLaAPof7DJB/KD2tPuiHP3OVSp/Fqv5mToHQ7hR
TNMjYuUVvct4LgfkhXQdmXNIW9Zg3whiv03gM0WI35dot6Gx71nr3RFNF12p5wrTHLJdkXSFQLnD
88FRd1FQHvjj4Ur+PRXN9mrH2l7nqD96LTPkJpdRtvylfZ5HeMAGTidAWmGQk6EDw2e+iXBpWFcv
ZframyYMxjm9uTQ4IFAr/pC3p5uPhoDQt+gr9m8w1GWCfYlqN8AAvlZ7deVwdDBP8ZP5ECrQCc7Z
g3htHtzABs7gUlApyVwfBWxS6GcGnIjHIs1xOqwiENstAlQcWxIExhsufSLRplDJquIggd7Xp1qd
ujzJzb9aBvId64t4/bT89r36BQRkQZ/uKNlyHZeEJD6N8emPEM/qIHmmlTrDj0tztldPjkODRcdy
5DbhPaKxwDAJ+jlFg2dxOcFPb/9TRAQsHVesi9qmI4We3BvUsRFYJOTdOAA7/mogd1WKbbJRz+4l
DPfXyF4DqQvDlysfOtviHXfwmx4tAkblmCa3O3mMbQJzw3Vf/YOK76nMjddz2X4r8yewZwwb+I5c
F5XB+gYCw71REtm3WTravbf3luJkkcndVTo2yjdGvkpQIQPng0ua9djNbVTWx82KAgMRUNJGr/Rc
3SKBPwa6mIgcBQTNIGpkY3qhKj6K/l/4jxiIOXpxDVJ53ILiecp7gHiP/sJ5Lwxto+o6emAOncHY
tD10PKGLmixLAgMpisseUfHsc3Y30KtBj6nzUu+Q7MVoBR9LbNRKW75fRhbc/Zi0hlDf8BpiCfI8
bldM0Qcm/s3GurOVbYvIOSa+d3q4uTsArHHNzGiKQjnindcAMs+D/oORDvQgu8/b+urgS/b0NhMR
7j8MaN/bE5Hj3njKqkTIFVlBbXDKM4bw1QaHwstScqNJnoAR2yRx+FLGu5TI42j913BYf9k5ttrV
G6mVomQDHVjuOQF96yyIFdnOSStro81QxKTvxNH8u0nW8dT4ATNsh2TMMvGJ0Lo6hpzIJVU77kH+
YySYo094LTCQYLX0VPz1HLQuQecj/eZ2Jzxos+eV5mK3SmKnQXCPMLdcv3maV6xAmMdBHGi/sPdx
P3g4UdrDFsAPre+HyLAyihzk73+bADmCVGksGTRLwdZJJsuVS49FjAq9Kk9f5X3SJly5d8wBeCX0
rp6ma1xvv8ed67ph8H+udTzwtQzus8wU0tvozbLeQxCb1+Jzbm4e+9r7OiJ9r7K+vt0LHwfYsimW
+nnTUtih//lOyxaiSP3Fty/KejKMsIVwh29t1zSujoD2hClWkG+usFUgu22Dj8MQRHEH4tmQp8Lv
DEep9+YXExQO3kYoHnESfCGRdfhsz562XjsirDXYUmKqx3SYSkmKJ7YcOKkt1tprcHqupp4YQWDe
vi9GulkRo4+WkJ4QJCEaXCL8qBq07fAxyIIRPXmbopd4Nz/6FFU9KRtDATF5a6KfmdtDX1ld4K2N
PizrV0doYFpnAf1y+YG88dnJgxipYQPx5s3QnYnEScnU1Ml3TDyTF1TgiXjbMh7acSxaTe8gwdTS
dZpwz750dwiSY1/aE8Vw2PfJvcZgijgGCW3g9pF1TUW5G+/x8RV1AFyAg+fm2KmOXfrqV2nMnQhs
Yi9pW7JcE4EFpBTY9VMDI+xIp6syUTN6tjycLu4PlYCRUkZ5PPKXYj2M8rFTptibCjL+RNHsA4AJ
DeYwIAC5JyHbKxhN3maBMgSg68gAO6A9x16fA41ERee66pK2r/rdbkx+izOmUWcJ+iyPfEWBtEMS
dFzTFTJXSeioqLEhiQF5uEE4PtGvM78G9f3hXx7P8hy2+FrOh6NG51oEuiiV6scwC8DSwZj5q6Z6
8aBKfoA3x4HJ6dJ7bKQC/KqvuBUA5cFkr3ZTPw5oFvOh3yj23CajR1AX+mgmUXbccsdohathbb/P
Red9jLZ7SCQoz+ZtGY55LV9GKXyIw7YqDJAqshL9Fc8Q35ylhXaiS5Sp8QCjLALFHGJhs6TASOZJ
pSUBbLEZimFLz9v9M5W3myCBn0m+Re/7yCqLbHkkoI1cX2KW1vDMXpOWmLuN33RRMrAzLe2NqtnT
CeLWiWcFZy8EqsNkQFfYxFBWZXM+0QUpTnYWjNlvgmzIo8H/fjZ6LYtEzefSD4P1ppz6boLU6GOS
DvsBtACnAM6OzHbiIqpOemZYbv0/Ri9uABcdjaIfOiRlT1cQrUSrx2H0mwDjOf2jScb1mE48mwBG
Dd2AnrFSu7N66I65a0xgDbLZ48sL603JnClePZfk1axxkhQrZxDzG4UDAK5zRjtKhc+asGFK3KFu
V29pjIg81+fdMQKt4U6eZ+3mYbjmaAURWI7DFDsJpTn6jzoVdgNbV3GU6OaeujBYiik/wy/nf6kv
2dMnjQ6fFRp4KbQU7twyvhC0pQAJfLjwtzMO/cjZ1gi536vESo5mkdvKbQM0DY9U1A0xABDjA5vo
wPpbL8TMijHx/y7fQV5mIZpxGXAXizqFHJ5BuIGGlYVWA2fkBvZcb5XXQf4gtdTFG2KY/rQ+EAOz
bl45ngq4fSR/E3D/fxYEfPgIGJd7Ev12NDe6seCpDYU4Ph6xxXlAFGkCDD8an6XjnbYDqmU+hbX4
TXa0PEg/+RHJypEV+xwcZNRXg2m3G9R661kM/yzHKg68dZUr2I2YLNAv7K3yjcWduZSpHmppWGtP
uiLaxT1B99R0qRoirmw0xNFtlgj5ZJ0dOSmeXNmnY5p5Ob4v6YYG1fWLG+aWy+xcA/XYydazT+cY
7Qp+eQ/s0ewigv3osaTjbuPB8quJd5v1i2PV8zV8TO/59o7NRZQaqdQXIGnBovQ+9cSQfaOVI5Kv
c6TSVkeWwzDp8poluj2nfV3K8xy2VI4gs0cCEveF/jn+Igh0eYDeLCvGLMCpCZVd0BdtzqD3SVfq
U9GVZ8KGq5mHMqn6g215FkoJuocWfmGShUtwRBTWZsLCLzqxEcXZbVhY6ZSGjrcC5tkJWE04B9Oy
nH/wGg9qkoIQ4unSCaaoaqSEXGbpWk9jn/Sbb8ow4Kl1pzlT4MpvOlerC7fI7JskJE+6F9ayB6HN
n++GboCITnBK1ldJfsaQ6T5hD5vtBqtMB/eefN3PLNgo/1+EUOLTTQp1FCrSbM5NKl5cCBpoPOqH
Ogpk+go3KrFIez1mKzKAU72crvd4fykUFWPbDh1cxYMY7u3zRlocTykYc3hd/7VdaDadOfhIgmtG
X5yEUaawnMEGd2Ia7bS+cAKiKVDylDGQf007UJMRKZoToYQTA7AJRXyt1c925qyVRXXubcew+lNi
e2V7+O4WJ9KgLluD681gnQ2T+usQ5/3tT8N+H1MbWsO2okZLUOV/k+bGRe1UoU4pYVjCI5XtMuwj
4rVTLYaW/oIg05yVsJCgY4MQaMHZL+nu/odJNVIH+OZiUC7QaEIE0tVgj2q1zXXh0VKA8iVKuaTr
92KUJZWzntHE8JRJBZTjjSD2t+51nMeyTI4541IMRZSE78wcqMHMPjI2PfF7nt1BPZkadw9AsC3M
DgwL8IjSGd1UanTCFyeCinWiVV7R+KyZb5YL1T3kSMmC/ui64pyFnODkcSe+MUICpXR+MbcU0Mah
FZTDde5eL+I1fsmLNVVcxaQkewRJM8MTKiFU3Ms2tAo7XIJL5N1Jl1UV+4Drp24GUzTlypblg5QP
0FjNMuzhHkfPeEcVy0JsGPPogDZT6QN2FjDF+0VNQrfxjWImY2xEoyJs0xgzB6ADbzPLHUsvwf7b
acT8/+8vp1SlAW/ndAjmU4ZWB4eopfYakFIiFwxj/44Ta/N94I8gB9jgKPGN6huSPPU8gREsSd3R
hVZrAGPrnd03HmixSSCXyww97Y8U1vV73fDyDvKkTDxVqMr4P0zsL0gac+5m24ui0/+ECqM43hE5
E6Qstgk5fpKOQ3U08SP9ZlNe92YonhXrBuw+hnyVNUnXmGR0e1N//TbzDYGFX73aBYEulC8BAwsy
8MgLdcIa9fiOnI/kMfKeLI9CHG970n/BoPBPdzl71SbigR+ZCkn9TmroJAYo8KnQF4rK5iisyOHp
+mWTVfHfHUTbDf+w8ioRw/UpjNeTVuc/hmi51WCp1zdoAdI2pF9QpVEHXjo7zpvLujiL6vUEXU/V
jceZD3hBjuBgjzTHNNUlXJpE0b42o7yth7uz3J1URkNXyrMGZlCGhE9KPGwyd/yGuUbzFpEpozYJ
w98pXzzqsro7RK/uwybMxvGnW8pv+0AbKKJf9yC4v+a65WG2IYkNEAsyXiYDC68M7f7XpLqIoTj1
GV96vxNALU87+p4pohefsXbMQ53eQQTCsoF4swsyBe9gLTpizDG28zxwEeNk3Qp1IOS/JUzRI4+N
FfLiIdF83mjTBj+NPuE8+nyUauFkG0vRWDsVdiMuvyVvy9xcMQYGwv4T6czkuLnKb66U528MUoOs
CVfptxSHo24uI+snOQQiwPgXGTFVLZjcKdmOg4jb+3RfawwcGW22Vg4hauMb7MNvLCku9GoyDH2h
8uQxJhwh7hWL4btwCqNTs9VlXCWrsVx4u7GWaWIH7jwx993RnqumFqkGaTYG+TkB7mZDwQq88cNL
n+CMGTHvHxXjuTtobAjOB2fBJFKcUHTPN0dW1NXbf4fPTHvly63Ik3KqF8FA0aKyWJVRRT18l7Ep
dlyHeufFSe84/EJx4ZW8PafxCfD4+RNZOW5pJCIfGHXpmPnjmlV/zTA4y9HXK81hBvP5720aZr/N
30Xsm82LBTrzEO/5r/h74Quo4cviIADWNylzgb5D1BeKwe0h3eFbxycc7+zkqBAws7dAypqiGZMt
vZzHhHtMq7RQOmlQooagBJtf7glqDQ+iutKC9uAdpbq4jiYi4RYrPTtTwtrMWBzh+S+lwtwI+bkh
62lp8KUJ5kMSykl7Ocvse3ueQXbtyEokg8AjzQ1+iVYpBPHBLA9XfBP3Kn5H/X1W57i3638XQyjN
lJ7lv+pXZQonjwVIKrSeHxbh/7A4tzwMEr7Okd4gCHpJa2cesQ593HwgN/cjhmsXDKdAMOE536HL
XXuDzJifsHXd7QA5aU2nWKsh8s8dZ7YdYfhwgm4IlZgBUSbZIXIEKabQbdCwFdNbCndzkhsS/2eA
a0ZSCxwnFog8eTkAjkCaM7i6vK+tVKJDAJC4AhvOG2y8eTPvQF38pQBPPU7QIFyVuA2zmNvLpNHK
j51hGoXPJ8pAg+jy69d3AupNIaN+vMw1Az3Dz8c1IvcOYq/WcGhCZ/QNr8vV9CvvPfz209s0Ocs4
6pNt4k8mzo1jVCyBDpHUjeTkfC4sCmJv+3MgtRquba51f9eP6XU+ufDqnFCYBWqsWPaVh12NF1b4
TDauUr/cIUb75YVnxiymetctMc0wduU2ri4G6LjVNAQzQ2Gsg7a7lvlpshXrRpdACEAxwtSgK/xg
gqDQQp9g798rY2U3hKgAY3pI1IBUJLZA2j5oyFk/5EmRSdmgBXzUwpgYBO5vgIQzVMH1ZzRDR9NT
pyqqa1gjhJ8fmvWMbAFXmZuAvWjwlMh2euRE2KNhKxuj6qoir718E6+reHG5W9hZeqm33M4zup1H
+QdbXJd3MZw8fKfBoaw6IMqxG285/oYUzsbLWKU9zE9IsCOh+zmRyR5WkTj6WzR1WwnaDmPFXsW7
W4QdWQTnIHIAt/coJQnlu70qcSZkZgwMRd6axuXdDxeYJ8QifCNYc8j6bu3zyGF0Kvong1Jo8FzX
4XKrmbNsdgIGvyrwBw40fc4jlI3N6vcrltqrVkEsLUt4ERAXlAOvz02jUylHz/qJxaHkxpbSqNlt
xpACY0zq+j1cH1+DSCVyVrs2KMoQMSrRKDVrvrBoU6zaaiuEwsK348aBAOiVG7eAS8JfDxLKd9pu
GCbk0WarCqxvycLZKQrF9CSRPKnPXucfXzCcpTvvgX8F8xG7ImMDZ3zYjO3RaeDBt3PinjuRt86C
VGGgHsXjdvN5hfHX9p2FuRtWd+mlampe6wrPiAYpjB1sZLPFXwIfot6vee1ZY9hyxCBbKcMi5ve1
1AvVxRKrtQpY8LqLGfFUyqAbG/Whp4uIpxKpWtMzZIKgUkBSleOLULOt9zbc69vXlsduB7dIqBFK
QgZrd32XisMNfpfQEkaSzvFYohyElL4y85D0E5auNIWpgT7pMySgSRTszxlNG9TuZ1EMZ7RSdVPn
YE6n90z03XR937wL0IKp0jYExSwMXYBf/YZux7cUiP2+mRN2PQqRUcNday3KHpApaLzBhprUsWmr
tLF6U4zPSm6NSlkHIq8NiYjHg/h9SENfopV2nLO9KCiR1pHN8I5yv72ijsjWmPFmtxbDRMSBRkzI
6BSiZzNuWzBwd7+g1H7j62B16oSShTEt8lIfBvh8ugUoWm7sPiHYQUTe2o/Dl10gqIMuPou/Cv5f
yes4qv45Go3X/Mr8OA9IbyiW7T1E49GWniDbj1ZcNE83g0pAzA4/IQsPAisMq43LgKjyMA6diqyn
tGFBQrLOl2xYNQPJoj50/hUS6hefXXuK2yLJXmPWEpHhGWoZdTF1IaC725o0cYcnCflEremtvFoe
G6E3xcuTxCDN0HuuX163pHBfqGClYn5sL7gq9USM5bDzAT2cTU1nf9Lw/eDOgi3w77MydjxJWNiQ
ZBx2yxaWP5Jegj6R/N9wawJS2hfCQvO6scnZUno3g7ejErEQYEcZ0hpty7yVZSPQVbc77eT/m6Wp
fKMuiYYtSAngoT/TuCz67js+HBBwRi9/3XFEAnGH6Mcwvgzw7Rw3H4K9E/8Y3WutsPiTTbJ9CGWk
k4pChroTV6E5/kqzsrip9FPnYTOdsBz9lXWXOyPr5F7adC7pn0YjvJhbfNNCZBQ7kyIPp2yxcwFn
f6c+NQUweZvt6Hxz6k32E82JeDCW0FlUHuN25io+8Z/wWyTHVQm1BbI0YY5UDVFQo30GCLQg7QSQ
z7dX2jI51cRPIry7aO47bEAKMHL94DocG6wNMIxJ8BM4pP9GfxaSUX88bVQwM3w07MGIxh/zaP+K
23DGiQa8Zr9rnwDa4HTGt+fXJjl1lwBVFXl5jH/ihBD0d3ILuvJUWULFk78eQarCWdGQYajerWIA
jni0QYTXq1UwhQtGgJO/PJFHZcUlQrpc1m/++Qojh8terDbn7ev5biwnRqmGtFvRwzyJ09bFqamq
4F3gsLabCBwJPUQ8dLwV0gnFCzIz4WfxY6A0WL/tyX9ieqEi69JtxV1snyo36jFqGCgMGHcFpcnX
z3P4J2sGlUnnA9rzJM6vsz/642aLs+hNsNQtf07z1vMWtCjzz0RDaFyinxoND4Dpn5lUF7IVd6ix
Zf8opopOoX/PtYhx7+kt5ioqTvaKbm0Hw/4UaqrE/1zoI46giSGPCqyIA51ooE+NihMo143QLchT
MTvjaazgIo9DS8kyo7xzGUGYxGSmWc992MqYcopTLGcXJEFcp5ZZTGrFPhSt3Jqa/Np3niL4V2bZ
WxevPRNmu+TkEJ025dUdt81MUo4xCdFoBYSzsn+2sU/1EoV3NCCmY1T40ECnYH0+1QKPjCfZ+f+p
GjFoeyaAToz8Z0lZNuOvr6TwBUaloOMWgqu/PmUE+R/Gv/UwrFfscSqYuD9HmOT50NM+/TamC9KM
k2kxc7gtD0yhNZackM8Y9qO8QtsQ8RXzKqAM1suD47n3mOz5z87J4fsZazCWqExgYwf0PbEtiYxB
Hzt/9lYoZ+yyuqyrG1UVysP72bnAJllM7wIbEv9qwnKZ4NvQqLQQ+ujqalQQPTOpG6AyzgqO00OF
eVGGriwg02Uns9y/qOaA4VAFPSucG7w4ENSzuEWEozG33FBLVQd3qzKaM5r1nXdPLN9iKtpn5PCz
AXx5gY29FBs2rJkMh5E5Yp9W0hyRh61zivXqHSIVBCujwrxXrLhv/ABhv1MrAGbQ1+2/XbAm8WLR
BEoAqJCIvk43jwEiKEl4Wv+dF8Gy4fwZVPdTo3C5gVD6TKEzMlq6vTwfpmejc9m+PkXOEa+m3PsV
UGch9DuuwmQgXZnCGEVNL4CoNKDfE0OOEhNu6PxdRgCpsAdwaJ4Q0bVQ3uCSnr2MgSz5kmJwOgzn
jdMdSmYPplDzLb/uNykFjviMrqpyz/KV+PXEQpc19v2Z94GcKl0/awDpfLkMx4Q90ArI/nbsVQCO
eoYF0d/RPJwPhUoRUeRbwhBXIZm0gvlIWLkz7IXWZJYACAPrNpHxKN3RLIPVyxSP5G75jd9Bzv9h
t0zFNb36QLyF/7BLk7vXSPMMQlJkbq190OqV2ZOerC/Yd/ivPDXscE5RQOQDlFvuwUclvuAcAZeU
7LL+wsvUWTVsKI8QaNbZMQJz0DONfVT2NYg/G3TwX3UPUCs6E0xR9YysT1W93TL9KOYdD17r/MMa
sePrDJiINgM1DsdF0zbtW1wd054AeAKcODdHi7VS9x9mDjq0G6wbremBAQR9MpreiRMtlPsQdy52
QFuGSPgZyJDRA1hWRRMef4946EKRmT82mUwX4ckII88EEvwB4XZGtGOZMYsBCBJu3z78PgkHg7/y
UT+/5cC6ipmDRN77+6iz/zlUsoJhhcOjJIN1BkTwtJ69s7t27hxoTXKKeiY6grxGYc4vcbBOB3rR
wmPdz6Wuxh+gajX+22UyVEac3E9is7o8TZZcktB0w1FLHyFXAkLlR829acL2J1Hm5CAzebjPs2bC
wmU+Y7ZFJj0jgM7AJK89T/mNGoH1OEz52nLNefgi5NRMUCzYU0TFg2UQQKunGND1mCiHoJF7nAPY
XK9uTniBR+ArBMPoj7uAj9pn7o5IbdWWYFewjvLpxFW/lC5n9CayMzxw+y0gnrbpeK/uOkBJQyjS
anmknMgl/coOa61MwVvuaQvtN1pH25WVlC8QawumyYiqTAIWME4FuHll7GqpjRFeRGXrmU6ZvxpF
8FBOnizRO6Ti4f/5B55yb3oHyaOgGB+kSUyKvoZ64B+ohDdLXiOseBLYa4V5dbv0YQuCwhTsRew5
SwJhZLPVr/75VHxjwBGow6yQO9fhgj/tdJEzzDIHzYdPFGmUm0EA79p8ZHkooQu7VdmR4XhDPSoR
Vs7u15UR/kjZZ13Z+rwaR4nKGfum5cpObBzxDwp8Wfy2N8NgdZWbqYEf71E2mNBIa1qdaOCnTg+w
Vc57+lu9wHxFWyqN6uPneZiybdEUgyS/hksrjNlcNYcjrdYUzzIUD+ftYoAzZbEROTLxRLf6gU2A
yftE0EUirjbs+nk3Ovdb+gOk/d9ghc4bqbvMfUic3rcqwc7+b5hjhLmfRGaiELptMcunIDMtwshh
+KkIFu8CEYacHN8h5HbX5ID9gSZbHdrpH1vsfIgqZUDZw39rlzwYGJbVWdumzol/VbjGwrUxjXVc
+Wud1XMEArHnhc02/WbsJdpivLetQF3wDi3HRAI6KuuYxokSiyEwJpLJj177TJpjtXwSwcHdBnbQ
2JQINEaMpud+l2SKR65wxIqoS7PnYFmfyhdwMfaqItLiRHIFjuONul6MxKCeJlpQOIJX9HncCz+t
2NET+tTGkhTrzI96R8RLgK95dCYOrqQpFUVfS+np2Vf6wIZEVWZ5jqVcxfoR6Cc/VRHWNjazI1yb
RuCFqioXzeDSqr3f2uVF3PB+ukWZuDYHvEDF2/cBbsof8VwG8B6BNyfHNoZPe7xgCD6SWETII3PA
JcAFB6U84S528Z9iBx7zK13UsxQriK8972q5n76MI3jmHoSjeqSVLknrFFhxC105vjc4FN/LWfSs
6obRzYrUKQN5RzApEZt+EHt/OFNSl5ALf4vezH1lhc+GoFqa+XCSD0RjJB9DXUIQ0JpX6R5oR/5A
CwbmKx/e7sSGKAxMhqnf6fa+Qch9qjNFJXInsHtW/HzTNTOXS0VdRzjFxcB1urbCFAtPmenyebRX
ug5ojZSv0WWRZx3yJjqAjf0in4x9cotik7/gKJuY5aCKd8ZQOUbbqVbuh+v0uiU2xjcdV0Z30Sld
dQ4RVt6ceBKf9d6fRV5RGOh2a1UNGgHu+L47PC2GHPGCORkpujWXndMfC0ISRZfZgOJ4Sc3CZ63J
TrzSyDhO5ZkAY+qfhsFomLTBqApyLlrPS7Jpbwl7UvEP7S4FGrftnqJD3fVoQ+SitkKVpyF0aZ5E
qZXSnQZg2x+h5N90EBQrN3Qou7+EzACzIAvq0lBrdOmMleF13rM3Cu1dbHAR1qez8NQgO12AE6Mn
N2W/AhMy1nkg/d8CxZ4YGPQL7aqOPxASxOw50YnBQKd1TSvigGxStvyePBj984n68ZTEIbjbJzLW
UeJh924UwYynmT9zR0pphhjEDdztUHCfD2rwUEPP4DesDONOAH+oBKb5Cz+vkAdcB3txHzAzGMDa
sNvCQjENdT6sxYR+ZpAuK6faoCFjOHlbU5GuauwKaH5LBCgqTipUrkAAvOngeXqR+GlNGc+sXyCa
DSGAAakDM9454l0PSxLzIQS8BMaIkg1Y6p1H3BESKPUF7hLV70ie9K6XVidrjOVDOxt9xMnpijEw
h6WCxu9YK8QXN5MTFwaIu33pnwVEmF8ObhW6AzPQA8GL+E4uTnRlA4uMOf9gC9xCubaDyF8YIGKU
qgTRK+8uABoT0XPU42U0ifnkzBnsZnf4KNgVwe8JEgmqXU2SyRFawlPtwmVg8z1wm07qYvMPYHoK
e3A4eshYonbJoC4tl8xrdP2g4zmkL80/c5fDRy4rkHMiZLgKzNUI5jdZjF2uZ0yTRWLCkbA15bZK
LwUPdqH1R5Lv0MEAHbsXbqTQiQIKCWQc4/E6kD5wCIAWtu0t9UAMcEp5gQohZEQ78xWJ0v9xZruE
y5PQZaWuZrVPoYhFg93wGkhoSsIabwzfw87PNY+CL7PHsdXB/mxYd1t+sI4C9n+gbIdmeW0KrbDG
l5/vjf/xnt3be6MCLdWSprUvxmTy38678t3fnPkAKNkMAAozNKVatraIvNOE50CuFBqJ9sdplNmF
pYNVvO71QjJze4goCRoiiDeg6E/sSWMw7TPqL1X6cjrDuDeiqWT0of/y/LuhDS73zQiCsu5OB5SD
jDAsM23z+/7BSmkzcOkh2EFzX1dOSJLtAGTQoDA7lnVTluIAytuQO6RUS6vVlbVrplMKuOKavgpX
7dnUfrlKETS5ZbG8x5jMUTgKb07uwUMWU9rEiHxfSaeW2SlelQZjryX/YcuWrMfqLNHNoyx4nqZb
+QJQtABu8qqmQHePQKpbj1fxEQyhWFbOhnPYWUQuHiSz0CQNDkOcePoxpbsjX/MA4Xp1O33OKWkU
kcBCdHkga9ZSjov+byEGO1cwCfsS5XND+sjWjB/XLKLwcblgwnr5Waf6bpyIuHBs3d3keQJZ/HLM
FyMGeczjOx/4THP8EmZelZtyj9236Hjj8dv2G+5yDM9NHbU83atOj1bKWnLWpx1dHTdNTAfkD/TI
NLGyPMpxan6Lq19MZJqbv8LW0VhS8VmYhY/vogyWDcciEmyLS2haxy/78oTTjr7e4OGc2kUrQs89
tPQpVahJxpuuTNImG1jmoaqZVTNsyceEV4K2o/G9rV8B/PrDBCBpDemomYAI3/F9SfuX1XsgEs9s
JQU1W2THXrRrznKe9NUzqXx6SjGzsCj8McDnj26BOi5R9CzPAqpVRqmdlH45Br9/iyw3So8q3dIc
Ny7SyRvS4ExQpYeGKzpISBj+IS6HwXQ9BgmfcPwICzbVNviCf90nxVDIMRMgdDcc66X59EH+GI7r
YLVgV02Nx1fXFRZ3G8MGSt5HjaC54yi4mbto22RImS4CTiBWQf/q6NNI3VbIIPPc8qCg3R1mbNAy
v6GGBvesErlInCaSJgXmHDSrvdGJ4Tu5HHJmm0DyRM9eBETa+EB7hyF5LtZ2THQ70oDy+kjHp4Jn
CZjCxmt2U/yHOWdiBXBe37OvJeE2eOj2RSan1bc+/oliQJ/RdJFzIJMvBJdBfry9rqhoxQa11MRV
AdPmsCw3MvqlN33MPvqPNs3VBG7T/4zjKsp7C5376iYH21V19/5GVgnyKz8khNjT5WmQVe9rCwA7
vdMvekLxGPpPoBhIxK1xFIqI+Tr1A1NMhmRYCTo1NLm+N8Z3UkRT5jWS4uQgBS+q1NcuLPAtAxM0
XYM7qGwSYuPoB0iTn7F+NiFcFRND7sb6CpEaRWd3Iv4m7rU0AnFfWfzPsQ/1BiquuhZ2fBLzTrWs
qDg6LRdEQKMQ82hgDceE7UWRiwhJcl94siMUMHBBK5WqrHqXUZpNsnoyMVTtQyDCIOzNEER5Jg/r
ogQLCOTsQmz+XVrpTc/rsmTO63iy/ZPuyxapYr7fvoN7L9betIPAneduOenGoy6bzrupBzuVOpF7
xw8zJBjgcwAcNLjTfvbMWcLmHHgNCuMZlaoUjjimjqpIqO8S5bx/4Wv4o7EKZmC7Wr9MVSGgDE3D
tkdzZrATE7WHFOFyaZ9bwNM2KMGFO2+RzuTLAvoGJCrHSsvFRyqCADQl/ONkDUtifo15ASw/hwpI
v3Ny7QBpg5IINNWjYTCyW92k8x7n1xOlqn1FLHkh5OMCy2PxiTResPpGrWt7qbaTDDIZo5gHyX8B
PkiCqUYvJ0WjVJ2DVaxV6El01njp9cfrtDS+gzrcLB95vsVfXlLIGwT7ACcaP1SxjI/D5d1tsGGL
MnTXFurynzTvDd1Ny7Ol5PvWGMPWcd6tl9TmB7gYNHJMmEG5Fkt+kV0iI7QbU3Yu/+LD8l2+bitq
TM0AxifBkPXmsihGiiyTq0r2n6wgn8VVnFv5UrGuKmVMF5mxGAVz/v2PeuzU34jP6PuXKTphFfdg
tq3+okrBeHhFJmdKcEhBy83UeLJnR85xMLc5atHx5f7XMf9gO/1kbcnpUDjttRZk6WH04UyuGvG9
kwf2o61jcaePMQrWcCxdb4gJWZMO6z/uhxJvJpJuHivv2vuCAM5G67xJpmSwlm061mEeiAKluogu
ESaomLxeKKIGpgjnyccle++kFZGNxpPCDcoqvTbO+x2SRQd52s3xc86glk7TY1fsexiWD6hihLhc
MbJ1iw/xjEL4ZzlfgOkXnxoT8O5i96TuYoHpVPynjI+eyQo/ZrivaXuHmBFupX1NSy3SuAWu0jk7
EboONLaRL2HIh6NneDN/Z/1Ts+iUMRDK1j39oc0zafpiu64+ngCFEoIhBNGqkMG7Xk37NzpY085r
PGbA0Pq+32prk+cLjcuaweioZvHS4cueVoWbV0WQQMZ9QvLqfzU60MqorauzgfXAy0WjFcBdAwcj
uM70wZSD9Edr6nuDEAsIAbfjxi4aFuXXnWrZr8F3ek1A3Wrgi5dVXwM4qaYenQZO0f3OccDl6eN+
MJEut3RgdO1nQoa4ymI5/9Qv5qLq/FdbPUgiOPna9k+uy8RojVkh9nX4A7c22frt0PrNzrUSlve8
Cf3wSlNOQH866wzh/zPKUkWglU9HcZIjVi+Hk2yasWP/6fPLTRTAfZn/mJnMuQ3YmNBjwEb8ZZG+
NNXjRAAPWGBBE9kgZ5KMYclPwKfrAcp8iJDdNfr4em36Jzua6Je21+pfIxGMDNv8TGXnbIHVr48d
np0QmPEFG+AKlq1FZygnmzq8olHPGiJN/XyrsC/CtVycHDBXsbIS0ajFtgsMrzq4Ll+Hydbo8lXq
sPBMSg6mcgOam1D9ns4XISDHxe/jHj1u7Bo/VO+gmwjV6PcFCOEwdymAq2KY7g5NUTi3kAreiEwl
3jh8bbDVAfSp00hO74OHK7k7EF3HItufj9Kl7IkS3KbDD6Tdq2G6qHavdsp7lCRs6erdPf6HanvA
yu62bfEoAOW/o6A4b6AjevTkRuzvBzB7GjYbZSkVyBwU2n09KXn9YJ6nRfEHALfMsfG04vfIOtR+
QfcFdAOWHpboByfjJlObtx755nTWOHVwueNxMkuBjRmLehBf8ipa3o5zo3p1ORvHaGDc7PUXtEDg
tti3/nHXA7fUYu1Uy6V+3ON5HZieVYydB294quNIbwRqxOnlhg3NXJSArgQi+jecWJjnRkFNETvC
S2dWabbHskLcu/vtcnmLU8etMBayHOXthJnFp/L7/YjCsplDYf9ZN1vK3yppcHVisT4TRwdtqGib
WYGQwHJUVWmXmOpVx0xM3gPwPAhCQH3cE18H1639arkRoJEd45n3d/UniYr3R5zMYfC7BDILjJx3
EoFt3F6PboZPweD1PKPYiAplI/KHBSFQhf4FKrQs6mGVL/+ONAgL0oYXk6I3ktbl+X5dvc5/qwwS
RWT/LknB/7Ab93QLUuuumu8jwmMb0bZRfWB114pn/t2LX1O5Abhhe2hnsa13GFewsn335sKj966C
THmdAm2UAzikvTqMyrQve92DrX2flVAf7TnREfr/5DnIqz3syo1lUr+ccGIkFirSAy03qDuRLTTl
zAbHcprbcRLw6TJjRpvWP3qmeyBQahmzVlkz977rg1lib/j2x+DayHWr1hjo4IXJmUH5AxTm7Kn+
HjkDYeeZnlIyQW/RLyUOOPJ6YutbsV8Eo8gGi2JdStcKsqr4w98se37ZcgM4nFm6+dZizn+KHc9x
VouIUCg3Yejs901+o0aQJ2C55YB5eZWgelN0ELOEMV1EPpm9E1G8qr8IdNF4a6hjTqi5zKyoFNuW
5vnjgfHEMj53H3DPFzNZJZcEO5gFkZFpoekDSdKv3NYpwX5ICOakzfK2jzkcWA0O+qK3zrK28SJR
fnq1wzWKtL6dxjp4bDLKmw0TegRoHLxnlqk61+znmscV7362N4gxP85mgASvS2ptx7ukGEF2bEDO
judlYhwtDu8NqVNpJvt+XzjBIbuSpx6PXWJ9A0pG94Svd3nwVNQn6mZapu8OWmPrjot2cRLYblmj
aMbSmPwfia1BKAxbRIpEok6UhXKy5UEcqZUdU/nvxNwKdPsdKO+xKX9mPmheE+dmON1Npp+Xfmn4
A2c+hE8A+w+lL+SAODzmvM+ydPSrbIj23RrdIKFwKYTpLN1oB3rmEYMvqBVY97bQXia1YRryIK6Y
SuItTg/m0Bh0iQ3dBKemOjWzxHwJIuu4CAMGFah6ERCU8VnJdMOrrIANDVLvC82BSQ5fuSI60L/r
c090GmVE/RJe9HederipTkgQj5BUbBVxN1dHqz8yrl56I2RphLp10m5Z0pPPJme7DlWZAAkyPsBs
x2LTnNEu/GfmZmhWcmT2c6pxDG674hynxyJf4kHdxb72Ggwn7SNKk8AykVm8r/v07/a2lzKxyWwT
a6rQb5COwesEH3MoXpFyuHWLHHnezQxLsXmuGcQoepKeH4ekVfs7DX1D1ZFZjLFzMECN9vCrMxSH
ORjvP0wmJ69gzsLMMFy0FwmW7c20bI193OCe/sex5kp/RQQVwO18oCksIq+uqjD1rwlq1+twPwp0
rUp613PC82IdkEiUToF35KLUr8FgNN1ezSnrIOYOIoLNlGB7dmN2biOpE2ALF3/qLWfm5eysh8a3
H1Ssb8mcW6FOL2yfh3bJ3jmcT4uGeNtmIPneZTKrhkFPVu0SzNGSZuKGEsZq9xgC8I5wQk8bog33
wjn/SLN0cPCWIU5SchlWy4pctx/dtOL6BmRaPDzAURkGbzNGho5d3BbUHJUfRxqwvDqQTbs3wSDE
GfWGxwx1/d3giHAmXc8y/j2buedR6egIMfrbsFFkqZxhJNefTKAYLR/NlERMJeVaxlGAFeOs5jAM
AaV6h8NXuyA55UDn0ZDfvvDUjHLSUyaUlo5lxNkdSkm0IQBr2BNhPs+0xeDNM/U/x1ajM7THrPvz
SSYsy/+KkASYK5B1j/5a5VQM1MnioEc/r/Q7IDp5Sxt6BncOUinYEGaDasVUljoNn91HqQNHFPB/
trPOm4StLt2U/gY3wzc2sIA1ovlMa0qTLG+dI6Xr3LTOPBnlUeJmaNUuQM3JkHkhEtizCsiumD2R
95Y+vqkyAxSNkzJuqw+jMSs/a4BriKgh8DMqprP0cH+RWBAXfI/DA1UATKrYuicmaZGeQZClLT03
Z6w/ZjWAzfJdOE1foZgDccsh1aW7xfWRhO2U2PhK9Hwr8aUMl8pXilvWKEyMF/fF5Fbu4/ZLt2Hf
c+FVumCb3iUmoQWuYeGGz+pEUvKcYUuC8Jh0UUuAvLlWRGT0PLZIR7Ttfdaf1mUNQMzPJjmyOXJo
+nezo5SCIQ7Dkawtr5sPWCxRuVAAxVscEiPgKJKJxLGhTt/NASTV7SDtcSocDVht6QZcY6pLPhRQ
wQ7N0doMxvwFJFn39koy3pSx4TzXL6qjIL+LieGpA7L9vuGR+WTTBc5Yo9o2u6X9yLTXSN4chEXq
8HUl6DAa/HJ98cP/19VxcLs546u/DITA3vyx6jHULk8KQvcq4kriwKlQdGjkxEK/II1X58CAacgX
xbjTApCkHAFNanU3eizdVTLkWOR9ZZgEYLZE9ITG4V+lITUEZ3SlpWIudMHwQqA2XENax48dpZLg
inLzd6gKTwLGudxohgMiWzDsfHAf3oFasu6KLIEGX9SVcMv/ooYD3DhH0BqbopDh1Oj6VzyIJvGS
Obaj6RUO3C7tMvFCCfD4G1uBvhmBZoOL/m3azvZoB/THqlqt8v7Hu/wu05nt1xdq7XEAUZJV6dOR
zjdnNZmV9y+JGrTh1EWU6xofcFerNaF685xAjyp+3fV1yNAhWC6du8FNX/Srf6GjXErMN5WfdF95
A0ytIZ9lBsltpozxZ0/VNoVo9HOF4fneYC/AmmFfaOe5KPJI+gT8cV2DFvIChr7CRpbWSyBJ2YYV
msEp1b+W1+GRMCHF+WK/lv+955VcVQAkhu+PmT8krp6avd1n5t9ZsYekvjkdphIewngsHUOGy1yo
xHXAz6ixnN39hi/wgZhtgMytHM0MeURaRoEuo+SRnOB0VXV3sRLjkUMTz04VARMcAXhmLQnuOpVb
pGjt1R80FTdnQPXIbCJ+VKOSAmxts30RDQMFFVp0gPbKT4XhTQ7omZwPei1kTlnyQVJhGSS7yMzE
Zzt/86QHsJP0O/hQ+DHTptSp7FPEzIgLPsWlPBvcknABqW4hgDgRPlYziKd8uNOQpxkSi/RdKU5X
1bU8h0M+5nQmbPet7TPzXNpIw+hV/qt+/H7uzOQqNnkC19+FTnJkNbiWhrmJzx6h/P5b+yNmGYr9
rk4wSjThajTqNiRJXGslDSEJzHL3uVLsBCou4rml1jm6ksMqAyssQ4ltLKl+57/uHoo5veWX5LX+
Fa42pvSLxA6hNDkNgXI5H/VEKkpiEwWpcdbjIpQDk/yohHZP/+diEcoxpTGfRZIQcivtFwfs40dv
nZMck3Dz32aZriNvpZap03nuBZgvCxAVw8VuqRcGzvf+ET+x/N2Y0uPawM6C9xNVxTs7FloxdW3j
QqlIx7/OB863NShJhBIM9eP6OLWQAjh5oWmwuFD8chgH7wQiH1XdBp+OTjcomWejIdZiqFZNJS1Z
EqGBh1fyeSwQI/fwUJps1b9OxoYxlfNIWCpco+Sle1KuYLNhnC+WV0/k6m+bwCWp/Cj9IPa/NbVk
+1/rhTnjIU7aM1zT0hpg6TEMZkVUo8FLiOpFCMS+fJSTAeEoZ2pECxz/4mIVUezZqFdHubLatLM+
ZF86rCPtJw99DOV1wAhDJNuYbGNAuDjptCjNf0C7JggnWCoT0Jj2MzN+yq6AaOp2R2QlgkKn04/c
sMyCtob8sdvgbfoCp7YA+s+AM1V+hlkwL/fHRsLLUEJcmJFp78tYtaEKZM4MGYDgvZVBoX8XRH13
JKfkDhJTq1Qa/VQS3mAS6qcP6U37aOYUM6O/A8QAuw2hu62ghJGEEmy33oiICAts3ezVVy34IKRw
nQvkjccw1Z6FrEd5eMlK/d26SngSztcyh0vtgzHTq0q4L2lVO/bSJMGSZKoMqYykUGr+Q6PeF1if
GjbKVDc3PWbA66P5fcBklZw5q6S21LR1RjndPk8583km4MWsSOwKFIZRyO0BUMmu2bcpcvHnCbGA
DVhWZKXe8Ny+nv7ZhQCLJB/tP8qbZOO/dU5gs+mJbGnzuwxZTzaknXo8HlPexkZtMEjjNKDS5Nkd
9ytq+cqO+l4cCWF2Fzhyv9DRvoMajdZmM86w0wOw0uKtEh7IXSYi8WanzLoCL33irq29l8s8dTSD
SENP3EA0GV2WCJwR/+v9qOs9FaFLh3KL2a+DY7Jblwmq30M9qRz2NJhZAWo/GStCyMmQxTz2x/lY
iS+A9AybjqYrXts6UgE5ShJzbh4yapsEEnu455CfcUWM5cQ0L3S5zzJkz2O7UV1I+pkK2/y4zvFO
xad6YWhkRft94O3wuyUK071ykswRdAUKikMvlNVzhaLJwoMpVINtxVaNzdWaz8Wt16+v/miZRG9X
W/zCMtXN9jAGcvMqujo/lttmFF4/38mHeqhXZC7kovlt63665eccp7Xg5ujQg7Dp0yB364yjkIZ5
u3A4ZSl4GnL+tO92FVCjO41UMHnZpEUj0tHqJKhziyKn+Mgs99i8OOuKSVHOwTyKhpko5E/AM3u3
YsJWWACSuUKnDaQDx7pshnxSkhrUWOMRk6tUibh6FzV7RFCNrBNq3fuNG/MWVHyCsoW/SpwQ1TxA
kVNIveUKD0j2u3Kf2LARNl/w5tIelhzvmLMKs5zKBPF/qZFWae0g+4hMHy2mMtBLxavFgp+oOgaf
Dveli4ZnId+HnYNhy/+INHKq41KLtzEgFQDzFSLTIgmkx0t5S3WnSsTzFZkYskE5fmRLNRDgZjI2
HOPvFwJpMeHgc16GkKTGAmNHtYLa+e5WwGbCKZfVIfIsuGHGu1lX6F5Do60R11hWooQLmbGCR+aL
Y+/HTFLnJ3Uw1cOV0AaYVnccIGiSVgsWmiiKikAphLoIlHnFtDDDzwK84h39LPeroVa7LBjTyX5y
iahUOVOGJtnN8C1Fc/h9jRlr1cnrffahfoTfkwm6jiUT0oz7FGpG6+uycXsBHQFvl563eWVYNOHA
jzxRrY2hgdm+LblAUe+WqTq5kCzgRLC1UvJfaODAITX0Sd4xYiEZvEwlOng9ptZFifLK3QnI4HPd
zijMu3IIZ2PP0P5KgL6O0n19EqdFPybCuR3xHGp/tpcfxyhTcHD8y1jYBYt0Q2TJSO+5X5er7F2O
gOQU2DzUJMVvWl/+5Ox759zMVabRiXyO5gPWYf/fPkRedDEuwzZNaEPk+XR9s+qrlJ5/ffD/A9Oi
zEsWqhhmiztviY1hq437Nrkj3DGrdS4fM2MNWjZ2f0VWU8TwFDdcs+EFFxZGX6n/X1KuU9Koy629
xkYvQKUl+Qz9SHgqIjSfKN7KjJ6UHwiGravElpJnLxIq25Eht8TB2z+l6f+zU8eLPU8kkDwXzCuA
lWHnWQg6e1aVAdHgzgxSXbN/AShzBeNLO4UlG+FoqeZXgvISGADpAvZieY/zhFyi3v/44ia7q5gI
4E8vVRVsAX8cKWJUbPeOZFWn4HLM2icZXyQRm63B/JWQdMm4hx9fDB5M+aT/QeXIl6lSolHfYsST
5Icb3vOGnCtzNCRXFz3VeDGLywusXpMNpY39XzpVtsYlCZ8VWIeypARqFOTEnVD+xmRtABb3HtJP
w/dk2XWWG/aPX+QmBUaSr9baMQ2XuB+Kv54NQ6lCO0iLM4cg2NR8qo5g060Y9mTxt4lDXqwqChPo
t8vnLJQv6/f9yCEXQXby8FzvAJg8VB2hDT8NylkPU2kpw6tkq0WN6iWCcAIbokCagUbtWe0gB2nY
WVPxXrV/jEz8qFDywBy2QelSlcEkyDdUNwqoqhZJ37dNF/EYTg1GUicvKuKWX5bgHDWbrb8zjymw
zvi3ONzJ8OKxb4GDQ3TkRH7UyGhOZCqhP0uaKi4H6Z7aiF7qSiBmOrYaCcaInVh5v3ky3itBXiXR
nQFK4yy/ZHnnYpZwIbhG6PylcKgxzVj18OgIV+N3SQpV8R9VnUdMjTQ83EYjhO6Yuq/1Jz2rBlR9
lossNm7rmFJoHWQlW+GXhGewDnOSPywakZ+IQZjLa1Z94hcDegan+9y64beAr8qTAMWdc4cv2mf5
SGVMjlKXw99ODey5aYu4tv7dpFzByBjB/6ltzL2CQQBOpNrNR/AhlNrJDfsATiOFmmw1ySHync4W
A6zMvWWv8bVYC+rOxosE1rXbhlCEB5DXZjkKCwrdG/rfoRcyfZngIffA6wh1yLET/3sgey8acsus
2NoQRLNT5F9gr1cLapFBzEW0ZMHxEhlkgeBlqQJe1zxzdHHnyEd72XK0jLhymCP5lm0QY6qpsW8i
zuHkubBrwSAI7YVO12RkjA3JRtcYd89n+8Y9O+i/ZGNl/EOynEWjJCMpsjwOtpz21K6/SZSmLkNQ
BF3hnNw+5IXZ1bSzoSjxbSkzWNGFPAX2KcC95ae0OQZNzfuVEjESq0EPSI4ddr5N27JUestDcVkC
GdR4011IHzq6bV9h8Yt0po1wWsyk8NperN4/Ed4c6yW2D7E75NDq8BvwducbDWHS31SPYcag4dF+
4lqpJjMXHKZlgQuDRa0Lq/mPwCOrVDqA/llDKbaFGbeDj76tjl/IEEUoJO0FuSXOIcqlj/cDUzqV
mDJL4azRBeeeKx2lGuTskoCQIKeDNo2BxrLsRQeHO54okxQK32in07bf0V1WT7rcOL2Z1MonFBJg
B1rnf0eDo0JoWupDfEB3oQ1ksNU0P0dqEvh9kTlwoPI2t8lw/aYEIepAmmoyxJ7HZGeC4G81wKg7
jtfrcNmMmTAdZd4oSZgkiQK1o+57gMUpFNCrzVbfMvcria7TAw4vY6qtkU1YWg5xSp+1roa+1fQY
B4JpXLBF75zy5NsixH2+nkKdQWPqNbtZzpXO+2FmUaN/gxfWr6Wm/VSGrZCKRvNSUQtLSKeWUndd
pSqxYkm5u/78cIOVaUHMixOcq0qMvX58MM+uTLdTGKNesklOacAUGrmQB1TXDFeWLG11XvjKslZt
ja/0CxvfCm7kpGbFUUKAZpxUdwBEckFmfa/wo6RyxN44KkWHmWZk9SUX3phBd+csBNJcUabo4ICM
7likBhNetACWrbaKuUPHzBTeAdbgB+Mem3cVDmqETRznjgxnBLIiv3OYwh4HWSxPDWgEV7fwb4c9
/NirdVtj6/ZcW2cpVfFSJ9TjkBUCED7e9TTYQU78J7ptbibZetrRjLziLONIKnT2DznPILiDIZyl
BqkV5mK9XVzxR4z2MMQ8F7xV+3nF5WEqZgrbrDnvZqPWp7tlUbZxmEc4zdLSzusqT/PUn8Apr7vJ
dKcy3N+wInc0bNt5aaasyo+nuvc5DOgZilALIbOTWviVMdifcMAuPq05dfQa4eUB7vWFcMfX4Ykg
4B+v7/N8zpWcG1YidnPzzJx/hYuCTr+AXzDfwxXdHoO4Gulu0TCFoiSJsubUoL2sbKzuXilc8AVD
dAWsWO6pBg6/hsLUlbkmB7jIhlpt8ELNPvw3HTbWtf9MmODjrcjvDtmg3wJVXkOD5k7tV3iTD3n4
3qQD0q0ZTbWiRO5UNWwLKkoy0M3endfiE9wBInipZwFeu2Zk2h7n3ERGPliHZ6fQNnBDoHX/gGLb
XAE//FraNxhE0qQMX50KfKXgzby83pGrQILastuRi3QFNCfMYVaJpr3fqC0CF2+GalMQgZMQFW0J
qNAEUPpNgVMtMhjtGBARz7VnLV3mt2Ot17Xfj2HLRur5wFR+d7nXkwQIn0PU8oUKVSty8HmMC8Qw
44ibB089Rd7Eb0p18wvSc43YdBCeV/6MJIaRYduaCs625oYliM7dLFz9m786KY4//j/nAcCtYSx5
Rh59rUSGshpcozn9o4ZY5HslsNA1JkNRLZDeRdr7Ngk+DHGbkON+lgEND1vluekLzjHllp2djQqU
DyO68X/7CSJgKYp1/oQjwVc90vaYp2hoRVNWVa1uOEI+T5cpgyKsII2/k9cnz1JDa3ZCTz1/sFf8
oioRNxNJh0mVw/xJLm7PA7Ll+CAVlSlsOjlKVw/Osm9SzpUBBvAuS8dRBSugVLboKH2VLf64jOdU
G2D8i0nJISdSAabHgP3/bmQYAIwrZ0e/cpiJWXdUpnzNCI3NA2FaQVAF1bSInZITX4Ney5vrZe6S
Ci7V6OZ3MyUymV5YLBP5t6lyWqkcG/6cwekuDJtAMp62ffh9C1J8zGsi52GxK0IhvMFa4fH4DSVJ
1v5wkIE7arS49zVA7WMH79qJaoSQHfYyCGAm8LRU36mpktP85uSxvZVidq2KfaBUiiz/AP0rdxoT
oNG2EJEsdcADt6B3lSV3rGLULtGFN+lnomq/tOGt7rgMJSmwEiN3oGZXm1/GFLQP4Xy0gdpnN+iO
3Z4WnYuyqcTRf9xHmdKe8BJflibeIh3I82x/38IPULAkaVY7FBUfpH+g2rjQmBR5TlX7lDbRaaP1
qeWeRSRZAr4mCJ4IJfnpnXeVCKmgVQuB+uHgGL7T9qjuZhszpiu8bz0/pEQoYOuCtehdhcwW3wMp
+7LicTOv7hXdlv2Bj4UPDaLraZVdKxQjZPGKZf0dwmoN9cgHSd9E4OtYswPlVmHCbxdRh1lfp0eJ
PX11BZeL1uNkDBBY//rhRe6Y5IOAPTnzLgFLOMCu1LeynAiNELTqQKFDvBBFUNHgVE/0EXnWZdYS
rV384IujyEU8zyE0lluAqxinvR+HtxkhCE//ZpwNDJ4pRIhMO7zRpTMaTnLCsZcxGVH41UMWDEIA
vmXY33DZPDc4J5dUV3oN8pWROo2TzFJokC501Jzf0QRd1ShO0+67PnI8pI/VzThBEePgaXQ8P/me
oDe04jKyrVzApDfkQ8emzp56EMt66hnxBsG8Ox0toyMCGsM0HIhb/dwLoo7oZduxxoTAN4f4rXfd
Iiq7V2y14eJ3J0OzPXmg7XLodKUpWzuAtpPX1FdvdJmn2UP41jywuYHYvJNURT2WlxR3WYU5OdNa
pX5seZo90+MLpz9HFVKqdNh1/8jiYDt6Qre7YVjsw5c64ItLOX3Xq5WKbu30CNZV6KpHql82hIlF
4JgUIKzY/GqnupWwouKvmfSYVy1MFLPyRPhLcD3fmmUq9yWPl324e80AKmKeQhZKxv7OkuUcIwdM
Xi08kNVqewWLdxwAJo+SzxL8LGoI6U58WGdrQ86Bv+DkdFT9/PF46QtChEnDmCSoM8OIaTIbNdHh
zgJsOA0E7i+3OhLkJpXSuRATtAbRbxO+RIv6uTrbvIfVmeUhMn/1kAk83KlHsfKVhAiJn8FScAE9
sSHZpyWASubcjhJuosPmaYoHQFR+y/n3aptQD9xuCGAk5szzCSpdaAOi8HB1WvAjrR4JU5k4DSeN
q4dTwnkaXtwr1RqE8eMViJS2WtCFUIF/z+9iPEzzmpKSqj6TBMge6/fe6cXLZtdTQGTKWdaBPMfO
h4+NrnrxZiyDi2CZozYXlh2gHwVVC6DHinfQt27i43/NGHkifvEUyTZ1+vdyrqJuhO0Op1TP0DrT
RwjC68j6AXAyViyHJa7/QdVXVehmBsBkDx8QsS7DDAKfGwkMFpTSPaGG8QA7dHqq5JiV3bCcs8j9
8JUdulkNRnw48zM8PvLWrCRPhql5JKlB/ewfCCkyfJ4uPgoUO1Uy65cRgOmQbPwnB+21quKmwr/P
EWDNQhw17QiKSMs5wdOv07a+zs5ocw0Vj6m0K8CEe3y8s+clsy70B7vCpK9gz7jd/Qjv8jmI4Y5a
3jBcMBImro4wICUzW2fDd5PBmDixMf4lReTY4dn/dFvT3lCvN3rbSkj3H7hLBUwEMrhXFU3TYyPF
LKL7lRjGaylsLWtWpP/3j7spj96Ukk/vXgRHQ18p2sgLjzA3gg9EMzezlEQ1zqGPdw4xyGk/ewDk
EMx5x5fvIJSEpS3JLjlXC6YewU3oEw8Rkq91ESkD3CcBEuX/OUtG/vzP63selafl/mzHNL4X+aAv
SKmCrw9xJKCC8DKv23tZTvNphBPN9QnD0g5HWz2HwjqNPp4LGgTp8Cn2rXZzEi5cB0Sw5R9u68p3
KXJbfEsxX8k5bbqYzCOfoSbEv8hl1xLofEhohFkYOkhXZX60o9iM409Ttki9lu2rs+I8rXDaRaGK
PaNPNWEySPskV5HvtAGMPfu2rYJ0rH5z+9HUjLqK7LiGSUKE5065kLGG7SOO+9HUaFNdJ/rYrdHw
9SlPtMN6VGzlMtaQuPrpn4PwhRAin6Hy0Z+I2rhNB9pjz/44LR3x0ULEkMHUUSWGQ+7A6+y/zIUL
wXm/LmHIF+hzb/M+yeK6aHpFPNRn4U+fWUu+MPca60MKcNCuTYytXycuqLZc0J7WpJi92rPwCGgA
C+PingE2oGilLan/JNa7t1y/BdlwLtIWUJbKg2bPSsFiM/HQIpbn3X9OuwsuyrAF8Bpwfz0K8dlm
R3B1BwZgQ0awmCtqJhHUJZO3/5bvroARxC2wTWf51QVIzgAAotSrYEgBdmqUeLxOM0MsuVChOcpS
6qrJ/TJTPVsR+Xsft1/ODrTRx10KuagWfPZHiLrElRjVVc50mYJS2jrQUqpGGnomOIf/9js5kdI2
JRlNLWwqZ3kSSu2gOjirKiZ8wsV0hnCSA7EAJNfWlbIkfC8VMU4OLRxq0RWEEIex42e3qrLxvPaH
n0JK6jZ77rWtM+UZ9omhxTthzexjch3Bho4EHa1wPyq0b3Rb7nf3+/vZoH/tjstzma0jkyKhiq7y
aQedhCdAh/w3jI4RgtjlnWKk+2xFjCMNDqlYQAWnxUFL1lQZvnmC4BUJyJGNizAlEVHP6+z5X9xi
5qw/CTUqdBk9aJ7VQLXLVQiBvkX7ie2kSxhP91TrMDefKyp/rPt2NhKPwx+r8Nw42r/UhdMqirR+
gLDIAnUDzAlj7yoEXMSvJyjh8b5sZIUSY7Q2J1+nTCx+U4ngsY75D6AdadUAZS4AVnhOjwg1buhy
0qCeZUeH23fh3fB06SxFBEEf9BWmMJ2jb50McJqkO4tQElWh3FRh7CXu2dcdcMMotEIGx1aL+pym
yB6PNFA5HmbB1BIeafK6V/KfDcPPaShfcfF/r+sTuVclCaLSavncQB4ixKT6dSmmBM06lFXd+K+I
n83nmLYjq0JVGzj/UmXyHbvJhpLM5KXSDNJdqAw2WxR0m1R5SwZljidH3ijGyH1pvikKmZdMy8zK
58luz9YmtwtSOPuhFovvJlD4Gv0x0RistqMFiLy6V9OwD85XPjnLC0Ff+Nkyw/TmPOh68ZUS/Mn9
r3k7l8lDROOnzwpWAvDWcfcu/T3CajSreKRKTzDba/zKLq+ViQ2x6SQDhpPCz1G8HA09jjN15sj4
IoRqX8Q5mFS7DMmeukgE7Baz6VnAfRj2ZOeeY38YVmwHnmdViQRYR+TERYExJtvVQZwdrKEiVJ5T
F4yuJt+6hqriQ8/d/niSyNYcf1dYQPSoB7TXKG49X0sWCKRWkcAL3837Dn//pFov8w5Rjgw+M9Xo
X3ToRl5KRRY9EC8GbLS+NU4dZvEcw4G1SMIvT8j1hs5YaWalbzjtEO5QRFvjz0yTqDDBcwKyTDu+
qjK7SxXeAkARjiIZ2Rw0/Ja4sMQc+XFPjvpt42NS5bXqZCjssAR3uTWbHWrwb7b6HHoTREwzMKN7
J7QAhfuJ6LIiIjOUfyKV4zP/hT0ccqOKH2ECtxID51jfyI4=
`protect end_protected
