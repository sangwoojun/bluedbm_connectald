`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
m9r7E2C4m5Kv4muOcZ0HM1f/DIcqeF0OYjRDXNZo3gvNXUCKXcrXkX+/GGMEh0D7LMh4xO2RCO+3
IiHp04j4Lw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H8XjI3Yko7OWF2rxLOS4CzY1b9QCbL8RrdLfBb49UlY544dSqHKwKDFThay4LdvV4q0nn/gubLqJ
gbS70MyAeVb67eaxuWSs2gNtlOsbui2jlWighqQ4jvlUQCuJQcdMd+p/4iYCqVTOA33H7/DBTB9f
OggtPnVvUMkcGVOirvs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V30QkDSXhbO9t+xnaTOm8HhCzIRwGjmkjB0K0qelGeupx1Oj5Z90aYz7Ti1g+dmQIIv7d/kCcoH8
V0diNpZ00nO43n/ijjeevZpEoGht4JnUK6HtnL/ExbZfN0b2UpB/GjJlYegZPT82pr7dZKr5kspN
TzOKBsTKVjMvWpoNCQBWSheeqnRGcP9wa53wm41U8YaweMQo1jd0KgUKn+mjHIMQjtkegnJXV/oo
V9aIlXtU3qwctlUHftBPCQIs2EOXng+6E0hVwWjd8jzfL7bmdTdaST7rbi3gHBZi2ce6htbSzrFm
93QlMXgeI0jQvMvqzlPsZCi7BFMQ5t30qtU3HA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1STAq7Nds8UxVdwUXOVdWZwczC3R1Ea0CBS2ZRlej+vgF4+ykRc5ow0CLl3B4AYTTFLxp17AYgPN
TwV7gcQD4HKXHfAix76zDT8FHK6mPrB+F1XKwWEqxmQ5z2g1i3KskWOwFshX/dUb1BS6LcO9dfk2
fmykF66fMJ1kqEexe5c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nF3J+LFDO7zOsx0eIWAVOPBat42+rOw+HOoi6+Sxry9otKO6ib560XZSLsQuj7NAuPU7pAYUUCC3
pwlkbD3Gahpk48bTYuF0jEElrkXhxv2emOLJp4qiyVo7Kl7nb7kG9xb0MgS8P6aCAHvWW2rEFBnr
Z8aJLRdheHhnqGbkBYhd6cYvxED2sAVt9ToTNFxnX/DYPkXTbTSw7MPZVnpFffOwaVTer0bRauMx
VQAaUh3F4HRW0UF1Ge87/WyGjmNRboW6mhjDMvicJwFsOpykfPfE3Y+U4M411snODHiys4t9JyGO
PaWI7r8raCzaClltX8v+3HVJX5DjRWo7b7RFZQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 66352)
`protect data_block
3NW+cjCfmJYbQsRfqvkqG4TceNheMRaxYCeqdv2jkqg21hs8xGSY2wduTKoGb9WPh792vg0U+6Bn
Q+Nz/T/PPZmf00eeHd8B8DNPpVEIXALsT4xqu5ZQdA0ZxWzbFIIuj7GtnsQMl8LS0n51g7Ij38mk
d/lRmUAo8Yq4ORXE6awNSfRqgRSe2oNYhxUcZuyEXJJC7cL7Dbi8b9O963FIrg8/Q4H/l+FYwiwu
L4FYRzhMoJ885k1OfH1on6XCPo3k1AGB9eb6371XBp/vagG3AsQu6QsCLINIABN7puD8o0HZuQ6M
pdU60nY7si+dLWIBqfWz+5fDjVSZ6tUbZGl77ZadYwIxXggBRc3Z3o3vQhrneDmZHMJuzo7JKGLR
eetTrTPWZGrxxS0r+Sd9JvZ73/vxP2CL1aveTDzJwg17Lw6FKuiUq9tpcB8gAHD+7IjyvHvslhK3
1zgop0H9Jo+HPoKoJjB4I758pXVawuNyIf/poN8xWMdBoaVGJpDk/SglxxV44lD0Tyu2iHYwsOo7
oly4pOS2nnhdutSAJJJ1+ybFQsJC45MhmbVkP4OlLBpwms815YPD+ZpeM6FP5eJ6YdklovLOjFEl
Zc3mEskT2zEsw9q3X8kDpV96Mo2lQGty0DcV90+zCtcfLcWg+1PDwARzpZ789qBKYtWUNsCB1CLj
OzDaGvYc+C2OQywFmwysyZ6CAEjr6lzwrIm2Ca5k9cMq0b77mDQHrqriKPhfPHhP87R3xltbnytK
dfGX8Ic6H5Pat7LJ3FDinrsG1IhTGWTUs2oDCZv3Or7J1XCnZx7K6xcD6SER+qbCkJZZFXoby2tA
MV4QJs0YTECS90P/0/6HMLW+Qz7i6LeNLeQv8lJx1GulAJgCQ0KxNQqD/9nyCJcdd3jal0VQPvGW
A347nBs8ZDbQRG+ZIt1jPk7zGiw78w1iOuVmmNbJ/QxUlraWclaJKVCW9eD9hAP23HyutcmmQKED
vYVr1ft3sdig7gPeJ3pY3XHAMHOkQunOM7s41487++n9QOTfU6BeRHcOD4f0WZCzmYegNHGeMu6E
zrMDawZRS6dkO/l9NB3GFrDTM8PsusSITMaLu1aFdLeO6RBhV2MF4/ZelggApc08E+Z3oyBkJJ6G
bl81C52tdYph/A3GZDDbMmqxbyqeYJlsU08CrV9n9WzgBBj27OtQ8Dms9D5tBtoumvnIiBQ/p2Ei
Te9Rl+lpikjkGcsCW3QUeGVq5j7A11mrXVVjEXL3PXW+D3RGw2w9T/OMsQD2V9awocoKSEztLaov
kRY6eYSAfBc10T/aF711S3yMRMHd5wTqcBJyxm84DLFajjz13J1D6k7nGnJp2Gy89xxMhbSm9wlS
nn41ZyBrUYeg3XsHoFrgxQQ5zlNW/R33NIL5Fbg6ooCZPudnSQCSIIn+NTiD+DJRINKCCwRFm7lz
e44GpeaRVFh0rvQJq/QuVwjUf00wyfPbS/okiXYUUCXZNALfNxd+QNNoq9KL7XWr5mC5a4WGVnvh
KuVAlj0adx6jEzv4fyuV3QEJF3JRD0LVEfPiCpsJKrt2nM3+lwGxHKa5CcMlrgyRdgGGtt2J8Q77
ci80DKxmBYoBusqWanc+aARgphZ+ukBvLoyfg1nQRmTohM9i2qc6GcUDhW9hxlk2LH2fkrKE4JDE
8TG1D5hRLphQmbf4nQZXgHxzlxIKtVlMQFwwfIEHzpT8sw944IRK0H+SwTJ6YUQSttdol+pbzFlb
Hv+8tBh8Yg7FAO5sBeQt6RMnxheUT4wmBBveaetxWG8mvKjqmSmhsLzDtI6QMhyhNr71LViXqfSb
JzKQ80QeEYcm4Nf3a0fpTK8MyNx4jeq/bEgnfxChpyFdAi/YwLwO4E3MzV3mHhOA2M/CF1b2H5+Q
D7t6e1Do+VWHQSRVSBHc+RPSp7jm7p0f9r26uze3AXIm7Zyyr06hb56eeNWBZrjYAxpJKwoGnsnR
fXFAoyg94q5QP8A5CMV1YUmw8vLL2hw6KFy1cAf3jLZ48QmnJeOO08YpScJMROln+ioWumXZzdg4
X5n7CZcPGYLYKZj0/Y9+teMsTpkWx7F57wx3G7KM8sHWj5eBu2JgSievVIUg5KLEBrSj8iZAa3+z
D3/W/fOALCWBGMe6lLgXaT89sGRq5Zd2T0DhNOQtKhe42gTMa2BtMN56V9ZxH2NZzPYv1ETBwhPA
//FYtxrJaJilwF9M/kQxRnJIeazG23H6UHquiIHaiYGQ610SvQRZ+llH/STPOi6pE/Eayr+dICNQ
sdpqupCsaIi2kktWdKVBrOskbJ4XRWBX3793DSU2HiohGlEsjDXptLnUwHJ6rpdFRAtNLt7XpoiU
9J/Z88q6Thl/BxJ7AdnSY0Ppxb6dF9uqqIl3TzArN8M6hz8DvDtIhneud3fIXhIuf5RlufDgxreR
lGEchi43ubG9iikAu99OnomD2vbNvOCy1DsMuJZjWnecwQj/5t/VJq/CAEy7RKu6Th0C16MbHiRK
Fq+85bKYxt6pGZfGd5YP4DExoN/nutVF9jrKXG0g6J4QShYu+S+CbqG7Tq1g9/UnO80ed3iXmTXX
iOWxRJiCReEFJd1D/HZO0o2dZsg5NsLpQ8fBRgpzM6kwlNA2FV8kgjYER/yUWBfq5N0bFm+psAh8
tIRuIjTF9y4ptrIFbxsmuRxHEYiOQTgHgRBAM19iJOPBfPJBGBfIWGfZw6Q6s0tCY3JJrWRfFuDf
cwxsD633Cm2wZq5Ir4HeUWHex9CTg3lvBnc76WpmJ2qVg8y0oC7OQH/weJcjGfyNhUH1lB/hHcsF
7DWP2JUi9VXVa7QmWeWMI943o8E57K5VfOgqVkAg1WNdnaN1E7hUBMF2wFlYMmzcdNuTbHxA7Pr0
S/lQphicCYJxlPnf+BVlCvwpdRK38+PJNrkAdJN9eCCeQ0H9XNqcKIfw3bOafwQJH+7fB5m5kMBL
lTcRNgxCoE17JnRu3/UADmitPuYkbRrA9vmd9b509LcE0THagGn8fqCWCQweQOKCE6N03mqWV3SK
1jgTh+on9w/9yOIGB2FzEzO4QCjK2d7pCEkIfvDkEiCUFdp7+Ax9mjw3YMaGFHH6RlSfkCW3AjBI
5jJD2Vg5Q5noNPfjQlwXOWWTbSQGzX6wFwDxsbz6nTfc80RvwKVpUWHe8DgGArZBlnP20OZJVy4g
Fs6KdKCCwmSxOJ1xavdgb9Y7FRnl7PPOGyRqUUK7jeaHpeKLTATmCFdMLNcg1d/R3nC3A1QCDe11
kCQ199X7LGVxAKYcvv6499CKF9FktTTFN2WYBraXEBAy+UMM8bph9q5HVVkjKKnzJW3qJqeAwyWe
Vy6+y7B0fDFU1EudhweyOgrHqKq0G7V0R5/uesTWFCIVM4bq8xNjSVgqR2akaQswqWCE6UzwcZ6s
zgoJSXrC4+kQZjees33J/bY1YkS1Swdl3aKsjyqDy19C4+XtKteJYP6SZNSIiSMVsm8PoS8QFdQs
qGGFz3MK7SuL0YwzHELO+gmJJczghtY66KEUc5CMEpHWQdPdFYd7VKbM/4UBg2e/LXz1LyGbD9eC
n1eyBLGqfpun8IOxqYvySgBpQm8hfqrWgj1rnZrSgzRgQ+F9ZI6+8gDKC1M5j6rt1XEdUAtkmFG9
/SKvUCNZVN+E5CX1ai6Ag4Ch2+9VeOn1HgGilMrrDlkEBtd6YTuSRRQtdCAlB7IvoKf/VL6eesgf
j77Yusamr3t4JPj8tw8gFdeDxYSjr6t8u26SdpnV/6eC5VvmWa6hsYwN/7aWaqlxL1sSIR9Rl0zD
5Wf28kBpl0ti7hTVLCubyHRoZwqrqDBpLxvKOi8hAklKUTcBBCNNvp3E3Z6RvIKSBfdcX8drB+jP
rexr3yK7+sMZ6eWz25f0Q7ELlD5PEBBTttvbmtpZGjsfOKCVmMCZ4wQFbX0SUfy8ZKoQC17UTp3g
5t/KwnrIAqCqUyFwIEZZo/RTortfVkF13slKOubBfWsQnkFLpqfh5KllVMBgYpQt82D7SJUJl8Vy
WGdU0vR5K/wqdTmk8MU/EFNFJQNo5QAIehQyhyLpxR944z+nMWGpE3D0GAHxc4X9wvc/rmtaF9NU
bX4Xm5T8+LLV1iZXNY26w5fbHNjvxk3pB4ltONZmpHC2XIkK6GEAddgY60PLtWe0QuN20PZdoDJT
ioEleZcxuYLnMciwsVGye5GZdTwgXmP/FTG/1RbjLv/W79lOao874d9VkjRrbJE4DGXuYOEwuQA3
9kKfO7Mwc0kIVC4fN5mi5hsP/ZdyEwPS97mGEZJ2OLd8JuIKfI7pKX7jJhv4Zls6OnOQ1d481smY
DkM7/6rqC83yG/DJMO3aA2dWKBh0nwuWd0kQZnVc2yu3QBbvCuF3rVTFGZbj5fLAf7Jjvqmfsxax
gzkGjlCnhRD3dnXmkaOyhYvlC+XaNPWLxZ7/BTTPQTwwPH5RU+o4hbA7r6X2um5GUMoGy4jiQ8YH
BBBJEabGpOJXTcVmm9tprG9cZTkychgxn1vVaVfv1Dc2jbqzGC9i4nEAsiVCXGkhtCTQjOcfWpKo
OO/CCMchiED9kxuamofdgqvfqysZX3NoxWxC22DzTQ6/QLi6s7ymCuPeMry2qgUBQOVOPNaMwmQ5
9pOMgBGREmCcz7OVZX2uo6MhyR4ypJxHu9g2DRc/iaKnD5cHaLw6RSiUv4sq78rIBy8qh4QKrnus
VXNZr6DKnKvLN4WJkFZ8Tq309AmWmJygmUIr6I6hw19fKX0FfQqQtED1yhBVZTtJGR5Y8ufnUo0N
cCBbS/4hGOLvgzu4VwhVpR3gV5os6WWoMMjrhdA1+3iBiW0l6umMDwPXm268S9EpTc46QVq0lojT
XlIu4zhaIXFKbR33bbTjPi0nhBoXqqhSZVQ56ewFjKTgPtjBuIiReFH/1E2iqW/5PAgfCkSTrcxn
1jxy/tYk5NLcAqQwuk+wISh8jkxYsFPAKt1X2vGmLjCLuQPjg3gZ27xU/YYHAA+T/BeNBtiPIacv
fhMMgHKhdOhy9mZaMOeM8EOqx5gEXZBzxmnGcBquRI2c15sNnzTuMX6FdkebLPmlR0FAUrTHZJMT
5DfBiX4GIhauqgTM3jtkHu3pkpVhISSUyJvV/qe1pWlWSOpg54nEjJmp744ndGXmUANpRpTWISFB
fvUOZLZycC6kOxoVrpv/x9M9SJqx0xvrkXrOAahpCf8JpX8rlBlEQivUY4aOADYf/nZm3ns5DAOb
UYdbfmau8Xa6o3JcQwNr6uvmfcd+fOL5RteTuFgpMqJpp1XfHuvjQHgsXzZOOS5k3ZLBLCOrRgrF
JeNP/9Y4eM7oYEAZJ25safjbv2fOkPqn0Kl3nguifwnSwtDW/67iTTI9Cl1j9tfOHdZx4CPHd0yl
BvdVsn+ae3OpzeY0F5SJXtSK7paYSUGSz8CACAWOGGzl3ITLcUUOR1kiuoRV0Fld/A7ORtxYEe3l
KxP0UhbltuXi/ZypncIuJiU0E0x1yu3hAM0kB0shzS0JHV0msTc54WmhWkru5CzX4iqeQoLwBq4N
BAbMtVV9O5FDDHgHyzsAoWKrb00rrQp9ZTXLoL0ouEzjlbXNQinigGN4oo7vHFUnLen6jkpQvvxG
K2diO2uwzMCaO2ZvTu3IKnxmVeXhErlMyNskJ4mmVZaxaPY0mDNnAKLx3Onn4GuJECOxN/MK62Nb
BZ4aBiXFXLrhexNhBswUywbHR1hzmqguMcs0S4fa80ZP06QeT8W/TH6yR9va+W29E0TQLJd05ebq
6onvHA4E0E75oqrvAlFbsVQfxs5lsHsw8PJakcBPaBSssjw9O1zjd5sut2/2xWWzbCY/X/TlIN+A
LFadfdAmjGHIXkuxQujJAEMWpKeXLNV5UmTZZ+8Add2v6aXIAIfksotEGGZY4rOHUGIjwxjTuyDf
PWUdIgKyP9aKd4eT48assUIsqc5eUQge3eqtCArAMQOZoCXpiI7OB9LYOZA/6UB2EvMWlCYBY7k+
5Ei3joWe7XF4pFegkqYkGwyvPessprnlAangC2g/1syOv7ns35AVf6YWDPIEPThKbAWgXRfvQB/0
pDKWgpZso/mMj2gwvP+talArSfReDhWxpIh97CA5wnJl7bqC8wXdys7+WX27Sx7vEN3qtTqAER0+
rXwcMyIHEbhbEl/6XOg234rpyt3s/Lfmrwn0D+Bvkp23Vbtc/OaNhADGYLcT2ZPLIrGsEL7kUk8X
VFxRr7xvhnnjmF7grjg5PjW6aZjwPKUMrMXeJW3mP2dc7xHkYlogmtpXMpvq+fMjd9lFvgX8azjR
UCczpkM+CWsfn5rfv35E2Zjv3v75AW1oM25M0C1nhqi+S3klNzuAdMONwEJ+CDnzD5jAumu5QcY4
j4iOQp9bwwpM9quktPxkjWvEor99a/Mecc1CZmcWno9VZxAgEV9H5H0J2hT7/i/6KOUWP2Z6Xgov
oIm/2MKiZg2KR/HVvfWGPR3ORumm7uFE+iBUbcL8YhVXyasrY//2xYP3tUyCzajSCkrRYQ84e+dI
MhWphtRHp0CONoLfBvNCn3TT5h5rjVNaeVPKoiWfXpxzwb6zRo4kMUc6IKXBOvuU0ZbNKk1/OTTL
tQMvyjmg76LoWusArrAxuvcUd8SpkuhHhxsKI3ygxpI92w5y71diwCtn5lYaYcIDjyXU71baY/Jy
nm2fguf56aX/8beW6+rx5Y+f0kGYq025ntvjiHN2mNqnuHWYAmwPqG6J56VDC6P68TBLFQJ7+PPz
mztNMwCjbW++/+YZQfZ1AIbv5snmbbXa1lWlXZ+Yfh/5HWoPERtGVRXTOADxD2suHfi537E+CI42
MQKsU/FxaHQpZOgYbLry5fNkrFWd/lAjgvoDYRI80Vs1uaMMtTTwNKxOCbRQBaxyzRDF8UWMF1dO
JwudFgf1v79hwhEq4+H4HHFFQWnWj0cQn2IjxpSWmnqmZwlc7L88KFBZlmncDr+017QpIG796bsc
gjWSdG6zEgXwOJKv2ScFty2zqyoWRCg9HFcstEiz76aTuEXwY9zJtWkICplmMkGuHb/Cy7QeiTm0
TmexhtySIpDp69cxa2KtK7reCWMcsy0piz1j20cT1WhqyMFuu7nxu0RNCaRv5jAbMtwgmsg0B9HT
1R+kYqfRirbv9+IGKdPHaoifwy+Rhw3cVvVZ/kY8r3ArjWjE17wvOT+pcH+7XS81AodgEW/vuiS2
MnfPCyLNCzosrBw9MFy6VSj7Zl7JvsJ06BJBB78qW/90YCdiVHuAoxNAySRleh/tMpBYbsayVLgL
+1aUuv8qmfeC8Lw7Wt15Um/CSb01PwHzA1fmqvgMJdS4czCjiNFXJdBDF0jHeQm70iejSCovCL1o
6kjSyCAWRiHC4GtBT8dJPYbkgX1aovYcnOazK9XjuRVdO+9NzYBDmv4wGaDEuyUYkucW+jQboDnx
+m7/ZeUGJjTSMnQSU/14udrzS0SFpv3iWBs914SldquzYMPDzPnJ1K5+WJT0hAP0khV9H3wJmdwG
sV/9E8N8fWGBsQttfaWAs9nB3g9UeOc57TStyOO/ghE6/SlwGoJY4OA4wEqUy3be8Vg40oBw7rwj
X7IFdwSErYG0QY2Y5UcQJ6AkSc/kGuQS1ygjYJvJrAbcC2bqC2q/foCAQRS4L+HoBgd+X7f4Kdnq
NNTa20ozeQ0QfQrV1j7oyCI52bR5rsAgzDNeJtLDQKQ906hlFnLWDm8E4GX422Do9JVkoHj1MaJl
3SdtO4guF25GzBUEFo3OL0aJTCMhXhfXlQg0RsWR0Tvo8AHZERAKpdbWoMCxB5YXAMipE45Tdpfz
CC+oR+BUQYM6SBRcpzOOSditLQvycmeuv9HwTqIFFKQ3Ey4CCJObOLHUHwBMyBD3uLWXQy2Q3p2b
6tR6SNMGR8Lw8z7uib0dZEDyM5A1uI8XS9nVR4cm7Z9K65wNIw9OIr5010Iv9NG46mdDo4Dm1aVB
42p+jGxmn6bZhc4jOUod932r24GNdQFqRRAnSZqAnGNVNTtwmmg7adLNo/MrQB9WHrqHO+/TOGWN
i//Nk/whoxVugrUumfxR9+srsrdR2wpXt+gQa2OwWCK43HTx2uDuw97BVX0R5R3+RwTPklKyYxtH
HoOMes7xGw5aN1ialq87HG9Fbl0LoScOgGPOiHspOGr7+PO0XcfZMOGD/A5n49HTdTTDlbzki6yh
SOqxpQJiq1lgoDcnS8DSRLfOP7NFNSIvotLyLLDQg4CPycZix+TYSdXVQY71aAQQV4F+2oDLHIIz
PqMWjnpPkZAUK2/gYck+ITbE5NExZbMa9ae2NtCmEX/u3PGwWZruBH6Xy53CDOm7xuiQuu5kGxaG
telmGlefSizZ1prEGSuYbED/MYwTRrNLThk0jm3eJ7++6tzMOWcRDwR46HHdZsNCbQ5+ODXYwzI+
66M7SnF6HneCYg5lzaXr1wHmBSINKTiQNcjo+ca5ZPbEvllUqPQU1xVfo3UrLJylW4OYkcBcj+qy
TzV32ulQhb2HtpV9cKvIakJ8s4n5B4ZgPTckq37/qUT7LXMMX7NtkOzTfGb8oybOnCED7WQFWhX8
ok/cs/eTN7ZKKPqBuWUKGBgIV3L9UOjwwnQdQWF7vbNoLZdP4Xh1rOAYoxU2mw4rbausMVeumawY
6/l8s5njvBEQUPaDLyElMSVu3hMPNhJ4MhpHn74tLm5rkKLCcjAtjoUT0dzJQ5GgmQHMteOJsyHV
d6VC+7yd616mezMqMj2CwxHzKs7BC89JZCEhRFE/nSuP9NWzjbUT++L8Wtnp8Yjp8jHb/ovJCa+J
Ccgp37atuJVwySsmccWa3TaZd/3R2iA+ddNVgG3jRIM0MtIWeVBzXwnj+xRZEPpdEgONvTMTafHa
NbVoauLqIPkaS/vQ31NlYAllfT91ZVf/KZSqnydQEexZvtftUt09waQLS19r2XPQ0NQQXcfgo/Pl
7oA5Styt//jooyPTfv7yHLyjYuBjWMCdhR5/e6HJ27aG9YqFEbxUHDVVEuVBY7w6PxD5ToL+tBk1
iO61Xbbu7Rp55VbJEuSh4h261j7cfEamBvQzO2NL7WAD1KNZhfYydrH9qRRMZtEYDYh/v74D583j
cQcqHxrefdtQnYwHEY/aQC4De2Ain8somOydx/1WhjxFu3OdzyeBm9ZZ88ylDh7VsJU9WOhWwxgQ
WwAvbTjdp6LAEEY2vpl1LkhWgT+vcZeFqHgeOKUIXDvWUpvsYyUVA3hR0dRv6DozrntyEVf27Yf2
IflOxb68Xb4d8PGIzsVHOUQJXXIsHh2WA7hpOKC7uEOS0xEyi4jtLjdPBa6vMbm7yl4X3h0PxNRr
vJBbMZb2MGYu8QblNc1CfF0Yatkd6XOv6DqM/t7tL6ucvKnsJ5uuRbMjVidIp/Ziq7kQwaAVczLX
ERPX5bSd31rjkhxxykrsIB6z7WiyDzGPubvyGx45mdqqkuh8/brPMgYJ0EqJNtqfefhjdLx+W+nI
ML/rPFFrBFNrdfPTBDV4kgceKaolJ3FefAhyfmjiE3gxLa/IIhBfDsFgOHb8ZdO9Az66FcbbmFDn
TQp7BO4MMEXfy5aqs1rl2cprDpCk9dDokfhzi6mVA8R5yxX1RbIAOofJYW12n3wH+GbiFsYa0ak7
X2M4mYVMQ3MHY3gljTMnNpWx0w1QvExbqJGIOioiN6svMl+fDoofy5yrcJYyF318oTNMSv5+LK4X
iLUdbYLgbZDAmQJPMmoQxKPQrS+MC6RAx1+b1KLYHNv19TnS+h/8NJplHtHosdxNfe+eIts1MB56
r9ymLav0fB31UTSTVOll4muHfpqbZ40N8S9SnYeJrv6IQ3jVyhj8F8u58L3IZhxn45LcfD3esP7n
zgzq/yUz9/ZzzWee2MD16ksVAGef1GTk8tUTOrGjfcUrZj1qsZH5mS6VJHLDq5tCXwIZF9r5tXH0
08owNO8byZLR4YvHcxgIQ7s7lRhfdzOKDKf6KuEHGtL/tbPWqM0Fv2FwFQWmBEV+kxZ7JSEi5yGq
k1E8oj6LM9FSknEZigQOKgBQFEsDl8vhGOAgLn4nnyuQATTYNkemgmbxH21SRYdG2L6eAraVbpkb
mncdshIp4vcrs+1Be7SEBylPpITwrV1s1x2CRjCoStkC1lKINgTn9Ry0rczQJ83UJjAUwJDZT3B/
+AcLcmeTdXHOwKZSMf8zTf2lNLes06z8lvXW1APclwex7fHLi9FS0/+bBuLoYe9a4PSekS4pYT6Q
G+IpZaCvo69cbdSfoMlSSxOftXl8zA1KLMXGlWKDb6bHD8k2QoFY7TD0/4GGfliqk84bTtr3mur3
ye3MQ43kNA0jCqO3Toojc2flhzFCgliWHzdo9fItU+Kg3rHKoxmaTRb6Geu6w3Ou4bhr6DIbS/zc
6qvSlZo+C8rcv4VjAik/Gn9DED64qtrYI1BBdNF75RGSE6kC2b3l5xmOTN+/hM/LTdAMCwdpFmT2
4ngCIQ23jUuxvzEhJm8CeTwv5NnNPnmnYhWjuXFNq3KkBqISFEd0VeXqWWVnTDFrFUJEaPvRZ16f
BQx1ejuZWbORXZPq0/aYLWbN5aumrtIwzaWE+mNeX6PfH9U3tHHtkEavxv2nFD4SCtW4q2Y1fVda
DiyDndNwhHaR8VgPv9F3xls6xL9uNXyyLiuSw29EU8DYFS574a7KruR/lHr7ck83rjO9DsX/5Dpd
Aw960Uw1XffmylVBIakR4GPPvE1iAD3U/8uESK7KJZUX+CDoLIC4nq9a6oNV1GPHtwNEBGfWo4Ca
sxHtDg2tbp6fjQ0zkuE9xEy9tQQiirRfEFOpq16cbYzaqaIcYFh9fj7tgySMfzNdqHcxnPzul7+s
YOOc8GR3lvcPba4pVOB8dKtBO3aKv9EwYGI0DKLM6Wxbv7Yiiruk72LgiM9DwlX0TPYyvXU9Nulh
rWEh8vtJs/6cDUYbWaznXM3F2M5H9PWkPaguXnjWb5RbBqqSPHJui02CppPbmMk7Ua+iam6Pjp6k
cvO/Kza7e8U+hCAjWHjSDx35GTLTEXzu8eovnYk9Puvi7MO1DMVs3xu7zd9vUEFWlxc6quM5QCkn
6sIebYUr3CxelAA25RoS1fZgI5Ui/LhVIGT6rAa10fhtAXUlYy7w8vV7aNreOfvhyFtuFyVaI9g3
xJxgdSZc8Ye8e50U7dv/49lPbnQcrfc4S83ilq8RVFUrxkeRLRnlOorbNVxJh2baCUq754SEGt3F
8LBpx/Ev7KS/uG6ZQ18hjeO0Xp62Uj4iBQ4eK6PTxzOTaAAbQltBSrkmRl3VAu60J0b1d9xkdwcB
+syi1hYgZe7icb0Rye2KbJxOQk3dN6A6RJZvEoIcZvMV29ceaYxQUIB/E3MMDzvBxzG/ILtj/FP7
DxQcs/fNihduGUMGHBeWynbop/TniAabrtSa4LBkXcsdhftNyr8B3pSvi0Xiv9C7Y3a5Zup+v32F
7MKAZTeH9rqAFtoXiJRl7dv/JOO5cn47ODJOC2qDJjHpBBEfCmD/g9JgxCdJjRiYYrbi0tYJsRDO
AwDcnDIcz+I27PSuYYcm5C2jTnjAwTn1uGOJZW8k3DfJS4JoyPaxPn5KIWbPKyd35+iHvm6ICXNn
Wna0g2gGwQEVysKnb1wj+yjW1QW8XQODbCseCzxDb940BmtUn828yRXKNln30SgdvrskxytFrw8S
vDcabNIE0nKNTOikAmMXfi0p25SZq1pbE7DfsieB9kALLTzhrTdHQibl0jTkGmYJqX02iWPooApv
zfXMRYS2t1U1p0Xz7bN32qzt84XfEhMzNt/IlCmAtwOTEQn4O4dUiE9GSItHo1zaQXbewVXS131l
u/4JV+uq2Nt4tpSP7BmeEDSaWKxEBPNlcsRTHHBy4gMPEFgx+iaVdP1hsH6UqJ9FvP7yF6MmwscD
1joUTHlp5bAHvZBvJKRUALNpj9aTWzMmyY6eKeeJg/sgzDUgWQ5Ox4u4ogrZ9NV3P5QUZyMdvzOT
8XFuv4AunqUbXKCk5oRXrJVX4DQ1/AZo+xBNTxZ8NwTbwY8NDbB72bln7A6oYcZjcO4zW0Qzl6F5
onvpTTT4O+TMyG6FmhxV6LVzCvgZZG1VL3ue6ve0kYPheG3n612tbBZ+LT9eEe3aH2lpAmrKu/sF
JgctdFwJ0HRYoWW8jjocX3KBrK/erdtFbqJkrGhz+EniNszzT2qnuFvAkaSPXKI/uo9jXNoJkiBc
aZbTKQJVZ/kcuSwYtgF8ox0hWX74m78E+iGZW9DRLCM5WD34vDH7PdhHCGHznXRGcQPlBaNI3mNT
CMewYIEwOMDpGrEoG1KOw8ScJi4P/tmi0FmDT9+2v4IAlTyYmCg2jC++Xt6BW+hodTssg+sK/HrJ
s5/WBwWipmvfsaFKa8cX83N0f4ngWWmbHmYTMLgcm+ZZTpABEEBNdkuj74jAKQ7HNWDDhvqMgRHc
l63vT1S3u0BgF5O/bmXhO/e3Jb3rNUUH9Rh6+kVshQW4t0FTsTaCfRVZjdCmMd6WVvzS/ccfw7Up
hox+HlmUggAE+SD+DbO6oxGY2KxPPxiOk0Jt7qmeJLSmiHPmFxESqGiTzYlGCws9RRS5kMd1rTNS
Hdw7S/rPAhpfAfZkCGkqTEn92B1bAjM3NvZyHIv0WCWLiHF0E+Hl1CX7ICxlqchWiADJtANKAmt0
FStb8aVgKY2ns2uUkURzKRGYwTX9/jKqEq6tPpwfRwKU1NZDne15Yygl/hr3pvTlCG3TqYd1kyEv
9hI7ax3o9bCIeNFXGE72vDKa3kudkjAEOwh6myTwmmM5hsxFtSouVrVK5Y/q3VhhjDKidwgWdxsL
7SurZDUyHl9G5nnP7sNZMTX2y2pHWpnMp7Ps2WATrohFBWPOGDTlH99GKgMxFSagAKUkrxR2km1X
u4FQFWhGbrVpmW5JG8Jd6hzxPz76LQHiZ5YKBVLTHlMvrbNnabbxd2CwS3aUNXEINCc8gAhzbKhe
pFvxxqRR3jGEc8zTbCy6pXJzXGTMMkiWrfMRzrf9kLXb1KCvuh1xBx6zET466piHjZMb49NQhM1C
RtEXvRmwqQX4HOVo12MmnrN9DqE0cgGg5a6xNfyYbo6QpyYGTFyPwGbo+cNsbQYB5R/DmvimrOos
Luaa1ojf81vG+3MOJWpcSBEpEOjqybZluTCQ1AO11WjqybMGntlz1OFqfJHfSFwGoloiabDB3IGB
xz9fS37Eg8N0IZEdXzUBR16tJ1/paaMMQdAJwXbLFdkDQ4FbXSRLui8jhJAIy6Zom8+L6NhWaEsn
ZTeGFw0ZJHs3VvQ919WiAfDjQZfEcJnLRTj8P0N9XLwDPpTJz/sw0UfoQOXQwuA6FImaZ42bWHGu
ImKCQb0rEuan2PSJcQEl8ZpIZeOB7QCCsJ+AFLJe9a5us0GzdtNqaaFB44/kTNgZGLuoDPlBwDpv
1T61D2ylOmoGcVE/dUe27EZ++cqJlbEQeXJ/ih4vNkCen+xaP35kLUwrkfQLPph72tFcQRUr9zxJ
3ZuBIvXSsKBO0VmorckA7RoVk4Bdhj1kB5Fbuf3gBsvCMsUR2fDH5eqFs2ZtJaAzDvsdmOgz2a4c
U0DL1QI4CI7pli+98me67nSZ7+tT/0XHEEtZlr9eMlFOKjjBSDnKXmZjpxfG9iOp2/Q5JbwNPtix
//qNadD0cqE6JwdETDJtGNpADcdcjjBKlO074cofqJQDYm3cjaN0sEC3mHg0IeMHN6QSpnFq/YWy
Cu+G7JTPAnXiulw6rPrHpHaLVsmv35ubrXkpjv1QL6ZX3fUiihXm9Vj+8x3l8JkGGkYPqpptfQ/S
cFmLpbpztEI36eH7HyH8LcUOyPov+sfFIdGQ8Dsr9X8soOTcP3k56k8iAQcF3luvFDrGIBwOXGIl
RPRsU9uaFceAFatgiKtGALnZgISn+hQ6RFWdYqGWtPqFZAeuxeTdXC/AyGXWDE6yIKaPNEEd4RJl
ATIgzZzNYVa3ljndAdQLG2lwaICjozf8NO1vHl6Zl3+GqdAB2HsgHOffZ+vbgTXRPAaP9uB19XRh
6u8A2vbA3B4eJQQPx5qK9Ta1LWy2bPolM/En4NYdO/XY9fv5Mgtw5v1QBHjvgIgWKGFGv6yOOrvM
Qrdl75J0s7e31N3w2yqOSnkIpCotYs4CVExkOsAJHRK90X/2YG5ixtpFL3obYqiVu79lujh2uXB4
Ix2qyr/t9qQ+LydaLF/kum1MSeY9mgjp2MX5DvjOmuaeh55iqu8deTC6XdoNbSnrc6+ulZQm2cZN
77SMjjGMNcWScyod+HTg+7ql9+fD7zTPYpFUAJ2UL1A6TN7SCP8ik0szor1ok284gRzE8mbmh+aN
M1oPulmVk993eYbNUqyLx9OWv4drSf/Yf1XYksRYGnIIsoXx5IvqFYgiEpUUiKtuAmXuOse4ua6h
2J+3sfjvELBrtKmt2U721F5YinwZ0qM5alkvPZkwIWuEniSqKgpXgqJyZ6KpCbqmeeheONR1CEJb
7e65/im/cGV22j8vW/qMP28FOveVssY5XphI2RU3/J6Obs1Hi9I8dGE/XGN7hwrFAzMKgadCZVBY
ryYdCMZ68r4t/knyCWPuXV5duWc3EooeSSvHjYu8XQRArjDRugrubl8QPcfz4a88S8UnGiaePtBK
vD/UXUYUwiB9itWP9fxZj3REfrj2KPv1lBbf80/P3bkz+se2wip3tJ8OUoJUD7s2cZqkUsjEa55W
XAfiVwa8FgEFkAE/yaUPFkZsXr3XecYcVgJh6ycMwq1bxDzQ35DOH2zEuAboR2VvoXsqRXgPQ+il
889PS5KRhan6II7zgYiMNHZROM5eaRpc5C5N7+eT3xjbZY6e9P/tthLtE1Dz7OrFXp4muuDvPs8D
uugh1gycLX5+zDr8ZfXZdcNLiQO/1fZFPEuubMUsMjnqOuElyY3OOjp9VeAaxynNr9YZojLlQO9a
gwTBjC7n1KMQXt3IEemMy42cFaQL81cPgTu8UPbzfq4vA55hEn6Jq4kcqehKoIkEcxknW+jjv6by
Dd8Jn4KXP4/aJrHal+OA1XtEjQ8bhBBYML9LpUJpClL1TL1J2U4V7F+x9nqDhzRrXOIcZL07ttqu
ygAdsT08cNMg7fUqAyZdCITc0AvaLMkjnG6BL6XY7ydHjWcgPUoOVcHm/gtAqz1109GqvtW3qXcK
Pj39CbYh11jdOutgIE6h1xhGYURcnG7e8ptjyFm9M2atRQHXC78j3E1cJGz10VxviUEriZi0V17U
PwbdJPPQqGBdTXO2FfBiyi5urL7S42UldmxNV/sGU1uBPr8p0Yvi6c8MGuAd6gkwvT3etgUFK5IF
drOSaIXUuK1SCVjbJRUJAfLRQrjvjgQ+m73ukMbLpiliQ1BZJnw6agq14R7GEOKkcyAvNqzHBL7M
h/bhHpMK1tGt0+lChKcmubXyrlSrwl0E0+f+D1WkSj1QCbxWC3BMErHsHcuGjS//iIVe5t3H6L6p
+dK6dH/pkCYQ/8TtRzBXwSUSpRpksKLwUf5FrkJP8SZMtczolV1JV7pGmTUHgeq5N49sFO+c/Mvc
Ncx7SR3jz3EYLyHcLfQY8+APrJ5FFFLiabxDe9wEcLbwPLIUqSHsl3kKWqSwdB3kMkCt5ftzYTMN
oAh/bghtX+mT+D8JxDs4Neri7N3YWJXI+XJYHjUSRQUdzMm9FMkfyUh4HfmHchheoAFqxBYyCzSq
nNM1tyqcSVONeTXjzwy0QIDEygPoRh1QDNzidq08qaabcZokrZ/zTmSsQlHNav/y94aW+txYu8w2
lxfD7IFLxbNK2VRNPHjhhJT8Yv7l25RLEoYEjrRBAEBm/8wY14A0dqpXQG6Vax+8ZzSi2o/GGQuf
ig5GsLt2KIcC4GiKMvL5tfAJG5RYl6sbvSOVc1uKQ+ANNXA9Evoj57tWCrTIWtJkdhj20TWCckzS
XTZDMwyh1T1mKlGWObkJWiD0ixHTyyEHSUUROvzh88TXWcDz2U0cK+jwH8zkhAdgBrGMQPr39g7b
AS6StbKYWdUiM+1kxjOwfKSLuVJCp8Yx2cgWeEcK6ReSHJreJGk+PCRN9RFM8QONvNB9ezi0soTB
tWzz/9RYqjDfzPMtqRwVYESIo+lNhR9bWVXhTjmSpL3EeI+hesNPJt4FpmiKZBEaFNeUBAmk5huU
PSdCK+66IBf0sVkCeBzERCP31v6g3CB4eAGJMk+cBL9AoCUWDetKgaf7ELx/bbu8yNTWmcdPhdGO
VmBagVASppzqx3NzvThINUO/Zs7TmPXPVYQGU+tUGeKbfQjvIUkJ1HMPhbX6hpiBx8EE/THhzPys
KXFRC0XHROR1zM6QFGX+kiiixazGsgRRAq2dByfSCe+Z1CixBIZdikSAblzC6qaK9Fd5FKctXXqC
ZYX4M8XSabA/E6KBePh+YWd+df1+y14JP+3H2PgU83ZB0Fq0xR5HfDJK4xxxuWcXrTg4Zy/8wlrQ
d0RokKD9mXfjlAcAFHxvC8NQkCeFk82vZqK3L9MtvcFghvofrCtStqIaP5XRA/eWdI4oE4B1coOT
gS3n8dUMaUcjcyqxcZWcsYR1JFc6mzMIqtjmWl5qzAjFf/Z2nCWHSaSXpRmTyNHdBdTFYY/Aafll
k+V7nd3mzOv4korXER687t1SAnEnayPqlnEiwDAgxs8LL4wrM6XQFIXIL7pfPFQAn5sOx4/3G7M2
zIYZmA7eslfIHHPOZL5SXZUO9FnDbIA5cf/gENJWCO+RcR07IJHddgDiU4qBD4nQVW/3OKIn/pW1
hiBeeN3X4IMtbpQlqBvG3dQJRfJs8we0134jKhIQq8iTChlaAVg9MTa2koJT923Ca8xhwJxMPFzh
9SCaec5S0uSkz07OBrgEmcrpSGccVlU96qgdOWVKteoswWH5ziWCOq7E/kBu/LyW9J0v9cto3WpB
ctZGz2f12a412ReHBq6jT0uAfrjnjNlSMlndtXObLboYDPg/RT0DpGj8heKOIB4BIlKXugWH1cBu
Z7eBSXXSELNEyOZhZNGPeN0SQuA2PZbrL29fObQNfMfe+4nY8zZ96AvFTil3XEokoUUrvFlM1ETW
tAs+b2/QC5GOCIzJi2jHtYo0SfM4myATAnB8NkhHknGMtTg1QjPin8nQ99uvYATQFQ4+x811U3mY
xQJ9J7yOsAtMxDutJYXFpFKa3kvw2VRKJBZ6pDGfMfmfoshhavrZe3rkKBwTrUYrAnXu0PVBYoDg
hVHWa5OMi2zOjL5agC2fUYP5c5XGY/XbPNuDfXGXYL1vDz6lyPNzcR5WkU1acPBPAFgh6NyPKlTf
kSSt/aM0hNJ6xNRHYwA9Y30JFmhje+jdmBmP0DwbihEtL8QbSqPBSZDokCa58XDQAPsc4ClLLV0e
BJ1CJZApkR8nYdOFIM5I8+Ipom2YmmtCuNS54W3U1cVWZZUdt8imRXJJPesqx43a0/uU08SUZP9w
pMJPM8PgmiQlAAb/MTPzCSBXz5J1EKdpIzL5NrZaXTfY+h6U6g7loV8/csr+nCPg1Zu8zAbm+faB
ENR+3i4jU12/AHRUhZuqLYOleTG46gchgrpAh33oyCNXNaQpQVmhOApc72KM02ibZuKD6yVnxeX7
4oeN3txrG+0okSEBQhQxq/8aNH//uF53MmudtT5/r5GHV6L+3V5tOWtTVvEJGApUWA2sQcKGB73z
+Ki9pEc+uTZmfIvG48ybVn73LE5FVCeDhe+i2zNdhNSyUbTDRkQLyJEigPD0qOxcTx95fap12jg9
QwzhkvbJf2SYgrBOh22Xn2g5/8Xjbm0mrUMJX1ngaJS6fanOeZGPAi8JJ5Hb2y6PXtsMzbzMFf9X
zueG+4h3HAUt0Mho5C7J5uawywbQCNwfC5towUE7BJxKJEofdwZq4HZ+tHEbkj76Mh1I9enYrgit
7HsFBqIeqaiWbXHwEMSYwwmiuZjQLmWCq+k7YD3dhJQUb7uIyR9DSwNEPZVW6kfG3QF9ks9AATuu
yR9lOAofd1HfG1OklWGTB3aIBh9qXD+RF2NtiyrhBWrG5QGh/ryRS8pEJuGRWUz9BaMEp8QLRa3p
cLvLdi1cPKuYi8xDml7a0OdGlFZKCHjyxu0ZmfevglrpaWfEVu4YK6EH/ICmK7F2qVFrq/nhzk7N
cOqx4xNW52Ji5Ic6bA7nexM6p/DVs9YyoEGO4C177kcTesNj7Y0/hYXh9FOfqRJV3w16HO1BP2MO
QGXg3FAKxi8XlvyTLO5nBuHghM53Vj0AlWcJ7U4QjZQraYadoGMTrw4/YeXwuUGJcvaeMNLVVXNM
ZWgyPW8G/+uSIUI9mNkmcZcKig5EtJIlUKyrQqxrT+Rn8r654Pv+fXmyJLh8ld6hyTTwU7+RxvdW
y/wYjw0J4EedtKudt7//LSn82DQBRf8+4st0+rEayGWctxQyhO4mWAlJyeteL0yGwHM+pIB3JzJw
71YlX2xDXNyJEhfV1h10UDjImqaL6bK7cPOUvTqClp34s30gE0QfRahfRpkFmse63hsws26Pb98+
IVEq6rzMgDqHqlA6apn7h8cYqzxxMs3VjabSztfSoBHHlB6TqXhCbaWbBcSNqiwanN+IdkSMqn4s
YwcQbFjAXPP1tnJwYk+usMVPgaWG5oBrIt2vMfHS0J94BnDMVg92AMD7dqeg1UP+geZ9+SHWyzvd
uyLB4rAxDpLyMDUxa5P4ArgnIQW8Oi9qoNtVFcnDjl9j1UwOjsmH4CItljrK+pDXVOex4gXJc6RO
lEC3idmbBL7QcXdyNxwV0HA6xyb5HJMEfz/3DDsHr1TJlIMSSThiS6AniFcIlaJJR//noMyg5ns+
njvpMcKtw7m5ISu1PK4vl3oXjudcogV8662LwwrwMGRHDnH3VV/Sb/JqoyDEyLJWZe89EViSH1rs
1y4QQJHMf9fwq5cYnagc8ctQq2eSeuKoN4yPTD92aNhG7AOncp6sWyA/vFzmBZR9X+bCa9alULXp
JE5H8VA1FH0hPQigjOrNAlP6L+XKMC97XfeJmS/QT+uM9sTtjts2/jnSnBWjqWJ+30J2orhojkBR
5yGGp8BZCREo3VXd+d2X93XyEStceKojxdyWHIEv5LYBVzs/LhGVQUCVDA080pYyqK/KwdNTVqLA
wpHaKMJ+Neivc2CAm3oIiuJLdKseIkQlbyP1lOEFsAOn6c40Dr4wOYMqV1h3JYf2gchJQ5WtaiHc
amkBZMy4BPGvjIOyn+EQPUQ9tUPHIkvzVANlGpSLdsYDaTrHabfbWbDavYVsJWmi4E9ItqEWiJX6
CIjCRRl4+QAywKWZr+PGKubF+5EyWDP2lZTLtHsxOxyn7nDiVS2M7DPKleLwFBdTH4kPlN+3y+VU
iXQdHa1/bsGlfdgUVsF1xUaNEnkGwajtpoDJLc2T973djoJwDhFvjBKu4SrgO/PmCX4hR0F3xOzK
gVFXyjnn41Gnl7kelux7xMN6HsBw0gQpkW8zZ//Ftch3n9RCMfC6ly6pW/EMTq0QlKcMpb8atVOR
X4pzucq0m0xZ54ebI5+i9HQWO55OBJC0HlBqMAcNjkec0wLX5Fqb0IAfDv1BTbuXIe/juB0ZVKJS
QTnufXK2wL+okH2HZwcksH1ZgwkxHFEG6+9JcD3s/nsvtHFS8IYSV9LoVpb11Eo93sEgIxryO0ei
H+o4Y5d/zoX6jwr+aomnGA0OQ3TjsRBxuCPiQoyKqZrvoO12er4xiLA2UvwGLBGr1vM8U0/zgXyW
Hho9ZRBhLaSwpkJxB6h2lezcX8tSelAGSL92XF3uDPTeQX6rtXvhhVo2Sez94ysGu9FZN779k55z
/5wn6/EGqOmXPLj/cIm5xvRcCUNf1D5sARUbymbbUeTTiqLJMwMdDNaaR09qs99rBQIVC38FwOhu
HzT1EDjFJJs0OnK6g9sLu+Pt2P+S9YuLbZBOWI3hgMNjeWS15M7IhmVhU7GXBgdRX48NccXqHiBy
pR6A9t+wWNndXQEJJs/IhSe4Hsu0DZ/qOO68WS3enS9nUymBz7H+ev1pJmXlf1utUn1ayruEJg29
kM7jLCmuseyCUbs7/CbOSdfzMAfUGOrJgIzdoUhJz8ulTeCNoPOfi3k4wk+O7e3XLaZElsSjwOoB
xh2N7Y/uKRvpo9bBdgry1QM6bHmY1s7xybCru4MJNX+WU+SpKVDMcQykjlfvcDE8tJdrhefgw+Nl
+mxLxRvdnPLOEGx7pdTnU5iEL3b1T93ZdipP5IxG6qmwvMsb6CnmxBBQoQpH3qpvdSPgOwPAt5Yf
5XB1vOkRNumsBWEeUlM7kANLKEnRnnpiVFOKwNI7IbSFN3bm72ucIQ0upCZiLifybHaFDwClU+gW
GMilU9Osme1C/P3CW44HMVhwoZMwuacOxjX35W5Mf5J9eGfMcdxAW1L8aCowE5IXU9OpQZsfHZS7
cxDslDjsBlV8s5376EaWHUmANPsRKhusQvmlKsd01CGtmQGSx8SYakkNawsfP5a5WnKna2L7rM8g
bhA3QC2Eu6cI5BPe90u0IFmoh0QglIBImC79d/UBBCRo/UMu9nzkICn+1KzWci0z5vZQN7czHGSh
I8gjRvLuwBMopz705REN4yW4wPT52kM6Y+wIFooCU/gaPHWRaGkaJc6mLvQz01FvakRSu0FuAjQr
UWYNhiLKZJUwJHaB/Yn7TJOkNfXHFXah5KCILIQsI0AtcMbBG7a994jDhX3gTOCO6Bf78tMx3pk7
Vddo3ZOT98jCThG10ojK6FPMjDLnpoyYEHe3gXDPAmZO1ifV+4NCfMPbcuFW7HDqeL5K/xzBCndw
WjGAhI8Ez/BmbXxrU3drc2nF3wjVGA28foXg36NNEE6fpvNqAJQa7DNhOiLhMth4Y+tF2RmUBcDQ
EUgnRakSCIWQzHCd2mQY3OWIR7WZFUaILbvg/Ew1le2aQvRhOXMqD//j0C6i+bKGBTXjwdldyL1s
v2uB9+eWWuT1xPA6AhKhNbd4zgf+SjR5uJaqXnE38PD1bAqRNqI0JjKkbNC20R9mDuNAFQmEstJL
4EoQ1SKO5sytrwlDbkGebpGU1kZeJM90P1qrjns38oxUWLaeOiJLpYzZE9nqG3bopoFiILEmStPG
QWJXU5asFvhLRiFX2gPOuAg1lyg+u/gzs3KNIdwpoQDaEzO9yF5IU1pcQCyXXsWbUcpq4vlsrTAJ
fQ9VnZ2p//0pLwsceBNVY2SE0j8J24BhzqeIyHHfy+4Msy8PNp/DIFF7eCYpSCZMvQkB4uQUugX/
FR6HeYSCmAjlpnerC84vjKN3Ml+8NUVO4+X66kDFPdBK3Jcf2kCu5YkLXVF+WFiJMpbTOMNxWJjk
GutfAa5Zj3RNslLvQM2NcPCPovpIulHUBjsH8N1TQF1AS3RRsyewx2MExqiN+vkB7Mi05AgUp9iv
TNz8tTVEynBiNUm0SsBLo1CgD2qSDNu3iSHcjJ6HKdorV6joxaEVqhXUbCGS2yaszuQ5sWEQMwWr
N3C6TeaOimMdqGgQWlu0uzIId2pf4PC17eoJujqZkfvEQSb5OfjzbtQW9g+6Ql2TrWxTbShXmMQR
cjwrfQNzEPJoo1uRnggJm72n+tU3qI5/aaIcHUdd7t4WIpW0IkUFMnZeocTwtb8lghfrVPrePDy6
HDHzwjA17MBm6tAc0umQIFk3lxVcEDuVih9B6X4OlR12R7/plEDr0DuZ7xTiOOHZmo2twpsRIG+3
pHGyxk8+qNhBpiWn3dQBcZuAwp9Up5E9lQbaTpJmpgFVj3Op253hOVYs8H0pUgQgZMrToY70paBQ
ixdQRXUvzkqORlFWk5kYfygVvb22k9703Z5vRWXTOdJzm0j+x3LvxCE+JvP/C04UGHYFW2Lmtzq3
ULxMSxDNUSXxd38R3S9QczDrjbniLpmEPyqOAQw6LU703fTBmvHK8OvUmErinhRn9/OLKAL+fa50
6bRidvPCFh2jMT4w1aiAXtc/jm/3fDwHrg8aXLyAGaH60cXKGbScDwuUCbnuHbJCynykPhI6mlSo
Rwo6elhHQbNsT2q6EO23YtI+zvuVudunV/xZhNMfj0XN11xuUZgN5Nv8MRNYkGfYanRhNRHpHIIN
Db675L2zt5cbuG6w3VNz/94y8VmLPDd/LbUNfbbuvpt6SiXJWJSuJj7+a9WsjWnsvN1SnIjJraTA
8J/VTWTg4yqV1NKP7QtYbrGefIK3U/2mamCcgMwbA05Qnyjs32Resm8njP/TKp+aEcO5ahQypfIj
LYd4Q8GLx9NM4emUFi7Jj0kXiBiyIXe9BGfFU60xtXR03Ce2ni/OAXTJG9cBftRD8c1Eg3foscAQ
xP0era544aa6pEqXT4gyR1D52i4TMSPe9b/lEQtOo2sntmCTbDdN7h2dTtrSpc3o5eXqEke1KChi
hnxvfaC394mofSHV3pXn6AaUDCRbloIRH7JIL3XvQ3bRDIflK/Pl4pqK//QFaAPOy/Q0P6ZweUrx
/6J+wwnL2Rn6KUGBVnLNELAiP6HipBFdG1nvAS/WqzrwqBWM/WxDMv57tD9LGkqpXurjewSfCnFp
/pPG8X0da25FIezxPRb3sLELSir+mmzrG/n33CENJxz58D4L6OPkuwi5e21sgkSNJXT4SppKQb09
4YO/6c5rzSvPlLw0KOA64Dom55gxCBvTwVFq7uAzXwu8ZVHtuqrYxncPqeN5aYZUCVGnnXS4+pr9
dhhv47eaZHdo06fhPDPzhJlyydTSG1CO0XSgKPmvA2uubWnHlxFtPK7ftKeKZNZRNOc4j3ehJJ4P
SUPfJG5ngcpXodP1OQPfNjhXmZGDZ/GgMZq25KSG/dGekUNOgCug0Rzqw/1MjxwcBl3M6yArgYzS
WUHamkxSDBHD/cNHCszoEYzczxTTCggCiT8o0HQGpPSr0QmlLnd4dDFFqEYSLAFdk4SPHQ2neOcu
/2bN5Klx08ySvZDcMG/MBRgTVvkg8Txu5QZy02qYkzDaSE5dxU0UVKJBgVkVIOtItgMfxQiuHvS3
DPQNyMsM/z9o3j4Dxu1uH9A5+BsmKBzz70aORgy17WAVxZ3Ze+bT8PJLNjn3sKdlTxTjiamxpNK5
giUPbic0CUpDvVmYJy+i8BshTBZ1VoYxIiMLqlH8iVDpO9ldgJmRYvxYy3r5BRzrhX3prvsZZDx0
gChYRVTWj/jBtOh3jcMXuUm8EYws+XlDYkRZKqTC+SvndBdJTBjFZXn0WatoLsQAV7OkOv/IGowz
/lh/0lmOfgREOS1LmJItt3roY89mBv1wVBBv2aZBPNp9QvPQfJMwrUKKots4KXs9Yr0RlonthhXA
GR6w0iilkinkp7O2PF76RsqA/EWDf54lSm/RMCSztDBmfBNWWwqyUsOG1tEHg6BtmDN+C26epPuC
2hXxoPcWd3C8L+B5MZ+6iFtneo8GyY5Txozf2c0KdeXaucOXXFZXL5gBkGQjqw4rkcb7RT9zZ5ek
w2gNCyjnX3pMzVatdJsCID9JmusTjfb32VV/4gtlfzdUtuhg26HSjVSb9Vb4gr4DdrHScOI68Bc9
Dlq/hx6XUqCoW6Ido6AyMN+0mGM3XG0M8EPDEvr8guvVsYp3wqDWYcvj9sd5C9EgIVZn82HOTzlm
MLCfvauUK8CWiVudRJHzAQFnKrRpLdbcX7EGyIme7pxnZsQe7GtyOHdyht6tyrwZ2NsHVZwJIFpc
ky9t5Z5hKzZId4fJQID4rizQZSuJzRjZ+Ch8rwtRyunNRflpw4T8rv6NrAgmVlc3iFQGG/3lAty5
d8qI8NHgwjvQvqJSJamnveai8UEyZD4Ml9s6lowIyuDm7CQ11HprgwoiNwTSC4aU4cMd8EMyMZIW
fxbTZJLPmwdrdmVJX4zzp7ahVii9XXk0CzjLyiAFVa2a7UwHQtnfk6QskpOYiTPI0lP4Im1FqBqd
rIV+gqRiH1p6xamCMecyxPoruBovaQ6t+WwVVR/lUevVBzG3gAq97fRY8Dr++ueUe4qRabNt9lcK
Q/GGeXDnPmZ+K8OmkaV6IVxOqk3iTz5Av16M0SIgOGglb0FZNsyr0/zOeQT1iuHZwUJ9OL4HZs6B
kMrDb7gm+6BEl5LIFOawNAm/bNULciKSsF8+dA98XvMptyzeJEQ/Abt5QmsY+RDa+sORjI1VSz7M
t0zNc6gWkqKfEAUwDvujHAT8k6BN5E61zDG3UfQiAd0mb9Vg9h9k92SegQ7/jODgy73ekN2SIdXl
/JH4S10xXe4GMp1lHu9rDbd/b+2tDL03oGlqNvHz70nyzqiBr37T5IZ2qYbx4n+rz1SzKGEuw6jz
NS1ade35u3mMJPjE92EANZBE3hBQJTKs56Mn6hPW4X/f+d1TV8Y3uIYybXe7XUWqS2JpzSTrKB3u
j/IpmV5kUIJsgD1foLu0mXqXlTJQ2V70RH8kssFLkzwrVykIvpliZsXW+RQ9YRGVDoVD+TKqn2BY
umewk6v+d6CDq68Lx6MV3G4mAJYfjQR95q9Pvd4HN6cv/XCHNelp87eHWoyKUC3LBRUwMVIQEJaS
1vprWv2dJtoPIkk7cJWCVh21ytqMDguZZqOMqzj2M/rM/btV7bNHRnN2+4lt/w26Er/3sOUeVKJJ
5lg/ZUvxLfjEt7PS4d5GnjKm5i5TbHTvdXxfcWYgr/hWPsfcuDo8mHcRlMqw7WSuVzCIpXApiy3S
GYulkj3G/gHxnvdGp9ACZp0L9vyomPxa7ZFs4r3UvytuzqjDI7xl/brOKeyDBNLClsL2VAJuzHKv
C0G+leXNWNYVj12e723zggVVwiYbKO+0zynjpvP0UIAGMnCPEkQsBcEqxdq9iO4fcuBo+WddUC8/
+Xi1rg3gz14spabw/o4ZrGhmq8FzKvJxQrM1yrxJfH8bR1QbV6itUEYe29eqyHcUsY3zXEvkOD0v
oeGVWWJCQ60YpkYtklNcZQIGVUvqNcimM8A0d0SfeQziNxdDqd0Xan2Sv97oea+GQTZ1piiQiU+P
s35moTguHL1WNgfCSlNqQIBHzyXqAFRcQSDdaB1HqKFCotspN3m7cQDLz9V8phhri0OVTmkEMnwb
EreRQcDDmX0YdWxz+0fJNkd7ghN9hV4vHgq5TJIzzSfVER8zUYU0LONcO/4WpPMBF21kMS12+Lap
QN7AhiN/HhrHgG7ZWbnVcBlOUco5EsR8q5gn/bkzzqg0PL74iNimpcHnbsneBsO02R5P1HIMl5lW
QkV6pwdkIGUFcJU5Kd515H4j7KIUe5IAjJdOfq1vpiKSzi36EsQroJvNPyLgNKyxtxW4WArDjBHV
fCvaWnI1BCu4fHkdubQNqmSjgGZZxzuXd2dr0JS8qUf5ucjnfUNb7FabEu0KBusega21YbGhH1Ts
ndWcq5UVr04mVL7L2cjv6xDVi/QfcXtE7uf8R//3gxSCFpbGK7GQkOYXA8hh97Q9WYt6Ez6gOJZx
3M9y2PDapzymF2TrHVYKQ6nZHDq9D1Qa0kgZEcu4cE2HGfwJ9V/e2uTSXPJ62RVdc51SoADssM43
2dRPKiM91fA2T9foWE8NBFFWTHDz+euig+MxuxhcppEYU8rLvhKIvnjA3XcYi/Exkq0NYGdUpf+q
BMDhSnwAtu7noKGiSxP0kJisWPugXKu1X/tiIMK8i6O+7wDnMc9Cm1TbFAI5YzXWw0NvApc3aXR1
R59F/Z0Irsreyx5HFiVOLS4BfZeOTuCubr9ocIN1XhqttnDZnAEGgiJQEm5oio10QRJRccf67Zq6
Y+Byk7ADCBc57XB6717ycD14xMx4no8i9TNAonesXFK9it+k8L/G4dC2mjMPvehzWXVVzze2TKC0
GGkk4+m1VYcFn4Hv82mGQHFqtgVvXS+dJWsgW+fdCL57rHHSZyUDq/7XKrrlbpxtDyPsh565Cx2T
JtHbuymDvyYu10EuH7OhED4j4FOyvdukqAy934qiZbjEzqjKYKnMLBIgu//8Sn3ZC8yNsLrJOl5m
VhdjQz7Ln0g8vC43rOnODBqbs8iu7uLoYrb+sBK4g0FzjZge6qK+QKW0EOTI1XjzFmFoD6YKLtOk
+9mpPcIav0huirLa9mj1XCiW+nXulCzOEY9R7CipYFwXcc9utOI8iF7RrGho4u0A/PhPlmxibOd6
00VhcYFYIa6BBjXVkKbewzNPVCKJbgk5pW4dwirLLqekiPXousZbXFIbmyzXYtEhcy23fUTPddzv
QQ9Bg7urSD6EshaB+o6wnWvyiZGfenRzjkf7YRPtk5M3ZyJ4OOfjFYCUFXyt1jhMfGoPNeMWv8Y7
8RV30ZP9fn/5O+1eryvzaT2TdC4gk76ScCltyxHOtCDQXAkwNmtqhrJjB00qAzDGMaedLzn00gji
/ZYE318EmXTObj6atYfBLU/Y53ra5Du0p9MiAg/gyh5AxGASoYJ0GDF+majWFaoPH6dO2VhFFPiN
Ri4NSVm7ZLKxORxnUvTgwD9IbPWFU1GUCD7tEyg4f6g3T6fOFzp+U3BWoXoPVUURzhNU1gPJjIxk
B4+NaywoMeKHlCVIJYKAXRqUJQ4dQCA6VkjH0f5zyadp463KHqqb32J+Qrvzk4jKhyqtp9QCdj/j
jAkXUAD02xQLFwON2z0yrRhoDx92RrymW47GhTBGuRMmtcmaI7R3vHTA79Jxp9Q3oZCshhsGPJ33
UICicmn3GyGgP5GW99Imh34lTBLlEpsCE6Al5WzYxW0Lzo7uAwAJYD6A10dd77Y65kn8qjJeUWbm
tdCKeIhQ8X59U7Dq2h0mBtPxo+E3rttEAJDOm7R2bL9W3GaHLZfq9hLVkfh7QL2eiUWCjBv5nses
xvY/CZdD6Q2RTnbpvukmOTA/aVidFWBUwe+3VGW8tGsAsqwJV4cLh72mPmt4mrJLJZo1KTysAU+/
HLSD5nau4Jz/2/bDJwIzNk2/HCiDhIUmOepgXIg0ItVQ9JgQ3gg2ugY0j8VSwCRWBDo9rtrS5mQf
8HmXWH8jvwlDYh3Y8vYUudXbT8YgcsfKGfNGP3LWuBziMDPRQXCr9igcXolskaE2LHUvuYpz6g6T
3OafvCfSMnn2YGAt11caolwA7TwYo8Y08QCZFDrqii2rsiZw4i3BNx0Hf1BeROqLAIjYp5MxfJxx
/mJm+1UbNFMZWGMfADxNN/3VQ4ctCzzPe8wtkrM8TtZOgZ/GK2UNRBmMlUfFwPAW8BoGqjcvwL7O
m6yZkmLjCuXbmRYkq/9B4khJnVdu+YtU5+IEDcNsISgBQ2PAXyGtK39ducxsRGJKCi+SqXslXL3S
lkqdwUcpyGJl5MqtjE6ETXb7JYArw0AWLIqO6FNjBHZNPMvHDnkyyBtKcIKffgxasZ1GljTu+47X
gX6KnpcrR/zyXk0dWxozUtwoJW8ehNFQyb8URmelqr87BXCDUg7y3w7lXRVpv8UwCx3+16O8u+wR
xRnT5WmWWh8tUW9MaJ5W6flN5JfBdchgTW5vzI/qLWTMa1a9jCea3jpwvM6sM9IUTLP42gbLEciI
tYeNihXmRlnVXir434UHHlvV3OPg0H+9XVmsQlndHsYrthVSLgIz7fJVyLT6Orx06yXbEZGKLXVW
NEQj+KBwJL28SwrEXqhMd9SmhcUcR+zeBN7l87FIJAUSnNC6HTvGT2+Zd9rDD4f9uY57foYX2Y/D
A1SpKponKiO+iYG4pTtsnF9M9cNnQ4motownwO4Fe/3eN8BZLAj4oETdS9qHh81CBU7XNZX0QWP5
0pTROOMiF1vkDJzvyTiPho674iZsdwO2esjcfWBroTXFSpF0NAbvrlCOaikZEf1938tebLjbSbRX
dMUw7xrmnrVyHpzSCFFtQH7jIE23pi2dmOZP+E/V/8SelETv0sNDQnin2l69Bh8ioI0P0LYuyLjw
mtMyYLRSrIs+Uhm9wf/mVfWMOk/jEaMFt9OjvRZL3FPr+2TnCaYvRf9JBEdwtuamQYgC2VonaCWr
sCyof6/TtAzgi0O9rS9Dg/1Idi/BbgYUWgR3S5Fsp/ygt1AInBu9p6JKQYyhwqwvz1Bp1w+bWfvC
RjcjU4glxctkqkBcHVsXldAWRtpRkB7TwIBeFGzDfM/ya1PQgwJQ7+Gdj7JxWCzD3Ye47O3l0D+y
w+aCQ1LJ1eDxUreBijjSKVC9A8jI2GSoQ6hrFfs7LKy1Jf5auCctN51CQs2B0yqc9g9vaGiq0I2R
2OjlXTt9Io4FBtlRG4vF/raIly++Gi1BVFsv9RSS2ZU8KZAB6n8XHm52mbi3cQ9v9Q7/xCI6lnIC
EYysQpQKFZAVfuDYQ6+alb9T87f1oLzXf7nf5Uz2/NzEMvceyN5aE5p1FbY3zmbBWdicwZ+qo35M
ZlqIMY2x7uwo83JkSZdjkVLz0ZCCzFD6deXvdwT51jhGoSbKeO4Ik+yxqgwZqIa+OXAu45a2AP7N
auXV68b0bux/VHtFMndZiWvHBui2sUL6fdCH7vyF/aElfbRAT9+a9KB/iW5z1FVEhw6zDX+By8H3
16eyj17rQBU98rsKDq3BgZJvt8qBTJsKAOjAsiFPcW2Qm14ZMJ02tggUZz+EUqJpIsJ4ikeoPRTm
tSCAExGZoU+EYOUp/R7T0Wsq00Q0oDysjZIIrrLfqV1qSs8FZVpxnfEWVLTH94Iu16UHhBs0N1z3
q95pxuzSFFeLq8h3+f4UNzxdSfXHeJxriwoDnryLbfzwfXyIezjJRJ1wAaNNgK5a+h5W0Vm6slgW
2PklkMIyMydhv4LhUu/91zsmQnLoNVGVkSecNWpWr1ljoaLkQaK/JpEUGvoW/78qQDDXVF9iUwkM
FaDKsuErWNGNVYe6/J7xc7SFtiJTn2xkMCGl/2voolk2tZJp15c5ITMdVrnqdCiHy9GgeCK93rDS
pavy7Y3LNwZYoAANsC/ydD6wnwVqHAzIYjPdwvWd/B35AZm1sYcEUgtVq+ob+Z1aKwze9LAVUDDK
x7/tu/7J/HJaZ5eUQNkq3N3gpOFE+NAvj8FaBG2DEhjFxPqwk3GpDOuv8CgsnujqMv7K46Ee+xRe
VdBnvhcRzsgyc/LiIdy5mcWeED25Gkt/ZSk2lQMPoVX129IKiuJ40L8wDahP6wGctBVPyBu/RdiO
vm33UmoaNq0LPvtfmc/wbW5K9eWpVJkgHLDGpNr2HScxcS9Nz2kurJsDOOFPUEFGLc4ZZg0ecC1+
t0zIsvuywja1Z54UD6EXwbz55g8sH/PYy1pkGIMEZUVKvP9oVPjYE38K9mCtbSYN25FU4rRlZ38k
uKv+DyO9RG2vgxWkmPhIwSh6sYe29maip/Bps5A/CitaPlfeCk+8/bOFXI/RPGUpzCEamf5pFlgl
Yg/+4lmQ0zEy8Eo5vTo4e9nc5N8l5ZOiYX1PfzC54aLMNdxNhkDr+WJK5jraX5esyR1ifrJT0P3D
UHwlyOoEKVyHAoR6FxJZKPNFfmil9H7BwGYTwxaMT3BQuBq/o1BLLWU4Ag+iYxJJhaagIctXARvq
bUtTF6QTbUJMp4Era+nOA3coKe0Wp2O/v9S2iE2fNIQQREw2DmuTu5yFH1ySBR/GYpvL2fXqqVJ7
0YWM866Jdwwk3RdvksJbqyTJebf3V87CKBy8iIeGgWQXIeVtPvvX9mX57V8ZYSP22H4k0KRzInAk
7ESfaG1dln1trnjdz7/TK5N+o/3gFwDA/K9cOTszQfAOArMfqhSiVw3esSgff3WdDUPUMXpmV8GU
dLIgVosTizns9cCotS5d3tLj6OFLdK7HUapBpxIJCHi5m80YEe0Mx7VxRfxV6VY++e5J+jvhPKxx
P5e4Cfhx4fX5uPISruiP/LRsbDsAePwa1rmWF3X9hsuhPOMT9qSVJZvt3gxGBnWcw5nl6po/+479
UD9kVdna+9HDwQePrtziQ+7/fslyDMyZclJBYgJ/MlmoqSOCB//qFKAt91diZsIvxx4WOoxyVmWQ
tWunD3Hrr+9GkaVhAtXzUwB0nDEClbCTBkyCcwSFm+cIyoxLUtHjC8idfZjagc3ebF/NM/LtMPRJ
O/aECBtwUnLaJUSxiWa6oI5qetLbeukL1MeJ/svCaCGXErEUwN240PyCP7YWCBgsQytCLUypRSqu
9quU3L9j4+T6Vze8lFnvuH5Jk7B9XLDVymXqeWsaoMnsXylw61l7TxuR9WB5lG0nNY/W+hN1tStP
TRlgmo0BuMMgYyrXuZwIw3a5HEsN7a8V1+XdS+aer+dIkVzmEXzshsdLolO0qxMf1muoGrZc7IPc
mR46KDTU/gpohTF1sTf59m4GFK6gucPViw4V6raQb+0pPNRc3WNWOpEqsAsD48TEp143sELCXvjo
8gWwvMFY/gflL8owImOF1hRwWYa3Dt8EXqIP/N4VkhXxv663SzWd5goHztOwwF786ZllDwWNVNrQ
Ad3QTctEgyB+0Jsz7wvisacrurn/XeXnI72WP8ikvjooeVc9kqrUYUOXP8BV4vddf+7leXKmbGdO
W6LI4dzwLD5JRd137v44qHjtk1vpDjzFW31b4NRZAClNMFk9kPjgFZ40WNpGQmOHiYRc4A+oHVPo
NlBLKn68lCWCteprIM37+kPOMR5KLQZe5JtzBJlLRKb0vKEO09VQiGVberVwaeuZ2GtNjEh6aY6U
4jtAfHfYfoE8AyWwFNE0DKGaI0El0DfJ8YnLhXKXAWurFj82QND6oXwyiRR6p9yhHQTZUM4oCJnQ
p9fNnSQ0BLqlviUSCOYYpqo5DuN57pYXJPTYpiyqmk0vANLFVG2nfU3Ev/lQm0kkiyHrdIbJKczl
0XNTxgKNC7Bc5I5R1PCTdWurgtfPqeHd2PaBSmQLQwKgAFB28hSshf3tG8iZ0I/KgB0/swcHKGyb
kWB6/xDqG/wGE6VvJjLzk4pmCxmGN4DehmaXs0DEBq61TtixAzrZbOtMZfUAWHqweWBzZE7dn/tn
8QZxDfB8tZi8/EQKQlCVMil8iH8UGsxktMzGKP7+I4cHbv53R42wQ68i9CrZQDMiuuDp4LFx49Z6
m6t1htkTSnB+1Ajt6tOupIfjIaDmswDN4gnF12L7Ws4H5JRGOYdby4bqXSeSgLuRWzQHIHRvm+b/
kR1tB4yd31PPBD0HOldUvtauIVv7H7uESTQ3bdx42ZEi4FdlSEyeL7bJoll4mZioL7QWBC8ijM1n
tzafURK9hVvUFLUh2+tMcqwby6/dYIZYAQ4TGiBSANg9mTeepA2FgCB2ibAjvSYC1OsVxDrKKcVm
q2BzgTfIqudSA5Sl3X4rUnwfDFnhLL3yL1ZlhGRA6mZrtimhZ6OCHmz0AAtEO1/qnxQWEKSNbRZ8
OEjB+v2QWNFeF+gKP2fjeVGUiFMxtYFjGx442avLOqRCmd5zRNBT66Mbd5j0zrDz+ur0TA3QC64x
myIeV01vtLOyAAF/X6Nuce4MtovmVaDima7mYW4TxrqZxYY8WqvcPKlHZpT9K9iR8c+LMO3ExOhs
gSEdVVJ0/y/wQ2dK/JTYmDZSXpHmZfj8aI0zNMaUOZEFFWfHxlgrxiwLUer327I7bnX4DzjbrsGo
1CW7LHXULxKv57EHfY2btN11UFaq649W1Mtm27IxSfTkjByAR6iNHintovNE9AZCLmd1czCnAt3J
FAvLBC+pc+L0dP9BJSOc7/Iy0Swa1ss2q1FzHC5i98BNEmPkapKfD3aj5rHYa/AI9LoZQlB1Wjnn
uWAblVpE/CM3PEsWqj9SVTzeKIAGL3U81hOwI1tgeHpVJ/D6Tm3d7OCgQo/0TwH90HhnteOOM8Ba
XKJG+IRk3z9zTc/d0jWloxvAqORzxjY4+P9l+Cq9a89E8urgRD+BFVIHkanz1bTaFQZd5EXRIJ1R
oGGtCPK7yEiSKaJf6wPe2uhzuHp26XLBbV9x2uhfVrPwzMPmq0sHSgOa2sJQXGLDEWXsNbQySVJX
F1Lzn7yDty2oWT9/8d2nE+f228MtrcsAtj0/uq5sTwdZA+kjvGLVyxW701DYgaBsQBZrSNoc45gz
s5BNpaSojLi3fRbXPBX0O8P/PPLlwznZNfCtthdfmoU37U8TFjMpWilX7XB4weMWKiZQICvNHCID
VrtHqa5mzCVrU/p2zZypQsdrSA6h8tC6eQDSvB00bQK4Kqh8zelsiNtVn4dpNPS4NoA0+PewUM8p
A8VHGfK6d5XkPHtdVpApTX66WrByWKSq6h/TLia4h16c++oNNQXRkqjP6x4EQKYw9A3btk+RAlet
abC5PDwfu2IgKjGQU8zJ+Ww4BcSHMBnUvkOL/3pubEP0mUturDNiX/3x/02/YuHh1SCbjOUTd1zL
bg668y3jVOKjBoEWMeMcLhWvjnQKqmiK8u39Viet3+5TYV+W3Hkiodg/9TfxBCKhbd5bq0aqHFm0
pLZdoeGVVIxZCkKdXSPj+NHNfZZm9kRGYRhOzEMmhbIA2DnC0BrP5MWLjQWGfQo3JQn0bEfYZAtR
H/kBXQBPdDEXpmnmw4pyaUW6w0wOmspO4HGxd7DEJkQvROzYnwR4BPllDXJeHj558KcULQnCQNUQ
XDl5xcu+xG+gRpyDCB5mL7tsE1z2hgF2a21GRUHQ3z8zGMU/KVaxpC0pf2Jy6A8GYugPHP9h47mo
8iKVRHLXpX3fYIN2oDdeh7tI/AoOj9NsWWlaXs/smNsWRJUH7yZ1EXlU69YkM1p3UCEtayA8Bxr+
cb17MAFGvRnlJEhTDxncw3zbb6BFiRmqXZr8V7t+kLX2bQk771UrbaevnE9xxbVjQAlidP3cZNrZ
3A4kc1qc7q3DH1/5NWjfEEm4KFWr/ELSU8ub6fwMw92VwA5vVxJ81CjAXzNYcvWcWgOKMnPhjiDO
mJUvQMbGK5yuLagdyvldXoXRTr8sa31bk8ZlcPBh6Au8u70mduePYSBmQbuPY8b1ZD1n6XCotNP/
cVRbsvfBMq/Cn/MOwj9Obbmgz3Sb3fMWKt9b65mK+qZFlNixfgSQfOAnKXGounu5imLF2ea1p02i
XbK8hJvh1aZY9679QiwHw/xRozqvhhv5NPr1B4w5p7f0xEIafqb3KXQDvW6azzNYYtdWWB1oL9/V
eWuhv0NKk6IaXsYYA1SzYLD3Iruc7n+sbFdNj9k/GgPssF3vd2OhqGmwfpC7exYfexOwFyhp0jlr
ViQmB5tqZL4luQsh33UHotCN21mfXEFdORYcGfjGd2XxV+iTw7kWGTcPf4IhPRv/UkiYa4894XJy
eFg6LTM4VqnXrM7ZtEmHvJ6iBMVzlD51rw7gplLJa4rYwi5EfHuSR2Ir+kZvCQ0INk3HYyoIW8XL
OOiVypqbQCKXNSKRmwZWJEDVMJupflK9DVFTS+o9tMiUfzWJ3C4F1irnBsFUW3MWW7ezwGZ6MqAV
QnN7wTnEeIJx/hR0npUBu85hwLkqjsZhoNhkZ93le4MQkcNIJXjq1Kmv2qBqA0Rq+7lzJT7iP50j
O1ZJQmKtqh2FtWpicmS0x/vLu/CYBWna56SQ2B3xo7fDmjG6BC/iXl+1S0UNMMK/8LYPqc7W7FiX
mXqXG9H/11V98+SCTVRcO4xyXX/2A+rSoTzHd4Rwzgwpx+YXV+EqFiS58Ruyq1079g+1hJ0FxXMN
qVWLAHop+VMLx74k4UH1fq4Uxnv8Q/64ZgnGzeJtg1xMZYtsMXa1t/Ggzy3u0FNvEdbBs3vctNWK
GS5Ais6P0PLLgmHoH8KvS2laSXB/KETS+J5B/nDR0u6lPc1a69QiXNnxOCrkQGzJugSgYFcrhZmU
iRR/8AOrx4G7A+mlNbK43Yt1iSJ3+n7MJ81KbbZL/tMy/OVjXajMpj2nahQ69qyTsptgg7v1YJP5
CsNJrcmun3PM4R69Wa0IwrtV24rq2/tbJ3x0s21mjrsbAokr/U/q6wa0sT9S5c0mH3sTncxvIDoV
Uc3+f8w/IL+rVpCTnRbmscUq4LUsg0/gcavGWKPe5itcBwESd2DfnAL74G3MHn7Lg3Xp4NkhewLe
i0njba/Qq71/Cr1ldJWPiZ8jgQJ6gy+fFev1EtgvX4LQTNQSGjKJTijItNB08OQ5rZqroh6KfzAl
i6MEMwPLm2lGc71RisHXYj8GhPViU2lsZTP1tX9nC2Q/EM1mjgdlQp8lxyobN315Bzf60dMtc4UW
5XdtEslMo05dHGOj5gP4EwLkzwQ1/l/wYVUFuTrWRWYY0Cp5difZLjslIEE0O5Uxu2bB2NocwGkW
VRSncZ6DxT4ZaWPlscJxPPixweSUhyTzLnK+eGPT7TDNxbe231eP9fcinvUVJwYp2hPjWf7eBto8
sen1Vd30OupBZkhR1HS3igOnTEKtS73k/bvTx69iRXu9j7aN0yBHC/qBfHVy0d8f0qjb4DYOzo1p
c9qflZEDBdNvnMb8NfuJJ8Bw8pS1dqeKeQgC8AKw/v26ePGT2TnPv0SODCq4cKNsOhlqpAfIMtb6
yAR9vLoKtXCaxv5ZX76NIn79zkORv3coid7szDc3d1jZqJ3GXciUdMFavbrlS5eUFKMIcEN/tKLL
ES1fs8vcEDWoFhq4g04vCNnsbyv41EP8/VJKR79+OpgfyByuOhyTLNCvvD2ibxOe4rWVO3XXxLNk
iBDeEky+zPymYPaCGlP4ALCTED3VdeD1ZCPvYcdXKLD261M7dq5v+99/oWkKPtYle5khG/S3KShq
NNUblAr/F7VUKrRl6H08LYlkEzkJ0MROCoZ9SkxzCNuMFBJD8MxctG0JhL4g0NIcaOC/NsfThtFF
ykOSF1JJ6sfvSuYeeA9+eVqL5WOAqTisrI3rSZJh7A2bupMGLe2D2eWHuLW/msuj+HTnGRQ6boDx
nhsLq+2hLOYjEoFQnIwzp6lbd8WFZO9op1sdZVaZh9bhUUb0xazcneWP8pf0VM/RrwMUoeAjDpqx
VV8qVqDeYqd19QOel/P4Cr1ClNXGBCxHyz7o8zI2XOkZcQZ2oWuxPuCOEuinN7Fl3wSLAsfysvmh
JoS1A3eSUwp7HuG8A1GW3SHcpYx3R4oYfAgPV274F1XBbSTbyPYej2L6mkpD10iG0ZkL8psudigg
DlUkdoWgyYq6Two/JNQP8w2A/t5DmYmT7sBsPVstVGExhMwFC077n0qujr/9Uz9DP/nKDZjkZs9x
uIHsPJHqtRZ0d+AAF4BSaohIuFVFpOPQapVybt3237ILORGEHvPzhErrPKZaoA8LcPvRr1guYwro
3IvDMxuDiNprJY0GxnjiKYaEVrpHq04FPLdxI+cXBryNxGEDfF1OsSX0FIbgmSyL6Twb45Ek0AtJ
l67eR6Fvq8iiTDky+55qSogQCzrrL32VqVMPZ8fQgPeJQegEEN6NDMcRmVeVLAATNIff26iU9Pcv
F3nvZ7E8Vm/sLVYq0aTiz4QPX2A8aDysnJO/0L2Tdqm4htdviRzdp8+urSObJX5HBvTEpbrBC+8p
Mn2FZxWzjj2QNhK4U7TzFX968lYNklS1AIKpSHMgAkxSi9Le5anbcbek/rwvQsmMKRNRUh9zY+fY
8/xl4QujTcJ5Rcj1y3jfdWdy8Gy9XdA4XmsQu6u2MopKtyziR0vVRucwVAs7+n283Wh3neY2wqHM
J6mQGE/T75/VP5Y3QywD4YrjsYP/ynJcM0ibGbDSjGOzkktjEZ7nWku+bEMa8gdsMEdg9Ql1gMvu
pxkjncYQl2/nnTeUCt+ZONVS4vqgbdPwgy5JxhyMvX2WUYPrl3GpgV9wUhNfAH3K8CaCv88KsYeI
duXEumwmJxPSgOD1vcQ7HvAqI/Le0gacNdUT02yHKwqoQCu97h5bXLs3kx+at6bR6WqVi23FSBtj
vxpXrput2yBVhXN2wi/5B8Igwgm3EGWC4crD9gZ33DN99Upv9ZnrpLoPXssA/bEAx5K2XBI/g3n0
gEvMghngSqIUtz7UD8YgsZ5h+FrmhBVenpRAq+ylZuzA9ACgWrFrSVNN/zV7UNAiNw2UcKaS1aro
BqSA+He4pIjoEfYe6DrWSpOmWMQFNSQDnfPayhGdREovMLR1rE4du8rPWZJIRcrH6QBQzisM+5QR
TZ2YzV1vNv8Pv1RDM4W2oY5fQV4bWJmPQs/qiA19EiMOMbDdCSrgTPR/1S4baUGqUw+vQpyDyTtO
aaaJF1bXS2Dz2d7ZnYjng/K4XH5RY2bY+mM5QrPwqmeK/ydOKpltKTSc6kVeJijJAACm9BXq1/+0
FMA/dYZqSxROopSDT+ecTMah0a/DSX9+hy//JKdNwLQ/SJQL2yTSMLZwNWPdph9CWSE45yWUCoqv
/6xQW7imUP2PMmgw+mugNgjI4UKvQyCpqZO8BQf8JQ4gHC1Q1G+QtHfhNOV7Zc1zOhGFMt+2bYUY
XuH2oU6l5ykQJuaGGJuAWRw0qiXjtHxmjYx7vums1bYEwsSB/pwEkbNSqYjA0mQAyp5OcNyBPHOW
nDmgIapLXypTMwVxdS1RaxeZ9rInMbZx/p9Sx8D2QbcuXRN0X7Hr1efTNcP9BMYEMSp/zrcdtI2O
jUFDfWbVRrhSnE7scTo33FPj1CIR+UTCE4IXkmKHjzFMQ+jH8pryPhkhsc7jD9lfubYVi7VblXgP
x4MpbxoDtx603NSLT+1IU90G3wgcZmDtvtdQR0hy03yTShWjRi5ha6+HP2RJHpByJ1LyZfIWoO79
2UYgiXLEeJpCQPP7moZkckDITKWEf8UNjyi+/pcvxnpIiC6RfIwRTGQV5n6DSdsg+mQ3brwalBNU
EOOeW7tGh159v6V9TJZfXnlia9yVllqivoWdm/d+gmn9t49T88eNW13VOKXlTf0cA637n30b/ZXD
PHfE7fqvj0Bl2rnT3GX1CIxLGT5kZZ0DbWsunOMxVhoV950lV/qOZcgsHuFQ82J5mGnh9hwWE01D
NDH7fUcwehJKvRQeeZg1fVUtzGIEYz4fwETzbIh+Sg8FbNcjxclS706NcYCxm9SQpMW5fxNqaSkg
f9ssdq/mLOaokmf2Qbchcp6cF0bcV21rOSbACYWbAK6ZMi/uIPJmcKkkTflXBYJrs0xvKSO8ARl/
/7qmTjJkWbmSZhTZ9BBHTjdhFui0o7GHVeXn/VArwE7aKeWVUm1SxPiW/Fse5KmyOJIMJphVFwEV
0/4jYeUa/lVfSUqzxlD33lcBbHtymwhocTsNyv6kJg9WhibgxQqjdG90uUSoL5d4OWX1EkenFd6m
b3PW/XzvctKrzrC3e3qFpeqd3rz9V9nI9cYQ3qYDnf5mgFR+K552eZyIilbHKbuJ5x31U5isYVDU
PZgBiSQbXIkfcrYSsBllKPkERGUz1V+e4yi0vnv5SXDuVvM5X2HEnBh5jVxoFn7zd8hEk+2Pcx7B
7h1rm7aa7QzJI07p371b5BsefCuYUyzhHrZ3ct/TswyEMg7iShBVfhHM0jv5yeDasHDGi98bnxoc
ebJ6h5zq8pTOVuErTaoGokaKh1APsYAc0LWNTMhVSZdwGd89YUu8YQUF4rjWwmbj8+5ETq1Ak6t1
vJfXE+kJLO2vqtWQunADXuONUWXBhfsJ09DAaqsKxrXkz8Wa+qbcq6hI7FPKMB5fhcGLZLcwNU3n
9HeGKtVBMaDxMYDhqcFNUVy3cEPEN55Pn/cTmPA0c6qs5bMAqL2E03NIoE0zQsYxt7Z6zDdnltDU
RJAweHI0fNZQgv8ar9F2hcVy8p1O6pmxhisW6IdJMQcP45Fufp6KuK3M75pzK/TkIKjtIjI6ogCO
rvq/JfonJCSqPofuED2wDd5W/L3UV+OkxDuVqq7I58qJ2P2WvVLd1xCdc/pZdvZasxUL/b5I5L0Q
XKrqvmZRv4np1Kn8ESaCzz+FbYOedzEM7S+JRJMCTMI80LZM1y4Xb2SLO0WsXuvIRf8j4q3nzr46
AjDmkSWNkM0tuH8/ddnjw9XUcbzyTxh2Q1ihY9R4S8l2l3eZxIET+B5Qx4kdv2slX0Ec5n1DFeKf
QXapbNclSqU5RPZ/sJtZ5tpTKxgwvHzsomlsiTYUNYngWUYG9z+FUxsFbnQXOaWObvOQV2Eu/3N0
sZiuifHRWQyMCzqIG+Nk3zxbkOMPA1z40l1jeNSAKllP/oquq+ngQNqsypnpQPOBSO75Q5RC5h+u
JfOLwmJWRXl/JC2zIylIFX3ruA07DWNHNvAoBle6i3B8VW7iHuVogvPH0iQ+9WZLzB0EWfxUwhJ6
qdeHXeBwp/6CRXBadafALKo4NDE4rfDedxsUtN8IBGy0WpIzfYrLoU/1ewFY+vIX+KuTrspjkykC
xyOlG6yRco/fDTVf9wI/howlwftghrazx1Zwf/JJuCgowJm4J+s64nbCRT5E8voATI2fVKpQG6L8
kVG+xCSaAhfswySwsg7rYC1JXhEg8suIBXTf87ZIPDSIs7yVrzR+a+mxMcwH/5Bt3F565cU0/x87
Z6rsl4g5in++70bMESYxqTGBfZqY1Bw9Qo7oNJZUyiB4qNOmlM9syypr/cWRrRqv2NGP1qt76KB8
iikVtP/8LyyXQjke1HrmDi6ycIbCH3I6KfPlYD6Gy06g+rNFQXm+E2CnlmHex+m/wBXxpt52CaL6
m1T5NDa5DvauyhPdc4u05HVv2v30pmjLCdFNnbxvfj/NWnDQbssnJJ5vOf/b3/1PYnEYNJaGAi0J
E8xeDsgxdFLvhnbFm1iUeVw9JbMkBwKSwkjOkvbRDXOFaWMl/lXm6/Xd/LrtsBCiVfv2bODwJ5nx
zfdrVm09kgmS1yIHhcoB+amW5+ItbtvGVYR6CquxWPKOLD/Yzhhv5w0sHwDz4z+t9DsCR54Tkviy
svB0x3pG/aKroWqMEbQV1nckuP5p9xaTgl9HV6UseBmCPAobemMM9nwctzgsttEAkXmo4OBme0nL
h0u7F2n5rgIEYa4f8fkqIKcWkV2inUx+ptF0FTY97e+6lRHdK5uPFfvTOez+SXA7MptjJzQKmiTQ
XDZsJqenM4URWgqVFS3fLNfsXsM8/SQur84emR9/X0l6v6myWhyzJBQpFR5bDbBaBY3e/DSNEtko
dBJ2dbIs1RP78XBd4NmHCVajQZI9t9wDbzoMVmSWvLN1ep66IIn88GFmils5oIPWMwtVFpgZVJ+R
tnVd5XQ4ruBBlHm0bQYp5M4h51bwtkn3SNl0nEVXDeuzspp9IjBenKlGkszfL0KVSR0+hXzIUaC5
Xw2dKdDn7vCqmqKyUlxcCUOLgUndam2uNtwp1AWK+no81SN4OyDTSQlLI7bt0KW3a7K++egyK9GK
XXILlysaahv01O1GiwcpRn5X39xzgWKPfvbqRWm7NJUSFaeqMpDmjmLtgHfiUI+MX0tVEPMLVmdO
UfxVwZ8HdGMVih38qUQl/+/NJX6Oe8U8i3xsNeWi7FhKJ2vFwLUcJqxf/DfBF8B7bsdSWfZurVTM
dsXVvoQGz8WyszJU1W0eabdunilAXdcJ/e3Oj06a5iQIeAhyCoppJpIE0p3QIl+E6YyY8nX+GoV7
bKVcjfMjRfx4EkNdZ+V3vDah8lWMnmdhtS1scDfZnJ+WG5NHO9gxYo+LHn90TzdaxFF20H3Fn2+x
fYBpbnYuJA8snCqoIClddPHntVKaZZaEG6rqnrmuXSAgocSGQc1UesXGgit0nQBR0MVPy9HOsYlz
WO1cgbiMenUMdqLfQNLrkXYSjT5r2f1a3uqmfKjajRXxUW9mH1LS8o60xw/B36u/nwIbL9STrGpu
RJdEnFLuFAvmAdxN3DC6UM5TibWVZviRN1q3FZ8NDRkOwz/8byeSSQoTyG2WeVL7jmZP8QYhDnJD
y5LbodlS3zd+n+5SXEfodOmeS7JifSwjLRW/mBUysy1PSCuKUDtgddD9z0uBQ3V22Xp3e3T+yVBe
xssQ0xgJh0lMMOqYQjAlkydaV8DKKbh83Zxsxm/dUNeDosQzFtV6AKwK1GMnR6mXgcVX76Lu0FPX
wzASrzfNlyQHeRqs49P42rG9vSAGyUf3zQiRE3vQhujbwg6b5CYsljeJe25Oc/HjSgONwLnYOHHE
jgs8xq0eIgmbIF5yXjRox1ULb4tcKQLnnhL3xUXw7iWV/5dr2mjaXfXv7YOmOHjdeicz487ZqKFz
jDopv6ytT+YqPJ1ZiV74/Z6kaGsIrHjfYGy7yIObA8wD8F3abKKPotgtyiDD8btTMgs7PvykRp1N
+2fe+VuzWOdGCDZkGuk0WY8ErvWl04bsSaNTWIA30x896Ju0MFUSUujbNOBzCvduYmQhBs9lk6C+
ZTVot5Qozb6Q+omTOi/+FGPwLLyWTNvpeau7WFxRNVmmQAGBaYIYhtCqXWmSxGyeLN7WQXthZKym
db2TKgIjlmsoNWqLTrO/7wq4CMzXq8ThDXxa9Jdr0eSMZLz+zGoUZSJso2iffiex4y6KdOIfqrgE
hJTgqWBKKQRNi/2d+QGflxMgwfv3sdtnIkc8bXw9CyLFLXp7tqjeGG+Jq5DbDeT7PhrZxuN5y91Q
2T9Y7HTubWYouKBEVZs0j1eLeDhFTBhCwFEkVLPVvuXSDq+HRXWg4uFWjbM+0n3u4C7/sGOdx0vx
5/jCFhT4hYmpsX9vBZMcqepf/8ND8w+uGLXs1TXqLL++H4GOhW5f9a/PLetjztuSlW54zoUVS1EB
VgtD/p6kMaE0gqrV+ggRN+r0GqZZf1c7ePCm+EMMZshIm1BSYY6ICKXUSek+bqopf4tgw3j1OFkh
kn3QXViXd0mMoVAZD1lFRXr7O+fAAXYFYG30u2nWH2VNCvzsDIyhfWi1OqAkFLU/YehGmB3pb0/U
ZiRJ+6l4BLoIqOtAbdpDJod3co1UsUACWnWkloKGTXCDiGu2XrPRhZayr3yk3W4MfzaOx4QT1NVF
AkiSzgnvIv7DrlTdmG1+8KEGA6H2iqzs3BAvDA7s6RoNjXIxSWID7+W7zx2I28hYUCtYsDQIrH11
ckDzERngsr6shOg9dr1kG0Zarqj/3zQMuiHLMaaoHmPiqt4zIAPo00aR0OqK8Eg4PR/8jpbY9jxz
d4+ZvELjewu7zZMX7dpqVBQgYwBNLhUf2qr7WpPUH6L4qzc1lTAGjfpc6BmziVoVVeXN8wzwIn/P
bI3Hp8581pgNUBBLhDgKy5PbJOjRlJpn+K/fUHz+DLCZZEzcanasU7Mhqr86voG5JbHWD07963Ip
nSJolfX5JdkZET7Z+Kk2PwyRyQ/FtwPLQD0wLXhEs+/3qOFmrP8vrNdY3tlAj7FwKPoFd/b9AfQ+
zHwjyliNHSPs7MceV42XkdN1MoCQCtnek3QKgsy3OG0sYXHQYyVkLv+oGuSDSSLg/jtoSDCfT4k/
3GHW+woQdXyFY22MUkR5qpHyae3py1Xyfpp2s5+kyLyBNsb+0KCQKJRD1Kisio3uuWXIfGapjY+w
+eeKljrBd+ljb0BXLPXowEwOWyQRlHcXfKFFP0l6idUD1NJuZ+fS7md+S1ij3ASjoBC0MFA5d98d
qxWXKwfJMr9jTzu7jcaECDYnFyMEJNYdWd+QxAUFlZfGNM46cRir+qcy8zEwOz56G3jHYfCQey1I
Yknfz0Nuu5l3KnbDUAzqwhbYcjn22g6TXrP9bOJ+MMHm637HcDSxt5+VM2gypiyd4rXKyCptzO+/
0MfKWV6wthmYn2an0kQZNq+iTFBNnmBezofm6Z0wn0F5qL3pafyplrYArvyi0QegtG6GRJb+kmD1
COcvPt927gQiqaqRe6QCtaVBcbZBDIwvww8nUh4ETMXIl/jaYCX+YfnTUy04/nEeDXWiTOyQp+A4
AGDLcE0YdgNTflvVK+L8fVR6SHPAwk5qvaFbs0a0qRHVGtq0NCfg81J80xKMo1LBXkgf5/4tYKJx
ivNjol1iIfaIDiZhgJLzZPafqUg1IPhJM1Y0SQGIZaLSdCQAwzOJApQPYEWTh2d7jk+VqbNRaZP6
yMLk+sKc6SGJgyPYO7ZQYbjEmaGDKCIfqrlpk7a+1JulnOcRPZh13aF1i/EZFqqlzOTlBMKziImt
HfnYHiRdRqWjGcbCxTKaQU3v48xJYc98y/ap5Tk+m/pySs1m7kJ1gr2PBmHEnqu+D5fphXxnzUa7
cpIw2UpVtXrqH1lfLpXxcZ/5MjkiEj6/OJrNoSxx8tZxN/2eSd4uFJr7+eFnh/zbQi/9Nrk+R4/4
cxgnHeb8wfE8RqMtdff+G5v7k0SVdyBY1WCHwSooOEJ5nQMnRYqjXeYy2lsR7CqRihsUuUnPT8e/
7Qyrl5g51moZow4AW6RDMRGAxTp08r9YmxWjAi15wmTFN6PMqbobQtCdpYXD3y0A5C2hRKxWWi+g
U1Eq0F+VDyEdXofqFqnSq0fylve2+zgoiuRO+7Ji27KQ6J2xwHNUOzHcZwStDLrpleWIhnaCZX+z
bThKjq1lWXX5B4jSXGQ2xSKF0Ln7v9cp4TdC+cPEnXEVXNVADNmqS9FbkFCk2ONPKpdbQW3M94d7
HsqZF9dbhved5PnV+mZwyiw4VMLCTqzoSpbf6bnMxk1IRmkFCWfpGFbJVulkfv8orhJoOji09Bd1
HPC2Jj9VSPvaF+737FlaPGeln6qHZj7EIli2tfrggYd9ialhSS360V/TXu5yCVov3cMFGwFd0xod
xQE+7m3lNFgvFtX1ngMvGl+q4ID+Twqy69RrlQsx0MnlnD0MzJ8lTwlw5xQb9Sdf5JU0ktJr0biL
O6uzlXf3k9+St175ny3eLaw9mbLxKYl/25zNsFJrmQn4jG1DoRfEsdTM+xI3EG4SPOMKnHhq/0Ec
liwAnT4gj9bfrjrZ2aA1Y3+5EGy6L+5o15bbOEZhR7bJr3LD5L7OJU2a89rEvqnzyjZpf5wqnlWH
hA6Ez3bIyH6I6lQXef8z0FoOVWdzCTrIfGTh/EWn/p0SgcGcvJKqsGqYUwsSbzEgt0M0JiFWf4aO
xySIkEnBupLRLHAD8b1A7hn0+4dc8sSvg4NTL/I8/4C14B2XJTxWS3PO8rr5OZcQDkF6CscfNOkx
O7ipIEAVaIuyJE1KIG+dkk4AcWjn64fzUZym6+BZF26glpzUCNL0irj8vPgiNlR6vfuvaGYWRKT8
PcGww5dcZVhfCZd5rupeZCZdv6JuFLQcghyhcwooRHWhrT9H6s1GB1sqpWHvHk/oSHOBb5ZKPjTM
f5o54zAfOR2V9GueFTfqQeEksTKMSzy7CV08dEWWLv3MC+BYgUWYqYG5DmBy3yXDDi42rRpH46FB
YbYS7nrGo1f5jAedcJix2qpdTMK7PRMZvk+8Zf7cyTYbaENSyhUwU1gbOnQTx7Ahkt+hAPy5vEGS
BX7ABVL/giZ57aiKqyH+EpH2UxCFtR1pQnMzQe3wP+Iaq6LQc9ihlxP66o37kLbE9vT8FlFPDxJO
B/3KKdlIT1gkYKNgl7bCif7x7blHKLG8TvueHd/qwSnAOeBiBSam+u3OHG+zxAoztZ+vHiyXnJPf
NQMBz0N0TcOkr3sIZWwZGwTuHlL3TPzAi58jz40XBe2FFYwZhzryYomwkV/HOGq/UM7rXA36mfQr
Tv7D7oI0rCRIG678p9teKAIgLs4TQnKmRv/TVSZQucGelh8g0Ye14OfSFbcHIkHn3mg6ULVuqMuf
f2K8REvbZGSyUgSL1yqIixOSiehWEVOj+mNb3klTkKhRUN0QzDOtJr4OqNBzPboKEwxIy0eoGXtz
BUZrAUl9gsGQsN1hYCTCua8K0fMFZW6tGsGqqmFw9vwkSXJOjgNHMSAHbBIjIygtN8dZOHQG4EUF
8b7BMslZkaecpIQsBVqYac4v2spBATm++LopVRpwBViTZ3YbBxaN93DJH3wr4L892PLYw5IC0irU
8zc6L3fVwBUwInAO5+yOHXgrudCtRzpY4qes2fV3PfIqSM/huWqGWOtnHrZI8NGFGOrKIFqrZ8tI
pu+qbAi1hLewHeEWnXG4ArAvcCwlukgWHjy2bbbFIBKfBX+a8c5ruBIsS6Gro4x+00atIAvcCYVJ
r418PKsvt76d7QaTKvy/rW4MN/jNt6FUX5P3pmJtYygOG8y1B6d2F7pLPCpqBPwGX24MvkKiNflT
jg9u5XR4up9I2WkxA6blUTWuBSFddKoV50yDtIdzloFa7DhZBq0TSgc044uyROhWTx6bcRRlxGsN
mM+9+XT11n/qUT8fVEb1hy5Cb6C3Qfdn+nYlsAsu2OcZ92MniFRuD9MEpjYnAVKZv+O/ARpYQrfA
01UyGr1d9jzfSMvtSxXYvvh1UliZyZgHJCV0FOcPpVVui4Cgqs/ma01qkKFSz6UoigV4v92u2eZ1
TV4pTG5WD1vAKSex/1VFWJciKfZafwCX9p2n7PpPVymuZC7IE4np2znKpHx42QpY3lL7UpANYKCI
dw68vM5y72yTkHFm5dT27w9dQJcWk97X5I34vPxAfp1JxONLYyMOn45g6+oZmWESEWcya+JD0I5s
AEm979IywzPqzVbqqb2sIlQK3xhStdu0VFxf2LoTV7797gKX98mxmt8CRidiU2xuHBop4TxNyAt9
RbwbgpXd0u92T0877JGS0VYvY+fl3m/Uzkp5MmBLxfAANngM65lvRPSnM6p1o5pEBLlgpM4a+omL
2Hv9PB4AxuFTlu5U155TuJqhZh5aUKVrTueT8/coEdx8s+/5hB9hg98E4h/ocgmsRBybciYSh+DB
I2qrI/0DigHS4Jt/u+StCRSrJeDR6EeAWjo8wZZA3hpje+/ZygJ3eMAMHs5ilq9UwQykzpZyrm+L
IDUoWcv+nIKbml/gC9lT3AOZocfQYsjXEbg5HH1QcLmat8YgZuhE5nSlwpUkiD09IYIta10jQQJL
NREiGK3myuNGyo756NWh3R9W6IQTJ8VP55ewb48ure7SwWs1D9M07Zt09GktOgKq4EpM9Mv3Y7v2
ebokN986bz5apacwbBv9UZVIKZFHwa47ZIZt1Yj3vWSJMz4xkncR2cc+CcaY84hetdDdJr/u/0zl
OURF71PtYVH7HVbOa1zFxxoLXFq+0+vLB9PdoRtBJARFtIySr89Ka4g3QiqBd2baRps4VREyoYiQ
inhUhLAwfc2t1ZLzsmab3jMtChEn4SV9AY7j+hr14EfQ7Pc/s/o9FQSfbjEFkgYrv9SCakaqfET0
g3xlOicbGTMfPufLf8GPYZ3YJ79BmOCYvtC+JcFbcBj5TPjoHeknsh0jc0nGCHw4k1FbWB+HtRPy
NQzPO5mSnzbWzRH+XsGNDJSB3OYVMXGlgfn1FjZ+A/TvLz2OHuDvEzKPoeBv4RYalSrg8jYmq4M2
UyqA0l1K0LL8OHL4rxoary3PEsJTHI0zm+0WIb7yuVX0mB9D4DM5X7FuQBY0YWk4WoQ4V32HWFYg
3Pdxw51qY40x7AC/0pOx+QD+yRcaDem1MW2rhrXyCCAMko5inhMZueSi6TOxIbCaBcLNj9yCab+c
sL00GnB2Z02873/63VAud+I62HK0AAClKUEnqqW9jXIRr4NunuJfaKz3kWaPmG5R6ketyhZJRJuM
O2z1cQ/Rd5e118Asr6wgjot3gnhI8OGbTIa1fwbTuZ/H/MrLKbXoNG5fD7mJXAG6orO7bJez5zZ3
axYMRWsltC5r/Mw9ERE4NTg5eAMUr9KHUI8RgspA36YxqTJanfVOKZRAnnlMUX6ioAM4CMjxCv2N
SxmTqrBeK7ORDTQTNj7ImP8SJsC8RBrZUoiZkHxInbPLMxomlI0zXTeKseYoi2kxvQdm93UGNNPj
pTeZqUgdJlV38Ip9Y8BCJXqRmtZLMGPSNWJIXAE7SABPdnTwX3XAsZHhvbbyfL0a+s/IWOODnJcp
mWL3JHztvvFp0IaYdgz3bEAy8y5Jv9xWvoMTzF8n1ccmcFL2h9ItCt8to5Ne13gGgGJ0Dd6Go7/3
MyZFin7z2nZzRRJ0zKskICl4ahqKyZXEBascGRWK1J8+Ch4ov6s2Obyfjb7BlTLEO8ZXzgGsjCQ/
hRGCK3XBJnW7nJjkKVV+tJx8FN4giOJ60yAD5WsNuw9TrgN5R8PwxY5x6eWcvFcYJqvK3q2FLFFm
2XQP47oGCw15INpXXbpsmnBzO7C96byyYCx85T2q1iWrf+OvOG8UroY6rDD01TjIsPd2Du9aJg4f
bXoR8WEt9KBhcERgInYbFmD35QpH8+K6nJXeONfxe9sRCgBug+sz1t2iLziLu8w3o9IUVnXLu00O
KVLmCvGNlgo2EVXdU4t40nnTC2hhtsNmCi0BdNNarZR7iGM4+fKlaKtJNui76QwmheXPqkTGyXOz
vzI0jn/qT3qaPAfWQAk+o4WoTeO7Sp9HzZt13mnozv8nVMwp4OO4e8xd1bf6PnjEWKDcJT3Uf6QP
rqMrw4t0IvYNVO3qp/7dHRew6xYV2mx/aLCcJEr6DygFgRPCbx+Oh9kB4ih725YLDqykKI+6VQah
o6L0G3iugy9/4LeLXAGyG13Ah82BTwk/wrv3hfoCkbPp++nMOyRvFZEk4MHXpRSNiC0uxittoVwu
9GiG4rx1Er5HNwPef+xM/sOrPUtaLVm7wlxBtJZt7iyHGA0KcJhdFm00koip/yO9liSTmfv5JVFi
Qb1TZleI9ZhuXCXv4KylM/fZqGxmo+cSIcdSi2cOQPMBLgQdzISeb00cDFo2q6wB3a8otytdrCM6
bIYhdVyMfaonKpRcGdZPC6Mu7Aa2HTOcu8/guc0CQ2KATyLVml0BP+U6/iEAnnGjx7+4rFaPJfhI
QpT6CsfcexhCkL/BEXJioa2qCkfnddTdLeK1EH+2tWfVNPHLflsT1WTR7gcte90dz7Ju9VA/RVcW
YxWsKHQaZ8DBu5cWzgPBlB4dJcYHJsJV0CtEyykwdOf/4mrd4R1yyTNOKgyxWvrfP/vPBuw1bYO/
tVC505oqZQwNkuJUzCNBgb0AJOxxyn64L5a+wBrYjc6icCrpsTmOmx/tZrcT4m4OJSbz1wQaAb0x
PG79zgNmTSrblthX0ihB/dbPsV31J1ePUreP9xTX2J5ZZKXUzxee0LB3acxWUwrSpr9l2XtBE2g4
yqnma3vivKHPz0WvW/0sGpzdwxzGX5D642CVgDPLzBGyOeFUH6Vg52zVhsQPJNGsjc2s9u/ifjGK
panPLkegMV794xWYwrepZHtldvrPPlM7rXT0T2y1C1KMv8htygxqpSBvJQl+89uDbewaQ0mwxoNg
EWlwEUJi4Kch1lgCO7qVL8P5NW2vBdmsrEFF0a+w5Cr85GGpojHk8sbiZvAa6sN1fP/oSl/klyi1
ey84+Kfv9vKFpmWuqUyo9rPLIznYp0Jf16N3U4QhzOsPsJETq/RFDhAzIsIpJifxdfUtPTwiqZML
O0ubKqI080N6VFnZsbjZWgEq7HcSwQSkhoLMRSZ6hHzvn8raF3f5IHEYiqYrJKtfuNqTyZlKmzLu
j413mKYxTu5r/gKWhn8KYIxIMXkUZcZ679MqSHIrt0VQSh0AbGZ/JQdb42rAtNC42M9loo/utczJ
37b/vQ7xbEk7KdcGrmksKRPrhzYsZ4Sn2jCb44J0ciUzEp78Q0bE1O6PEX5s83z6z7QuhgWwroJt
aEf3PtdB2kD1MW+0bXwHQTGfKHGtDxbSwsWCu0ZATxCBydY4v5NR8mYyUbdeU2xLavS21j7J27Mh
gMGjITqNMjxdk/FJhjflI4IR8OIaZbl0uHyZQSGxTdorc6SHrz0Sy5yMCY/Pvaj8lYJZqR6bjMhE
nnrwSLLsZ87/7XH9qZgpQynXvdQ4sz9sHF/OXByXNDItqoCJLn13RPMoKcFUMyKHeE5jB9KRXfL/
Meb3ioLRo+l7AV2zpuoI+0K1z08a3q106JRPPAZKS9y2uU8eYbaABh25NUTPPndnWyP2MGbRBQFp
VLsGibIDvppdTNTC+Dr8WqTrKzvJjAUgbxD03sW/sgLwrDM2uynkzlgdAmVXQhAq7bZafX+KF7p1
c/TxzQx/TsEAR996ODVCDPikSAt40w6ITpa5XySRr+g0oMjm+VrMA1TdjC9eg/yP9u91GPHXAen/
0KkHgsz85xo8/HRApe85DwBx/rcG1K6VZa9MJxuxQG4tkrn5cKiiVxKjX0R3Ln9jJP63YrpB0+4z
zDuUkow2C8Q2B98GC4NN1stxiQOmRBfFQ89C5D34L8hqSsSf5+R2n89ZnqbZ1Y0shag8jAEy8l6N
wRDdVIDerW2AG2Nb481rGFWqLDeaADlXwCU/fXDVbG1qSQcA3daQ7Cvimchxvy1mXJQUvGSjUAGz
nYWHSxxnmVjE82E3QXN07XmODeUTk9i42f2nnxzDjtmN8vc4pRIDO+HF9E636Q9JFFG0N5Hdk2D0
5xV2xBO1BWnFOpL+FdIWA1gJf9DL2ZTfx9A3tegGqrpt50Tct48cpZvnbPftX0rY2aQiYH2Tfei+
pNynW/WfKOuw6o+/nq9p7d2jl1hYSVxxRvA2ERveFxHEF7ReCIxhlLa5IwSYsPHd6y9JkD8No48V
V+ATP4hw3bmkaFyuXZ7Meptit+ZQnsx06jrfgry105Qmgv4/YF2tTGc4Nbfp2BJmLlxQ6hcA9R9e
zoUT7QJGrOsx6dOM04K/CWv0DVQD18ZHIs/3qBXT0aNZGFAXQtXAbuWUsfgvVZYm3Tcd+LMNA5iG
+ItAlD2QUf6gIfjXQuqHOwYzPuBA9VlrWDia1O+40MloGKCLRA3RKtm6g0u86uaRzRANsFAMeKXt
RaZObi+UNh+ljMrMt+sOkMZb3XamE/VP4XxeC0KvP3Mn7Noj5p3BbDeoAhd/w5Z1NSRy0JPOcCtO
cRjyBOcZ9QQDlZEZAvv9vOE7WabJkzvONzpWwbmqW74TfWQC1ruQdi26fzJtKRNi8L/JO3oDoq+B
HnK48xJIzd12GQMzIpUoEXDy31zJHd/fwqRpQXMKlEsEweLiGrsMvqlhZteAbG4ltxNmTyJlhNEN
osTJ589Z4gjIhDZrjj+8Uty3BRxngQskXxKbW8pYex1iBD6VTiZ2vwCEZIg0rL1yks/7UDM/nufc
QxpmE8Y1AYXHbatI42aj+BJqspa4/B6i1+ncJXELeiuotGpZbSS1Pqp7QO6s3OgRGSiNAFAxnwWK
bAhjkC9IuCKNGWMAt6q/RnM+/70X/SQ8SkeH+6WiLh4RI2ne9VKMsXWwnDgIhgGH8gOdK7T5FD4e
CAIO6OV1u2+kOjAj9cb+FfFKT7vDFtUzmQkAhlU16F2pT/hiVSJacdco54ehiu5syb6/JN0SXXiu
Gxcod+a1A2xnULK9C/TrGe0C16DgX22CpajVqc50xv5RdgrtsfNSpTzwomQs2FbQagSEteIe3EZ1
2hvhGd+wWA4COtvYGjT+HyKn36GKKrkIMIYcDXmPPVGhcOXUZ6vPYtBPSgEViFr5+RJvcURBt6dq
hgu6YMrV8CGll985XPfjYZtJM6zezkEYCJddnP0Gpf5PyRLD6uW29k3zX2kWuMRpzQ2zqFW0QEO6
QAUNvjKm3lZ1J1Hf3Kkgw2iUPfw4VqFZWL3azH17/U7t3VMe8pf7zLQCok6ypqq4tUbfa1r9sKE9
vS6dhy5o+rF0faMogB29otd/rVQtjNF5ukZiACntLgnfnL3AbXPJ8ukCZIiqRRr27iVikdGOTuIh
ZJjvviCdd08GEDPxMTQjznBuAp9wiVUHXSli8J+8mdkWum7hqEG3QOVt4GzVlCoxdVTmsy79/NM2
+o0+CPUMqPOiIngPEs4BHJN8i/Tw8jyFfEIKy3dhS/TDO+6oQsV2oYL0HhYgne61bStqBMVs7gRV
0RAfiWgd3BE4M393dnJ48Y12lbXuDITFysyBAJeB2E43PBjix88kN5V8ytxqdl+qyDbeshQDSAoX
YM5le7ddxGqlOIlevGwXqskwkgVAKnCpOuxD6u3+axzqw0W4Li5/cjYt+fr8QCIpjGGPVzAmCUky
0XqxEYScmfeELZSlWONeEQJ2SLLSz14wrJbQP1KSR0pyRKmGlTVh35jvFrhJtf7ja09wx04OhXJ9
/M8HrmgM2HUnJ7iDUSgmeU6t34azw41eiafcozb8dFQuuZ8Kmoe2KVkn5T8myy3Gj5zno8rFzBoJ
R9rbQ+0z3ZwzJdJGjn9SFFjeKffOVWMQ1SyOSb6aDbJAjMdpIF2AeVFbljTdF0oczYXaiBJbI5BW
VsjSYeQceya77GNKYDic5PJc05x5BY8r5U2JmUj9BWVb60PuTUDCMWnkPGY2ceboP+j1J+kD06qy
x6sp/bewluwme+BMyLVirQPkiW5vHmWdLpsPS6igafSSVltDw2p5N2bsICt/XIzHGauUEw/+DIsq
wzM9dP2HzzYedE9M7ZOpNlnB2HySm0pYP7Pp+02Xm1L8yS7bDwsoEbcfruVjIL4e1vLqOhbnNeDn
wzDTeJ2wKc6B0fp6YrPE5QjtvEpjVIeK2Tygyil9oLq1Bmr/IhhJgGk/5iLKMb5HsufolZmd9/0J
OL9QuOCb4SZAlGrCgf9L/YOM6DKtSBS+1805rEjZtpjs3hmc2Tz5BSXPK0rYNDe2xH6TB8qDRnHE
iFmbcqDHv/f1T2xXgdxO5Ok3558Qtl6IPGvVF3tgo2XuXuDz+/j/SUvSXFJk2CC3+oNQNofIhijm
kXszZbMibHSGG4B+SbdlMtIPPj0MqNobTKtL1Y7TwmtBi2CoVcsbUp1o9fTD/OT1Wb2pL1jIIZx1
QI2/2umaH1C+b6zfzrPVZWyH1RoueouoKRDAf3p6s75fFbvr5hO+0H8dqAErhsWDnyvtKy0+zZAd
umn0DtQyRQD2fqljpoth6/Woyxsu48TGbrzShwm1jM1EJNI91k94fkQg2A+flKNe6Q4rV2q22sWN
Tf33vTAHrbwiyNStWV5jjHkKLxBAQbT/nMpeNrxQ9bpFH4mWzu2Co5SThiEsn6PMVosOi9uaQy4d
CCWqbMrdMj7cA35o9+Y0qy9GzLUXFJ6NUVTwvVKixIQa072h7WwTqlaqsY0Se7aIc4aqOGP6ubGT
kYPZdHa3W7WxZ625MdoTjTYskCmDRxyhd6vg6Cdrv823BDD+MwdeuCS4eyG0oAM4/wOwVkt9E1ck
3J8hAg+gLN3KoFbUfUKyIogJ2Ebu7G+eWc4Gt7QLDJpa9lM8JIDu58i0soFRpX0Z8rNA1uL4ZSJd
xrNrlFxQB0K9BS8/BXdq8AaS2QggT8lBXt84VqeWscluWnTAnJUoLYz9QIm/P+EOynpTOMncYp+6
xjGJ10kJ/kNLOjuqCbx9uP/zUbAGWXZoOdMLm7f4eLNdupFaeYRtsziEbw1M6f6qDfRtNKJTKa4s
qTu9RXmQrUH6C7ua5HFeXGYlc7OU+VGKcuJbLEEAlghzZCsRmk740uYOSg12it7YL4AXSB9NqoWs
/FgEHZewBOCFHHonytRTzgNqA8s4bFH57zFW8TZDUuO41d/zqmj/rh7XLxX2P+YEoGlX/CosMBr+
QBQeSQRvTVO3ox/izmkZTnnSTmSy0NznquUCZh4bB+AJSnXFL8+F03ytoBRuS0h0E4d6+I37q5hZ
vEDwRxgrfsV18lkzwhha615eBagV74CMzEUF7ctbdKJbnsl1iMK2x7ale36odqJEHTb7wt6GWLxy
PfsLepBIvjqQwsfQQVtlP5jB8dxF4RxGCnCFGT2OXp/NqQnH0XaeX+odrenTVXKX19xNnDb6uLPR
Xnue9Frgi7pVKmVmO3Xs6/yYQPPcsgNU9JhI+1YpZzVdVjsUvvsy6UPvAz78BZ+dOfTQMmRTa1aj
Tt1BxdEkFtJmIQSRVHa9th5IQ12E4+HGGMpMYvYEjENtgzYSlAtZNhXOTFrlmbn0aKzVpRe9cOGt
l86K4jlVxopeUMu9JRGtwv8rgzXvJ2qeNEZfuV5fQAaXWRc2HJ2v772l6wk447l7Q0Gu1ARIMa1k
7fp/50mQYxow1LCg2bgOap9+YgxBIpyOrq2qVzPkri9HEJdPtejz+ndLQ2aWJ0jt0ROOWsv5C2ip
F3i+RTOdfCZW12JjQNnaI0hJ+asSippAOGIywBWl+P+jN2GlMB19w7sgH1VCoOfeLPO4idZISuvn
DYl+NtiYtl5cWSd+B6dXgIouKotZADX6UU4zvFKB8QLBtFt0RnOPutlIvHzkm7IlYss2WrChFxgF
GECQ/gFzvEdvRAhPHrYEp63pqnasSp7A21e7ioko6Q9Hcsu7G7ZJaBOf82yk+bwzWNRbf5J5CxlC
rbaDMVihfhniLS84qJFFmLWOQbn/Vcntci5fU9mQu19OCdidgkF2Co1cP33c7Aq2zd+hkFMV6T7W
klHmM46v7mb0Aja+AM2krwieB1YyzgabYpqsDCIgEgEopjHqpZJXSZn/Y/JRF9OZ8B0tbY7Mrcqc
gi/9/Js4zSG+t69pwqDM2dPdf4aQCDrryEtTd24yUsnScD0arW7pruGz8+YxVOIkA0strBLIzfxb
2dTs4gY3zt0GX5Xs9P7oho5lm2yD9ULZsJdpBi1hBekdy0i+hOcFIbOBsmVQGk6j7nitk4HAivXC
q/vVurA9i/4F4+mVSyct4Oauq8zvzADMJbdh/iWvkVG1Y69kHQovwmjw7+9Cy4pWGYkZG275sLy1
BSCa68mP36r6kEbQXnISeAkTzdtgXNzsAEc/sdQYr7L/+j78xNLMUU/+31LgJTslCy2nHqZevPBP
mR/dd6bsJ/PkdL5lsdty/cM0JuTL+mEYjO45w6uLhREHB2QewN5SqojfFeTPF8SIFOd5JJRmongx
Bj7AFKnNWnmQIAPtj9XJJwWbcd3WAGB+O7wL71jxF4NNweZi7lgzZ3KWZ3XkGdVAdZ7JjIT+tGS/
MTkTIfWIYIYBDYf+GzJOKhoib9SBFD7bSQAIjIJEanKi+hoQ0JanzVPUEqPYlI2DO4+a+EAdsTAW
bwboSGpN+gp40IuteUOpoj0YhWQBVRvR5DvAYTTvacRqaLYt9cxwXIkxIxqoK08O7mC1vpubTOpk
c/aw75pXw6WeKHJ23KwQ29tA0PmTuTZ73TyitzdyPohG8u3s5ML6WmJtQZMcCDoPSPTJV9LV7TVB
zcjXK8Kri8eWQyd7yL7QGUP8p3zEKHXusHXCEWW7cBfanKVwSltRq/T6sd16HdpYCxqil182bd78
tQOedwmZBEnsmk1D1xi9d+EGHOhWbO1BlsUY2c5i78qR9VfIn+wjZWeudujvDRoeB++nNz06H0vZ
fC6Qxg0Gz9k/7O+1gTGiOxoGwX83tzPD8x0UMsmelwAHGaMEttYU1MSzJeKsCGLoicOeiSiDTVT9
5R+hVA/jqDVzVAyl7L27zesvgPHQcpK9vCH8zW9zhd0gIJCeQ7Kj6Sqpl/6iQdWGAubE/xmOBtr/
YcqHNeMmgxd8FQoFHJ2Z93zrmZ06JovLhe9/SYveZ58tHLXcjehphUfoZi58rR6vxdTaNXQmEaW5
VdDRz7HsPMN6PrmDdzc2qe2MqJEq/uUw1Xi4Y2ifQTnk0CcDY4qNXPQtwc9aHEVNb83SYlgNZoP8
BLOX6pFPaKPKm/oIMmhs03fNWXlvDye0czCEIpKVrGGSLjVwBYxKjq1o17Tlf0kQCmNvdQucDuEF
5qAicTdbVr+aKPrxlrK6kHLMWRWyTidlyAwXMMImjfoh9BGfGxEIqfIvGtiT84QFkQaAzl2++9nS
UWZO1NxpSik/JWzqj9bjB4QUKgRl9wyIe3/KV4MWVmn94VmI/MaR3UiwoFB7pmIgmzZoflRgbjm/
9Q9WBWa15I4ZNezbl8pWuj6d/3RvaC5uBtQB2SQlfmUyVB26ztf5fc1FlU4E15uJLkA/4eDDCs/h
r6qHYptb61GEqzkkferpTE3joyPjWR4Zpy5hx0HGo/Ajuq7uhPW/OM9PG1kGAx4sGCwEH0n/O0LY
hVs0M3QnNN2SXIz7xx9FgqzJBqdePEgNsZlFlSw0n0En2gHyT8BfwtmURoc/7JCvs+74xWI01rIY
Ykr/ollP6VO/hprl0EEgxsgtjOXXjatSfJ9zSlPzYKNyrf6FZm4SvRUW0x9zrHmB2bJDrH1q+np5
VC9Mf59j8tzrp5bpqPLG0n8hnqd4B8712xXxBxlIzIx8t8caALkhq28YJ0/ap4JkhTtllDbqr6Og
tRs7ig4Gy+LzH9GLn/KkUmvHumPQJR5r3Z9Utrk1B7TfmMbqG63HrscHPomldrC4mZtKwt8qSTCC
0T06XQQOeUhWH7ak0zaUl75DsQGJuFYavNE/Zfutuu3l2I0uZ1jZ4SlRgRGyWdPTZombpb0QKY0z
QDylFb4nU1GnK1aMDNerEjWJmTNXkF/Na1Z6FqlvdP4DfTsBNFdSAqwsXn5Bfqo8g0cVAUEDZqlL
bifIRkmUxwDtf8tx7jdcqA468cxpAyk2As9N3/RKv3VeV7h23gNc3Mf8wUIOD8HZgqY0RrdVo7OD
Z883EI928wJT5hhP/Kr1DVZyExNw2gkC5LaPIHumcuxaFOBY/qzg4/emWW7z6SpOJkneWPeNjMz9
76rrVs0VGb9FEdhyzxmUPb+PsYUpG/JMbgNvaoRgqL1Lp/LHohHlNnfIkZcyAgcm9igctlzmFBWJ
tmGlbVFha+nQr0/M8k174v4RjoVsk1XyoSb8SFNwK3sa/+COHJhIMcfUJYJqbAB/JfMWI3cnTzQA
oeRsRTbAzQnDT/Za63FT0UVVuOTROJpwFKrgQOYI+Qr7K77inJoHuPvYmkccRn65e1Q7Xwl7woQJ
odumlPRnERrr6IA51GUTY1Mfcab0UwlXqa4CMbuzgrszgzVLWAkltwRRnh/XQSEZfUJRjyUftDq2
pUyRYaHI6XrhDOOqwfXboX+vgP9viPSbqG+cPMoMiFRznXAVHt1zQgTJslh+ilbNxt12yHbagMns
NecncwuzuAr9ohZKkOzaoDdWP29M2V6bsdInpaV2SRaYxJgtNw9ji52AMYQlcT0W8x8weK6Mw9nM
GCVSUnnL/M1R1vt3uoo4Y3LUw/y1Bwg/tFd8s5XVfQPy6JeoAkMLjoX3oRWgfqwlqpv3dapF31Xd
gnOzvRuahoakPBq6A6BCVA0Fhdj8OWc38s6ieIGx7GPrGKQVi5MZ+WAXrIWMML+2+ECkc7Vx0KtQ
RsGyTl5xCjvA+x4rHrV2dK5WJQoRdi4sfMcHNKPWv9aDi29vyx1A9/nVHey314c8/IVDi11ApHWu
wxdJ87tvLZY4Pe+Vfi66mMGmaMcFv/MgN9rra6Lpyd9aMSrPLiw6uU2BxtBJO2LwgqKnPgh189Jr
Oc7enLXYbWx03gqr7terShYNjSVLhccC3mh+L69XAZvuMb1qX0dfblL76PjBdrvf1QsYxOL4Pn0n
yo3DJv9SXaoeMRVEStoZub9SbKH+A5SudIiSf7TEJPyYxYYvQyVndo3/B+0ZiiB6CrrSLl21RFQy
Sxblop1pc/EvlQPZvM1Ryr2iHBhC8fPeQeBl2WGrbYULRLdMAduNm4lHy55o4b9IyOuO/Ju2//AJ
9YVZU71Pn0uD4ZrYwhlOW2WoeFOXaaBn4x/dHmgdVQKQmfnUXX0ihlCVugbnHN1qjyWdlblSJWuL
ffVyeYzKFRhY0D76znMrESyyHjcCGT53/avjNNuHWoOvCn5S2lHEW3cLw4OFiNV0nkPxdf9+PlAG
uGHP7nJIxwSm8dcFAEK4wVJpTCxspOA43/DkDciQAKPu9Bs6cN9ycjNmidztVu4wZksf5mRIiBSe
C2Dvy3y+ZyesUBqbqcAetJpN1Dp6sdiOyqu3G9UEPtzLE9JQboleTk0YbVeTf0ItFKL2lqU/2Swe
i/WMIgm0K8LeqnNPODuTwMbmXL1IxPB8R7+rx27jNQwusEfRAlv8UXNjel34Zjw80Ybk/p5JlZRF
N9JM8LQy1hAV0Jr4G5vIcwg0S4Q76NE73eQnSXQ1hk9iI9FM2sImNI74pw4umqqf18eNmafq0Cuu
MZdg1rdqlH4PhQFMGcflXmPtvyxOKYwzfGSP8eECYZ8elEAxQsx5fMqo2h5TeUNVm3dSUezkKmCW
90ia3BloAKr6yS8LrOs4acclfUEnRGbk919V0UgBzzafKQZw0CtrcHe+ydlcMTJ/Mufnn09gYIgY
ciTrDhCdg4Iz8a+NXhFH3SXWIiCfIXoXsE/RmXFvT0KzMQxCRGhUgZM7C92VWWHR7lbMI0U7l9u6
NDFi8tOtIThq+Jo/duafJ5iZxp+znI00xcbDk4hP8d7FS3MMTAkHzIa6rW/L+EW2PqdoKATFVJAK
/MxfuJuuELkMCbGbuyaTPJl3GJx6upyPVOVP8RzZO21ubsDvBLNeGtj2DtFhmRi+idouWy/i+zUB
t9zYBXH+fzXm6ejQtLD27q75my7c+GTfL7GGRXYcW0pQUBXRh4n3I0F7sfVOOxov+s6BBBzrnIab
KInJEgVAllTsPPkVo6UMATKmBTxIxCAiv2ZNnTlEQrPdKJsW4ip9vR1RqZLE2gMXpSsGd7uXhHbh
YdLLWnbXgpRErfWUvhTKK9pjSCDu2ZcN7cyolDnhGVDSEDDxEGA4fVPd136g/OEpdM47+l+qM9oE
Ut8yIJH9Os+JUihdFNn/z97f42aFM7wMzULV9qO6PIP2SvfI4j/Dlc4jkhIR44Vp+E3GHlpuYXxm
m2UnKJv8WslWudvDCWpUoYScLXuFFvtZz3WAGUY8+TYnfbiheVxJHn1Yd0Ae363HS73Iwb6BaxY0
ugFJF/tL47/aCMlPFrtGbXO/U2Cm1MnOG6+EkcmDJOoDoW42/SIjLM5Usuo4zDRjZJAR8AKe2Rli
76FvhMJulGNazTn9PCGVrv7S9fZCR7C0buYECcusztowPgLP6Lqch0ZpA/uS4cG1AVL3znwspmWD
y9Oz//ZhPZ8f22+VWaFbwXeDKlHEFaXyYnG0agiRdBnwzhZYMSPRvn6UTkdXIWu1sgKKkwqiI4lD
0iiQcSmefq+GEyJzfDHscsWhtc3QdrsLG9aSwFNsPWcbzrmGsl7aFHWkrnxnIssHQpnQ94AFwgD7
9jx1mcBclNGp+SaCse+2sOw6603lOZLH+QhYL2/NaNQMC8HCaBBJkrXrcm2JFJ26gsI7Bkfy1xeK
iObxIDeGUR/DcHSjJcnfIdKwseSSN33rsmnAwYGaFzToxpoCFcTpTzBpScA+KkZoycYxpojgNoSA
qLERQ4XYwYHNZNAIop1cyKvyA2LV+YcGmhViAscY/gSuqEsAakPEicDVVPSZyyk1A4K4XAfxAsNR
0vFCmq8ZWp/1OJTGrCPNx6+nPINyrXcmtRcfXrNIADOmFMBOqOqetcc68AJzmdvKoHhtWpzZvKqC
zdW5lxmG4+uKbT8uootFfv3HJKsPWdEuPM3KceztpBY7kSfNmbKVGZ0Ai0xUtLJxEIgXVTcuJzqC
A4BXhYAqPsGovx/zl3sPAuhBTz3c7z0+ej32fXQUuxbDKQjq1jMLWEFLbjyVZV4Ieo051CpWIH63
jE1CgWjGWcfF3ZpUnPiZIwPA+rkka8pkgKDCGZg7UHkUdAg0rCN0fuuN1Ld7HJdaxGZQFg5q6ZS/
pKqDjxEKCzhHxn+SViJXmqI3drNRfaI397Jl/KUr0NKB9gAES4Nvb+AUliXq74tl0cCwcZVzgo6l
KBVh+I34MSra81XcJfmNKPt9woyWgvu4Yqwr5HFh94yZCJoXR/FeR94Vod827dr472fpBzp41HdE
JM0o67P6gCBtkOCTmyVjj6NWyQ8f/sz/FaDOTZiYBGurRJxlTlNz+YXlaZ7SR8Lsih33h2AAKeun
hmZ9uA9rc8nmGCQSNMIlI3FMW1Pmj4VOv7OhqI1ExpXzXMdue2lnrEj8coFkBMPnrLMCwPqBP9ae
9GbQ6zVYAeoLb3KccntG644RiLIf7TajcK79C8KUS/HsATeNMuBHqTy/XB5u0QbXLb2uijIzL2Uc
6MuoacI+oZCVF4tMzvU02sr9CHtJB79KUgyc/ly2fgbVcY2j6tfM4EIhJBkg7FedxJeKOneYRhqQ
JgGRw4Pz+uTDw1vMCrxReEGlE8dB2A322tq40KRtz/f+sGmyhw8tFq2NE+knM9vsmIK+toTOjK1E
ugrXhf0+sKJ93qLCHCY9aMDnjkiQ7VaobicUCp7AOCyLVA/MoB2dlQS1WsHrXdka/eT5qRSND6ym
V1iyvu0m54hNhFr6MIEWb+md33RDBfffxI4NlDZ73Q4jnbElpsszNuA0KihHWILbTv1XGqdAZVPD
/gqWd3crpI7Ta6Qdfh8jXlBP0u+KZSBytQu33o8UqbIDVQL54QPNCbA41/eAHe7IvuLMEPNui/aU
IIWUUjbeFpk54WQhjvSHGcHJpNFLmcHh/TTRLyMZuIbot4SlcuQmjSb7ukyBdlTXkdhiwwMhwvPM
gHtCi+0nBQuGsWm0YyJ2KSd/rbJznIbwu+xanfW7TsgywkGNWMqQX/g70JE+viA11IK58F6DmRTU
0KwXio/JeT897ClRZxXMUcdPXO0ABLnKaps0WLYmPN0JvkkwydcyAUts3B9+cNjiNBIb8x0+IZM3
HAkQrxeib5gBIvyUi0MMGefKAvl/zP2jUJW2Gl+ADDmANGij/XkOc9r23M1wM0+l7QMD9H0Vs7F/
B90VzQEu0oF2yX9wPw/xCMX/nCmF1saWQLwCDaxBbNtnA9BBfTcwxNiBA0zgPxTx623lcSLO21eo
i7GHWBrNDirBeZnwHjFu+zfdmVTUEynC3BC19DE2QxlEiX1u9MHlxU9zcCKzbmIT4pFDlRB95thf
d8rNwntR0TUGEXx0HQiX+H6GsggVKheb47djzWGLz1d0pR9wJ8Pq4E7UtYvGclI8wZozGE/hG9h0
lNMuUvqEGdHh/Ald6l52V5uL3aiAR9II9eZKQs3cfv8xpSe+GnU7Y2WBsnoxxrw6Ab/bni4dFNPt
56bgBKrPYlnZynTgjTLtspXaP8Gu/BgA2nNFm+oNbglPky3815L0HQ8r5G4606OwKviHcDrRJQLX
GLg8VCoFGPPUPTsd5IG4XQ/AZhbtbd7bKt/7mHTINLgfO3ZO4rdRLMvGGPCXn9MdmChg5+DFR/pC
Ne8HFO7Z4K69+IezRHXFT/N2dQzLiPN6OPH9yBKbM1+9sOd/8qCGtH757bHzp89MJZTAFRMhaVtH
uH7ZOdDA4ccV21NVNLnYUqfJuxP2e8h5aauBBvzRojEBDiAqLW3QRzXTHMuOgE+/tWmLtWKqGXMn
29U/vxuAvhxlbzQXtPLULGoS9rKutbl84wcpwdHGjBOHRAfJ03HN+YxkrHz9AggRp1VUGeSy3l3h
RaRYFfzUan49fizmJUqLv58bkHkDCQqXIFYJrV6NM0Q/Yjo4GN9KARRDrDB0Be//GmIic7KO60Y2
xmPG7/cFF6NNa89zgzX6YuoGXIOGXPMEUx1nAKB3WWbdfC0U6nc0mJR5ICs5QcNile9dqIEPivcD
r0u1oVZ9eiNvlRiLmRCEXb+zykGDJsKb2ebcUdJPwEz2i4Os3+UHVqqInTKgY13VgGmVOeAHet6N
1BEIcjy6ahLSK8nIoux89+q/K5wXPO+3JVJCAeCPScpN0GCKg0UeRLCV8KC8DJ6Ur7+GF+zJ0FFC
45HhLg67kAdW2U5E/wRXoDdn51SYBw99WhZNqmaZmLd9+/9IOHwoQrpXKOMg9IN3k/lpJLErVx9I
AXAkJqcyxaefxaD8NxPahUHvnsuRWYQGXUbiW93VtlP6UI6VfVWy6hRnK4ICTeziqUTj1IKx6/FU
TYTGz9VpWofiVs51/v1rOdnJR+ofM1Fwnbd9RuM0ssmJLC9ZEnskpl0/ObjAQO7am8IwjJUNujnh
hrjcomNYa8sPSxx39mzRnb+H3YQy/6ra2nvM3WPIzx6GnEbyZAFTO8jNHsra4ggi1PqbfRduQToP
tXAc69b5FTdXgg4G1tO/kwEdG2onKHtBPL/bnwWk9n61mp5VaYOstI50krcJs2MWg5N5CGY4UwAK
grBFL1mwRkzo5tV8eM0jqV7WUWCWKD2AtHNnmse8B34JFZaKPZfIrM49ERpxZzJCj4+sT8yzVKhw
4NYGtHz2O701csuPorxMoYbgXZw99wg6pOJLqQ9H8kooLHtthcB7LZCppqOYfh+YVqZunDlZH3CI
6If6TyXrHC0bQnifpFYAgtz7VuVeoTwxf7GO9H5vP/b4qjRtASa7Jdy38j3llyRuiueg/kzj83CH
tS5CxabBFbpx86t4nRb5p0cQmy1a7klKhSXJl1AgBlyb9QVUUR/c5+ZbHxegZz32+gaJ4FvGsJsv
cSYvVh0rchYBzD6/yW7HAfQxplIplErXfs1azyIGGXrIppAZ46HOSrSVnf4yE0T9Ph10ArXuHEq1
g1Ulyu60x7TyP56U3wDpsEHrg5cCKs1nPohdYDsURwduP/1hoXjpx8pWBOsvI9kfSmAeLsU2uYnM
oxQ+JqbdCpk7Zhk49WIm9wYBSU/Srd5FiRqBRWfeIlVLV8MTIpDPFx8Tq0C7c+E/sT6EhxkfYlks
nWydT+c7JP82H3MgQbbir5uIazFMVdZlqkTwuLwgJk8h4esKfXtEjC33D5rG6ah3gZ3bWrFfFF9I
QYqbhGimVCpIOnEjpiTivzJskGHuYefvzbMUQLF0RlAX2EXRpou+n9RCC/+aFQjk/bKacf6DSd7j
wuFTzVCjMSTTQq66LEob2M93f+kcHF4cu1pQJnQqTN0taotglPmxbJneuMvqY25451IDpEBSyHA6
tP+FeZlsDo9avrdMljUgJk8zBLMfilsAKxWbeCHEicCpcyIOABFFGvZRJwE7LhfNmp1pSGfrh41o
Tnb5oeA+kUtvi9F9fIvm9gaQlySpLDYX99pU/8tyNp9qwOdGYNgtU6HYhazlBz+BuSMOkiOrNso1
5rQQkdJg7sshzJOwp8ta6g1YKEqDqOzTc73OiO3p6FMk1+debUGyLbouQobKOB94Bw6v4dtB+XiB
TGKPG1rxXLR3p8VV95bIJk7LZdrMbsb4ELPOLli9RZx7xmRD8fnBNCeqorpKdaR7BXAQHMi7ffLa
6KtOTvmEyJ47DX6I3+HiRsI2HzvrrRJP19W7jmX1K7uic8WpQtNKNITdRnQ7CapOvkVtT+WXl07R
hjlc5ahBXCbbblBf6p0AJREUSVscTyRXaNKkXD1bbzBqyKSPXRmoFfEF3hEpsN9vw+HhbjyA5M+f
tvnDekg0xD96Dzd0Vf+WJFagnuALuFBu4IIp4WsxaOV+woRxnMwGpnFFumLhUCISFvtrtnt53LQF
Xe1H9en++V4VVXyvteR4HCE1kkQWb/YPytKimM8dET6WpocX5WF17+FG+xaFFQ1QWEIRKfb/Y4oi
msilH5kbv35e5RaIthrEF8VEs8z/SWKoZhEuth6Gb1rMSIZ9rwp51V9BGiEWeTyKVRz8OafjOcly
0LsipLA9W0FLb9BZBS1v8LGs2LoN92yzEV0IHMUWpKCEdnhV+oXflxFyhhMS8hngLGDOlH1+D7u0
b/aym3oj46JUX59UPvYQ4Oq0SIoXhjmmIdSxAfpsvdgDtupBbbzbt0JzrQsgh5SS8XpjRds8mLMv
QldfMcccdo6q5IO1G7mGfVH2U+7EbcV+KOfxtCAfNRLd0k6oy56fG+yFR6Bm2j6brW28p1GDtIDY
J7esXxZr48pn7MDryWUhtaeBba9yT9IQeyWz1cNG2JvgH/rBDG0Cr6Z9156x3twDi7MfUlGZhpew
Dnah8vmQS2GakOiXcFTb0L7ZEyVCmcjXrvgj8BKNHyp5LO9Tm0Toy/PJsZgvogy9Bs25o3SZ/icB
D2pV20b/+3ZFMYpBE2DVPsaUNrahqtyK8vsAcVoCXzP11pcmTvePsi9XWKz0RynFMx4MUxgPTuqs
/CuAB6umHCELLKAHHNssbL4WmmG48M2qjAmjO/uHXSi2zfQszH610hJIkxOIyI6ESwJTet1j6Q0P
CBzN6WOXmOkw681n/X4W5vbROEnRXIJvnuF8BStOZzbzhHtnNOB3AYe8qgwESsPq9JHK8JHr+AXr
cnRTIxpts4z2nNeIQN2/AcJl7mUWpurjgY4ecGa26kscmS92DkJFosGZo9jgWaDfyz+RQsK5q4rn
jM0W1pchoVEeSOXHD4f+Up1jRRvVkbTUrLi6vAf+7W6+ivUoFL4ChxnZ3bRQ+3FyqLZ2+7w5EcWJ
spEzEbYh5X71Yg4O5YNo+smdV2K7+qeGwjranEh1TZOHf/DF0Ay2pSeTvvZ+7wM/gwtDB6PORJif
+0P12MuFh9uAv0M/EgUoLfsO00so/aHqt9gAnfpB+NeHTq6cq10DdBVXb0pm9M0t646SI6wuNg2U
92/bIMNFm2O8bOV/lWO91hZ2m4zO8cff8R8KSlrR/D8fRI7hCzl+klMer9zn68WOty4gaYx393qB
vqcw2SQyYNp5vU/EAlpte6X3wGcPhukOQNlDKL9hnYzK+dG5CmHOphAck3QSMRO8qDV1wE15hAR/
nEvACV1IL1YNFrsqnmUe8b45p9I3A83UGPjSwMz0k73GeKUHwhmJ9+dL+WMasygE+Bcb1Fodwo8Q
Z2Yn5mByCz82yDeSBjJZcsFQD/eLaHYWhg6Cu/lJSGmPyEs8Lz79pV/pxZL0oMlIU2Im9bLunU7M
VXsg55LhpscR+x/qWQtlvoS5UV4PG54IR6CdkomKVRFRP7hloMfJQeiO3yi1lXToWpNKB1YjED6F
5I3mDXFxdW8z041U6xWANItVihC7lRV4M9cVBRjTlGBMUe6ET+nGv0dUp/sAUS380oWfp3WK8f0G
dEFeF8iaTil4MCd1CoTmdQi38IdSbQgDkHfk51XuVuQ4S5IZ10nrrDhaZU80IAL67SlecllgqkXi
3JcaU8u8Zhm+6qL7SgzWVVJNLxIdzxRzf1pBP6JbUQfoiON1AURiihoBdxSbIFvm2awm37bqt+Ck
CRwbhlhzBVR44YNEqOBo0RYVCXKr8vWP8DDSac1a2jOZyQwoVmIuc1SRZH90jh5rlJlcwsl34O0w
G+W5PeHa6ZKkrHwvDcvBupNmXZ6mawA+XT19N+UA2NEPPcxnCkKNFMhPtqGfdCuQ/BMX9smUDLkm
r/OHP/S95mKg7LuJ9jlooQgLY6XlfH/gRA1gJ60x2dnXRP1odqE8eIVHKfqR3bNRl/GBfiGMLHkr
OwAMhJ4uB6ZhE5hkRQkk936IIu6qmdXi9nUYWg/uP1KyfHIzZL/yyS+mxXaa4MpTadXAsCwEYFAP
GCQfXj9BTWoW2cZ3ZGdwY+poSe+d9f8rp9muEI3AORfuQuO2xdhfRhtLy9TmGA/v0k63W2jeWYgd
jXeU7czkiWR+57E+vuR7leRfsoJv29zqIh7iBkoNtamL8i1cN1iLjdQ5OAUPfRV9XTyMSgCZQ/fh
aKSAOORw2bRLUeUnUzqFdwktyQKuawgpoSy5R/+yWdIVl43lVAT1CyRFfpNk7Dkudc+w1NVPJIe/
do4fmy2seAjIcswxDcSDA1N/ugPa3D6Lna8IP66DEXN2J65F9024E1tzI/lJs9ty0qH4wyIDYv49
MnyRmiPuyg9+rOMfA1Xs3agq7bUjgAzEsZrL/rbrKpGzb9FH93zcJj5FTr9ihS2aUVy2uLo82Dyv
J4wml/veA/T/RI0g0NR+sMssf8XLjVoKWG4mOdAzpY+OfWt702in96vov68Y1FHP3VSgpDPQePOM
Vrm132+SvxBI/MiibfXPrXM1Q9ug7rM27z01/Qoo56ARr6pNCJHV43/dXV0lLbqEkONQfVeAOpKI
Aqp5/UJG22oPZht4wUAFsiiuHP3dpIvwHPuMfr+Jos5UMkOV7q10uEoXNdMd5yIFTnMMPCVKaFMa
fLs8SPvgvFxu4GCz87wBPGIirEWbSvg7P4miH6tM894KIvJ20RTGMZC+CyyX47hoSAfBKdZhZlBR
J3Wcc1E00ZOYjQf1VTECoQZ6Lc74A5JLdFItY1lOA9hdwbgwIco6CKCwzGhvxBfCZfRL1kdfQkmM
1ou4IfeJUf9FrmV0uS35gFBJuEcdSun1L39jiN8T5m8eTHnHVGBSiuVtcvGWE84XK2QYqueglV0t
SQWy/SpeDoNJJN072074RpX5CYraEYC7Lyr/PheLXolISK99XDWx8XHIIuxx5wBZkly72WlIgSVA
1cMl8A9GBV3QNUc0NYm5/wZ5WYk5ef5XViuitXSPlt9zA1f2meKF3hkhYa1Rw9WXvuYPihPRKco3
MEQzYi2bR0fPNxJpE/J0rWQ7c2krDEnHJdKcF1nZy56k/J7EfLlm7sG9lNY6zjnTlMpO2xiltAX8
3aFb2rYDDlmTwoDqZCY0hxhWytbt29WL1xcjcp0lUKUnUEz7Vpe0whxsGBqanBlTOX2eB/2u0Mcp
AEcZCnjJ6cMcAT10E1EnbEdYxiUnFpCDNF+RjcsMeL5pI7x2sPoz46AVQKdkuFaH97/lyYdgPWHj
o8sRxRvF7HhHOQX81xv5SAeXTvNQVoNAh1tN+YJ7p/isOYtEtKFh+rRQH/S2Ya5U1lu4vF0vwM9g
9VdWwe/bQO9Z5oB/VzqYPlZl1HgK/iwr2agpQGFir3ylEPxcaYR4ZwvObbihqOlUdHqGS97Fvlsf
va/JHxDjsaCBZrmdEUXPuy3Zxffddf9GnCUdsBnpsLMuhKVvoxYzNKk9sJAUhlImlR6/SWvNP2Dm
nv93JuCKeEcYo9g0Y9tqIfUuFw5lXncVa6ruf2oZUO0aQCA6uP1cVXnqmXF3JgL08BflfoXl0pdm
5ThaSo6AHAbYmbLMKZWZbx4u+OOaoKJqIgaYTSEx2KYKTM9k9Fr7pn4nf60LZhcwqeKy3EjPwjJ0
seNe7XSZ2jSbfr4hh3sQ+xxpgfFCB/LiTeubBwmQtT/Fo1PNO7PjG+Az58Cm5UQx8p88iMRu52qO
1C7nvZrSdlTIWriMICoOpmv2fD/d+rE0/s3dSflO0bS4RMX3MH6DLXtndPavzn/VUw9QKNeQVfEp
37tPPhfMkfHkE0ikTfLCRjL5MRyS0W9Fl9u8+kL67dRJQXSDWyuiGNeiokcoCFHAlpG7DI4vyMDD
wyGu+3Z4UapLq4BTRSh4o1MBJ5E9aNvksDtm388bVUdbjHCy9lif8yvEZMPjijRJoxxsyqvFeqgG
gNEMHFLqYX0egkgm8k4TnuQb9EqEgY9FrM6CwyKzWvSTOswkZ8wP8zdTrRJzmSiFCK1IrjkVet0F
OHgM+2XS97Dr3McFJsu8M8vNeALN1QXJoeNTqy8vTmTo2AHsnbWzVOz6QNybsRObA1dbJ4YS9vKO
m50xBXoNLx/EnX1dSi9vmgT83UJURG7U9Ymc8HgwUZv3C0xLm7C+bBg2D5a2jyOS6i7/zrvWNwfe
ewV7x1SOeyB4Rz27bKxo5R7MQEiSO+TNoNOTak9oMtaXgE1PYndfet7SSplUtTqqbq2iN/zv6DkJ
01xXZ515znKiPmhx7NpA405vdpNh2ovl2ANH1g/wIQh55Z6v79KoYP1t4VrPxM4mGz5VWxZvqTe0
ljfv7BaAkbL84T9jWHL8CtSec0kdbT+784tcLU1/2f6AiiFRCJm3pWuqHfqaUBiUzF3CN3tpCftX
dLWfSSz4o8mX4N/96bgHKb1BTannj+EJ9qQ3MYKkGn+vPp2zk8MIpQDyrTroSRVUaX2TgRfB2dGq
rE1HrHe0d/YYEJnMNiRjMEFJDR7/lwcOBKlA+R/8M7j1iikWODm8QZEl0aFiQKJ7cU9NYgsaXYFU
dPmI0XC7tavPQ/lhf/frDt6iKZTACSQrwySd2HYXy5P9iD6ppdNLLdavm3aPfe1x22SBsw/jt+A1
WuV77+3hkKTTbJkGNwOFITynJQqPuTe0v6fQyzmaHkRXNuqeZUuG/whz8MFJsls/lPGsrVHpk+mt
fHpsDsC5BMukSIbIB/KtCghsT7SDAkce7aWQgeZba5WLqvnPDyRhSCp0suKMNrZ8vN5rldp4uNYK
6VgfnxfqEtcnUVj5ms44pBg6H9AaEdYDHcxj7hVy1bCv3MMMXuaBVYW2BirgAcvvBDWBIzhKF1OJ
aGBUUSX249V/QybnM0xrvMeg4tLr/22dul6qtNtiMzieEhr8zWz+tM8C7HeoHLgF4E8FF4TMh9Ta
pMVWIo77FoLazXXaMD9ypRqy61YePsz/uumMNkMV2vaetupotqqloUbjnu+Lb38mUrpBCQvgYpS4
3yzbItsg3v32hho4RBtUAR7dZ4ACBLtJTpCGzbAgDQtaCzNICoqG15AEQK5iEgyXzbuxXkfZnun1
mTQY+oHr+l/ER+V7kTIrjpglxPk/17GNg0V0tI0oNf8QIhUECQqnPdZa6ObOEwhhTf0KFai4f6Tt
Sy+tDcNs6EwIEmRoRKz1IJLPczXSdWns06l/aReaLcAStHPu9QtVRAIalIIegHrYsxHLxN68s4zE
OXqRWLChY35fXquR5GkxQIbAqlsxoaHOR+5k0WsIk1krhYQtfS6MxQWhAdC4dnrsNWhUDPYtisZ9
pbwLVy3YZEEMHBKWA4shfL5H7ImTIVM1+0/L0rSW6MOFTZ1DOCJbjhdPeoMyg/KDbH4luhDlkquS
0ebgMb045npnPA9b5Gd5FKQSLpvnYP5+FQ5z/u4/dIgMSitrS5aBeRYbmduikHuijMUXm9rF0FN1
rGaunJN0TCoFvU/Igva387pGcGfoAK5p5PX4RSkzUDQgUEDdsGCPyq+Gg5z3HQICgCwKzFtWUKuH
MB0b7N2upiWrVH6PFNbxQR0Oi/z8nn8LxZHZOs1MAwI9erhZvPo8Q+BRdd8vBOOVqYc/JEngqBdk
eH9V7gKbUZo8xneoyzZZjkl4f29MZht9cxw6f97YITeozQKInSN0/htlFk43Ok+FRrSPatxeoepv
k6mOFwDIxUzbxBBarCFMNQEruhmr39I8XFdChKDgQboD7t9EyJ+cpxkgR6YWNAdI1tizvIeSIQ6B
dgJAOt2ON3LaTaTlYwEIPBu+wRNSEzsFVTVIMYYS6ucHjAOzzuk2dfj4d6ChNfc6t21tjMTE8QDH
n7BDWtCiIh9l4wIPcDOF8BB/zMfazlSaPsRKcvsrkMEOOC1ez1mKgFVg7il2KwSmIf17LOgnBER7
Q1zHUdRPq87ZixUBDXboub5g6QRUrjQoPD1qVsI6PfLjL47JMJsSiPddCx10SPxVIZ8lCpMvVZT9
b04U+knOkOwRkwMHmgVEg42eWR3jBygIr/nhGr2mRwtU+tk7rtW5hNuYueTIpK/bysW1e88XkAbL
vDhDjsPVMYFHDl0cNp/wWgmfNyvFkkfGdhwSJC2pHvuDFq3IZ4Escv6/5cMAYvfMbh/TixDhM9Az
VQ5oS2pzdMRrMqxIyXvN/P/crZBOglWsz1tuYykCFPITCiDNdt8cvJ+MelSjBj+wtwN/0Dkl3ePH
yU1Ae0uf23h/Diykk0R9qpN38H21dZvYO2qHXGH8mVsR6u9UijbKUCdI7BIqfB//ArbGTXiube1P
fVaWSODbchYfwKI0PLV5AmwdhpKGwB7P22PoDGdjaZCIA7lyjN9MPh68KVvttVT+QvG5PUGrix58
eElL5vT+4QUaUH1q+NLraNFT7wTi7EG8RvMx1UWoGlZCQOVQYHdNH7fMWNbMpsAfbnC0ZtjLBIFN
frDlhtuqK1rYvYB9kZBs1zbsOsHXKH6uaZgE53xI6TrsCdJ5jqOz0WUu9VeDKnnagxZpsWWWp4Mc
kNes0fnpGDWk1ZzO6+AKIQtZTd9RCgYicfox28pTuN1PE0a5rS7sk6033yYJ+JykK4kmettrxXEb
fox07s/BH0yR17jy6EpTmY8068qgCqClNpx0BYSta6CzNZlKVPHFzsaf0qjEMU8+yDy6XjAkkLHC
0TvCLcq0lk/Ln5FFutPlXiIVJ/zUoOZr1iUAkD6POHW13M9rtAqlbgQAQhllO8DrznDAx37qJDGO
NdOHqcKtlzPROAijm6HzsFzur0bJnBEOauF192nDzmNCv/UgsNxe6dGL66hr2zFYvXqubEF+IQ0G
2AvPwwH8gr4o7YDH24YxBJtFQr+4dQvJn3uJBcJtOhLBOyMwj7+LZNWj/8Tz3FYwjFVRn+Bgu8pj
olAQV89Df/D/is/+OTOiQLkabc5rQTjEzj72AZU98VAYZ+2QonFHh1MTq/Z2nJhjc/jLnPUEeane
2PKGnZdQN9yvQkDr+8MoutSnWRoQzKr3Ovc8ovX3RUvxgdJ+CO2zRfl+Kge6SXV9/Og7iYiunowS
SKjmW7SxUkjQEYUw/LHu62pEgTlaTHh5Idd4ar63M76kOuJ/MmOQrF03tDg3JvaoKhKAZHN7TJ0s
aPqv8jj2OjBqaVeOsdt4iILrZLh96V9gie9+/61yembD4Fvr0djjR3MhI4h2f6lW1dlGoNSh2VPD
QmJBJEACfzfVo814g9fwjOwXewkp08j8MkjPgWhR77ei3oq2TJ7sisn58RV2mBF3L4X5OVRDjm45
+zVsMlQ7rfPdqzxG3u3S0sQw+SOgpeN65GYgTD49eBUYxyhtp2Qnef/nKrPwv4IH7i2Srr8cRiQp
+XbOCxWa8iGJ/AW5FY8CM8Oh/+jTS8A3kbJktxLOcKjEgPbtO1M7C+wtRdz6+j6rE+sqV74ui0Us
olI+fY8fR5p3i7He5MJSdMGMCfBxtw/H+wc+U4mB5Y0z+Wq+b5zgiRhUUu0PkIj35Ivg5OWddvMs
QrixjY3ManhsgbjEjX3oNgaAaVJa/3WtRtxVlHAZX4TpTadealZAjLE+lEUTkia8Rm8gGoDA42KM
6v7azjUbCz5RiSOz1TQpzASFUtwhJgNkchSiFa8E20AekagbGN59qQdV9JVNKB8PchmDz0kAvw6C
AHYLBJKd8wavanZ9xKwtU0a12Gr0BDOslmL7dNWYpaHMCrRBVfD5vUrq7D2QKz14/EmBh8+WNRIo
lCBBOlkc84EMD5UZs9ZoxnhA+Y1yL5+9zSwwH4jXIWSYxC4r3YZSaQbaXNHrdDGtXEedQYxA2hJq
aIQILRR/JxO7E3Jew2/ItG2Adh4LYrompL6kBNwNFvX7LeajEBEyPfIW9KVYp9crv4+jufdvD8f3
h1PQ2PtJ2UuDaRhIuuU7aetefYnssGIY8M74vAvU6nOLJLSWK+1e5MriuYrJRcMgvQZSMTsq6brH
kij967AeUF+yGOAHp81TQb8tZvhRaoYe4o4SfOzGN7E36SoFRMsXKn2WF5HQFDhBKh/k6EQf8hgm
39kr06mDfJoSlbnWrC/YBS3PZi25MQu5RgPsLP03KdKhrC5YnQC0SmZgyWXyFTzP07Sz9/WTUk9a
TT6cUl8fvFz6EghrncNxnltOTy9vNBY415vmUCMkxsDEBHXAI+EPrR5YpQPCZjuYODUBGw5rwkWx
zDzxlc5g87zXomLxOLu4grJahNGb5QcBPgbL36YpLuH31HRxtksR0H9CR1n19qu5+MgWfpSu36KB
GbbNLpXdhEdyT+AYCuEru1jxyKldqhFCQUqkGHGSGS/4TG+kpltYB5WGJ7boR8vbM4skIahcx1nm
LXboZ4kSyTqpBDa2R1C/OWFNLQAsdrOVUyK54qKKiq4nfJwt0PwQbFWktCgCDCw3yCQ78L0/1kWx
kL5EsuCKoWc8s+iDYkglrHD3SZhRD+ioVogpO0xuCDM9ASv/N5C5WopGM1VbQRDoHOPPCLltnshE
cEfHQriwQeQA0UEABBY5JZh4ignTnEJIiSIEphQUMRSAyzyISHKk3fBkN5L+l/0G1YoeHyICMZ/j
U1Xy0INowi3qP+FDv8AXFYOSUmOoWGlJ0FMaVmE0Abpgv8c0zhw3b+0qz5zk39or9vLcR0jtfFrw
zM3Yc5ft9BwP1rcTC2nG+BvLn3dg8rKF+S2S43rEBXB7Kab+0TFn4ixNfTjqAUHGwSZfFfrrSABE
H7863ctBe2y80bC8FVrCg9Ri8CjI84MJBi5ymBdCbdoqcNLMDNPmjmBkMg7LthhhZZaFD1WLwGrD
ZHZxSPShW+iKS1Vjt1fBgXd0M2f8O/jHayN8rFnvegUNiXqBDALav7/dewFbgL2FFfLt5XO76zsR
i1/zGQa5/byDUcAEBPKm9gUj3KhN+Clbn3fi0yGLM+QVKzNspldHGzCq5DNrtl/RZHrpfU2TIXcH
jpbHcIyCy5PAQ/l6c8YmSFcnbicDkFYWeYzG3g6UEbaIVgZdB+gAYn2/YFE+ksOnfsk3iU32CJzy
AfWTw9y9PLJX0fgy7OG9kIGamc25P8mqzwLwHPmSw7EuySRY6h7F6LQMtHcllrohU7Jyp3x64/D/
q3mUIIUpaLDyk0Riy76aCdTIEQcNh88lWGSCPPoA3FbLWeGIyeEuofqqfeROKJQFcwLLyOHCv+VV
NalB3r8s14+yoWfLySJ+zKQdRBGQ3ZWl5omRHIwK6T5geCYdma8zonrABH5FP01aQxC0Y/nB7kSi
PZZ243APWp3fPx1E30tFTYz39LCaPbHfxNoSHhtW4r2seUYoTUTvJq6csH2rVPcTpt+LiQaHki+J
1ot4SfPySkGUo9BlcfDfxbkj4N1P83bYoPEhRwDSfgu2zAQw0NYaH+wkb3oZN1BfJDwDJEVBsMZp
kADPm6RW/P+s8vCjrkIOyMxkbHyygq0y/FyhroH0ZcMrOJTplikWQh1eRUfHOX4vzkw87/0FsQ5X
wg4iiF1+gSwRuszP5qnbLFkp79M/auvxLMpIOmis5V38z4cFFQLNOGqwkYpEfajtXWIi4o7088jo
COpPprUAVIaUSR8nSDLXw/HOICC1VhpYG7cGl/CKbglb80V2Qjom38m4TwgYJmRy3W4hhBYiU3nh
EUzBP5u7PNWdwvzAluziUVG+AMo3P5NZrtJazX+c40BMnkEz2msm4Qo2WapN96inFOrbxZ91ZyVD
j1XXUjhmP6v6qTsUTuiElKM9lQ3J5VyTR5dEbtwN7w5srzafvCuHz0T+1iHYSJQ2t+JhdBwoU5z1
bB/f0Rtp2DlAKjXuJsNJrZj0ZS164hos7073qHSVGVIWkbI33ilFCnKboqzUgKfGCEeuVBXgwUCi
DfFKXGkiRbDHx1B6l2CovWkFxGUA37UDj0eB9NzZxDDLcvrLBCbA0vgN2/k9tP/jyojSopZUEhnP
T83+xbYdZo6aDUKwL+GlVdfhe5hC4LBNDEbTlk5umY5nQl8LfsQXWYlghW/YOuvzDP+n5xcEEDtC
t2jhARnvzrMLPsPU/B+R7GkA2o47fm8Xx7AQovhnjEQNlqMJjleD8RT42F4jIKrGdm5b9hYHmlWt
qszgX18yhRWUo6uKlMq6xCNJbb8lqwXp14NJJMjyxvPJUVfUQ6tMhjFRARlWnFweZbzoDjWtk0wY
2lIT7Y3WZLwOlF1JSVL+VBmKT1Dp3v6dc7RkhxPJRmJ1K/O1U17TYI0W9YH01j/0765nyIrLN5Kq
ZoR0iAc8MXfxnd5g/f0WZjTg0WzcelklDL873l55/X9kACGyVa6fZy6rkgYTgx5QvKyqwDEFFx1m
g+QsJjouGV/eNus9AcxiL0CxYWNaGeppGCK8hW+A/rS/AiaOrJRFE0oEYuvvque/xnWbA1Dwf3LF
osTz8l5rS0vQx5Wrr3N5uw3Bu73o99TdRO7kDDx2bRwSjecNH5V7ca6OvI34rBJ8sqGdyCY4B9UW
deQ1+0sGI5eZnY3ycsfBnBFqranl1KUpUhCkHvcWYLgOxpvf1LIEupK3JoB1Bq9je6AIJk5oU9No
+BuvYEGJKQ3PjQiSBcJC/lBmq7srD2QIw3G/N5N2Z8z0QdT4EaApuK8C1rNNGRF5Gy18qsmXQDzj
8cXtS3rEEjWO0gcZLauCAO9nMKra6c+vniw1nc5clRQQiFj+k0/82/XTvwzAVAvOGV1LytpqtpFQ
CCzvxJZzM/VywyeK57UrJxuOvFo2TRq9ocAVNTrcbbqNtCJXIzl+vCOgNX8GjzFwjykuXGWWr5iP
CLhsrnHbp0xc4KK8VAS1GGy5ehivyPFRSejtSaftnlL+C998+qYx0nZWUADetgV9WblvLBU90+ut
Qw1QA4dquuuumDxTUe63u5X8NAvJ0rKsjpR1IsZsd708jVKRQngkZ6cBLfq27UawkBXSrQfHfGHb
QxsfrjSt2GbjTd4w6IOPTfLnPeH4O+8f08dF0m3BJNYqOehHQiN0xB/586BisOIWvQZLdiozWmPn
Z2UbsG/Ppb09ayV2zI3Qsg58iNlppIob0IN9vOhP9lDg81zMqE/mnyop26QwK0TZKfb0qWBxgBcE
t6NJDDZ7Iizz+CU9H24hTBsMLal7Mz6tMuOdXzpzT0pIZR3mw5xsRJo5OAhhaM70lasSt56pWY/L
Y/zazNZ/UEa5iZ5F+STTQBBpVodINMSK+QE/hbD9Yqvh6sgiGlt7bv4YuDVEwffvV0i7JZjGF3oX
1T55E88FBpRvv/KNdVFwos1CPGoN8T7jZjM32sQr4r/uj+QKsQDu6yYVNigUkQF23swON3JDnzWO
Vq5tmg70p2cpqWfdDxR+cxnIzDpiv6pg3ke1blvXinCRSec/HhhYsYMZdrP3NUNCaJNlxQcTNSyz
QGYcftL9hJcvc/gWa7kNOM9GJLzN5mL0Bm65KFZg6O2da5Yww49cYJM/nKyl1bhr5K4YMLNsEPrH
Bns7BBbDgi5iP9ZQD18VgsvKn7XpYVgYcijZRE+n+FWwMDLVrGmV5DPGvdYoNwy1O1mlc//HNNCT
K/+TWgeXjoclE2/UZOTWx2QGT0vcwW0FGpNdepiwu6Zfh6C5a9Ako+fCyLc7PhHvOtQ2/XCiJdOj
8MafmIJ5x57H2Y6gVui2DyLMhJDMpFlBQbQ5aljOjdgHXBQb8YxBzGvA0vC1ItBiM5s0U+xY6Qzw
bfDO9cotzxyhQJueu8Pt7MZ1l+BcKj6xkKWHfzY9PEVLCfhrzNTkna/4L5eJFQljBbO7V3W01u2j
T9gTSLouG6T8fCQTFuWf6pDPG9FhWjb0CX/XLyBcoPA6h6QZbrELE2QGzjMcwK4epH9ngDmibiaY
Lq0sNS/fyhlUdcg2tN8vSbL5WL8cf3S5UgbWUzaGTSSzT/lp7/14EbNR40h9SiYtzycIxDVmirkw
8d2NjcZWorPkZ+3bUDp3fWQ4nhpalsvnHQ01eLe7NQz3l2y0zJ50InSZvlBVsBIC1ZNR1PYP0DLb
bD1/SgXqF9XZbhM5IiczpEepvaJS18p/m2JUqeC6VEWUzCNHgTo4q/jteaGWvR+MBKButGvSwOn+
t5EM8NEBs4VhT8BTmNNAYwM6niGrL6rW9+GVOKJ/jVsV0qL8FTR/zFeJ+efZHYUOwBi0yKh4Y+FJ
v0CXA70A537dA/GGmPiCclf2QDBp6KOE7U9+Vku4XW8oGSrF0d09hLvxxUEwTz1sRTkOg1pg0jin
YzT7EOMBv0LceCnJzUiwLjYWhphYbsCuLzlBRUmGzvzdf2W6Tdzs2BFLhjdaMiOPFHN9KTgHqfkB
CbG6/6vnarO9u0XI6sRNTbssQV/6elxXkGmEZBq2SEHC0unO4Dx/BPH7BH9ACYcdYv5UDkwALUlS
Up0PAds/pSxrKHLGofiYcjXpp9FiG7xKjGsCu6U931Dy4kbt+a/xpnTljx8KyApPshVMymM2CSKq
+axqvW7gwX0DCEKhlVpySR2+EJajz/9kwHuX5u+SN0QI1gXK38rTPMJkxAMKn7a8aIWOtlTxAcCY
p/2pOMlFPqwd4hhcULuroOSV/25FdxV9Q49wHbvntxGjohsLMfr+0FNugEeO7z9ZiNg3/m4RRJFf
DkwQG9lhFBtFADqqzrlUeasbqN9ylhGMC4Qhj/JVMnBG/vACLRuUqVITgexHSWM3C+ZsKQX5C2vi
PjNX+Z6P2IJBC7R9LQ0rpuCkwMWfBTFRemWW35hE6uuabEbZCwOco7icDp0h0Us62ya5aRZvwA4z
diSG5K8RW8II6lQCeGePW9sGJ6HkMia2hlB/owOLngdQ3WTM0QX94FnGzg+MznQuQAZ2nGFEz/ff
7FSex6yKrjitK29v/qYZw6ZEJAeyLAoaxlQaq9hftrr+6RCcZoQBkPTm3jDT7R9R2XxtgEUPLNNa
o2SUkZqesWIR9mBz2pgabCk8D1ZXBCIF2EG8UGGxGsRMsnHlK4TNOxeJVIibe0E0cbGvOgNfIIrh
6B6AaihZxXmw1W4UWe1gvcG2H+SlbJbaHDMJfov1igH1JdzPpjudyf8b0jUOt9utaKCDXfnstcR9
dknaePseYbkIxUJK1bg7lrcvJArWwyY+Sjb+9WpIXZeMbhGcs7g07UROV06XZ6PozgTkLquQCwGQ
fTiBCB6jaEGZRvEj1ydrmvEZLY2s5iSGSO6tX82YAxSLUdgSHAvNWi7LsYUq8hxS4Caa02vs7VN9
UHuIIN2h0/Ma9hV0z93Ju0oqfv0AyIyQUFy6QshJ7LDtX0p4SpYD9OuPKAACutQ5oMQVNYx9Nj04
2WDZtzdSxyl2aXCyodA34/j3aliB6Jw9qtlJQmrJPhCyvYxQxfrBXidgok9u+aBTxov5qhxdA1bH
rucG7/DwNKYdJ18VAtCQPq8jxQcSqdpymK/JNrXfmoJG0mB+T8BtTAFftk8nnwTo/5tSMICnJZu7
60e5ULc6QOZdtblRtxnCbhODOG7DfcIWmUCPIbPqT2rL+jrHRlI5jddqzQTRneP1ybUtXOIy4wX5
8iwcP7BbTdgLJyoR+J+B2SCeIRed6vxubp/E6qtyuvZ3J3353xug3vnNZX5nVOalOlgJZeqmaO+s
BU8Ya7ViuDGKEBWGeJO3Ken4VKsOhDctKppsYx0uB73y60d65b45dAdO1ciE41h2MuwattrBkQIG
HE2oP7O/jjOCWr9RLyaIJtLFrRhwPnphStFp4A21CBwkrCbSVGGQoP+tGu5DDAsqlCpA7EohQXgh
tpQwj8ogkxu2C/MEse852Mawr0Jr69qeqtjL+D6rJ3xCv/i4+FmUdnTHJAiTzswuPjp8EczzRN87
j0WdObSTMpY42ZS/xW/N51C/HpNSJyApN4zCd0Fys7ZHKLgFhNWllBW15ZfPfRH34tI/NYyVC2ZR
pK/lrsQKY29YYFPT/nw19RtyZGcuTnHMnCc602bFlcOGV2WdGq0tM9Q2NkdPmeLoQ5Pj/uJHhEvN
G0c6S812GS+mCrcqdM9FdLs/sVgaaMYCAncDRKDFQTJSuN323ib2YsogVMfwGvnVTNdZ9OpQ0/hs
yL8MzLMwAMmLZQU6n03m27toQPQFhyCUtd99M5KeXbCgmXYpjMSlaloDvIuwx7fNK5RW0CZGhChs
IVXO7/1XYwoBlb/Taef3pP8qFq8ujHlsRRV1dP4ErfG+tywK6mzY8Z2pxUCZ9CJr9DOlOwx8faa/
/sGnH08p/UT0X94y8NArFok8sPRxSx5K4v4Q0kl/nYTo0xXivTHHnR5waIYywdrPePw95O78UYHX
g4jUekoEicCmWhSwwKYthZJwgWEY2DwY+ebdsuHdONjpRY+ZlRR4Aa5prBth57iwQ23fB7kZLhaI
yIASy15mrfLxi3QRd1REnz5KkCK50JqwCK6WqEgDM/j3hC9YmhZQrJitPOQTruRxkdJHc1sxu2fs
AX1NrPiPHVESvu3r7+wolpXmSNXrIYlPk6Dr//PY+gmrVNxbTt3PbtSEjsrvl/V1DyNmdqqscpTn
R7AMWjE2tzUFVmQMKE4oZZ3H2gdChLxHIiauFPwgnNhyhjPqCtJ61BAbeUKPuoyoQbKmPdCwjXvX
zabOdB0I3vm4boY/124IhSSp2KPwrIRGFbOnWvS7e9dSFpSN21eRdWGOHvTia7jJuoGyu2CgrY0Y
s4VpCKOD/2QD27PkExKPqjd7pjHicNt/W+VxQX1oxJHZNjhDty2CiHuMi4xrHIOtL4qCOSCXP5BY
KkoS9v+oDpDXWr8dtTzbXb8GIcwfady7KQElNtVhqjBVYO3r7tTWQqXe5kOySLqlodCXKzjsL1Am
UJoBdJxkjrI1wZwlqVdAAtBhPTXbRblb0qTBXywpMXnPKvzID7p0/2t8Vmh0ZcLovzTcFqKh11f4
99VCIxOS312w2QXNZqK0XPvmGUypznKuKWpnjc9ziBXfvxoRiZTr8bbBAVZ36PmZqzK91P2DYoUf
Rbc2x+jgVlYIz+N0poetiXV/vTcKqSt9OMvQNb6U1Oo6f3SEKZau4ygB0V8Dh+ZjQUIwmITNUNr3
CMosAn4xTmtwoP0GXJP0K79twJuK/aWQAaeWFNXI9tVcdowJ6nmKJU0zy0tqmEfon5sMRqc7bXyk
8J5xViFUo5v1DDwcdIbIXJnCHmgMBrqR/Xdue0SqWoPZW4ZdCUBJ2iFFBgdLkS8VW3WcmLaNOUtU
gkn5WwQS/I3JzDlvS+rqUrPW7N4KmS8rkec1dGcCupmpWyFzeYrze0Azw9i8OV5Gj/+6H4Ib28UG
bxH8LDnmPx96bpbe+AQmmXpB2Pi2ub6fa/MKYM4km5XHbgO4eA/3bOucB5r0QRPqafrMn2FcjxQn
vVXi5nKMIIrxM5kFjvZRrsbfm8a5Wh84fz4MzqGjVdpysfY7B26INrxsJByxRXTk2i/d+fvTlMQH
jFCYAh9PNsA2eJMXgFuOM+jVzxCyPz1W9D97heCFkZ0kmUaD/q+gFRJYqJNrNEJJ8UysLh4zRy0n
k4hLz1OHw3q0k/kQjElY3d1nv17gB3ScQ3iVtFZtbec5lFhhDs7PUZPhd8YRmWdpGxTSJ0qa444c
bxyCr3MNstj7DT8SZ5CSt1bRs0TJcn/w9iue+IHloqnZWIRz+CxcOUOiAO+1lXg624fDy5ilTkFL
sav4zIS/bl9GNK1bt0pBDnaId2WEI9VR/lwMvRVGPK2CG6wiSTYuWD9jfFsPHFC2+9RKNDmlOVtn
jgOhsJxr+pAQXmx1bR/9pOzA8SNq9f7uPARG83Ma0fzIoc0r1krhBplvICR70Dt8vxjWDJQnwEQI
XwS6a/Rm8eZCQdvgZucPYJI6Q1ax2M3d7VxLHiTwKwVyZdI/q5e3sN7fkIdFRPJz9qWuf4Hu1lH5
DkgQ4+HNhQDFJTLmwBhUPgMlhUNI4BwB7TeJYrhlS/59Sz+IwkHQ6EnfkFu5LE48ILPzTfWKe+zZ
/lYE+6UGkZqnZnO5iKmyNmTduXkdKL66MCgQdv4tKeVZMbV85RNxv6SFu8ukTVV+6xU1fxJikVWJ
KMbysYwu9jaTtzCkPrVUOiYDKI595lN4ICGBxVmHteNqUIjnAr0d1mK0LW0YkYT0on9KoWvYaoN+
9YLDpEcjgnctqCYXPLHagsRZMhE4cdF/LgdOLIiJuGjOLDpjaT86KQCstV//vYqN3ZuAyrovC6MI
iE24jEwv+IfJXYO8XTnajepgN8Sm/Dnxhf8KSWDdbr4oUsHRK3C+VD7/B/MvdC70Gs8NIhywrgoa
LaNXUA9rGX+BItsgzpWqqQY44R8MUtUSrCNvnF2zyT0pgJZZXjIa0XO4zoTVtwbadCvqaYloC3yh
Gg1os+DBLR2B8EObF92X+0/y1Mfq9gqE8/neClc1HzWUl+W3ZOU0n94wc3gPsgTeJROLNB7E68Eo
FNt9Gy14vqWULguBm3a0M4xZW5EpEMyq9vrDKTJq8uxUK/GauSX6KIMJ1QH7b5QWFxa0HYeqepbi
W9s1utxulCgdZWXV0MqAYfhyO5AolVyAHkfC79iEnyQpsFAGsVpcsAEGQe4yEpHxzvHGZufUVvua
Q7QGsSCkB86+N5s2cfJfrJMYf60AzSkQ+bqWrnA1lKQt/ItNI2VRmfkGz33YWkR8/mZO2qDv7lho
FWUae6UqIDtSbA/SNOtbWOFuLE8Tesi1HeJnI6Ve8n9TZJdpKFgmOIAbvqNN3Zwzae2OsVNIlzHK
/wqhwTz1iD9axl8iGPR689iUC9xpj3ZMSYiek+o4B5xGgL/fP0gz1KrfcJBHvb02v0eSp97d3m89
Tu6D9iaB/L2zLns05pdiQRw4MCFh96s2EkyKzF3qPRDvV4j26TfyRi664O+L4dNOAD0UTr4LxWNn
5g7xS2aPw+0UYUcNt3pqCMBtGmi+VYS8L9MHrO9M/p6HQaSQLDepUoCRC1Hasj2ex+WM11eUlJRb
YOaMhgNOWc7KifJhF0MXjOcpOuRp6TiFMzlVmRi/Z911Mo11IcXYLPkPs9x/BMWWD6TpWbe5ORxl
5drFZhEOU9bdoUcUg487DlMptAkEO6Ra/1iG1nQ6kQhA6MHGtP9DHm5zcJYNd4++BUnFBE7B49D6
r7KicL6Tau14ORfT1WwD2Qi0ubQ5B0TsAre9R6ZIu3hLzvCbv7NTjftYGrx8EyZ+leJUAozZJ6rQ
F0fwA6YlRFHJQtp3jqEmvjR+D/HHItDqBGTwOwebkrSWR9B+dUg4FBNzzaR/Fud0JfKaK1Qs7rAG
uJCCG/W7xj0FXftFuUnQuxonHO4OTYMhg38s5lBcH28okR1eqhybmzgJEr18L87Ckj7bv0is4hmn
BNh03TOq+Uc2xmlntTPzvTvCFMduhPP97TLAgOtdm+53brLvr+3YLeivLUCq88lVK6fnNiunDoXL
AR3vXB/gST5oJ7qDzEOuUwlGLAq293iNXS4vDZ4j/Dn5u0l5NBQqMa3/95XF6JNVndOaoGbm9sxt
FLr5jCqkaRfiOwwD7NItvVi+xEbOp8xaStnY1vg3E/L2hTTlVmw6mKG0V26nhTPvvS+JZTy7+YAr
qrcAxUbyhQAzutrcUlWpTGp7wGIvTZ7A/f0+SrzffE2AgLR3GEASlOSJJ8iKfcs7oSlssfkIY/ef
Z6X7bEe7LfJ2a10z7rfqjMHw5elsIAHg3niio4mlSjzNeRBgqmk4aLwgryXiEkM/jyPynY+sGGu+
xORV7VgSE8EtHBZkQLUrRQMHwRiNTakBB0AQJsZcu4NY+uNPh1kt3lpB8G0+VvF0nZd3kjWFeTjh
26y9SHNCrZMAlCSKFHQxv82v5tGP2h+Qgdt2RQybTyVW+ka5GDTfaRrcLGsmJ5BXYY1ZJZaw1soy
IY2+JLAlNe+T+sUT9EF29jzJTzUBMqOkaoPZlEKAgRft0zK34QNtXhu70wixWvjmE8U188caCvht
LLsZjW4MwfL1YyRUreUfTRk4t97j+7vR/K6XBTZEXjYKDTecknXgZpnUAthAt6RctXAMd8FyZ9Yn
Z7LP5z2r02/03nNHlIBCLZtGxrWvdEaAw5zOjTLozG2RmKDUKQC1O6UBaBr+Ez3DcQhIrK9C6wSk
R8oY/I9rphFYo8ViGmIogsUEO6o4Qzvs7cP3ehPAv/0ifaeAD4SXbPyr1oQrzu1dFB7UsPG3wARs
Q/GMp/PHJQOXQ3SYMhDnJLTyiutiF1lI0nyDQo0F53wumdI/DBSxC43/RtHlEgDLeMJe2jZNmUy7
Cm4mMDR+DpUmkl57MTSHQtbEvN2TDxA+lqS+Sbvdx5hbP7yxFWiAH3yPfN9iBs29fVxo0CyAzBcE
GajuRanANTjQoNDm3509/0fFXLSmw91iF7hIOyXhkSA1Jd6yWJflNtRMYA6eZ5MbpZYFxOOxcZzc
Ei6sKRDT7gVqkzhSFMSzNysNzs2p5z8dXm+SAiPf2mBODQwrnG8CHcIDAVVXDG/VuUO6oq0vxoRN
eZvc+OG91fh5k67b+Yt8UlKqeN6tmnY6sCHD6cRLwKzS1H3VxEjJyIkIwFw5BWa0mqR3tP+5QKZ9
IeG8ohIuBIt8AVdhXBflAOE5S1PQ4yO8W4aOaQgDULcpaLWE9Z/gPf2oFRlk9yvQt5oT7BNvC9TD
PRBOfcbgd5Gmk7ULF93NhC0fDkSyscUDhlrlGHvf76tCdWuzts0mtTICUbEBt1Gi3oAaw3WpBaTN
nuB24Hbt0MjlUQL9QmHXgXxYPYTTbCtuYDmE2a66VcwiFFsiBszmB7IzHh7ue6azxluvnwFA4skp
zQ3aXyvHYoedGPV9LVaTSGGym4waOms1dHm2sp8jsbG+mWUv9DTuHRuLaVzItLLgVA8giT7EOzKX
8FPCsN8kY7r6FnnBWC5HhPWxI7rwmeoDB5CmX8MosBSAPIXemNP2rpJHJOBYFi1Z0IJYSFf/aPgp
Ffx+3nP/iz0ini4xEpVYCenEMFWaNap0k5eEDhxUCxBGIN7cG6FwyMyoWMr0niI0ZHHa31CHlDKt
KBi8E9OBffq3LCQXWL9gCFybUMVB5uvUOPyaPv1Deth/nN5fRWjCgmk6YRV3uUjC7oBtZZ9Oiezn
oiCHOM+5QimnrARza8VdkW6ch/9+ut4bmlmW5ABQqVfQ8PLK5+iM16Cq45JVx7HWnnpDmnhrgJhT
tbOkDDAPq85cOCzTYw4vdtg+HRdplNB97lIgOM4WP3GexEyAqdDKIZDgdMyo0zmBdX0bJel0Pk3o
0MKz9iMfaDCYI2tFE21V2RkWOie6+6dpU0uVCPdE9a4i9I/5M9xPRSZFdt8CO3sqePzeRCiSJcQe
1AjnrhFfCMdmRdztNGhtpzE2NZ9R3XlbPA+LvLhB33jnl6ukmeA4zWQmnjtVEn7H14K2fXCaDeX1
Bt5juj9EuCrzqMnBDWt54JzjNZPKAQ/s4lPBr6HGuo0x1r36Qy97h8ZbiMZpFVFwlbJvkiWkgA/b
eWeOZJ5HY3273CD76DuTROIuP340sr5tH6/AzO6k+FCEH26kODu/1aZmzJZuCzaOq8S+zZv9LPuE
uOE0HERGdeapAhZS5CrjuZMBSwziook+In3S5CJkgVZRDgm1qkeLu/8AnRsUF6xesBCCX7ofzI0o
kdjVCs6aGnIa9aWC71dxO26z7PgfoX2dyas9kGKgHLjzxQ5ieHIXcCaHMTvb5vufGpkALpbqLMEg
O1dMNTQioYYUJJATXHADoX2EtGOUD1KelwhAqRJHjc3P8RK5kEaMuBn5zEeN72Ks3yjpAsGYX+Zq
m7jHjcM/o1zo0zSNddLGmzAEfBl3Tcdk1ZJSL9hbFu3Jt1J0xydxAdjOMxDpl/HV1EkG1bpQZof5
28FfST6sHpcLo8OYnXr8BfqwUnjsCA0bZDnAt515NoZY0L7e3r9F3ubz3AsAPRK53GDMgv4qjQv/
EkoGr/lkr5B4BgFgxbJgBvBnmn0gnwvu782Z0PxBGbLg7kBdvPcx89fJ9uGx5Ax9oY/AeWqR1WbM
ADEn5P/wk34iLgtv4JxpGHwn+PzlMBjKaxKLRTuTfQvE65JUxA6YWn0aJuateNPON5ESDXUdEXYI
NbKlJ3cNctUYqPyx1+PF+voti63dw0Jnh+axh3z3pCJ0qIOizwmjsnR5yonn83qXrlis+P2HzFGa
Y3TB0OShLkLvV5raJz2hl5SVi7hyjSrs3NZIWwxALkGuK51z/wunvQH/jcFY89w4uHiIaDubcnHB
Fzgzusru34o2rRBmepOVNShy06384NX+5UKrwVagXZojR9FU2K76WeF0h5r+p1y2hXq+utQf/XJA
yaBGabf30e9INBNiDueI/g8iOExIRDn3fYwVez98VFPyrZRweevAallBtnZNMjg1Gdo2v1KfSe7x
GWW/PLWcmZU7Sgd8KmEEubmORUXQ2F5OVOpoVYp3lVMhy3hdnIpfJWJ+din9Fx3BzuARXeCT9h97
ryuqrDLLVhi0R72qLTdMF/mrKziq9xJkgJhtz9VrUVDT2T01TdGF4N4cePVplHGPHi9+fsKVOS6L
9LY5mNuGP79RlavAtfAFP1XjcIVjhahNTYfQ8GHGBOD8UFCaJMHZWQQrEc2y0/3hlOaiwdY+Jshm
8R6v4vgzF2X9bV8zrX0t8iwqA7RP5cbRRAtH4Ow/QbuaYhhSygENeIUlZyoM6Em6B6+AhsdqMRiF
G8kyXU2ATDpA1G2BM+1vlCwBVAbC/u4BcrXQYKkz50raxoDOIOd8vcKcj7Z0ewlL3LSIGdYlwt3t
PEO8ZUrYLaJ9YUSyIy0IshWJoKN1eRdraaJ10TXBCnbmye/ax2MwOgLIVBcEfhLgIswVvSQxywKG
TvoirKe609QoS/Psy6uqf9dfVj0MXaFiBRHb2C09gL+q4Mf9uVtET8buobziy7/1qunv2n1+ItU4
P1tAuUsN1Zm/qRtHerQlBk+mq55KmL9j/1oTbiqStfc+rh1RNhjIbaIDstJt2pjPRTDcEvAMHB4m
BCrpd78oVe5lXOizXbomxgMrke7QJbvUOTfJg0tV7w+8dTWYZCXkU8w4ql/5i7iKk2o5UF/gos+T
PGqcmsbxgrw0eqfVgGOqhVkaE90HYRzN9CD8zWDU52ZyBZBXHnsYKraJ5axkvqFJ+Tz2Bt2/XHV0
jLkX8pQZbTG3f5Qj7fp/UT9+eYnsABYM+f0DL5Y1+ZjmkjNN7JKOzE0xSDQKyGXwxtjHI+s0OpeR
02FdrAY+N0z7hc4FFuGvUIdZRYOp6tbdV8z0GZRNPIZ4FZ4HrMyTP3CEf8BzKeqMRDzNaiZ8Unnv
6bj46u+kLszqUu6ZoNfMtvXho7l3pB98P0Ab6cUPWFGUiR7SoOhq5cqugCMYXUib3FUyvAEk8uDO
UMg9Pgi9vTMjXkd0V6l9P/+zY8n7Iros+erz1wHu1A/ni5P9ttKzvprL21GA0XsDAiwXkSAdGAtT
X4Lelvw7Ksx0WmKMa413Wv/CjknFRP5rH6l4uLIXPNguMqUsqqo/om0nx/Vfo/TrViCaEUBTgXV7
swRASYzkDDPSyO53JgNnLcE7Dkcxs1Fih4OSvyvFlXBdhVaVJ4WO3BPKntDoXy5Sn7LfZ8HjV/UL
Z46/87MRcBpIFvvlHgAtMYSQYNFTyzdACt7NzqCEpSMljzun+V+/p2b7QVnKWvjGZY4tsZW4V4sJ
FTgINNkv2cPj/zWpCtFPiSkbKY4prDn9clY5YfIigEZ2EuuS7zOC9xdaQYRFrKEukO5odzNWIpUI
9CaLm0o1lUjH5p8uLQ4laUL6F2AADDzRBXTZu2WcvNEaK3ay+UFHGiVBK+5URftIg8vxwU7fSzHX
01e/xl0x2WMjRNNbmwbHJmYKOhPNa0nw1YHu+IFsQBB0k9RLqcm9AxyIYfXlwDYFSxgh8BiSv32R
JKEoQWDIw25iCGzGdcxSvPSZ04xDwS4vmRK75YbFDE/QwYd80S45Di5ytSNJUzsqhW8Dq688Waap
Rh2T8P7Cb8T6WMf5GWVGA2LCY/8ylSxUU6ZHI0J1SayRKnq1VD2ZyOmMaVr+E6iAKGuL/CCR7U7L
vICFAjccMWJMi/jSyMMq3mLCSwTWrsncn+1QZZEq/fNjhZxBw7LiP2Z9r+p5XLVWYtVTStK20EgN
0pr1vlXloOVRVdkyK5Ce2467RvCOEo0xXFT3nDA9fZ2M0Gwg8OMxlN2Dk6EKvq8EQi1B4dqPosjg
qga5fqwD427yPqhnyvuYFs5IkyeIBDDy4+IbnWbSaGQIJ1HEf3L4cEE+Lje4189ckN1hLAMoQk8y
KQN17jKxvz1F3XPQrIW20ZIGkVOHHfiZSDSjeJb6LD6ilnaE/u2oYU+QB2UiYuZab0533B2oZ49H
nwmilTVyYb0GjaLulcSZ0/n7B4psLDAU7qBJslOLPN9MnT3HixW5PmMls2ctE9Z4vsLihg3z45xp
v4axpBJNZy1dVCwN+veLssugsuj38OXX9Qd+okAcWEwWbur4xXedUs7XeLMgKj/IPLcj8BUUYppv
W+PPMVYNxTuLY0ir1tcDUQt9s0MquCJM2ziH4hi9/rycABfeCTzpErsc5gbqFWV2LxdW5Re2bV/K
iaXguONWw8jMoRCsSDZJsFxyAav9i0XJeleXHKdJOXawLB719ev+JRkFgpSV+wP5oBHGhYU1xcgT
SKva8VSweEBI0fJUiUViTnMsUq2A6cvnBHa5Svyx95vjUfBYHIjqwtpkxmNlR+sveAUPMIjcOpNT
JMVCPbrvXJBHiUAUDqfMApoEwLog0H5qPG0UP6zNFbAStoUoW5POALCh+YW1AIWF6aYnRFBiNXFI
JHaWieYSmB/gfBwDTb3dV86vusd45ENP7ytr2eJ4xRwou1ijx72PaxHw5LDNFM//Tfsn1mtNLuyW
8+NzUA+5RAIACLQ73JoxnzicrYDyPk0eNubOgCXwPrbm7xqswLVm8UjrLexo6YwnFcJQ9ALeRqK4
ETM/bGY0SmDL8n34JwhpmhmvL/ouoHDofyue6Dy9SfSEsguufYUc3QislQDZbtuQOwk1RcjXqSsa
719+UB6OYIANXsAuT0Xcd2+RPD/9qm6iAvgX321cuotmalLoiCgNf0/9YFcrZXPpf3I9892VeTWT
MCfEJz4BpUQziuLm7x2UDeIq5pSTpiTgD7E2lcCMLYOB5DtcQjpEK32sFhoPd4NGwxkK9SHpw8DY
km5vBZ+YVXWwVH0rOz0sXc9+0lyxK2Hq2w15t2J+pZNwCZq/1poF+dRodmIs6D3ctmtagyjLCS1e
+sN/r9QA3DnawC+aaprjuPBBS/Jcg9X+FhF2HhUG/h/sGgvLoXNGiFRVdSwN9sRqY16yGH4mpaQw
AGsELqlGL2yi5/APuCf9aYbQ430uLHvYz0kIEp/gdqcQkmBc/hMY7fNz5hnM5C02omK6e20eHm0V
imC6vy1ULq7gwkvr4I0sG+w1ZMpch3kSRcj1owlqMbR7lTfvkGo5lPm2TmYGBKjvdWa0vhfBZLWU
yaEAah7K8xZLDlWLPyI5D+XMHTQKVX+YG2GHNzgwouK1VmOcqFEXSps2sBFS/Yu1BgScaZZV7W6V
6+/9+JLgG7OJJCcGnIEos4tybLRMa0I7qMxDmonnW8THpjyDs5tour/sC579eQZj+Vz6iOWyPpov
3FivOCeyUulePJvelsM+QCM/q+sOoknf9UXM5pq6m4bfI93QIXuub/SqPlqS4ijHKyToyY8VvjX8
0kYkpud8rgsh0/c/ja6ZYVuQLSNhE86gS5YuKorkLswx3tC57cvKs6Mlxes55xglPeuS3Ro+7zX8
NINwM8WcRLEmi0doYe+giI+euZ5aXrw9UfPTJl+Q0XD9gbOLRYulUfQVVUfPz8x4LaBaCQanBFoB
gBbArTs9lvkE8jviP5Ux52YdR7cRQmZtt96SwpFb6fu2G4iXmy3x4YcOkxuYI3ULsCxgX55BeUtd
KFflyHnoKXNMU+PY4h9+msgopTH+rWALyIlfw8WcqsTAoJEZAijRQQGbXwy8Au7sJuNtoARlIM+W
/8jBbGzd3ZoMOVcqOHrguG1kxUU5EGJITdtZ4qD9ZA8xHKG3EWXaL1uuSovYfu8+ThN7imrur0n0
qhzkpsjZveLWFFP2xg27v/l9j22uqOrCm6vmBk8VPMlbV4vLv4TH9qK73BEKZ5R5K2gPLh9f3p5z
fclTwh9lxgq8LDHvVN0pfJAl8wYjKVI7fgsVDuaUzjRraEnQNcAz41NrJzX9lZhy1f2R4dlefo2k
fcVmdp8elOLXLk5P9VgExOzOXvNQlhjI0OHkQXM5PZTp6b+AR/qaqYUYHxoqnUKUiEjdzJiqzXyY
IKV9QyEUhRt3a8bgetpub83xbguqh6Io7PkkWxnZEX7KixmpjWWh0dPSSR1EEpVQJl1vFf5QsV8S
10Z1wXKJEiZjiO7KnM1/7fc1Ns5VZTY5unCEF9Vupjni9A7vr2Zv7IpcHWYGqH1IE8a2LUMstf1M
OCcpguuH1qFFN8v9Ubrc/WSsUglaOs2rYxryRFo84y04HGtcL7kSrlPmUDXxU0qySD3yA4+nddmi
HPclqWwJMkWa0iqDwjEBpdoy6MfP0jAUcL9f+OiopOtR+HHujkTZoJClhPtEJoJKIAnihBzCE8s6
WV7/WYMBngZY0fe57NxuAct6+WgUxinbeHc6Is8JU57iHm/axxTg/Zdf+u8IB5NeFiISep0uEQuP
4SDENqSytGYovRaNzgZ4/As05RPkjmG3cXHBXIfuyynEyGUOWfYSLyhDXd5ITFzS2uIipuYJudjS
7oXvJB+3VXDkNKyd5BQ4vGE0tLCao2hAyvQHSeVnUrjTKNZqB934BWOuRA8xP0/QC/M/hN0IFHJz
yMUTuPMAUS/nhuSNYTFSzcwQo3M/NXq8MX1A+qsesBLfLw73+kBV6Lh9M+sAq04V69fGT4oMS8Gm
aPnfA7NdVIZ2x4uY6MHC/EZHoPgNXDW5SyAOIaocgnAo9SYokmNuwmJkmc8xVJ+PpFz9Sh6wz4Nu
KYMWbQ/wSAlOHbF5IQ9Grs5DMbrRpAjj18fI0C/6Byr+GBwHkYdLFu/a0IovIRTQfxiY/hLn73P9
Im5MKZuQdUz526AgzgXo7epts689yESN4cM2KaDv2wsqzIvQ5qm9ESsmrtyZE9MbqALPtQLR04x6
kiq3U3+usQ2ymUZ7g7J+1A62mydSzaUxtnAN9aOXE7GCDS+krc5PQHvmeZTtWas5uNYMaQjev8ge
e1xr3RfQ4GPL9wGVYbucjNnLa+OBTX1sLQSvBT0f2cdjcfjSwRRfYwB/ESRjOEIJ1Kp8Cd1Q2p58
ce9m7q3Q+cs/Un1PHhcJvpc54YdAkXjfV3nUPMxUQGme9QenqjtJYJUC4RO4Ow4e41TGK++VFz3z
L6ccwsktAAiacXVjiDXSP7GyMAZsMMvLhthSTLU1XaNN2oCBk+5ygNULmiQLCDYpTIuLgPOeoYhc
9sTqiaRnm9MhFvIOCV6nHyMjURugK9AkKPyIeog+DvnBLlg+ieWf7YIQplxBbLoHV7VKRGDEj6Ed
d1gwVMrQXGWZsyQnvcdIQXHDm8GAnLTEcVT5tadN8U/simKs1HMzbWG0kIzwF9aLHcwybire2Che
BWyAt3AbLIzKQggw7IUpRXYCPmzEVeMlyzxcfgjLuSo1z/pT+qdvhF0f/HgFi9jheKwYFpNw4795
17ZlSdExF6BRKi3uyQuybhUQI38McOAI+JI+30yIuZK/br8SLJrwHVNPky0Gr/3fS6kF87EPb5Kb
JhT24I54Z763sGp9kI9r3lnmSx+YpgYU73ltN32R7Nu+8n89GzUX2H21S+fY0fQQ0d/MqDgRoKyP
T7HwHskakimNJb1hlAS2LHvNcJT529czlbGF2Xq2x28Dprqe9mP3BrjU6kt5QGJ+QRXk0q1ShGmk
ESO6m3WkSUVkNdcLnq222bqe+WOI/nlHH5T2Vpk/Kmo+ldLg++Fw7D9OJC1/2a006p6SJzx35m1h
n1GBGzPxNVP5pFIsGLXrT4Z9+OrujF9o7qPplWmLVSDFSLWbCEs7ilPHb4DSmiw34ksZbrVlIsvU
+zuThk7jOFP3NZ5qbPkfVH8UEmqEjt7GESVHZAmk8RMbsiVTKv54TQHUhuVOAC0X0VPYz+b46PNQ
kzw2+2SoZb9Fy2f7JyeMtWk/xvyYfFECOMIjGvLns5pvRXnl31SRBPe0JWWktU45MuBvI9O4jtj4
6L21mZJJHuq0QCUroZNjRvAPNN0Pd9GW0Vo4+U596UH265CohtWTQ4ksaJxN3EGlwf4lZ1JzmHcO
c7fAZsss4JrGXVZ9owN0tG5J2dPn88ovwTX2HRbYImnPWq5/iRcIfeB7jaB0w9zKSuun1jwelo3P
nA/u/x+GzrlrhGHP7bT8vlnGXYIjG+2s21j2w4i02/xTI+29GdoAQwW8Z0an6eC2I/VQ219OUbCv
1uHh5WjJWP95YpCtdQJgh+w9a5BkG1Mv5ZmcscbhOPQWJPfl26lldiZxdB+oC6AufHeKZL+73ss4
dQGahFce6Sc/36N9v7MJaeGkTwXONIqLSyvOm3Bm3s2KIXFuuI/u2bs6KdXy38EsZmTNPj/w26PE
IzrzJ0yx6omNXoXavgAskvfRb5jLDB6l+TVTyTZRZwvn+Uv4zqCwaleDKMprhssMWUKNYOoLgYQy
A5H1RLzAbtayffhQvQw99d9ODP5RAUOCafRV2RZ2bCAMSkXR3yMHWV3uoOwjHMwnr6PiLvHdZPNn
qavmfa3pJx8Fn6PdYLQ0BFaglsza/u+fGoPuZmZPJcs9XtY9r6Ya4tvonFoJKP5vdL4AZnNP9mHs
5CA5ApUSYavE4FHfwX6GiVfh/X6T/lBuzWk4kZKtyh750Z+5ghRKR0BQXY0SU0vIL7an5QzHVX5X
4yfemGI/FZi7OdkR2BGriJbYWbou4QB26iApn5MDpHBkj1UO2esU7sEa98HGMrH5XVI3QwPRjuLY
DfPBST2copTBorqnuPfAkY8AiTSFyAjs9q2/cFNSJVcAbqdCulLcSxx9RgDP7DIaflVF9hHzsYCs
ms7VazbHtqb6CXV/PE+ly1zszZU5pKkk/XifgALbqqY4qw0FQYTnyKiGrJUpN+YB5RIOsmxm9UEN
dS7G4EBsjS9j7kfaGBdF6EYX5mRYCVS1OeAPNeHeiPltcmqwvP/L8TjhwjCbV+CPE2lvyMg1CzXs
wYRaF3AwDV8zjbbisTPryBLTXBRrPE7SbPXN1KkQtsQLyvlzNFCVEAQCJ8Daemhi4rV0JrQc5oEd
e8xsuz20BjIeYxCjjoPR5QARug5ZlGQsogX31nVaokTz0m9TL8Sl1LJi4Ab+8tBz+dyYvbe/kBrv
Q8PjdA==
`protect end_protected
