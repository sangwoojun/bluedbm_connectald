`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mHbrJohU1+NLW18uCOXXqnJ8Y8qGd1j7SK9CpvcO4fZzP7H24vxhSl56CC+ATURWdynJUxjHVY4b
rTOO3nLhsQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PNpBjIQ+TAKc8qR8G30piOQCfwcfKahW9HwFftLzKDGUg0a/kOOeaWrJMK4oCip8wxctccjaAJQd
TZqJZTZOlqggMrwNYXp2YMkPpzDtZa1/lMk9dF5FgC2hPG8VtsOGc+vqxIuREHRYGgZa6n4NqGfW
6KpHOzGWRZhD6D0CypU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Y+0AjYa+YDslqfuztnYR7KTgIyBeYjSpeg8YhneZHvAH+f097/MMjaN5dEKliWhWtbnMuQGpPGP8
k35WDwY3sV1eQzlTbGvPG4vXoCyVyctpcVYRKxC5W370SbsATGBPPTDGYxx/Js4ktfWM/zCRdZgZ
XZ2kRYmT4rb2vtk+/kk87aJUJTaARgm6CGYW2CVoRYXfMu9KwLxcVmg+hLsgM7/+hg/zawIbTPC7
sJ6eEUBPkcR5aY7N/hjQiSa/u3n8c1ddRe+5SPyn42O01lqQrMJvmD0Y6ff3xQFIAIxJpeTmkTGW
tNjib/gv8/LFX2MXsQOKSO5JaLSjxlaca5AkKA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pdu+tE/nNv+AZu5q8V6x6FVi6/RSiD675BBeSBpVXD7fPWOFT5GrgOb6ZkieZv7AkGPNFyejUAnO
mxz6nH/HuQYiXIn3E14XYuzD2L3pm5UYu9iJRanZbv2WtOoGxIzmwro0sk0iEVSaM7ul847xoKO7
iFwz1yGSVaOTNC9f44w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gzF+D902W5+eS1a+HKYRDmll/ZcALiUUOPwkJidQgzPa4yT1AMSdbO6FhZcqBsdRq3uTGBqaeh3T
g1v7mHyp0XEbFBr7YYurwMesI2RE2k43plFRU+lSSx27YJYxawssZuVMUKDfUT0ttMjeaxRrS5WL
+d2Zn3LC59xAyHqG+dl8WOSuQpWFb/1D+A4c1YlyLp0PQ14hgtSPVrj5dU4eClKY2oV/KG287fds
8+TnfAIAEwAYZM1Khwd3VG2JtUrriAFngYk4PEPoyV6qsg3Z4TAvINU4mitoTCctZTFxfuGbDzer
kJNYoYUbna3O+jUgdESWI1MHA9kxJwsAL5L+8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 51440)
`protect data_block
z4zP8FNwowCDDlDXXYm7dvutOyiQgTdjpOaPuRn5NGKCCqDN0jMDIWCNAKjUfYgrueEF9C13p5Ir
NqE6WX9w7i+tREjcibnAakpe23g4EBJ90DBYOODHbBOV+6I6HvQDOqlAqBNTaQ5m+HQYmQvCjurQ
8VsEUcEmWy3T+ZAYSsg7sOz3QtVDqsNwK5PVk0SMFRuDWoo53OBtv5hSXwPQf7TGYJPc4q3EwP3S
up6dhBUGAsbB7JtaW7sm/E5MQwJivUm4VQtFWDHiZl2seijYqlJY9h8MXzaKE/j7Amskcx0FDY7G
CIpB7e/VWL/XbnXpFT3AD5oJwVB6cJAR9d30yzrsnLuZvJSfTEwzIe/Go3YYYypSDZHAAeTmRZeJ
9V1XvwK0SMNWpowf83dp/EWLV+gq+W3v2kkZ+X0/O4iYtLjejPOZGp0tXm4NeHyRrk/o+G6HJovh
WYB1B00PV4UtdQdqTkeKMSVZsfPUyBPNWvIXWue6meBxlpI9j3ntg8wmxHHG8K3s3PqW7QcmcSAd
ggniKOVSe3gGjkLw/a8Y6CZ50mbk+m2+gmaxtdWWoVLspyh3niQMmHtTHrTMC6t67+APitx9JoUD
H+vr9w1XRPoB5ux5jTE0Tk01oNv5fiSv8ydckodChlbmZY32rkzh+VdviK7e4WIoOiegm3ZdudSa
bX8XUFqJ2gpt47OJHd17aehlVstnCxjT9Ffd/HcCq8bhnMYxtr/7cWPmP+7ve3La5ZHhD1JzNk9n
yZm1fQOrKbDRR39jX9JpuGursApyrcJryXBlYg1zu8gePxISq6mgh+IVS0GmJbLZROp9+wLD/VTs
Dq/NhU0j585MByKqdAHXJoe8FiVMQcXTFpi8/5yyuO2jrd8PVKCSSXs8KZM8zRjB5IF1FLOQ3wHq
H+cT/74GHVtnV8bmnbGRm6VO3GV+aSIijULODXPMSnbzNamRIljUs2Ook2yl1hZ8253iWM7wG5pv
STceqZIC/IbJUGK1r2h74igvPUu0pb8PVT0P0TkZ21ujSY1LBNkjZ53Mv3AKKK29IWwRqh15v/jo
9J/EG/Ne2BUPp0F6iU/cT3+Og/sTISitExOEF19tHSwI7Uuxx0yWe6DLDfMEhstpEfSiTO7LLDL2
wsDHj+xqGGvX4Cm2DfLPaAIPLqV383cRYbYvVJPzUmHpcb6/TExGzslhOx4lufgmKHvBRXSiG/a/
baPsk4n8VDDJuw/lvSccuRukuMSVts3c0oqxB6J/mOei+2Bz6mm7F0DyKxxWwYR3cO2H2X/oYskm
QxYpvwA4sxDPbDAExk7h+l03yR5Rka7eaadazOOblZETs0YYB3/YrNjG3y+0qSh3hGAhHuAFX3Rv
7kr8FcXPy6U7Nd117yrSS1pUwLHfaDywDGvZp0bI3JiO4MLoR1K+TfGkTLZiy+RuP2Hpl5ow3Ui0
XOQwVwAigQfuqBhsh7ZQCX6+VRAtlQDnZFa9cSPPhXWUf5tSdZOnadA6rIulWDpT8ZdZTOxzc4fH
lujTrami7ZEjMvEiiTbJnX6qAKvJTXJ5c7NXfAo5IXLmsCkqJew1cMhyONzvmlSWqQV4o+HXW7rM
VkCkHWiadznM7sSqcwTbuw/Lzdpj2Jfs4IymAlyWI05MWJp6ZHV8moRMQY5YX3HuHvyNPQ7jZXlx
/5YHEY3BcfI1inuw4uyoZv7wMbOa7BS+/oeeBBm+PW2uIirmh8BS2nDaSRz9LZlCjPJpdQkzRbVj
iHra6NnQRbduqG2TSVD1wGZD9UgYuuxIEPmqx/ccBB8QtsmFoeiGFQWGvPoDvFyyysDK3v3IwIvR
RAsmuez43ac1WyNVylQ/6xV/hT+LBXnPi8V/mD8+Zq0OUuPL9iKcKxjFz+Knqg6bQX9ARLx2Jy/3
3yU8eton4x/iFnQ1RLd35ToAD+kvISSqUxzvHXTkpqeekzpYJOW3NJlUgt5FpowoHyAbxVQSfuCz
JMmRMfFdA0HdVdtO4Ff76ZyVm+nR7WAAhqfy0ehlIZ2lkZbXw5BW0ro2hTcdvNc/wLMH8/wTQ01G
qpp8y4kV0tr2aQoEzvN6ACZSrh5T8k+VfZujuqq/9VUhuX9fuGyXsmtqAzAoxUypre88kJIaQH52
qWNWJ7T5LMoaqdZPBecIkS3xTjGDdunEPdTAn5vQvd9nWNJmghL/jupwJqMzkXLdNvX+z/Wvc0Pp
JLrvkOyWrP/ALZgSLRfCCmRFWKomzgJ60/t1E5hTGFuVv2PpNX7sfi9hSUGXR+KSiVDYk/+8JQcK
BZQB+9VF+xZWucag9nlqimwgnYnlqWMAzm2akUgFLA8yBf08hgxua+ouyxlKyxI8UiAXI7DKlwrx
shGjnQgdeCjIP38SrCmsnNfbaXIZlRzMWaUxmhtuOX7iiPO9afFJOG0Dei6X1vY5WdnZN7Cx3uE3
fTOOqC0QNtP1UNmOOAsFDNv/R26GoGl3m3HmO7UkIIJfrVr10k6d5cI7Po6aFkHqygzDKjG8hFew
fQ9e7e0a6Y1IbS/Byvj8ssU0VeGcTe8yluPpq5wjfPJqNYZPVFrzeRMKyyAwcxDMz3aVFI7BRoqH
3WAtT8mk6xRt2LccyP3NgRq1iOypNR5bYV7XKKGhXmruwIqCsLEVuFQTO0gaRyTOGNeg3Q5ntDOr
mMHlXFnJzJUn4CdaYyg5rWRlNqr7KjebSuBPTahBM9Vm2NgNcgfowsZemRxR/pNom0V4BJu8A7GR
/pdVktmsn01a1kUHB+2IWPB8TlHo3iXUSKxnre0KX3Edmhev5Da8MmzAtGiyaGw5u3RTa7ltuBYq
tbBOlgwGXb2bG4rCQKfaJhatg8U2GMgIY8fcN7cJYR/0GIRZ2/EStvYuHKGjH/ThNQ1DuPDcj3Fk
aqT5sYgwxOwP8uyJjLTRVaf6DtqmVSEsOPWDgTG4pZGY8+2AieCbYZkHJT81mWamsAzdMm0AK1wh
e1gfM7uYBS2u+5N7oIB3SXwK+ReVAC4qoTO1sgvmP2YaecZrT4C6AL0d0w/CV0O29bW9wRo8cKhw
oOCOZbzo0OtFIEU4Oe65nUNCD7siJuxyQaf5zcBAdXzYKmNZRbjU2u8TLGeBVxm2mVWyalfCepOr
UgMHfGvOKWWAHzMSXJWyTvPCOLC/3mPOGKac82ZJVYVv6B5eXtHuBgzuG75gRCyNcPH3n7nc06XM
pYS49R/HrH7SCnQwAz04kffQyRE3mE1AfjZpq1Wwa/T4FtwR1N4OSQ8GtD9KZAH2KKbedTjsgc+6
Gjta+rP00G1txy5lZDFnxUQNaWTCANl7749o+CSfpDBSsvZfYBeiwH69Eo6xy8OUpco1PNsvo7je
oqp1bFw4I7QdFDMw24BPjO8hPh/Xf8PH1JjJJlMZiIwGqQ7CihRojLKXZOawOVNZlzedU+ye1pjH
jIfVfCSTCobq4tQ7Ojmii7UcX2rl7/PSUtcWGPhTGjjsmzhTfstcX6i2v4iq/t8VwubCE42+IzA6
9GZtKN64/urm7i9VWezn1jRHgiolGuLFNry70L0+1zHvJXdsKpZo6hTKf/T2rPA0Kca1QPXXLWRb
H2itk/K8g8oakPutC0ad6FGy4tchUWe2oEEvvcJ+XI6oV5A2UeQs579j56l1jMNR7kXbralXlG3c
5Wi3hDI4Hrh9bDi9taVPxOcGYsBlCLf8pcP0aOfxP0chuGZ2JLN9vXSvwHQ0JKVYnD8/fyq/BLyd
HY/scHN2P1i/3Bt63Z39yZBAZYtTU0Mz5dxCJ2Ak46BRYuXJbRONY1xmVe5ABY1y8bPgSCgK0VQ7
NQgSDEW/wJKyLmrGG1o/FKB9s/f/jZtyJ1iRzPTUETXbTbM2WoU7SH82a1nXB3BXlMDKOGSYwJf5
qP7gvS0b8pVBK7nZlL7qgwx0YTTA1hhkV17Awc5+4MyGu82E87y4HlLr9fxSuKwdDv3n96EnMmh+
x2hKruZZjcda3IR11REOyHy+iwLMcLvALp3AibXusOo5zv7lNU7RqKUNq+QGh6SRUfRl4FUgoZ4s
VL+rXPEpw1kQxQezLfLc4+Wb7ZGlGZER0wIA3Btqf2Z3mjY2pbvyNaBmY5pda76FB27hxCcgdy9h
o/bmz569OiqJ3EXuexbGYPUuOXG05TRxiXDmulhHy3RIW70YWmorMDBtDPMUFY3IL+Tq0uJZnZPx
TcWa2JxA8a/xe7jozTfpdAV+b/tTIvNy5dfaQWMD35jyaQwiaAsmzm3KYt3Tr5LYGDiegghDMS/6
1v8Huixr2e48q2S3xGYQr3449zFVNkzcJ0rH+jF4fzZyRCSXZp5/X+TKlnV0YzDJYsXxX1fCD+L+
xA8m9P6Uyvc8glPyHRM1bZzP6/TBIVTXNOQGa6Ur9wTQoKCL5HJv4VbzsRtUHinasst6w1xYDZEQ
9K1Ou1TTNsF/vwPM38y6NU4Hznw9uKHYDM5SIsi4YF4f00kUVSe8xwCIDcsQbTe/CMD7+c+ZHiQB
+SR3BjRskV4Xa/Z0SwxurK/tN+EPLQCcxuqDJlYdFSuq8wIKaZ68s5o9mzsKbHJ7kS6aRSF8AOXt
JN41z7XXTRLZmzzcsNdfwwhhleZ7RA0wSmm317Yi6Zm4EJb9FmjsdIRze+QXnpFZFBTcjPrbf4Qb
RGgbfgmEzn48Gb5ZQSR4PSEH1x6CeqB6JpRccBb8SqGffNatyeVVXZyLkizogDiAvvIGEtOC8jEX
wvimURo+xRxUHxgI67+SVhAUME1P3iVLkbtLBaQKLMU+2+FOawNkJ5DXDWm6K5Ya5htW/fxhh0Xu
G9pShT1kKV8f8J/kjWee9JDynoGZRNN+3SlX4Mjge5q7bly3oua3itwTcN4O5d9SEeuwRHMdqd79
SPdpr9oKn1FyrT8Bs+Hs2bhzBHjO8oOOGHrs3aPgC6GTswjCCIc4DfbuWwWHQ92dnQ/gIV7DaF/Z
UdBmtLmLdJlPW9gwH7XWfSITB61byNrIhN9Pob1I17oPGhk60jsxLMJHZtIKDxuadQe8imiqEsTK
THXWrb8cETvHFmI08XjDJqABA2WqDZoNHmKALDPTHBRfbz7fStaYh0FzPl85kfv9gHGzPXh2i2Ls
megMfosDiJxpY1iZMzd6gJIjIyRctXFgE2A2XCoJO1dWRn14YCU5EQNmcQmIMHgXc/YHsY3G8CJd
8560qcldnI/ym3dd2vffraMdsfWPvxV3Ywx2Ns6W6FfgvejFrHZY3pZGPqeQXfm5rL0TwTA3pxxj
HzcmDX5sPb4YYPPIz4kngTqnrIETF8yz8fBr9VFthjpbT5j4U37JDFUoy5NubI+VWuctddu5laT3
cVwiqDcKSAyu37XMeWT/kFBmS9kGZlw33FUBb17T/+u74SjkIcBjB7Hd7/EZ/+/Ldtg3cbduC8we
gasR9n35f6umdePf9x6lOEoYXFLIoU0ERla1Rpa7hXT6oNuHXuFgbPUk79Inv1YQitKD68cPltEN
8f5vhL6xCewB3xo6gq0KFE7M7fWubVaPTSZUQ9zeftz7ARBjZVLbJ3PoAvHPFSP6LZ1YQ12A7jsI
64rl0jvsiOdsCnML3Qt7Pn0tBURxdeH9yNdyJpfEKwPl2nJ753V5HBroEb3kKvX8kaW8AhNFuOq0
pqzaoYLMsdZN3rWhvQ3jydtZ9Ki6RelGn6jRolkag7OV/vMguLyYL3JS377+CPRNbA3YtjrH6NoX
L/deCqKYESIfkuT5MKzZ8/XHFIKtlCka4+gn8kvVoeRcNkopMZbkUnkUYBtXg32uthTD4J3piEJY
vl9YE2kxiqC/S7+CvOBDADBhAH19rtxtliQiCtXQTideJ/5rCoeDFWvKejPUbF4QGIRs2p0ZxA4k
rPMpdXs4hf7GaSf91F/oAhi+vQtClj3wBmT2NAqZSlFg6fiKy5F5sVslcNg2CJX0h60OgENz0UzY
sGruOULj9P2/K+1gS2GE8Dvebk3jS8MtkC4Y/vF/2hX+R+6ZFnXs8zEvaNlu1CtPvEFhFx7gNO+3
fhxoGQpNsI55xXZ5RSp1cYPwPLsV3vZuTWx/FJ28MEsTqwysDr8FX5Jb5bPIkd2RnvcytJouMajp
/wfVOMhaic4muMRiDMwibFnY64h9+TT5CxlUrFdOONIj3GErrzLZrrWUvMk7yZE6y5uLcRm/hZf1
+zteJOpuPAxfKIEQsyJESKKQDme5HtgO/KOY3H+LDlUwydyl7EbKLA5kKaVlfgqUo93Wm6dg7HXK
nNI1J6ydwmXO+yWBLcVYRStVIanXKa7SToSCe4NuYkufMQZMxHAcF3fNDMmNv+Eacl1A250w+8+J
6cKpE7piQnCzcFsKAu+41FftlpLfauGWUQIs+hpRuANwfG5coDA7gUrxYEhHTeO5qT30m14SkwDG
5aosg2+nZxrl2nEwRpNV3o633dHN9Z4KWXvS8A1O8LpbNmUVNrDfm2wZFnfdV6pFRbaxS5MNFz8Q
uKhQEU9USXOssFIO6ryOE3BYGzYT/qcxmBme7rkzuxonGs005Ddp1Ra/M+TBABdWFMNjFaxl5t3X
Hl2XSxeFqbzaOYvyEWBjl/8GSJ2sN87uDaWpZvk/+GzveGeBdXQc+KFNrrLkgyhs9Lbkn5QkItjs
z2LmWW58aVSFha3IOVYoTXSmowrWr+RCTSJEAGMw0xmSrtvaRlL161og7aJGZhh68BDTes0QEECx
Mp+gl3n8YZCUnxLfg8So5wf5dLYrc+sxD+lCpbItKTYfRvrDPyg25aCWph+aVK7NXKEpp7TxFXOq
nskX11nLEUNxxKUT9maNdWyUqUhXRuBSDOdqmWeseE1HxAxmZLlQScaENiTs0o9xykB+h71kxD49
ZQY0ckD++5ffvIcroPqILDwnoZt8qA+Wft49to5UZ5pw45VnAlXbvhYB35dwJ6o4xVDQTy+w0+lS
f8z4ZDSIpb1jp7b9dGkxa207lVYiHS1rRnRvtemLADdTvZ9KG2XdO23jtI7cuMSsj/D6ynYCKPXh
5PqWwRm2hUhtERdhOpX39lxyj8O2gOELMnxpYryBOQp5BEsqMaPTcFjKJJmxNdGOTCMBl9wiCeTr
JY23iRevkA7QDUC9SOTgUc2KjL2koHTpmSFtaBNhe0MFJNihikFUbqhpWVeucBV0Zyv+KuJ7cTme
22HHQ5suNLVpiHOmUDc6WEGYSzNhK1zR9umqyrdzA1cW1YDjDAF830bM7H+Qk9aPYCbeqyuQE9Zp
EwLMPxGHmNEXXCm2An11nmOE/ezQzLj17DqTGrFqOA7etAWVz7M3cdGCbIHa670nAliZa2yBmw8x
H9X+uCUZeDe4V+43iVfB1hKQZyjjhCXkhqAbS1X6ZJuXH0UXp2rTagiJXSoXv0aJQ76pj7SGZ6pk
sl6RP1ce8yL2FrJu+NpOsiSJ1GbENpaIUagCVCiFfh/CEpdy26oH/bWzPYdTD0gl5NE7BlZMxaAR
Y059b2bKE8eeTejtyqePOu9xR0dP8/2pRM8Lo0TZ+mxdDV8qSy07HV/75LMvMBYN1uKF8CTcBVDI
O2a5lfpXRrZvZ6HbQy2NRIgGju2G8IyK5/GVe60UcCtZvgJfn/VTeLXcQXMBKS75kBj3SDilHYHJ
ADdpEdVT3J26meqg1jQLTt71XqAj3x2OAyH1/cJefZDIM5ftLVPDiYwAqJJ5rYZS9KWLmTLYZDPA
XFjRJUj/2nubjT+qqML6gXVukgDXm5/QKw8ZaF/8z1sIGreh1nv2psVyPWe7WxUz//4lor2aVubH
qX6nXT/yS+SbL+tPaDfZ4i0WQGq4N/wqLr5MjzMcjbZYsFrCA97B0hJqg0eZuq04ps1voIuYD+Rm
Tydu5LQI4qEjE9Hd5IGDAn4Lkz5Mz/xAUw+vQdVTa4lfoHtyM1pMeQqz1c4VU4ZP7YkHBlcvSK+f
DJHLLT8SWCJ/gE2cR1K7fa6GbQY131O+brOYjX8Sg+pd1FMYmgFr/iwy0NRdSNy42vn8juEGydjR
nT9DgpN9uwGLxl1n53roP5QpD+B9Hw1DU7gFY5TahkYQEadAOr5FGfDV2BFHS9BP7Yd7Y2Q/4g/H
oPEgmJuj3E5jeG4MRUPdbHYhmboGdpQG9939gjYSzTfh1FF2i+brD/oS19eym3jDGrTvy8TykAsE
13n3X0rPwI0ANUh8ktZ5gItqgzan052BdUKjM9qT+bTCP3JVeYeQNpaIr+g4IDPo/0/YN0ZU59vp
8X6JnKilC8O6mgUV5G6BCAN9Mew80Myobg+UPcGanPqij4J5CSZf8D6ORVcKzlJpSQSbQCYHxl7h
mIZXttY5ylXZCUEJ4to+pI+xZI+7GfX+5gXE1z7YZtxUSRQvzm32SY9SpekDGGUOoOAKyZKivvTk
SB80c9Pt/GrpTnKjSYUy4x2UKwYpOIeC95Q7ZPFQtLDMcVrLf8wre91JVOGBh3OG/jTUm1cvgeyp
C7yPUh0KaMUretbwasVlNjTzfgkcHKlGh6/pP1zxXUuDWu3NwzOmu1xqpVSVSvJGxPlbhd0c03UT
Uien2GQLhNz/NNuOUxcME8c0+94UsKoXXSoXj+VG8C39lSq+dWgWHQVxTkvGzkwBB6phb5SjNguT
G8ba8t7oIJPKTJSO1KEPxQEFZfSFcpXUjo4ziGg70KpkrrTVqmVezugQIazeTJTeIqHngoptynZB
dEmas39IWX+DJ1bpFglJ1bOXBOaRsSgtbHTjeeYeJ12MRJ71oJEpcKV19FM5/VgZlI52RtzvAO8g
d81c9V6orbfYj/W6iloab5gctPgyFRqXvO8Gwyjc7I/9dnhxJNW0WiBSadj4ANym3QUe+YHlqOU/
j/mH6kqJx7WCAxBQ4XQ4QOQrjkgyQb+YwDTUe5o2djHn31Eie/iXlPNBJK21l1/qKYkghuY+XS4A
4QvXyVyixtxMygr7A4w5Bx33V08z2JQHLuJpPy79vGJ/XyJ8p2jTQ+R9k0jtazYUF0YDlFSmYrjH
KutB4nWakxfpz6R+VEFHlW1NbW41Ax1FWVQKlYINvp4BjUCtta0MM2os4m35+628ztm2aQdsURtY
4ppUwt485B5EYlVedXHfbA5xObNCJyU5cmouMbr02S5RZOJySLeJSMmBJWZn2VxdM0D9hBxtx2An
IiLP3GOZORfbfCYSpGpKqtIy+0ZD39ugcze7RUPZkpYeolHo4t6R00pYpVDVL/xEl/KXwxQM21Oo
b3zTiztDC5em2WvoVfyD0LBBYU/FHMLE7/Pl2xP7g/gYGq7BAyt3c6pfx3XjqPlWA7w3k/0M0ktn
9pOs41HgZ9Wj3dGYPlebs/aMSAeUvh2N1YL4jRYjgFFFu9WQ7IKuSBpzcJPmpTq7oOizkevzaTfp
LLm2mzWR/LJABMjA1LlGjuFE94u+tlkcSEHr2udHHgbP2hxLJu6LD21oHxY6YxxAx4Swh+d6hBIP
lrE2lrCua3Fkt5ZVw9Ifu56vznHEdRl45cn3ZLNcD0y896SvRNL6Oaout0YmOTmEYyQt9dEo5nxk
g7SG1K2Kkn79N6MWrB82MgwKq01vubx8A2U3wIZUf4rPWTxfRptzdDlQHXmZ11jl9fpasMdoYbQz
lDz9PrT6rBZU+Kkug9ya+b3+pQkygIFuR5laeERpZpsc8bwfDnT2WgQj024AhbRIJ5GmiI6Rnlve
srQDcZUtN+c1nMg/It8QGzC1/rWaZf5kZST/wI5uKPUHSLl4srhJLJkIKAeLeKol4fZ0xlbkYkx6
OnIlsBOVrZUHsx3no3v1RMiwTHF8PLCB56ld+DOIecqoahxNZ9zwQPa3kjMIJWYqwIVfa0BXIQ7o
ua4MT5ve+zuB/R50pi4aaR775DejNkr7rXiVfTIXmDdo1iVfTVJO49Aw3shN8V7oQu4XwFo01/02
63ySBk83lYPY+w4WR36xji9T5vn1UsPKQjGoKZs9Gl+CNTUhStP62PdxuKR9+r7VaFrIBpfurHMj
0PdJXf++NLZj9jBNku1vgP6rNl+2RLcsSh0Wa0XMKeDYG4zTEX1JD29XHXy14eiis82v1W3ka4Qs
E52+xk3LsjBUw21yg54elAYZdqEoH3YjIOW0o2vMCkwsyfy5m+oMS0vdpEVoImk5v1zr3BCgiijT
GKQac2AZRpwsBJT/F6SnAIXQR8LMRgEXxMJNOGfYukmju3PAfgumYoisFkcTZ8l47IcSWKFI+/dp
PWR2phczjiDShZajE8fWcujKfu2xnpHAbQb1QEBiLAD1gVCbKFB/gsjEpzXnAeVCCEZqrDuKORla
rJ4qORHwalZls5545UwyhRoHkSXbccRgb0EKb9S5yu7wsUpoVLozf+nJlp9oeEVGdfWc7z/Lo17p
/bpkl5E3fEVLl1WrmwsZszoV3uIHg+05XYx2Y/9XwqKhyBIoir+cDMgMQyDnS72+3qkh/onNHM66
XZa+6OGxOnz+HuawjeTMm5JJ8bxIRqPfhDp2WB3HLIGamRwUlP9b2R9lOxKbfu23ievR1s3kLrLY
aNhFI3QPyvvnDjE+Ecwn76akXynMWkGIzDfoIuqSxVn2O3wkPxNXTE22zLRYggZvJyZcwvJzTYAN
QeJ1rFkHU5w7EfPqBL4kDPzuyXryxsVBljX4UxcmE/0Cup3887g0/G09LX2HePTv9qNnrVj+aU27
sv7cea8rBI60r8KX2oj5WodaNoKZsCouTP3cv2Bz2Fb3Wvhc03Qxr6Fq6gVk25zeO5ksonpguAt6
WarmRrSEv7hxWbVIc4LbIm+nQNFl8JnGmgx1sU3ZF9FJrrvYD2dpZa92LYSYzDwHKKANmPhaTlvX
ukGZcRmi36DO1G3syh8J3yPtjeq4bDGBFLGB1Lk9PN9vNNSXzYbGTRKXPcDueHdAuBODCX+NH2ap
s4Kim8MENAqbgacOuTas6eA+q1gswAFRCWMUefyFqLdsp2YUvfJjzAb4z7b5WWM0sVsFHV4tuaf0
nCn/RhHe3X2N6wb+GGV8NGchz8B2XrxAZNDkSb+vOFFuM8+1hThx3UyFjL1li+n+ouNB6R28LLO8
yrhodUG3MYZ1+G50CSVu49Kfq0SBNp1yY4kjXFy6bxlb0ZdqO85iWs6zNqp5smGkO4Klz0k+EvpN
0o3PUyzxOawSWH9UlRMFf8y0immRlpOo6/FNiS9IFSSNJf5FF7uL8yMQ/4GQOkdZDTVU8wwQvElO
S4dhmI60WCdbaUUMp3tkMXbEUrR9eKu8V1ccssXPtFUfP0XiI4p2P2+mH7ODJ//KEOwDax5andiZ
u1OJwRKROw8QVQtAOA9sS8OJwADlyg7uzNb1Fvw72rcn5rNw4RD4YTwMfryG42uPOTqVOai5p3Zo
veI4vlA2nhpWSLLZ6Ji+/Tlt5FimhkHA9TqdFS+qmKj+NFWHHInpuFiwdgq1FHYg7XuEbSTe8yJv
XAZsTOdY+UfpnCQuxgsZ2JiEh6qywEflW+Z9ozFBHoO5/2052b3dqaimKap+rbZFraM3IltpGZsR
xcdoiluUEwBwbgp+z+5BP4tsQ49gVEpMD9NgPA3MJl3Ldq093t6VokvWlhe39o3LrrUfOjmnf0bO
dbdk67dqwCeia9R8ikDDUzbB/1E+/gy4axCDwtugtQgQA8CCXcB33lzy0N9K9FgJg+NqZpb+TN3z
WI6gyDYJFo9YmTA14chKrMJ5I992hp5jpXDYV5fr6t4K7vi1VlTitMTzodgr93MGhZl7FG+Ab51U
4ZVus/WhB2Sa5Y4onYDL5pwI0Gsc4pFILrBRYGOeSsJNGKtBjC+Se9OTAbwuy2aQP8gDhyglzh4q
qK4Q65AoJW260JVeEiO7rV5dmfTDnN//+y/VWUKKaywGV8sia++pQkk4KD8b1lbyvGODKj8sD4mc
PYWeTnFT6g+eT2CfkSWaYdh6pm9go6eTIWFDDKxrUzTaEPweoN7hoGj/DoQd8DQivE5IV92dYefw
pFC3kDoERwhdoPVkj6OOOVrNJMovFE1IM1hv/FUz6UGXrxzx6LfJCouRWmYkSaYB03YedaNkwWxB
XOrI1DgGx9/vESPjgChNEMW1wDuZnmwduB/Kc6WYVPtT7bvu4OYnS1fXo8Zr62ik3y2Dj5WPj0CW
7RRIGQndNDsXvG2p/AItusTaNCiwi+2JePV1+QzNlGzcC9YFGYfY+Rv3fynWPyxvsyjTkGG2X7ZC
VUfYbQkpi7AOAoc8gSsIHpOQNSJZJq/JxZ/PIa6gO0evcNrKkcgV9Vi7pWeYPn2MBW/rT/0hGUlq
CqEdG+XI6ZIoC+txgnxHN33CMPFZ2qa2Z8x0wA2pJgXR2pSZYBhwnDZfYS/AUUtddJe6DUqq/MKE
c6ZusiLe2gElTlvY5DVZEjdqfpd99HeAonr6EPxkpRR51R4AVvTP66qC9heqXlfe2St59nvPuSC1
i2eKrN/eYJJwz5jpwOvbUz07SbQCu+x/A671u+/z9kwM6J2N89AhS/esIDxjhimI1xs7jA+GHKz6
agPiuaLIu6uMnRym2ONtLzAGotD2BPNcvqi89nPuhd2VSwzah1U4o5Wv7XL5SD78qVxWAZwZkPfh
GoigDGxLHnVIYpaMYkIDlVvHDUh6UyWFxwsmIdvGHiRqD/uRpcrWaH7/wwrNn8604smNNGfu2nz3
0Kb+fK8mcSSAok4l03mCf5m2XoPwq+36/3xKoyOimv6z1YelaH9D40PKR213W4x0NPK9504Ryu9u
pn8Pg2AuwCqQhpnT1zU3z286V5D8w3Wt1JFLNA8eks9U33/XtPltiPcjqdMimJ9eNJ3j/Hu7N3Eo
XwcbEsh4cuqpEiM7jEbSC7+F+xR5vpE9Mcf7LbGqQyDkBsWJB1wZWWSHY2Z0JMEkExyJSaBeDxrU
a5tuWilZNJWfC/5Pt7+93cLXcbo/WyvffrH2wmU9rEDD/CyqxHDDWK5Cb03GPy7t5bg847RJ2VjQ
BVoXkdjzdWGC18sExKp7GQaoD80xMaaDiPV7bhQLtTYXOY30JdGjVKi60Rz5nuP1jR66p4tuXqxw
TsR46IUgCzDoMyEPjDkvPozAFh5YFwQva443Cm+dJAdYIsxSIB0ZpuK4QuVcB2W/k++r9lAF24fw
x6NtYOOWZJKRlxpi9BQMQ1ZbXl4vSPHOusZjd6ex/UmhoepO27XoPlQGsCQcVa/p7su9ZoQOZFWc
ZreBZNpN0sDzDFfwgCwxVaLQTIt27ynMOtiN0EAk1eJx17mzo+7N1xKqhShSCWO0sumF9g+u+hKm
9ZXr78Iv89XOplSX9n3WHTrbCjif2HK8ST6x6xMf7GEV8yF2Wq7oQwuI8j9vbcR6VBdxXN6zstZ2
m64XCXhriJD5tiZo/D+L4y6n99oCmMSuxLTFBFnkbsezjzXhQFf5PjbsgNJGN4r/fMw86PGInvWh
YVk+EFtwClrU+dszsNI6m0dDblCp7XCwrHayCYMib7CAIDhddIAiONpBSez0W4oGx+HtXPpLMflw
5jlcHC2+sh9hIcFz+JTlbxDsJ76WCPUHp7yCNThURl9QtRFAcMg3bhQLLjLxY/WiG2/8k7rHNjwG
nK1WuWTb0rgPDSHC/3JyIgEmbH70ZeF2XFDlXuQKkLasJ/Ho143HvtPKJW/cm3LdLJv5l/766Ojh
kkcUHchT2nwFvbsSoTyvPMSMcJzw7pxJq8NLEwTIq6ZUaG1xyWV8NX0yxt44LAwiEOBpYqd2mhld
/e2toFQkT7UAy1ytZouvJB2+QPBif5Q9I00Vjxu6JCUrKhsCw8Qh+cfUzZ7ykD4okxx4pBafOWEG
AlDie91k2t2cdKyCyKVCFClGnoKeynQca0gFGnUtD2Jj+Me85K1RlnMfQwX64IoWbu0FLSJ0Vp5W
G259yXeOQPRm7wvQqFyoxsrUyHfvpKJ+ZSzJNkpWCVwiRAz3LSBRLVws79BP6xPEyF0Wh5hwIqso
etJUulbSRteSZiqjOiZnBXpcNLClWUrcmBMkIWDTFZDxMyC8DkHJEO7f6d3Ei4I+Y91rCMM/phTA
owb7qmn/Gi5rr2m0HN/O0fr8jJXBnep1/dGpIODDpGFXjLM83TduL7DGTUhR0+OopJLkh/J45QNE
XGzq3JbqKAI9D52TnjlC6NZi9Hk4hL8UiTUhgmAxx0fhusnJ5gINNhlm7Io99VMCzmT12cj5/BKR
QmYthEWOfw9jkE+1CTAv6S+aCNt9Hccbq2FKbhMtuO4afqUiOBLRst0Cfmw7qgQMhLEDLTJpR6M/
M2aKb3cywm5CqwiRFOLjKEK/0nzpfFOU9U0gbvxKL7GWKS5evkqtNJY3HlNBsUPj477KMIRdh/lG
CV7gdpT4Vp7bLS31KEtMPLLyBbmkQjAN5Y0bQEPJivCARprPSm54fdQY4l76f6Fm6WY2CDKgFoFR
u83naK+ijZBtZRZmRnMpD1Vcm29qf2jJq9CHgw6GfUHvkSkCaw0m8mA1uk9Of8JDFcFRxoIQHyTl
4DGo9JrBtqd3bpi/GSRbuDomln2ecrGkUfXhrDzOoLSfi+yLdbc+vMb4PCDkhXOx2FZSvMgh/x2z
Dr0nssx1NPvyZEXkkf3+X50ZEzoyq2mVMfHWHR4JVilPdru1UpDPKEM2RUrgKYCGwTGWig4HRKPv
FdxzBHiwMMDcNHR1m58ob6vLArDLunuFhX1Q9LPqmlkW+XMJ8kQpR0gXJKEuZ6bAzziOYQTf9vVn
KPJY96zUNaNJxZ79NQiT9igNYksEfZ1dNr1kdE7u/V7XVr2a76D8v7d12K1KHk+6XtRBC7mE77Pk
6j2otuupQgyHybfBM8y4dwdwmktQ1QpyqFid9r5SZTgIdShITqxHfB6Yu3CxMrFnHoTNKoQLVvf1
aePoLjYaCoyORD9o2+p5kmVqn0prbM+9DGkMrRfabH08yWt/YVApq3FLHL7dP4dt9MHMnaCMCUuG
gsFyTTfd7GncYtym0Am5aTs4UeJo9lmWJGCjhOD24UoiMG4EMkov49hBDzE897d9PCHVnA5zsxR1
3ou02YUQShv2yAeKdVSSijAZ8fznTdqwdr/lKh0h5DjeXgowH+8bZUXPmk5fdsdsbvcWfDzl4QWf
dHWhprGPo/eMCb4kzCPUVynKOfDeaEeWESzVxbhTiRbs+Gpxn2VxnF+cEctnbHRd5TImftUF2KeI
1E/0FcTJuffszFTRRruDOAQMTa5pnuQjq+3uTwC0mCDgsvboeC6mZFfjtsfEXuOur0tbSlOIsuci
HuBzQZPntJkfN46xHA+1j7fsOLSDIisjytUPavxpcFi6R1zVJNvUO7Hr9IQ008yRvLwotyWEygxX
NpdQfvXqHsozq+1/EDvsWsSZ9Y5Xm7Mknlkyvo5qIJ0RMNCLBaCXcoKT7wP39jVyRSr1UWGzZXy1
/SpSn56fK5Q1cDJIoDKOX+Xh/C1Aga6FnD2VLegK/CcERGFjR9C4OmLb/7Vf+agiESJVHC9cEWyg
xL7H+TVzcmaz0gdakL//LTNqB68kqTcOnAlzS7ZFKmHB4ykw72qDomEPSB2EiOrzhk5yBR/Kaj73
VSoaPnYqgO5zSyj4mc5sshP0UrxRru3L8Q7++YjzGM0SbxPSgoNCFclMUwXPq0pUvAFpcLOWUI4O
rmlvu/LGUxl+lijzQD0JGBuM47fsndZISfmF2/3ZOFpwIAfR63y+coGoq5scta+mmPxRD27Pyc+G
79EbNw+PD//i5mJ8V2WZRlqj4/RgCiAgJFV3kWYsmhdy53XmKNTIIFr2s/heYPfEZMOx2tQKM8OF
PJv8/xynOhtAdgqywgdOaSixs+pelN/KcbO9AlZ5f5fL0abKlq20rd5NgBTpF3LQN6GtoZ8WIcxQ
MAfI7holxsDzBeDO2R6t6BSG9Z96J2iRStKacavk1y/X8d5rjYSqVgwPP11wNuNlEhtCyJ2ZGQbD
sRY9sRb5m6xHjLP4NQ+FlgR+AP/wGoYMw7LZ2nxpyQPGBkCLNYYyizlL/sTjdrUl/oF/retXk6PW
iVWYrioQPEAhu98qGvXvMsM/wNtCTtc3HotfHlIW6MzZYfjh5hrNwiLCOhJf1uGGEvojXHXeVZck
10qq9sqyVjv8uhmdKGqF8ki5tSqONFHNZa6roWUD3zBZPW8eQ/bD05ex3Oj3xcV4PvWE3x+g72yB
/XkeXRITd3lk+Qxkk0laSamOiGam08enekAA3YADkbdMqulZFS61ngImsXI+lQKJ9mF5xl2c/4lS
FRrTm5ZdlfYodGH7tuR/2K6pEHMKAFm8C9a371SYia2fpUnRJjK7WUdxRjc6W/PHbropdalVactA
pkXKTQPrmDbPSguVTGGATu+lQlFZXWu2DKe4V4wz+g3i3X8dDxYJPyM93bNPmP+SP5oqdnaQ500L
G64sg90Vz7/cPyJ7r/3RLFl2s+3RnfwpBDTE1ABxVysMoPKFucK05wFALZDME29fqko/vnDaZpJA
mVGjtiCvKLr+uZK1WTbVZyt4aQqpHsZdG4xDdaMTv5U5RC4eNRNuZgESkG3xexRB44hdVGRrf6WL
mLBjtMTN66+93MjUXYL7D+IKIz+5cF+xSbbChVQNeb8Q/egkj+HMUHJLCcQzYNtbhLOGXfM/Pdr7
/PbQI5lUwcOv0PEtWn2XWoIsfT7SX+/Q9OM8PxF6pA3M8fc7ZNIq3PAUSp+1Q6G1XVvH8aCiitp6
OpND2SnB8APyDP7ArXnDXZ7z6d8l6MGkxRUioNGqosz0wiGhiQqvV59ZPfA5GOqfEm3kghoexkK+
iyLdU64im0XW8uwzwMHvZvo6Db+z8Sg1gQ6Wl3qMi+dffLsvg3aQlawq9avv1sfsJ+xMe1dAJL8b
n1cQQQbhToLVZKKOScqLJYfmceeMPE0WzxotcnW0j9WZ+yV7MiDYAJVyRVjygL1nJI+U4VCEpVPk
pI1k9AxHcbdpClMMV8ABwk6PoDEo6MTyfewFRhSiofj1MnNRwN52idOK/hTS/FvzQuFMUuud9a0t
l9fwCZirOHjNsLttpnl6OeTPGUO9XydYJsojngKsvN3Zh46I6Di/VV8bsYT1d9RGLUMpyETqDtq6
/Vw2gL82dLixW1TCnrmdrzwMwBwuR2SCA23R/LfC9yRlFgZxb+cL4L9LQvUrvVORC75M8tnPGvzE
6SFW6ct8yE4Yl/hPJS/D0EsxprN9wvpz8ow4c0vYs6B83PIiAhQYFwCwOePL75kQC9uZmpCYY+7Y
MLE4NcI9oxj/kWlg532/M9tOiQyvEVSKAMfMTySISiwcHL3x5vqz2/Fe3SM4nxU0f3VpNXvpMFJ/
7L+gBXLx0bqD+m12mHO2MK7psPMYX/QkbMuuiCKRTqHvrvLOSYlcGWmG8gROMqjbbC4jIbF7dQhP
LUtMFT7fw+d3yRVosTToaPcfATPnHWfvFpev40zvVRTWMTwlJEuxcckgRTGA0eQjpgmhF+snowAj
aolL4F0m4APEsiISWCiJ4CXh0U8pwuOXBDkXvKFiMsB1fQDGScCJ7Yqy7wj+RjKccOMLRMjCXkn+
Kw5xsXn75TDacuTA5N4gt461gd1VWFLPeOgWfvtPjC8h7xlxvRrFg6X37cHFF+1NQigGzy6isVrG
/ixoev8/RR6vWLy9ZQ6pLLvK56MQy0fLKBBxIgzZhlYGM8mB+Xq4F9dfkm2IL7hAjlm7LKcTZN33
NuC7Ka3z1KuRfwHks5L6mBo4oVE+5RT5hPqlv/q4pGmDlV3eHf0z+Qxp6ZB7OkA7WFyxX65F3wh5
L4QsxjSV99COd25PWih0Dq1WXcXn4vEp0NDsyzd/f94ohzqVRHOdnByHA0OxQAZdu8KdsAtdvn3Q
iXQhxM754Te7tbdRXTSXerbw/xsFj7mPgyXSvF5B12A+JJFSgNoDiVdTLV6+itZ8/GUJCaFrKvhv
9Z6KTWZk8pN5ASFshSiMCqFA6NQNwuS90DdkeQh8k7NfHxqO9Zr9Dfld/wtpCuCL4UnuZIOTkMVu
NDQ1hXnziwM9BbW6StA3R1pZGD0X/uCvuTMzSN2yvldqvHDHsIMfU2GiiHOVrmYTFLRngZEXl4JI
PALAol/xqqfiJV7UcS3pLIhqS47G4qZftPruECbHKDhNgWZ1bd8q2dxoVGYTXCcvyV0TOGde3Ywq
8u/5TmvZC3Q2PjjiuICxWDwi26DMqIUY+aPsyV/cAmeNI3Dyf2eNPev5il4PPnuKIkyjcP8lWObe
IDmyqEmndXJamfsoOVvxK89jeWW+OfJlpBqzg+Hz9rzDOBTvMqDJJTdw2NUT7SKuz6M6n9MDuBOZ
8yDFlF9rBVl5UaJcoRe4AqM6dWPT9qhbP93kWVqE5vwYi3eAzuPcI8y9RuhHXDGwyrBX2ctLCjYi
Kc5t5yDwQX7LHqZNnD2GfO9rV7cxBoS3dfI5biAcVZ/17ZX4DMBVVIMD4qROaPKV8jI6PyB++3vb
D98UZKORRc9ZEA+ejYs9PSN7fsYGp5TdkpiOn0XrKH0yIHWCleIWClwtVzT+DKFYddeAYJamt6ja
IfkOGAYAPpfB/AUxmO8UAv+gfCXU1t9AKzvh4FLEP84iGNdV69va6w5jSr8ICL59VCq55ull3MXO
FdKR6JoBCWran7xaks7ACmRyLL9xd1V6g8Q1na8jj9j5InOi6BQRy55z6SzZmfW93K7aJLDb1NkS
g73RdjFVZhqxrStaz90s+cUftr1CEaC70FXe50fuFoJnJRF1uRk7VWH1PJJXiA8g0yDDZB7Gwci+
nY4nc+wX8EQEdgDtTvHZo6rqllqWLM4u375K3oLvrckX1WISXeS6/2EKEFt4WZAt+XZGQSQoGepx
hiETmKqMcwv3BF1B3rgz5kfnLAD267R1jDF/FY2ivQ/9mWLYw53A8u5PzmjH/tVjKvpJkBSlCjD4
m1sFU0HmfYSBcg22cWD2AxJMuSxxG1xmuixuv7hppbBhxgU7oJ1tWsUiMpr1ONCcXU21g8ZSczEU
t2zAHtHNhjlDjAC6wwZDHHA4ZA1X1VCeyUfcBqJ2Mdl/5ETIL6+b848w7I0lXYEKM2X/fGb7hCFM
FCMICzpgLa/HcJknBq8BzYqKAbwCo/5xXTCggJqLMQ3K84g3B1NnxkVdLNIQ/BdK14WwcvSE2fXr
wgF5t6j8iq2zdO6ERJnxYfTHnQSK8z/0Uy+SO5mht7hIMDs7+7HCOQPYTocTHplFcU/x2cosXgqW
eWH1DdJCB58WHFj+/GjLhaKz6sybMMyb4MoTtgUq0GRh4p1RTVpNxedfy3cC+ei8JS7GL7dtL5WN
c5zv66syVVwYhIvKF7yAQb9CjS8dT1xdMpICqBzCOr0++zA6u6vpK4tG6Jw/b7AShZJboMIBnHhW
HwjEHlUcLdfzncCWTvJJaDWzxTaYyqyO6In7ZRHO4CWLsOWulwCIdcacYHCm/zFs7wT7qGJuymGB
1t7TWH/pA8TAFRYhgQNvhotHDDU20TLvVVPxCVWYxjiVpQx3j3AWrvarlfrA6Uw5sHp13Q60mt/7
8E4FbuDxbBJYPnvbzIhxsmG79Q+UeoFANwEYQTlBAwD5fwn+g6Uqxxsk47BHTAGwfBfLiggwtYjM
XcfrTZxyHqlNK4Ulp/WWvzoekxGcmXWJd9wU3XqE3BijjoyHFpXrtEP7L1vZq6q/2KEZgBtjZq59
BBlRzxGqppU+sxKc1BQh6VAH2fRHPbTnt3A9OyxlXur5K4Khzy31SYa2Fcev+jiO/tspe/UNPhdm
JDTOKPpic4WGRAfAwzJ0c4rzI6328vwDLVMA22BPVlqTRAOcBXEq4AofIy7m+SLcQBYMF0G+ExFK
XiWjT/QK3ZdTNvgxYL3mtGwn0a1t3CFdYW/GJGKMWCfM9eV5GNEZmxOJBluVOhmF+nf8Vz8MAijc
gbPi6TwDpshksULy2EQxp+oelFrB34EIwtqF0qTLJyr64/dak8B1i0NW2UJVeB9yY7L2IfJa/RNA
cJJLYix/TxVVshkNiQ5mg/ClNLbH43i7TCG38nwj3aGXJrJ0lNKiZUdyycvaWcHDKH8kIg9xuKsQ
f5gUyySnelrwthZL7B/X4iDi1RameP0VtOIoVwdf4+Rec0lELyz2MbOAUBjEE49L6Zd8OSqH/2Fl
nZq07IAQhUhlT5+LO3Ui6s1tvc7auSEcMNTXvdjTippr0Y1XDO2V32Hhz21qLx9btdrrdpji6mDl
WfaAgj65/Vpcyrz2gyuNY1GMLpP2JsKg8tqNMvC/uEU36AfBpgpkJt3lTcVg/daP9BtMTqhcNCaf
mumzCgx5c9H4NhI+oeprpqBvrIviiZ8wAtUe6VeiYYB/ioVRqVZUKhX/wcW6FGkjkf+yA86BU7M9
4wFAFVoZiQ9fwNEPXELy2wzsxw8QXyL81IByu0YPO4F77Mw44nr73jZhg9RoDqwId6Bpn1sbc6k/
VoIaDthdPTOSFXzfKro+whj1mPJ4gKAFemUVSpYuR/PmjzGOlkFm2OmWoAINpJ5iov+SqX+D/JvS
twEU2/I1i25kg+7HdEg1g9COaD7PmJJ9jsU+l8URiiAyAlo+JeN1EyORLKg6gfDsh4gTgKfkYCSp
ywzvLUpKQlDIlYVXYhDHrRLYnotW5xzilb+mIo9sylazB9OrBM+KHWX20ApUKvQPpkY0wfUCS6lH
TRPvcIZbJdJJ5xwpZqycoOI3yhIRjC4hVeVE4QBqVKvTsUiAXC39HYDTlm+LtkQYtO+dWaUx5DOc
6lmCVbf0MvO+OJ4Eb/LTxy7DpXvhtZG5AKwCHAUhRfwyblOmFcNi152rATu7G/569Yijs8ZE0VBM
nEO5/t3WhWX1U/WTLKK45HCP7PMvJEk6Ofvt438wUtKDgbQQ16D5J/8F6DUE/jJf+5aQZ/63jxsy
eAmkTGgeXAfa+8JmpcDxxR7MRmh0mEXDX0TkuwOC4j5MTW0Hbe5LEPODhxRbbvBkFmO0TFXWhaB7
tHmoBbiiuf2N0uXF0VmQKAtMrTjrbJrNJ6sMDoJdw1ZWYtiqPguug6Yx23LEEp9JeUwt0eHZAzDU
MjiUF4iHhaaCF+pXfG5Z9RP1AxK25/mcNn1b0se/t3/kIu8gaa1XD31Kb+QlH97WxZR6ZKTZo1CZ
n63SNe2+COy7iA4nMx3av1mtO93aczeraAVj4reqP8fRjfLjNBcUk7OkVZqTe2HvujoyaAgVBCc5
fH5+paT5F8pgHBybxnLDrRu7APd90HtLWIVZVFaFNfx4Ld0Je7Z0tYT52gE2SV96eWFz/ARm8Bkp
kTwP3Wtlu8V2tYSRZxwX1oIaSLMm0GmaMoKfZX2mbWypjEcX5otpmCKBw3rb+ocFruUs9URbynvX
0XCXvy3w31XBvRYQtdRZWulVn4WBsG+twRUW1/oX/2T301ptAo/0J+MYLpzPmOs2q58q7BvToZsP
tRg5SP/stkImcKd7uJ9aDzV0lRRim6Ho2AH+8wubWC0mPXs4DuDpDss+F8DfhBhlMKmlC70XQu08
4Pe2TtdSeB5K8MgVsxtw5Nq18qlgkdKfVDWmNncb8EGH4HMf7XVP36IJkrH/9JyZoeeGXo1DNBI2
CpBLlJCX6W/MYe0wQbpgU5cvjjBxKoAGcDg091/TgSfoGit3/rNwXG59jPcTj7ePU1QYQsAb+Z4F
hc+HomO6VCWu/vp5d7F71ovvfD60llIlROD7kO7bvG7yKjtnrgMW1oUj2O1Ig1GEhtrT0FRFqcXY
48cbdDY6i9/bbSeP+TSMYPv/YMBkzkID9RMYFrsntruvwdcXHbEZDiFCpAnfaunBP+Z7LefWlAXz
yxQ2cQPMmbTlgaOzFPsaPJwEzIo7br/P9RktgfQip3tOz4Pc8cWAzrBOf11myWyYe4PlqNlnnTxc
SHZf/c9NNGtSNsNrjzbq57nFkPJrts9/u+brNX6cpE8zv9hpoFvR6nMPJWLIH1slnn+vWhii8vcv
gK+JDWliG6PQNskA/cFRYJW8yvPo05d5mvkqpLSoIr+pUtTyQdFLNNHou5sDguYDAUAll9Gzjfen
bd0xxx5zotwUFuE75sN+KjI/pexLecZhsq5TW4Qdg48JaAeyy1L2m8uMEBB1zq2jTSXVf4BSUOYY
iUjn2FrX4XzPDzNhGoLu49nG8JXu08O6LgGlB4Rd9I51DTs1UXcjna2VuF6nckT0CpkQd93I40r4
qRSyF/WQ0pN2RSJSqYXeZi6eaIgO4t2trqR4VXP3GVeKpPp3iU5JYiGejyZFftJNWUANrG+kODrE
+ARhBdt5FnbrhM0rAUCnuFdsVLvR21E0o595vOLfeiy8H5wFqvba/7dPx949qoL8rJQNUC5jRZGT
rY7yYiz0ZZzd9RhidyxdrHX8bdehjDDsw8Bq/CSxzHaMhv+XJSOW2naFJAvGz9S0IIQCJR/+m9qY
dW0l7B+CVXJiYGyz8nzHDnjI6X2J1uDDZBzqqTQhmEPzVHbg2m61w4ppXxSbohtMY3CfK7oWodY6
AQ1IoV56p6CNzTOF4rL5FIPeIaMNKGvYRYKnGZQFNl99XI9jnOYi4Y9JrQ3CDPD5GzBaOCVGsc72
lRfxb16Mc97Z56hEd+Tc286wayY5Jc61YMf9nf+b0av/MR3JfTX7tsAM1q8RNPkgP7j+vff5EbdS
6buyiqarLupHc94rpbnYWeQm98VuN/2PI4gXm879YxyWtJdmUkTJ+syrLIhE/VjWvMXEi1JNy0p6
YklKEbaSoyfEMJD1dr6Ullob8665dSmmspoXR9EhsjQbpwqumta89Sa2eXWKr5z+MeFer+1Ri9rp
YVIrKLZhTEQEt2Q3xtKm7Ktv8blsPNWfUiV3o5uijUK8YaeSWTr2TbYmWbFgpAYsCzRKdowDHcHx
dzgTJOX78iq9Hk+yR7X1tKn/dXH87RnJptAwQc8yu6YLabGXd4evgQVOpQfOgCMCArbpyaXMfI56
Nz7FLKSF9wO1cV1RKgMwU7VsWx2W+F0UMPgceTi/adTkouTYPORUgEbXEzXdh9woLeeAW4Qjx3z0
33VYqCbC0eeWabMyepWGBuJKgNK0WgLCZEQftGGCfPU7FVaNHerdzVWEbyXM4AgH9RL6ZQnmJosE
cEY/j2kwfcMnzhJCZEM+YNcjdVN47uLES9XAjRfe+OMb+n6X5OBL++jNm9XFYB2vsr8+JVNg9E/l
rn5bfooeAkuD+XzvB08zZkSQ8rH4ykLeL20ACZot2wA1h5QBGhfO0ER1BQeEFYMH9vgl5K+0wH00
zeRzoGdT0WtvvldV3+4F69MNt2OWXr4EVeLumWJ1Bk6dH/4FjDXzvd5KjGz+p2Y21wcN5QlrUEQA
KCz7ivlk/WAr+xhgXPMaTcs1BgzUrLwVd6cUNJ+SJC4Bx2+MHdmuBMrvL+Yx9LLpcu0baDKklL6x
wFi9RQQ+Ik5AYeixq361vDdB35nCQ/23InqyXukjWcGgPhSVBHIyFt/PxMABjarCfs4USxiXcF9R
GORAQ460VAb200KRND7+u94oj4JnoCjEkBCaA1yGMo3XRCzGLALL7OLHurMv4qLMEG3B0wbZK5+D
jn5aB7sSPn43lWwlyZRKNKyOQUm2Q3fM1FCrTFGq0etuwNVkGfgM5Hu9oZz2jMmG0rAv7csQZS25
9uMgGfbuYJqGyo9xLb2033+hvovGiJ5449TtCboMlszPBHq+to9b+qhgcZj3nvM9JwDdfEA47Ev8
PpBPrT9IoM86udjnIpjAcYiNn/o6vArWS3KAJ7F3q7bBrPdgP+PxEUQIQFf5mdl74khVIffcTAw2
2GhAaov4+Z7/LVlo0/NVJCBSTBBTdyFmK5tCuWjzk5ntmdGhXkrufoUPmeusMbGWZKsgQDT/COOk
UOePw6FYa6Dzx9qscxHpl0BDs7izXbM7wY7ElZIoiDVwlP0tawMoKEpE7jBOlaE26U0Lxo08fmEc
iLkzx8YivX+FkvZRhpNPWj96Hmd2MR7ebQJJugvKO8zMYDjVBntfoT5NBs+kSl3V8wC7qzGXrn3O
e8d5/zx9cuJewFtHUTNEzMrZOepEQWuiwibFzQS2TFYICggvLA+tg4um7ZiCDz/3iOkX434vPLZ4
2znPq+iXCZLR//sfwBPiMVRNPU7PwqwSp35S5jNTOZ0LyXM8D4bq2+0hCejh7x9x0ftHr0x7UsJI
4lgt2N2Igtz9tHEicsp3Pwqf9nnrs/B+WHdGTv9Ua/g4CUXuhJ7P5gJ1terf4xdcjGI+uU4vOtJZ
FAkZ5oAPwdlqgMwZ3MNMKCPZMrorxqp0nO96LZSYYfYBgzfUDs1o0nemT63+KDL7xtbIrcXMvb5W
zHF4WUxy2znaQluIIBMlMyHqSf6cGmKKB2MQmmMCHzp6wCscCXTaYlGWpVtrp1j6NEUJ6I0Gn8D2
ImzL9T4L/ePpm7AMhADayVgJSHXIOEn8lrCQnLBPM5Y0qA/IdrJb5QqRcBDK5ucFeSccwb3GBXxg
PE8Z/ie+LJBuG74pzUb9Ee/+KDfMIDuTQ6VQRLWQHtXwDN+f+7eyAknAmHVwpuk6sG+wyuLjQRU6
LU8O/xkHhvV0AT5dK2877ymDeemZgriWEu2Yunr/1Sw46upUywaF+iEpSuI0C2+xs77OQFIqv5A9
lz9qWaCk2b8NR5uMzdJ0ghuyQCZNHjALz3fXQT+534kUhbij+UMnVetd6RQekqrVLk3oHhtu5ngd
RT+e3HEAG+p4RIddpjM1lCZFAA4dYPC/P2C3jOnLHLPwR7gF7Vs/3MqZ+SEXuKdk5Uhx27GHDOBa
F+t5ARsZWM+9kPkLmeYOqLg7LpWLYEa7MNxsIBOjpTCpfI7fay3axOgtlKgqsUq4izDzorWRfd0B
c3wtZjjUphyBaPRyKqdmBbtDXZs807u1ctgq/DgacwE+bYmWAOgPPRQVRvp+yvLytMDsJWIjRMbV
qUoMjQM6H9eL4wtiBqZ5fOKJhuZuUNZT2ZyGeCo0/oxw4jPB7S+P9mUeKSgOsV/Z9T/TbEVlfImN
PjkWylBkOF8Fq/9pOpoHd8mr+pHIVNY5CLjmorBEK5bKr+GMu+SVC0tgJHyfX6aXFklJwtKrljy2
yTGTQJSIvNrIyeZaZs82zFOXfW0EH7CtAc17jnIKHMTZwRNHaOjpUr4QV1RaO3Bo6OkKBgC7My1B
jfWSmSkHNZ68o1/X1XgMiD2WogiwQsHY2TixHVR7l1b8IoDyImB5Iw/WSn7Sd6cL/LMoz0z63tV7
EH5kxaE3ifYdQ44zurzxdTXKJnYHxAKXGpZpaTO+2p888FsMFtUbV3UfwT6CjW/6Q+NY849ipEwa
TpitnRcWiAoJFDcBZATYZLt3x59Ao/g4yrt9g+VsJrOL34o9ZI6YtSgWRCVLqAUe8vnRGk/Cf7po
cpH1aAXNo/3rV/Ya93z+pF8BwO47r0SNqZffDbJ2uvuWFWvyKQqv249Yl30gVvXgCy0e7DUOku7v
GLOovNS34c8L/DMQ8QGABUUWQx1z47GwYikos12AUciqHUebsfuCyL/FWXi433ObpKiadjLg5sdT
KyjXkDT+8/JUkRV9t/JOVDedmh2WZjEv5YJhBufvZDO+HG/h4v99ZLNOZ9qf0WLICdKoXLyl17N1
3efLGYkEP7NPCqJ915ZheKDRKyLhg7Sb8pez0uvmWb7nEIOgNagYaQ9wPMRH1Mtn4kCa13d/BP+z
xoKnB4v2+FhVDuHREl0jTDT7OX6u58bNcnsob+uTOXIwSeJLlNAGKr4T+ECJlu+I87+8qu+y3WNi
+19s3DFM6Kxs0poa2DnOMs3gFgfMBq8xxtcm5mh988+WmBSbWAIQz4DxNIqNcay9qV3+cxl2/9DN
edZdlVBkOUzBMFkNtvP15BR56wMJ+8maNno/xfPb9eHo/yfdoRJX/vKyotnCc2MeCoYSHl8cIGjk
dXDYIg5Nd2/FdKXAjopkYfjVl2+XBDVMbbjOw8airTqBcKvXxxKhaC1QQAhh/VFL3ZUFU/PxqyYT
97i7PFfltBupYnKqHjNTbk/MkwnaIGMSnK3rv+GXgdQg4fEVvykfjB7ULUwzF6Lr88TolcjoUOFw
2biN//0OeVy2FOz1Id0qLSF21z63FZwXg7LHTHhjMsoyFzlkHtU6cQ1yTCr25gofWtdQDyp0Zytd
svv/V4l7V5uchUo5YDVUl0KZPY5afpPTazS5oNSsOQ88iuHPD8C6XlXul3EtLnZBRJZVW1gEREzy
22hUMIcWysjkDqp3z66rjKGZl1WlCuydfOGFY8b1Jo3icjO7kzD+gxZjqyLie2tAoLUZPXeEyVoO
FV95RtefgWNQm8x3ePzC4zE3nStDjWcpVoyG5TAhArajAv6AtL3FSu5rvAoYIVKU+ZTLrO3YKCts
GSI/2hmZUKsUwb8WpGODFnpTnH2/lLJwiYXrv86+LcBrVYJoFvzHo3o3Fj01G17px/FSy4R171vg
zi3sCc0Xyxmq0n7EyRqh0BveY0SuED6wDWns3nbBFUTNgGPSYLNPbgeiPTMSYK/kIv5o+1D+Vpwk
ezTGYkBm6r3X05PmHs4CSBKjLCW2XJVgR6n5PWSI7938bDz/buv1SCvp7zOrTKBRp1hPGoe/LT31
kKyjCFYSpUsAofyCSgM4MrvHhECACoGYyQSSy1KRX+rHN4uRhtnvh7T6HyAw6ixJFEB1FxMaQtDn
MFo9KZGlG37xKaTm1Fldydd67fn4CWza7d6yPRFoDciXGcfZzrEM7rEvT1cxkhuopTRdzw1ewyfk
JmFwm0gl3HpsYeP52dYcmLJoah9USOk1YHIgE9zZG2HtsCV+fJoTxxzmvRDoZM5m2oFBIyrqpVil
SgnT6mQPMNfWK+8jY5coxYK9eLjv2RHw3KnQPELwX7KrRfM5jK/+HWxuIB3QfTZ3TxL5Xyo1rabv
jW5kbgJ9UnSLhfsmBnVRcrbr++jmBmQM/jgTdC+PmRQ7NOMS/myCSI5Pz0fgujZ7ZHsX0cOuYgQR
Yg44eQXD48Xa2m3iwwcVpbzVUDdWLYoQdKsV8uQvZVSx4HAY1obTR9/agDXD3bBbaO1Yvaa2LniM
z4R25ATlYQkSZ8YqYNGy5aN3Vs+DkGZVkoH9ckI4JkYqzeXF/zQqzOOisnvGqpUvQ2+Gq2MhanFP
v3L/YOCzWQWJEBBUlg6DsUTCrgAuk/Mroyegm2FjUXtICqfRhXwNi4A0xKfBmZ7YvTQQbt/qc1rE
lnV/erT4PAJ7bdpjmOyOwfQm4nhrj4eYNC5eFRrYFWfz185eUiqGWbPRifSJZ4uT7EvnS06Z6cav
7ZyipQg3kMLWaVzP8Kuzux+/i6ceuBuhLy1fGh4YobMrj+jg32LxsYrqDWS4P8KWl+q9SDvqFRsE
KCPhlVVsw3rZGzjY4ck3bW4faB3jWIzwYgJBbw/YXKc2cP6tbNXC0o7/s4j0ICGR3FaANQrUtdMl
1xXKwAnWVTOQxVatp8FI/FvfPmfTnye7clvhCsK0DGxCDdqzli9WzlFFbEJO61s5HbG3Zusav9sB
9gRAsjnjhPRrQMvZmp6QBV9TMpVFxYNdlvQzy9M9YeXV35bpeMXfsZv+el3XQ6gzo79WnyVQzOE3
AxJFr7dBqL8EKAkfjhBv3/3F7zHLPQNyUJfpIi5DhlOHtM2j4xD/q1SWKJMEy3YPMUu46L0CQf7S
lWjub7SnWhSXyzfiqOYmv7vi0bXXiZXxtEz+ufOshlHFxsbiqqqE3kcmCp7HQIhfpmlCQKZwoj+a
MmcNxyeR0YtXFwqxnKNCu0YcN2mySId6937H8nl69V3T9aNT/P7uvnT7w0PVCfYPZRztvKTHTJDs
FwvD9vjf+u0iK8PADeaSvdp1FKPEsjvnLPUNY222McEigl+q3GWS4Mi+hpD0dd62QpItjnUS9zvp
i9hN0r12UrQBYYu2KOAJR5xnZIYpYT7NzxlUVU3hwv+rxtKKORIk65d1ewzvPDYIi5jESWF9QSb9
3gUXKJSrMmtMILl1Wqp71DUDg/19lrh/eu+1Y6lmNJT8aSkSesZfTZq5pSeINK0QwVGZeSWZdKsl
RNY6j0esUikpYk0b+4qvaj2MbD0CVsaR/clwZQ4rQmYWlJ/yGH4DaulAMEvI6h+bf2FIcs886lao
hkt8olE5f0BAYbzoUZWjNfRerEkwaenTywM2+905qd1BUP4IqCVh0hJ51s7FEocSHpMXBlVKR4PG
Wen4QnVKUMBk7AQSIZrXzH9zmQBdwZrHUIhtQEYXVak7/38nursardHyNRVYIveFxzknqxk6nCB1
YNjny7SaEQcJldJh1YAw9prnmvSLj0y4ChqkxGqIB3i8+hOBnza7QNqSf0nBTzviX85xJ5Ntte4K
UyLQLc8ZlTeY4TGdhuyQnbAbQHTyC44yCeznb2SpsXYQBXyIaalV1GZvbmUmgWAeRpv+kB0C2OmF
Sq4ZcNsH/yzJ64oLqtIY1IzPJX/iZvqO/2NxrCEv6qqMkJRiOYEcfmL5NUKuRWhbHr4G6JfgYwLs
6xvZsXSu0fSYinK6aLoEjmyWpSxfZnaHalLaqI/muScTzLaoe5JBYf0FEli73bf2RcZLUdXgtlEW
WVsUW6xvis2x6qZv6hmszyZ8ywpmT7nLd/+E9ysVIzRqWgAF+4HcQ7a6Tn+S0sFFSnN74epXjGij
74Y7BRo6pzYacbfdiGBTAHD9W6AcIWudZk8Efm+UW/LLUgRJofAVlCCJfvNgi6EhwszeutZxjLwv
KLi7uqtm+IRLlHKD/lV28do8FoNerWDZxpzZUwNwxb88ZuxeKFl21qe8tiDyvEtS2qOnb9w8lIqo
SJmqyOAD+32P3WgcBJ31t1wBH03vubDjUGf7q8DoCPHSUMdWQmBPogjoQKMLYUZWpYrsO/y5Kt5u
Ym6NTAitXOKF7ZvPGepTWrVAyXDV+e8cL1MAjNXobK0keOaLhniKL5LjWw6dIfDsySini2q060Yk
Bi/lS8Kx2UZrk4DlUEx8L1Ski4nu4D5H46ZCdLx/4tHXrj53Cxn8vkfooeWZwTybm/OtZH22bNbK
Buzd42JbkQg5oKur1FrSv2gV/l/GG5MyEc231qu540lopvNHdar5ba3NtILb+hJQl9EDpZBV0M2r
KeiWcWqzY7Sbos0LIAorQVam3LOcTCr2YM3w8l4ZWWd23NfZj8oZ9BgwJXVzgtJlcJmsM3ITKIx2
tbXQByVBntRwGFSX3cK4VCR06FxEGzQ47E4EvYloZzfkplpagTnnlCgBBjgHBDsF1ahJ40/T+33Y
QR5x4sYlAuypwScEKHzeZJQuzan5q69aMmHCvYzi9gIM6MNWFiRQqFFj7zRRCG6HKIW8+L+027Dy
5gDqT3pNdjDOEeF87Z3F/D9KwD3XT1Skhswp+Pe/ACEk2KZELvm2dIm/nlArNx4FRKj67VcOythI
AHoMNER/JoKvicVqtqU8E/uSXX12nPGphDEA+XBF56dWM2IXIXIifJTM6HZ/MISswTYUvOzDtWZt
m5Hx8BteG/19HeRgSrYrDgN953bHSPXnIa5fwL8Gwa7DbMlEpvwlbnOWwib8bFe13svngadGFS1l
YAm+dLsWRQKOtPFNTz+0nU16FzYhVDdhUDoTMXKA1qzEFHE9zxFPkiCltJM3R7DjJlxTihfC+1M8
dUni1BxJnNYJkApchFWzwSlkKsnfvmnQGcwFZCZFlzrVTd2dFUBKR4aJvIChfd58C0e5w/1Yukqw
SeWvuzh+t6wy+faCp8BLTM4MmNqtFUanbrzRxcdXGjI7/veWuPSY1Skr2lHfhbzmo4Hn3qIgX8x9
zxXU13mCH+B+EtRBo3EljNQ5cHaktUguytdffJbjT3ZAeFlh/rsa41fY3lB7bR2zDz18NQ3U7zD3
ayMNRYQUN6GUHmWSXZpyobRpPJ5J7rVhFt+upHznFR6EnKcmKtI/OIJJlnZ/fFsZn2/9uT5i27ny
gxBeYVzLR7EeW0ic6DcvW5EavK1E59+GiSLbou0YiFcUTFQ/hAay5ZhMQgt/uVAU76h2/T/gkef6
PBzG3TQe2em6yJS2v/YJE20QYbkKzsmkIeiWRH9UcmuJZh2tL2JI5eBuhrAJCxid9D5PnNUcj8t5
2MrSaqZmpp6KtlKAkJuRX+VG0be4qd6JgZM19rH9DM/retoii8/an8/ztGYM9awMX2yty00DcMDS
Wqn1nyQVRNtzqLksOC6af10D/KncJwm3pWk/Cxbj9aYqx2GtNpgGxajz1EsWFYB3veWJt0mFohN2
dmsqzd65M6Tkl0ahzNQQpw5wFOVMTsRisa0YvJSHgG1mnr5Jy4IEipRZOjBErGBqWmaQq9QAqhVV
b74eObCIL9BdGGRRQZCTsTRyQhuicoweqR1q9gSgwbT3YhSA+NsaIBky3LsZ8hNO5GDUZXj3vea0
yo2TOc9aOYde3QAITa7MkPVeWS1NdVmsASe7kOTzDMNAhY8OxyUSAKMeKzuCh8MA/7n97Y+l5TeM
mxJH3g0wqDRWnIAgXqNxhnU6859klXpcLKxL4qZAJNmQcB+Dct1Zbo+LcKoMMmG1PdXY3s8FKC4x
131CXxMQFuAF/sz7witCmOAK24vygKVhMgIsjVZlz3YzHCvpxexksNrGWuoEKIRb82dR3DloWtFY
432CU8B9iRwZyBzC8o5PUPvlmgZZkwG+8lIuHIwxn8SMVcL7OVWPhwdrqvdbgNi1q11TgrUGve6l
gEKqcRLCDdt+aWrbB6/ipjDkxGsMKB1Nos7rjGcY1oKh0S4rUjxlO/huZ/Drq1BEQW2n8ExcfYLa
A7bg8HHjko3jEU3pJZ9ekKavUSJ4sXgmFLelTDIv2k9W7XuDgdiKL3NRbk5ksS9+jseioPq1ikAZ
Fo6/3+0Zwk5kZoDJLHOz6S+eMHOzkI5ADahBLtKpNj7Q1yl0N2+eFzxh5yEFyO4Q4JDGZBmJemB1
TprBG+DiPoRQx/zj8uCsx7uz9OggFbf0Bebjfp65GxjzcSKelvSjoNXxPrj1ItBBLRRs+sfxKmTc
S2K+eq3OpB2QgCjwq/4KmW25btnTECrbImHhbXgbgbrQgjtETpQs14MpRrMV3n2n8F1+dKeZSTHf
UzJ8gr15zmEKkLjkY+GYf1LbAC5Ub79HoT+KChL8bNphQy/ythEyZCgssjM+hM9B9/g8qI+vE3iI
ns64loJFUQygC8qE6wNpkP/ubq9TH799KdzDLDOU2SBE4o8yHoV4qcEe92GrhSA9w5ACI4ng+aDt
dudtTyUIDe3Fx8tbwtOiBCrtpcrbzST6XqKb9mAE7iCG+haJd2wJM4cUI2XiTl/2bW6pohtnxIp0
U3WxS2lpbsI2uQhHTBTBgTIN5srxl+4EYheT9g47C3d106xnX8WgdmI1caxxpfKn1a22z1V5HLBn
6MMUq43w82QexoBULy3MDbhcsSfB1iCC4qLZEjebcvUt6JDFpq/kcMTOhCtmteKmpYJfVXZiSi4a
/KlsB2i1EKZIltW/zBlm/zGNZbyEen91NI0TdlfYmrZFw7DbRFME4cJ5lRZYOLfU+/Qq6CFANA07
XUEX5vEfiAjX5A6Lt6bWwlERvsWfY0NC3bNt6of06FzPwoe7L0WLpdHQIy8I3HC5rr0ea4H6zvUP
gzE9BVrDeaeafJJymmKIn9oC7OtyATd3zWef47h2GOXOhj8+VGdjmV7uDjNZA+4Xvf3ukIcv17Ms
0fC6EDTLSDo1N4ETZAIVvqwfaD08oKrXjESdytCrU3X8KwIhSb2iyxkZ5AoWhcxXvCzxFAHot9Rx
p09GiLWbKbneOgLbRHrAa0uwsMOMWWieJzbyPWNO4iPqJ8gDVLRFObagNGjV3gc8wBCKXoG7uhpM
9yer8GZtrSNSS/PHb3wL7hBHFHabu1DToSvezMjDMUQ00m/83zxil4jpO/y+h1YPZ+RZaK8NPLfx
sv9dfX7FXlCcyA5h8RyJqQhtDwQWh78km2nqrmjzWI2Av8Ihx0+040LC9PoPaXihTXsh35fPAUdP
fD0AG63fY0wHqK1muZ0xp4RI7O1mLm/qJ2oVtH+sRQaMTfWnEeX+6stIet/mOeP8USEcxuuC1d2f
G01RNKieq75p6CfNynrZea4LQBSPKsG7Pcwx4S4zEa8KSMZjORQq8GQqmG4lIkkMT4x9coScjY/y
DgnCvx42T09vyEneUTNMT+PSTOiw2OiXBbM+shp2PowvidQ7OaITd4Rf1RuOOFvmo1JeGIDW36Eu
xKDIQiHbAXTuS23+HjV8qmOhHswN8G9hJYZwPOK99SfZ0ksrwUFI1yrS1Xwl7HA4F//NB+mhJ8C/
SZTMdFFGNmoNEVGLaFd1c9K5CPNQC4G73JKqHreF3UNYtmTKTKlFRDmP28UaTKpU1el1+CTWObWF
WAI+nAxjhbXgBn0cWO8uvt2hGHwkRQhu37fQtiamAldIHviAHx2khVryM7G7EV6ifK6O5riC+M2y
Vzld+fZvkMHqhiaU+P8gAyiKAAWGB5xHLovSCpRH4YWVgxd6gbusrK9OL6W2sWwGccwIMb4fqAMl
nTQdYnQud1pXSOGDjJxPi8pzi3OJVsTHMPYIDY4hDiszSih6AgzB3+5PYNveLXBXw+pAXxRzdZLq
cnpzPItFAQBHMy4+gwvf9f8wQ9DXMQpiceBrCixHebZaC5hoNiTN1Nd6ah+03iiF1+avMCJU+Y/m
/5TxCSDtsfwc4uky9gf32P+4WvIfDa2El7D3lXvXqk4HEO9I9BevjJVCcUDXpsNjiuyuvj7Y/Q3J
Nvj/tD6TUv0yG7dq5wpoBiMQ1B2/0xYVidfWe7wkLxOrudgEDnSPmjbwPBS87t+TBELhZB6w7P3l
3h+g++D2GSAr8hYFWLyZz6/GaWAqZVWyl6nu/vnCwLxZpMWJOprOKjWRJ8xOvNsok+7G4OJnQqvk
BLR5SpYisIzt+qDfdamckx5wHwMOVrvTuvVOVI4wdrlDcIZltNLQNq5My7bbD+V2tiO5JnBDGsVZ
sPiOnf+JamGNLPQ7PY4pL2CDRcAbu9ws1pQ5MZw5w5maZULujDvf00BwBAxhTMSeqsK91HtKTNZM
3SyVbPwZV0tql/udQmgdKnasGOM0hmMSrgxOr4N/uiYBOw4yl2PpC2RwsXYRqW2Oy53iqtDQ/mP9
a5kAqBpOo/iT3Tja/Js6lzx8Nm4Jmo9uDraNJtw2/xLgp+9RdgSq1eBIS/BjJav6Iewnaq0EXfwa
aHTqK9L+eC+6oBk+1bd816wvWPTuuoGOHs3Kj9G3wY9x6nPrqXIkubzQgkwLhZ0oQDV8g46Sxxws
MEbakEwT8Yn2BZ0BnO3Kw5A3mxhRqXUQt/FdaOB6O1sGdZrnDPMjp2cWQAiLBExfEEPgVyeLKT9m
QEfjqA2NCUBZqHXrDc+f8Y7G43kcnG5ng4d5eGQn8AtS8xmh98FVHjxpUVjcRf/KxeuOjevtdJEO
I77prAZ8e0S25ieTfZLxkmlaRlHHeLbV7YePSGCZnAP8TDcVo+8Tgpw7Q0YAd2sHtZrL/FqOa1gS
SxrVTafa/xh5qrASzsMucx6c6DWWE5SUspmaxR7jz8CXAse5tHvNeiWcska5ncaGakr9s9v6Zeow
Sp/mUVfAlXw4DvuH2Mv9JjiFlbyqlPOeebN62HzmecTu11gyQ9CWYl9iwpQYoKscID5+ExpfiYDn
FkqNquO8O7N0CGzjSxddsrB/5W6X/L1T0EPcqsOzH0wT035XzdGP03nzkg92nBjsWFzhu7p8IgJT
yU15jbjmRL+pNBeK0EEgXhWVQDv0JEFTbLd3mJq6uv3fqVvFqIZSg6e8B2HiAa/rnxFObYWxp05X
jBHpFnJyawu+1Oo98W7C4TASCRzjV06AvWp2jG/ppvMOFAN9c6B4fEUXOA+V3K8c2WF1RQkiiq3X
4d9YfmYIB/MBFi1x2uLYOND2u5Mgybg0QJQ6xSqFr2g/0LpVa14rEmMYadRr7kEdqRa6tiBEvGWe
ug1E9u0ZWRKjeuSjagzkj1qsjaBlxzdhjZKGQ8sTENTxQV5LYnshW3rhxTaRISr85iXFFfMzRa0c
wnQJ2sAE2bTIO9Fma1dOTI6xxQLGYKJDU3IuJQQ5ZYdFmI7JKYoyT0cLqfcxbH1J3dSmtgjKAzUa
eSpEXfLoY/T0gp7ljJ4cRsGdFWODsc44w35IJJ64cIsNXK6fcfVen7n5yYu2ndqGIehT5s9REOZZ
iUdJ0hQoh6zJ96AF+Q8TvLZiObv4DlE+U3V638MHt6X9/y7VV3k9xSkMZR1zBcRXU5UDOaHjZaCd
48h8IBR5H4jOaJKvmnkVURVJgOeKlRPd8fFOMC9ZC0lXJO0+Apo9PYplACRf5eSHqz0GcBAmePgq
uQHLycKjF2BrxWnBxBTwFwzh+P+gHFrVzYHrqGA2Y6Pv1hjZybEqpsTGt/E08kvcNOCxYE7G94ml
hMuGS69s545JLOhFEvlX4X7zyXq1F+Qh5v15nTlS6Pin2psbTZm4Nd/6yx2hia66SlUd4rP9+zPm
9UbahRjC9Ui0orW4a2VVEU+KaLogZlRe36bc9By3KrEW/ktAtJoXawVN1Kdk36ABVK64VMll0g+p
MRSLPrQnCV2AJt9ZgsrpzhxaZmkL66BqhmhQl6PTQjSzDHAIqXzZ5yDi4mG2rCzNoTMLiuFwJkJ6
sQ/UoHUHD7TrPoy/8NLszRYbHqCMPLC7LdRzr4tFuXdlDSKcTwfEnN/UhXGRlyuUiKdnpLriQEyF
/E1qWTZinmWJof8pGf1V77+B2TAYWDFsadC12w8YKvVMg26+jO+drHFXYOUIGaj4MAitucus4C6E
bbwU2nxr7fJj/fZedl7dVB3jD6ILaeSyp/h3cdb1ECclLOtCl2iVJQU4S7Czb1wpeGH2pkxNF+eN
t/ngsAyzjU1Iwd5U/RZ3C4YRC7juG8V35XLIQXuTmM340XoAMHl6t8unWnafaMfs4MWd9D+wxruZ
0EkaUB8Fm6W+89CBw73l1SkDvh1RVW9cVOuNaPJjjs/fhOPfvZ1F1lrPipCyAbCockbgIGOCFbUM
zv/v2LDL84EkId1dz86qUz2psZY8s4Vee1mEKDzPOhIGitP3Qo7KgNdyLe4fGtDe8FRCZfY0qWx8
HMasFZl2rdifMM5NdedndsiDsewh1Lt/JiTM8Trxd3zC4ZjMdQLgH97gwjYu3a+vIwrKTMkE21x5
a12HpYuzQR+QwYGwaUJRb5RNVCkGTOX0TVXFJVN3IejVO+OhZGUZ4B8gVCvbDt/4wxKo4ikmGWgl
Ih/ZQ/LSZAJ1ZCOsWmxpRSq/DjHeTHWb0tpJ1L0byPxUeF4Js5V/sbwGq9P1BHfSFvF9p2sho95I
GR/TnX1P9D0Ta3YsRxRirx1Tkm1Dip27ifCqLAqNMej5xgQbj4aBTt2T47o2EWztvLrqjYyJhYmi
27K4cJ5Gm91HSyu/fM2ScG/ytIqbu/G9c551BuS6hz/r2JkBi6PJOHGPEQUB/xFGsvVEKupnZBav
wk+OcHVDv8vDlZ1BWK0+56BLUrPkrk+kd/MTNR+9AyDyLte2GR1MGcLBqEGWUtekFNLLUa/Qb77i
LIPzb+MkTKDFjYNynY4zhh4h+Jwdvvrj+3u1HA7umKb/plJ8KPHtYCH9r7yOBrSc1f5dsiR3lhlT
7OujXAxJk8P60apDA4EXlFUEZa7HX57BREipCIizL+Gi+hc/8+82jXqrL63LVuA3HvZAoynu5Qvq
25vtSJhDKuc65Cwu4NmDnTNBTvSZC6CAzzgvdTuIu0+G6rHXzWXEkAdFmPbwhjbWJcw1TnBLTAtZ
d6/rpoBcUqXxLsRDQB7znLtHog26vniZ02F/R+IBh+JdlrJhwj6lWBYxEv9LRsr8Yn+C0sKoXSFk
9QHv+2zkfFACIm2iJaBJ+CQ2vb5E1zcT73g9kyXUT3CuD9AEbaiRHxKy16oFfZS1POlbCctQbQnB
VfomsrvOlWeNlr5lufIy5s4sEdca0k4+5DfAOnwNbQ1cm3TPgX5TMgdMvrpww2PFV2cSJCS5AIsk
y1yzNrLBfaO/XrCweJZStIY3Ebn8Qi3htMnN89fv3LxFzTwRfk/jDhHQBhtJUdr94Jck6a71x8As
k6RF5q5F45MhZKloz1Yov6sgKK/WykzL8s5DMt5ydL1rjHSUW9axT97Zzy56PIU2fCdJPl9fcvY5
qGVHk8mJgTGjIPh0/q1hdcNqV2R6r7acGpl3yzlyeTUGT6zO36DGA3HiDVSb87LnEdXX3TSTmcN9
O6JlENxBtZxoOTCbdMa+9+xC9wP1nQGQPYV37GJ4qxc8l8E2DlHEQ1WDQudqZkP2EQy2Uo35KsZU
pibCHbVNt/gZxqd6jbMmEhIiyizXEDFxcL+3z22ubKvWlxGIVhV8S+CzMvwYABcBKq4C9qeYQUBH
OqEmyoApxPg0U4TBiJ+LTC75zODPHdkTzwS9WzyfQK4GlhWxnk/SfdtJYavrIvHIlN6uOKV2CvqL
1Ps2nvqnCV0oZUVTzNwS6qEVS+YJU3xuJOQzCtLwjl+lGUl6/pzy/4A8jvlImDMyQxK5Ly9/XSh5
qU1lHpOlNgcZeI0cLNwI2L32uOe0HozM+t6cF51RCLDIoE4L368NdLtQmtuE7yCaR23iCXqk3Vc0
trINNGuP5+QjGFbvGEQubLOAojzv23Yqsn/3fkO+P0U3lohvD5wQK8F05WynJBsCFsOFMOCLK6Me
biHImE0Lstte8B4ys4eDGc1FxUj0zJyTekqalR7tXaGi8zpejQRSnouvAS0aex0YjH0IF9SQ8wS3
K5yF3kwei+Z8UJfC6QhKWXe+ySI0Sv2SWwGQINxos+uRrsZn74LusQtWy/9SVP7118z7bFQQhOCL
jLvpA9IPd13pzhtMIAnbGrCD+Q/ZJonZNNWaoCYzWaK9EbZaJFg9Us1pi/sUj827OqfrgDWZmCoA
SfCN/g/S4Zr1le24oG4QD1vGs5iju6paGJ3gw9Nfhm1IHCDPh/Uw/M3TMQ6dTubZyzgDmK93wtua
+f5yo+1S3Wh/9HNSN0YRBNSPVlBRW9ubOIgt1Mfa79fgSz68qRmuE9LSXQodzuBzlaxzRzqTfQgi
+gTIHsf1RXB0S7wZivo+9zUoGWvZPWgeOjm2EwCZw4xVXen6HNc8FmKWCLN+pjMwYid6Bc76I7Hq
/q6yfBcGhitcxA+v9O6CGwFFq7w5w5RBQxl8NBrD9TU+OMOXiEJAH76p0KQRgv+UKcxP0hKYLwwk
bNsPPeeS7no3uS1Ng2Zl8knW6CspRY0BHbISxCUosZELlaRaOGPN0Tr5s5Q6a3nRLkfiuM3x/V6D
XRxE/5+csWBLm4O9FcNI84ZwocEaf8omNfBaCuw+9JFw8rWHOATdj0OZNtlI1roO2oLhHWULYbxe
M5kjPZ1OydvHTLoGQBXOeF8paKWsZQNBH8zabY+3HjnppMCYHy2OToy6LxaahL2+QGkioYuRlMvZ
5ehN8niE1eF1IC7cxdAYF9u3MpBEeXXgtU09z33Fk4ueeugfa2dvOgdFjUdXu84yVIaKKtp7a+cr
5qvoNbteYxMwwWsNIgDMmlsH1w73GcPZrFNxdquPs390bp2Nne067rkzzGBWTrlMWrpXMyhks9Zy
a42JR3yIQVGhCdvBQBLPoYubeaQINu6ujwkC2xevEUwDtfW7iDzELq6jL4XIzWKRM+RmH/0+RwXw
mVQjcH3dl2dt+jAWqk9BbMKwKtHADRkK1lxkSYxiNYFiW0xgKFKw77lM0zDM/sy9tqCfbAOUUswP
32FcNcJv9gMKokOUjGGVjfmHVWUM1vE4Iw5RA3y1WvKmTWnm8//vJ1lS4+FH887WjK8UUsjUPg7N
P5uRkEx/ekwCHLwBhYqkEXRzY1r7YOa479lDdJmTR7Z0r25q0eV2V9fluWTgZIare0efqKQczl7F
H/nsmpcnni9fCxyc9tIMET/Yy/870eAREbmtvBoLtCVGn+gYfBPm23fXUzXSPatJ5p/bZXOdcmqa
Xn6FnhaFsT35WQn+fBUIZP1f1oB5C85Ir97mPtOgE1wPdaR+QcefRzl/00Q+aJvscd1FlEZVDqkk
4uIeBbV+D/qPc1weTDM5EyNWiLSIhNd81bQLJGSQ32hW/hE7K9q2bp+H+ZP+FqFbHsSQfz8BXC5C
b3CdqNJ+hLaXlDsm+BD0xqAmXXk2AkL95C0OdicWG8t+U13ij9/7snlLbIXn19pODHboLNeUniMH
Lfy79tWtZsSYbPFMosj3qj/DlunSRdOBB4rMRJd3sXU8tH/6cMG6jZxyL8AO9iTtOYdvYPl07eUW
8hXAWiIbSD3rhzUZmXh+cxUgrYkzMtjPtzQkkmPPVUD8+Rv4SI4suleT7kNKkJAN+03iuLPIiMPf
hE6WlnEyWVQPSW0PN3sIzvs/7QULl70liitzUyaFxq4heQWYAEDkv1cDHt1ervAy3Kka19ckBLzm
1k+AZApOzc0EyopWsDn8C6kCMtHbU98xnOm48rRRqx7Y4LiZk4oQJMQZr9mUw4/QLBnu+3pNSUS+
I9hoW4Oy95t3Osqp6XzZZ2kffMf+JqDiSYfzIe/2KS90d0JgDdLHvXBFwUJEobEJ7TjM7mpFs0/3
5Ft1iHSSkFiIasMppTqNzgiBKRo2bFdelt8vZB2ZrG3W4bfLoFjtouyhUHPyJ3GDpESt4C5y7kgR
Jnz68OsEnSactd7y1qGKeRufQ5U1fKULaILtHnMg0zwRLZI2NuGj6kaZ5aSZ88YdPEG5b/WozCDo
woL/yZy1B5A2J130pKmgAbQTw6wswgK9udOCZLJhlSgsXzeJ4Pyb+X+cJ75USsEeNGfrNdhZslVP
UI3Y3OzYJlRgTw1UN84xdDgacMRp3DFbP5aOhCLQV8Dqx0JoCGlk1EOWjMxVtnXn5sQWRHEfJr5o
OrwgbGuSz1DaGb/yd4s7Fkj9az3AYSNd4P26tvurjybt40y7Zia3mWGn8pisHIhEp3vJSsOrMAFY
mlWI7/Bm5Whi9c3+jD9f9X+oThQvbo/sH4MI0SVViTbwGZ2+QhI3rZXmFYGDA9LDaRl5nMb/VD4Z
4Bo77jmLzRdouNLklg/yhdpgBZWeIWRQt2WQiNOtBfEZQUeaNgCxnewYRl+/OADvoV8QDCQm0sXI
7uM23MLobgcZx7+dZFJGWMsMrcHFfixkN+5AL1jhYgp3gIwKmR7ATDhxlQIiwp7CjWsC6/NXTo8v
eAkeyaDcl0UaIMJMh8BBiz0OyhG8kA4kvWk1QAEARXCVb8GSmL0XCsQcxvYTH73UTgAt5CuIoRHa
RvPa4j2WJ8T1zSxYA0MXIu0kocYGvzdRcbciL5WC2Gg4niHP2DLgIjmlv042g95xBDLBe6La9xHj
RwFWU8QTEcKsvmWCoKEfS0i1jv6yNpa/AwkDR3EnVwdpyl4j1ojgjboe+R0R1hSwELiYvQSt8DRo
tmUIdWIPHvH8IIdNeFkUBLlktuOWsP+u3a8ydTJopFH63vbMZ7keDX21vF+M1yGwIMtU/WA4jlfL
s0cyxRiICpEYt8E3cvLvwBk4+Y8VZdtILbk0QVfGAYSnHqLrhFoJzHITC40MA6UFKXGL1S9+qQLu
YjHVhgkfxJsGJhn5Zqvsf8FGaMMLb4ccJg9+a2QzaS574ALsFntXeTBT7ixv4cz2IOkFifzyFDz8
PCo0neIaeAWMVAdQRyHZFyDCzXKzibXa1Rj4JC0Owx6OQ6NWuUXITfElQRYxHzfUfdafjMSSj0n4
wAh/UdC9ChXXvrJ6XbALCWeFVCKT3KIpaRTzcOakTw3DlWM0ssRaCr16fVj1cbtmzaod6uyhbDet
7dyedWY3uCEi/Tt/96BU7DetccOy6BVMb7xgIBiwikaxrgulspUJTEyS4lo/tQDa5YdZ5i2LSmlT
KahDreOX3BLL8DwIYmCInpOPbNbiU85n3kicIounZm5NqOXRDzwKi2EH7xpUOFvZ94rabi76YZt4
Szs5uee5QGLnCsEzdL5ltNha+RfVWpOBqIEr3XJk9MWcvetxrQihZrcoMsa8CaCLdXcjWosJz2HR
P+aEMDDeno5XihlDGjZEm3jV+KXcGKCo4pBffnPeJfu1ldbL9J9RfyxdokUaLOVehfTdOSwFlcmd
hG7PGVo4bf1tqParVJeURK/6CFEfgkWwTbPe6QC1EXL6m1mXiGsd2ezfLl9axRV+0t+w6lThqpCa
wTnVLZvhpZEnQwejJX6ZYaLWY7rX/S8MqJTH5TlbHHVDFGP9VCWi2nCSpisL2gu9Mf9XZ5s8RI/W
B6qcRT8MaE0yspo9hLF/pzsxmjryrL84zit6wyIHv6CLkkKWQlImoYrVpBhSseshFN0z9CLUo3BR
OhB2UYr5DBhXhP3oR3XhsTCSnTgdi+Pt0hr9nc/f91i3vyaVLL5beVkf4KblAdjzjzIpK1x+ObOV
3h8s6yrw01lCdhTsf/dQyUCdDT4fiUyKuuegKLNd1ix3BwT9va2SVczcZKTYwYB5jAGs2D8J8V6e
LCP/5sZMHUrn/CR1HG73klheOaLYw9VOG0yR7Xx9y6YowLn9Lk8ZHBh6uhzMEvoxor4+UpC7EGuE
TQ4udVgBI/3r5CfuIrG7JxavJt/Nr4y6RSVPIIdpUrVlIFiBB31qLC5wT5zoRoRaTrWNCDOdNoyE
TYrTip+3TYpmUgOFXtTbgT+8VQKsmQslKKfWZ659FI+ElWGe1x0WbIItxcH0PTbCsXVLTV89O8vJ
+tiUTWnOTJ01F4ZDXG5lVMeogxYvmwo4RC2s/ibqJCuaqknRR4OPKDK0PP8kNPYfBlHrsOQa4hrS
/sYdH7unPakItuhNN6LuPcjl1ZbU8ahkdG2fo3D4pNQXOdDbiYfXAedbBFjaGdBoxqXpD2x8qHaR
VY7n8w/nYhc4SW/JPg1RydpcYfNMNAMUK1fgmTm3r68u+8Axrg9mqH+AEGwFr79i70tbgzdFuaGb
bfIrgDVvkmDdluruk1Lfa7xtPHxE9UB1J7Hp4xfO193bs/1dzWEscA66hlWiGMuUZNxUcjjoGY2y
sV5nMn2zZ6+1ZdTdeiffKdu6iH/t8ykD6tf3+zVYzTNeqKaNvYB0rKCvo+uzNSjwLu1GM1FLaK47
iCn50jP3mGuHrjYDGClJ8YS406EgiPeNUsD6W5IJFQVRh9cK5F8N2JDus/+Pk6lILldyjxhJyzV0
Q9ORIKgySaGnvXtf/t1rtAMO3n6pa24MYBu6zNomKgn59INb0jBR6cj33R6ir7iy6zQtwJdlbmv2
8e8rArRC3yHCs22PW6a5sRta2noieKHbR1ueKAe3rvceA0x/DwCAVZ11JxMOZbmz50XUtvtSSd0v
e8pUTJylpG8KeSrVpzRyVUg5eZbYztRHwDM0iasrsqA7r7U4+JUjVC5fKccARmrvL1ON33G0T88i
CtuGWH3Gyj5OhhYFpEGV29jy/oTMeoyulfvXQf9jERMlyP6lDz5x9gC1rVZnn8qrrEfmb0xuWal8
QVe46iCZ/n8+g4FeUj7LFIIHbCPOr3j8xcbPoBnuXiTgw3vXqDrVkd64MOx0QQk+5gYQWbAj0U3B
IDgu1+FpuwD9whBitSdGt7RTQXfm82A6fYQgx4Nhsl+/VfDddB6Ns8jWTCfWVWQLGK7+/APLCv0a
rx5lpfuC3Dqq15oM9TmRGzBfdGguONTzvwZLml3lVs6PT2MnJ0RyERvpT0AsGiAxd8h59EFp8x8A
b/DYwxeUw+/JC88fR3i0+DxY2wBOciFzP+bVAVuCTGmYydAn1YQV9NEDsbaoJi8MrgpU43k/orW4
eDGmBtBh+ImL/8klVgDoay/VDsnQhVfROgrHEdA8ppmLGm+roEtsfdXVg//82+oJNclMoyZ9GrlY
eLfcLDuL4pa8WrQOXdoGM5PGNGBUbEQhKuF5EWWtYCeR0+0zYDgpwodZrpMzNM6EUwvzQ/0WsYHA
0bLE1OMt9BHR6OxJYxW6K/cS3se7HUmETtjAl2ao/4eu58t1GRqtkfxPHUJrtGZwc99Y58mp4EPJ
hKww1KGVkj7G4jRqUDEzvMA/lqWoDP29jt6vtLa9eUNaWJoOrt/Exs5Yr6QopsoCRLNC6bkX42+c
1+i6PNHP+W+10iA4lsJFt7qbt3qO9rYLCXl8xOlHEpG71nE42297C79wtULFtmF7T/CP12Iwttj5
3YjolcOBQga52f8rQ8UkkXgzX0lDuZRmHTwIbk1xmJyIDFjOU2BM576y7Y49Ft5CF4BWS/3jj5fY
kLW43E5nksysSqF8dLrBzQkuDXEJIxi1psDOKRaD5li2+tW6UXK57nZEMEJnHWiIct4UkpeGDW+N
s2WRYD95eNFYZ/f7IG96ZmygMsY8PvAvRpI/6CGiYLDXjhpzpuph25PAfrE0Cc/CvwI62PDCJ602
vpOFxdrd6YSPZdhFVO7eXEBZCyF3mjIwRJtW6RaHH8q4yAJ7cyMBYugzgjQkLugJpI0FR7ft5Ac2
LPGVUW+shyavMtxQsQizEJ2ylkieYtBKT/oZ/aAmo3R3Wmspl5RNHHqxCwdVyxKMMqM90Tg6cn0U
BL8FWpW/bgXofMKR5mMykpZGbKFyq/uJhpPgiMV9pIVJmzbsPksNmpS5i4Kax+11Fsxdbx9dhVvH
Bn0eQGhYGnqZfDM6ogXPJp8TAnwj4CUNMhhbUURu6venWDohEq8pOLImXFrslMnUJN2TtKIDOmt4
F9zw1nT+MpxQk0QIe7NWULxU9O8KZQoFtA8YegMEHDGMeOWbufa/JjlzU1+9Z1a/u+DRloGzlfxT
1lcZTp+8eI8NFM/2s5znkO6NanBAFX1ol3gpzw5AgE+9x1FkP/faY8ROf2ZCRVb2VWi2nVPvakmt
ByCwSuGtQlntn/bbkbKX5G4Ej2xulpqYzOS/YQ/xGFEg23+jr4B9D+seopV4AXphDX2MAn32h8eE
JfWuZGEgoRiq13jYipvH6SHHob7Ux20QUjI951I/uROVUcXFRRtQ2CIdOY7oex1pKA3zZ2UUuWmG
7DuRjX2JeYzWdbSdZog+gRIPZR5mzPZLtdrF0CV15+2+m6+CmliarfBnr0I+jyy/oBQ5V665BeVO
YT6TTKGboq6Di4UuTWbbiBSsQbOb8nmF59gc5/CxbZ+FF2ETSG5imfG6z/9Ygl31ixitZJ7HxzQ8
fB4gicOtXNUnyD6wccrIPZJvU4qO/j/paR6JALzfgJc3En/tH/yr8b0F9BkXh84CMfC0NWJidZdS
El4t8p4q6c/pqDfgYhX1+fBb0R1PVvlofhNyXEu6hbWd9v7eI0EhZB9YYQY4CMQ3uOEJQQgBeddS
XnvRSBd58dYdcMLeYegLFu13w84eKStp1/V7GkDYjfIyif/BaohNdD2LlXMom2o0KZeBnEs3Gtzx
O/GEDGZ0c+jJ4GXWFDhwuD0Ihvk1YcpsVTE3pl5m8DM6EQ4e2NZ5SyQuKt5v9NKGFrdT8irqkf7Q
tabqnU/c92oeOWXr5aYG3e7C4sDTyDm1bJiaFq0LJ01Y7cUyiApdqFdWhrahgEMJqgluYQNA5CCb
nncPeS00jXKuu52VMrUsjTY8/oGeG+UYxjTyhpzEEMdBoztYFTlXKA51Bt67MfWgbsskzlvxY6Lf
0RXin9uOO2Vmx+VzpvZqldz4shoZ5XiD2BFOQwNdgEQ079DUSuJ3sRanximJVi3ovE+VYgjDjRw3
1tUPGNXHvrVgj5BzBA9xBrOvMqPiV6YwDcP45uviGgjtzzdoKxP6OwWjO9bDjmLEpBNTuOTI1yEE
jBFe8C2S56VBxxmje1mAnSj9WVIAUB75nkCL6bvT5pcpV3kxXDceO1z16UfBS/zb8FEcwAjHwJ6i
9aqo0GNy8dqVHGlQ+4t373LLeG6lPXrwNwgtaGN76AHOep4EcDTt2TZaYJ9CyMbT5DectoSB/yp9
AujyM/XO926VGHjdaW30NgvSHmtqYCFhWsE3Yvdsh+ko4kKN59xWCxyJf4kJg84UctdI2et6Y0Zz
SNzYDz+mQlkhhL4ZfBQdGpx6PZaqWtm+0GwDfvBZxV8tE/bwbqL/alOBR5S7Vof2gVLlyP7bcsws
Es0h5tPY6ItyoOD5flSfkrECoSzFB8+6bwRrpUgJOQYYeI6ywin52zFS2yRfp9jqREljEvbdDcnw
LWzT689afdK8mY2xoYxheP3taLXCqExYsovRhgCg6V9UvPBbnt/SKUKtPnOA5WzoqFuvXrPakr3i
xS4SnCMLh2d/gFsYqMnKWv67BUtf7/sUib3ZHbbXbknjFYPGE9SlzRl9rRvd/vOPfQRKhoO3G1IK
3SWDZ6jcCmgH5PekdC/IJ30EdrPuyLU1I2HXIG+Owncx3ibvDKaXvd2/2Bk86xkqfRm7d3k2LX3p
eZWoUoDQVuZNuSTT5sHmeh+VIl+ADoXiV5kF7tvNVdiRpjHYZa3rchoPqoOsrSLDQ0Vux6sayUXA
X+uWfZY4pM5DNU3vBvgXkW1NTuPkc3fCUgysLbEC6I4MLe/VPA9cye0Y6vIyIQE6oe+fpP0+ySPX
tf8svXxXovrKdW+oqvejpCbALfvy8QVBb5hRq0TEbTy07Z6cFmj3tc5vu1KBfA1NlG718KzFcOOO
zbEJBAoB7+f2AjkyBQfLG644bKcCTN3C9vZOZiDCIpyWuk7/UewL4hcducWN8d6Y1/tjfqk4d8NS
MYrBbWHZ9DWLa41dpL2k74x7Kdcv9VNM5Xjaqpu79Src8zsikePOQT/6pniPdE1jGtXgrWYwIiN8
VQ19X0kgHNzYh5urNYCQeQuP5ulQ+v4I7iFeofCswrc5d2O2lENiJrkSBJgejAXTAvQiomIgjCwg
B5lwDDBaZ1xLebaHWtoukJheR7hbkIfKr066lvIgeFYqnoGXnfBzlXVs/xV/P+lthRLmBm9HnTpV
t/T6sMhZQIehcQGdYHQsMUDXG8DC+Z/+CNuOqY0oIO/YoDf2DAVauuNZQWh28R3QPSkTK+5K/BZT
uxOhhXxFddNBwDPwE1FSL/G2OhYN5ejdeCw+1gBWrGdwivn3/YFw/Bj3lGY3TszvRurRmHkb3YXn
YBwjbmjtLYxJ6sPlmcjD1NNXwK1e72WnL4zp5gjuy2LdD9qQkAQjdyupkDVYSOj87oZL65HSyeEM
IFejJSG34XvgCXQFsYuhUWDK7KtVE46IBnUmjI0ZZGckhSDhzZ+baYU+/bWJpLK4bByKDPlyfAAZ
FNot4xH4AKDxsmMzM3WWJwgB3RRmQxfvGAxPbAaKUQLIyDp+ytnkEQvNUHcUzxRZAdcln67XGEJR
l7UvRUedSD/uGENlR6HNRum/UboX8Pb84WX8rIheL7hWRFnkyLZTXAKpsD7EPMOQLG+o09Kp96I1
C9d+ZzpQn/tMOfQ9vGVbKAb9GlujVK8kDuaAoIs4RdA+gyovWoFAr8/LX420W9FDYDp2w/58jog/
g8dACih4HvD7b6wP5gVugBST0CU8A+mZGy1UcQztKc6H4ugS5blSIgApN3BlG79VX5lAsEBMW3Xl
rnhAmVMHlWS6Yof0M+wWLVZs6dAM1HPruMTUa3Yf7kJVxaenE66sRWV7Ep6YI2pDbnnWtO+oQ+LO
hNzsKmreJO4JVXpNw6mMXLhSTQWZvGD6KP+rXrIFLaCNZLf9XA3aqhP/7BERp6AkUwHYSUWLx9dt
ifpX4iQU0Ymhe2iXLQgB3U/SRDnmLp94heI0JIMiI4wel43T2mZQZHTN42e/e793cCnIVmivu2U/
j9Bv/x4ZAWEhw3CpQhneZLG7nJfI2WUvHlSVsn+sjoqiEYnGl20YURjIYno7c+TR6CYJ3Y5Cpjjk
8EAx5vXuwuUpXk5FEfdjfOB21rBptsZ+OAgV3mpEZ8laIeIBuqZf40vOadyirQedS3gp0f90n7nP
CMkp7OYIPaRj6wlfrrf4dGOPu6n4qmNUx/G/rqJNgAPhI0WfYZhqWzG4FS1OWFfeHwUmtGM4+McB
UCdPGCEJkmM5s8UEhKqTFr1vyJFx6tnV/XjRtcgy5A47OK5LWGKT6cQSTRwsVQacom5NfnfIpa6p
OaZpx5VQm+5Luw+DlMZgsLmcix2jjhZdlEDZnuwhu/D2w0bbYe//5y9Ziv9WntJxw5Y99ZFaNmf7
NXlgu8kdRFepMvOKlaiGIGs3WD/3xwTUkFJg5S/+efiTHPU/bXvHXwhUYIjX/mF8taN4oVCt03nm
9yF9I3fY2iZ2ER04qzB+yYDVSjwFd2HbJBtyWa1SWj26eiR5fTHkt6z2Bq7mXiR8+ALh3V2cvK3j
8JNZc2S5Yu1EDUqLTSd+TdjnnXVjA6BiE0gYvKZvmhiX4TSZsAeCRPzk2mefBiuGnSE+uhLfAUQp
jfHsYCjLxdhZmuBo+G1zFid93+IVoIdTHkxO3w/Xm+8/ibyX1A90RSxM3yatFXQtmWN+ZYIXM6iy
tPUxiD7g+np3x5yojHz9mmL7HYtc/S7nhHltSjx0gvVjoqIm7cIh77ECmDpWGQyEMpgPst5qK7w1
j/gkLugFLNAnRpsdFYVoTTNwt4+m7vdh5xx1h9dzyE9VotpCRnnTTY8ax7slk8Eok+4Y8oOp9ykI
AnW9KFuG/ijDTjp8OGaiOIuaAuezWUzd2Gv4hu44cB4fBvMYt+ju9dJ3TWMFxN1CUE0IhB4isHJz
Ol3bajwi6KhNCUnl/KL79M+iWBriiszL7mo7jRYQg/Yk9Y93DmusGJEr/nYOAP+qMm98f/C9LW9L
dKTIPMaZHnKT2+DlI908RRKMA6w4MqlxX0NhCKlsdyYYKmNmBxqDbHADT7kDTjlKwqzhgZZ4sX4r
ZvyRqHyD2RD7MJoexzexmg5tQoF8GJ7yjsdOJD3wRJMNqEsFmgtNI/cANWi/enONhK3HS+kD+nR+
JWSDdsoO6EPkmtKsWxmNYTATsdkaFjINmyfo+vTov20DkOK9lDBcjZTOL/DyVqbpq/BYZnN7cRMR
7Jd68h70lnVVJ2TeAcqVRIEothjQ1b9bkpZD0ifKwgonA6cf4lSLz5OLlzsC6kNKZcfhEXtv4iN5
XdIreD1mqY4HHmUms8y4R2oRy1ZqCT1xtPODXt8hzXmx93xcc8RFfhLa34a88t83blIEUJ1MUjHq
XOgt90VpoNOgbP8filWv7Jv5Zm6Fxlc2ve2zBmMTw1Nyp6i10WajxxCIW82s70ifhm4z5MdBZmnj
TyendZmogZ2D1SXUg3EbxeqpsIB5XDQIUmr43ZPR5PrKSmMYN8VLitG54JLt3H4BiD7T40Csg8XX
Ug3WzEYDYHGaxazwT+ZkPGFpBkRRaJC1zN8kDd37f/ve3DjKYStCpUyWR2g0grjZmnNO9S6rNzrG
GF2vd9xw03q0dWLqWD4DNTxjkh5SYGkaLiXkSY7GdAPH1ifW7EaHaWamZtNpQGGpNibWh/lgZvh0
spCl8l4uXBD+S2QuH8jyOdFwfiiC58PLqIBSy2K9CEWcM8/dG5rIzPmDujUs51JxaIUK9GzTZfov
XiqedzqfcUE+YzVcjaKi9nV1mX73x8xMynvfi7KSxBOxxkPizfjDnLrQTPP5FEkuQNsV4yOHFWnw
IJufjmrzSJMDOFfyaNA+QMnzxCJ30Mkp7XJwMwA1d1UiFwFcNtfYthe1catx+SebMMATADqluLHw
PcTJQJHmNiqmSaplb18tNxObJtzEK5w89vFHtRdIQtH/zwemsJdPsC1bUd44WiLYaHuzLGmlT3uh
aoCfU+1GrScptdCBarD7OEJq7U3koK7evQBRnyF9iSVOHU5wX37yiSBFtjZyy5FHcHDJHqOg6iH8
HPpccPZnD7N0pMNHossec9jc3/2XLhkIG23udzJDOX9jyLqkrPmS63nS6hVcVg3E9JZqssdLeP9u
ytig246fqlpkvX9bXomx1+8+s3DDQSjoHToTjsp33kQ6DMEhJ5OmTwKFK6hEPuXir1HuRJJKprlF
9QP1hNemMM95kUcWiAJ1MVTwxin0qruVkDb8TJFbWgdBb930UwKPYrqjeKTsD+OhKuuFlYN6ztMX
AGNv+EZkAUoxauFOIcxZuonpMmkJLKg2HIpemu+KEc2rxrNyLK0UWYzsgtcTY7PDYzFx9gnF1kZH
mwoVkN/H8RvhzCoe934IIFIjrVmPOLpwXxf3jevJcCiRisXK1U/VL5aIp9pFSzWTfGXtHZd8E9tt
WFHop7CtpSTrYQY0t165KbBGxCGs1SnO/nN28briJce+DvHYY5xhHusSnA5M6hjcjSqKWrg68iEt
gJ79e1dDVeJeht5ngxGU4gTOFQVTMPep9BipsSmsGEKMbc8u5uihcqEuBKMA2eNdMjAxjVy8IavN
ujxGKdJ1FvynALsbfbZ5pUo9O9/TI3eRYTahy1tzffRVYwx/Tho/q4hBTu1TxIeVMbbFotu27kNj
0v9tVJvLzure/6jXzghq9dt8s6q2SaeGzIcs7oHHzfEqTXJRPWbBO9XQpoF17prtK4nmhjNe9dTK
pxabi7PVun7FDYWjqNOCZ4l6dBeBmv6A/k2TTmNzle1Om9dm8t+kg7m7Yee2XMslxE/qenVn/i00
mDyeZJTA/wpqlL/JQb+RtabhKxphaQ0uloLRK43oss1WdPjObYIHtLfZ2znXgiS++E6Wf0gjqWgF
ZC1MCeJGK8ZZyAQo1VcjwHz6FqfBfLVbhHg4XxCivUC7lACkoAAaPatsI8hazAIsBWeQo6V5HMwm
1Za0fUFszJWiTUG9e4U6bJ/Wk5S76n9vw/7CIjEqUrkO0prpiSNXibJR7Dk92Pn1vQymMd7Qk/9T
fGMqTA13cUOUbMPUgElBu+D7V4Xlmm0aloWQ/wpIvQL4mJ1VwPerxXefOPE/b3KINPENYIHGI2K3
nUtbzTnybFWkXtoYEJuL7CNEMr5w45LH0S+pnO0zM2PM5e7HKS2Iudk7PBVcHXqXyeA05uNJxWQi
4TWnZF43f2WZcJ4uv6mEsLVoU32Cjac7g/aD5F/YxNtjUR7964NVXvq2K8NGxSFSHKYd2t2POcWV
jia0VKYEnNYXhYIMbT4jrDKRXrf3AyhGdkNcfaC3twcS4RgPAMeJqvPT6xRmWzzS1BE5a5ctR8kO
izKRKQD3c2k83I3DqH0qjZIsDRRSuRPzZ7aUF5XIL6oeteG9OwB1mFeirw8oR9/u999Tsp9iXt5L
4JaBxXK9DVUlKUKZlyltLIpIH33+boeLD04eTnyZlRpuEk+2BDTQmKGoP5Nm+OWtZK6ouu49B4dD
pmixE9jnPpP+cVAXbQUKcGXY07U2l1+l4nSqWkPyzlyiPMLZlo3MG+KpVsZFMlh5SyXEucAJLEWC
M2bBEeKBRIntGDRbViBXNIUtMjr0iqiTkE0R3kae6W8oyYZaBYkzzrxeboyG7Tn7H2e9BkmfXsCL
bsYBmLP8AemZd9mUJP0v6ObrfPDi4XDVo4Mb7njM3K5nxDMr6/XWHlp8oWufAJmHoU15bTMrgcm8
Kw/4lAMtVfxhtGCpGeAjAKcbVmM/Ctd/gODGBmnRhPhU6/0mdeaqJz1ND2ZP2YttGCQFqeBsqGzy
QwmedZlVMxQwV/Y88HA+2in/quK6AHJKCTdQ2GIBbpQbAFHlkx87zUX/dgo3PdEgPu/eb578/3ey
asWakrt7iIJJ3amtJWBmXwOUYXJ3TsojBZcEtKX96K/fjLNS+g1lIMdg/VhdJz3/x81fuWLB/6HS
6Uje3WHtV9/AIB/G713+YRQkpKlopuqseZqVGUbQI1sy8NTglwnhuSoGcL+DxvMiRCppIvUKpP/b
rBJexwmrthk/vwau7DVGy5uoD3gQBjzLWc6kr7GQT+wH48XSraUP41GvoROxODWUNIABJHwMNdeg
iKp5ail6/ekwGHxY+hKVmVXnVKOydfJOn6aEy1cCKnJxVQ3LmZtVPbrEl9fya8y7zi+uayYIpdpd
lx941u+EfvTPvlQUnzX/HLRHpGMJSbmc9eiB0voH29R17vmu/NX2voUc/c2mFIp8n+4ei2ZGK9rK
P0ZYjpqwcyrHDOI1Z+MDF/uxqpSp6K5t3EcHcV0eIX9eYZ+GjcoxgYQQFYNcHepDGZe9Xny0rqOx
+R6cxwNnkuvofNPQLwdygvhnbiRby9SaiSNtR8M8nBlPtcSeT85bJkpmtHly9Uh8/NQ+o29EcdTi
nnZ/na0/g0duCHLstL3p9b5BH2w5HYh6YxRrIOVjBqvdkvc9/rRl8v0J2R6ROaO70pjRjCD7q/SX
heD2zBFTnAetAm7cZO8hCtg11acuXj6a9oGHOiVqzmB8fnD1bPipFJqbjvDHGqhbaUk1kL5OUwMS
CVVtwkV9udz6MJKN5xroLlc6jdYZcilXnab6udXHZfYSZ02jSe+ZdFTjdxxUVsCiip6ORDkavFWD
A2ERANjG+3/VxldpGc6C8NkCS59dSN8yGZUw5XWsUSYmu0uf24XmfQ8qJ0saqGq7ADS2JIV+EMYT
gUVbAUvcuswErIRiesM4RRrkq7bJj1lmusyKcADyf1yYbMF8qWVg/8c9t2Q7ZzIUeQ2lbn+wJLEW
l+BQA4JFesWqBMRUIrRNg9KEE28nbMeoM/0nzPFEUOUdtnCeBoA+cZVd5QmRSi69jFsJVbyoISw1
67yZYZ1tpuBGN2hwjCe9ghB40rOnOpb0Qr7hlxyHMboyjzf9iMeNVUBLJ/9h7vIb9zW29XPfIZLN
ZyH0n6BM79XAcOzmQLIkzOzu+LxCEDqPuAZEKQIj0Gm2inwewCJNyQGrHt0HtnYRH9KYe6CkiuDs
0meEKq+ZFGoceaTqeAD3oWHAzOGquS46spe2lQ9Z+OKMTrdYyikQGpMoW09J/Tpvb5/VSM2Kcbky
WBPekF0Nyu8tU4prrukZHY8KeJdvPpOSA7GMHqTB6Hx/4EThbteRmAyAKTeUHF/grQ0OgcX1F6hn
FF9XdY8PAQH2GpeLruYvkx0Io23Yv7DSWga6A5A/HVOOLjTghOORdzFTqY0XFHU8Ew+O+Wc2pxJt
4WsTB8pEjuXFJQbWwhAgSDPRmPJr56i+R+mLRPNyxOXrmuuDfuumRorrKNCJzq+nMIu52+GIcUT6
NtzMza8ypxn20O2rRHgkjDM+MBuNA0CL1D82LJRu2ZuLHp9lRRvg8QW3+ChCJ9HjhkFw4tNZtSti
C3ARPyczM+39/vBaye0+lZjTj/RjVUct+EpnKc2IfZ+vq81Mn6tXgzBTP8vWzU9STn+f8EUFu/4V
IShXHnuz09WaWIdWxJId3wCS6nyq50QNAXa/i2IEEakRESi5VEOhJ8K7lZNJoPy1u6Sn1PX8C60W
cubHjion5i4mk/xzpoYrumOArsMFxFP907VMEugNnULR1z0D1i0RVRGsOujnBpObZCsZE+/nyhHP
W0ARcNmZh275in5hYXsb62a9EXysot7ApyNcdbYXK3hCdeEW3VohzdT9tWg8KZPc54ml1KOPDrzt
BalByktjst1e6WObT6Zu1VpNAluvtLZuHAGTp66it3w3gB7hK2cpazVfBu9I45qJV9dAa6/9vIic
vl13QgdX4pdk3qHkYrdeWd2iZrzbzhpFMu2ZYDQBnch8e3t/jllURKo9Xo2cq4Qb2UnBoVlsuzRn
vSRp03kECwrqEcpJ24/5FMjRhuYNCOvrDUodyN9PguJs4XGpP2E/J4gHo0wWcTVuAdT/oIMp9IzL
mz54j1hNgHrBREliZErMixyTPUkys/2pDC/dIWXJDkAL4hS1x7jL8oFl9lC/LVaPNiDnw2y/RPMV
0mNNENW5Tmlo99D6koIQAZI7Yds9Jsta0J//hGX6KP1pKgY5CAsVMANRVssB4t90chfmh8tkpsCn
9KZezT2ZUx4VdjXkEv+H/dN5Q4l5c5BPHkRIOsyzeEkcOjNspTTdBoj+dM2fOwW+hJT0kj8AaPgy
GseDnjG1fP8xleIsThmABwEqzgofZj4yocMHP0AEhVfoAJHqou7+ATvxz8VpPIWdKuEz1wtNHDge
y4GkPvXB8hezoG1zKRwAYzreZ8iaNi24ZzObP1DGbV7anvmrSDZuLglz+BDTzhPGkEj9wDt69N11
KyejpgXno9Gli9DJWHft2n1+KAA0DH+S6BECI2bk9uc8sLvyeWOYY5/R1ORNcNTudCj6yZQD1OFa
yhLpvXlEufbRt8GwAra880xMrRX3NveV/iR7uaQuKrGGmNVnZo4XO4dGUMQ6GV3lTsJb53ln3C4X
qmn6oKr+1UzcGtp+UvjtWlIb0U5PiVm9eySsHy7XQxz+nFomCIGbHJyhaviPLnoxyI+TwQkHfEjF
b0ksXXSKrl0XjKy6jNituodkOlA2YfxTtEpHWiyAGwRlOC0RaNeagL5yR0px5M7dJ8eaeBMEUtAw
+x6AooGmfhfKDNMw5RnnscbGFuLFrMrK1WfALmUZkMK6tjXJa0Wv/MUZCQiwFVgy8K0ZPQWM2CV+
jgSxiROHhooOIaAyiGNX+jziL+WrlCBzWkbWTM4pUcJxOKNn1ys4Pe/HCpKO878hhGsGV6eJtc59
f6MpRZJ/khmq6i67wKMfTc8Ksdq9+BYR8Vm7fc9hf7RplZFQaHt3ua4oy1/WF2en5ke8MqTPU17/
VoLIXisYef4ld4x82o6J21MByAHwppkJrrs3FkFZcVLniL7uXTG8mROqniOXhSpiTbxhpb1iglxL
bf4kTbN1SFIvFSynkwVsg1a9pKVqhYQPlYbmcLAolNzlguxPrVI4JfY+4gH/cF+QXEa36UvpckOY
EBaNIdiWGGGztwbkGMgbadCWAUQ6Pqvg0EEKQt0Au2yp81Hw2PRX0tsEIFevS6J/n0bljqXh9Qmb
4AZI36w0j2dbNr5RTwGy82iBm7Y1kl3na2OOt+FwLWaUdVo9jNDhLaYwtns3kT/EOwgmIyc/GeOJ
qWWlrtXkGruf0EcTtiSWu6jWzbX8vEvLkPCJSQK1o1073Y6rbB6WKsPpGxhwIoIOD8kkN/gPpT6u
8xdJDPz6oM25F1sS8J6A02gf/hc4Dv6+Fm2cXXvLqTmlVFTGiwLAm/8F7Pqu5zc6bD3QiOkpg2Oa
K41hesbOhu4fqHCR6rfTKgKeb6hqAtx2oTjD2pshzwDCRKbnFKkdn5uCIhTEGKRHwoZEiTIYcwPc
v5lQ0k4jUP+8iR28QjGP13l5wqrYMO0hy+6a9DhMLtP6284RaFy1ErXD+01DZQuPskqUExG6EAY2
w6VLzJXjQH02lNO9YLJU2SWhAgAWSgT9M4/1AkVNckqul0abSSC5bqrGVT6TX9acOnvETHUKE4r+
cKBVRbbHCVGYtJ5HWWxRxbNu73LjV2pxmAR70OkO4nR4jl12NLObZKhQoa33IPbVXaRABga0W/tJ
zXur9MEPxytG94rkiM3bSCU9Sn8v4/U+77KKpiWvmxvvjpdpg4MHP5JJaFkWnn619uiYFlIhJfZy
GfRnY6H8vJJtQu+xz1Q6u31i5YKCEIwye+qY5PM6feksClTyVZH48bVGgx5RCIIe4jpkWLk1VJBI
Q5oTXrhO/TNvXVJEOciAoJ19+fuX2bh1z6Rx8ijd/hx2MK4sOptKBjVi2ZG3LIaGX1zGr38mpZbC
O/HisMWcUZA2VRyOXCTKUyyewHU8mQ00DWK50nMN46GKzmwBwh344L1zqQnPCqAEbGriOzzM1lq9
DojQWi1V2arw7yqOXUs2E1CQJ48dPV1mIdUA0fWxERS6+IOiL0fNKVXVBLaSYooePnRkTvbyJmtu
GivJJZyWn0Nvvn7JdGt68irT0v+HHpOxZRs9i/8zMC1SFJzUa1tyIzyvRN/jGYdEy00y6CiQUbIC
3ufQ58gb/XCrplHilkWqTVMocnk8TakUyLu96DuyctmtazjXhuREGuUiu02VHcUtT1w8qs80qceF
alV2sKpL6dk6XGgo6RIF0T8zODGrPgfVoqO9O42UvSMsOT47Sah9NYLT952kxEshGByaZ3YSpQAl
vqXJtGEf2R8WNlwlpTWiECdH6tcfnHCkWxPGIpSuXUFgWP2PMfckBg0ZE3XQoMLziHR5AsTtBwBY
8IXirmhSKUeekegkgEK5xmwuRrelayTkA3MCSsAf6DnxMCpPZOMTknL8LiDitC1Aj3QbhNLgoC37
ahomX0XBduZNna679oiutTFWH8NbIfvpfE4fozsBGd2E0hLF6lKWwXwUTYwlag8hN5dNbNCTOKQw
pFYUe12ia+BxmODgdolSCF3HwJMhPoOpINae9EvGDfDE9rQJ2TY8XH9MSkxZVc3JGmwRWbIJpP+d
FDPziXZydUY20/fkXTNyAMEru6ydPglznx5lfFKOgYTaqoWnw534S4RbiFzYyiQ1NyTCOesB0Vtx
CwVQb3pDFbMfjwafYmTyUMJ6rGuHnt8/gFR0JLY9tu5y5hx8SLIaBf441reWULtb8aTfDoiMYkEC
w4fA5ITrThORN2EJm75huJDn64iSyXvWKIh9ydkiWjJZv8e9molEFcz427XajV/GbbmpdDNbdHtQ
R24UUGObmfwrCqy2yS64Mhfx7PyfKT9K7VwlvMESKFQXLesDgW6jEVSBkzD/5EwNJCIIXRQrHyiw
kOJcbAq2733uF7YNh7V1HoaL2cpY7A7kAycvIrbzinx9moQ+SyFXFJvXSkkEOQfzRPf1lBaRvCrl
sE+1wT8CHv3iEGBwVbHZodZSoXZ/uxKBeKphLjvRw+/bpEcC5O+oJ223AARVofabzxmJCSWF6uMN
/51rhxmsnHKvM5bJqEegKOxeSjCZJqL+f82yX5kBImDj+WDQd6lvfBjYChz2dFYanojowK7C2eAz
90DQ3MPaHLSM6hFTlH+oHI7BkQ7DKeMIG9KMFpXBWoo1eGFYfYK+DzPk02BN8FAbVC71BGIfQ7oW
vmgwDx+b7H1PtVkH6mNrvK4x08UfDC/F1YTKM95dbbYD8qvqYuKrfr04OmWJv80Mzn5BLf/QM9FR
6diGa5gLq0MMLA7StMBsu4mBeAwBI5aaoYdmVXcFpfoU64GyrUKjNjuTKIp7OM2m1x3UK1oOS/iM
PFJp2dL19aeZqpyP501U8PwkRur6axfpgeC1jAR3mqLYYH24++/fK5Awu0I+VGauXRWQYIuxdN8p
MJ8SbqAiucucPirTqhBuFnMMqmeqiCWnNN3uAR382tQF1kZk8L+VZImuOrD79ygmyno5Ml6nqVjW
Jxbvvd3zuwuLn0kAFAR4goWYK0w1PO2Dhyt42pUlLn8BDujiWbgINX6FQMXZ/eE3H9DAxXrvcgpn
DGq0e8nNyuUH5H7NIWH8wEb0YjPH8t5y11N9jSWTQ5/el4Aq0VYQ8dc3ABb3PE150PEilMpGOt0y
amZ1hyGmew3De4fFWllEBU8hpcoO19iRuYQLEoYlT2qOmNPB/JXcOeMhE/lk2gsRHUrB6uCKDdRI
pD/H8EkrX4TbnACtJ6Ygdyd5kqBvGTRZt/j69pN//Jqxqg/efKoxR92W6ywad2/j2MO5thhD68u1
KggiFpRygKrY2DZ/bReztUYiT1pLdz+NeanMWb4rloaYMtfVrb+5jOQJa7u5OJR1UY1fMyzNDY0X
/4OfIubZyqVtlC/YctdBAvkqaajqCmt1OoC81ndMtiL2zvKPptnwTwdQVLOoWJP9X+BDlor/z+Xm
GXwecOm1qkG79+jEjn3/J2rKhBbjIZC0oW60O9/bv7MmfmiCe+/BsYTKxe2xHgW2r16+RI73cSob
eHLnRXipgg6eJ/yTKt7+/8RgS1R7S2k12imVC+niAC/dQJu28V+12gbg3rVqlRrgeoCZxb3GisHG
UeNvB16vkpa+bII4F3LGVvT9tz3kFlvN+nv3738dtdX6awlrgM8LwREvmpqm/U4Fs+goV+hwi10s
qIML+reSsg+9PUY+7WQrZ4TqPNhmlJ1egCtVoENrH6dT7+b1QnA1jRSM95egy8oBTi9W+sVe4a3f
TCw+uVdC8/YVtHKuaZvYXznV8sC9LCF0hWs+1uXDEJjNARfq3ZmjFbI4mHD0eCA6E9Ol9Oo6cTPB
0xKpik4XnKxvhoKIVoYIqMMi+yPgtQoTn7Rfjcv+QY5D+9c4oWEEypT+DdIw3+ZpmfhHAKhIN5+S
HXKddV2QB50KFIzUlcV4UVujSprEORMoWDYeu3NTdj9CMqqZO3DA/aonUMZjqDQXYN+ZJeKpGm3y
AybzkJB4tDs4w/jHaZKDZKH6OIHwik2R2JZ9sw93zAMqaZA3A/d+zAqUVb04PKHtfsCxzJCVfLJx
WhM8JPH8S0bs769bTeOB/U8AqZn6UmXVMA8rX3arg6yoT6rDkYU1R0temU+6YSN6ez1d2s32Jm18
Bpx+pLXz2MpDeRjEvUctj/Mi0Fc6Aj4dkj5W5oriXtIYEupGhfCfrVFGsAQWmkroyr4wOpQ6kZ84
eigeLiZcE40ivXyulQxqd8zrMS7lT+xnUkBSgYvVreG5t92b4oFQq9Rdcp+u7RGMnrTuDgT6QHsx
h7bbGkZ0zDH0WWoFO9+n6tAzCfuvG3l2a0ylsW+TvimHMAlElYH1yfj0pXCepK1DbYrVGSHMtuar
Btj6ulhoeyAF6LjXRWftqH/L64BFL1tS+Ii8Kz9g8wk/kbDgdbMtenMfRvaxgDVORqvbb7Fs2goU
AeN2PPqywr+Askv8Ce8yASexGHTSxzwdRU0v3lMPfKjukM5Udh7+bqrUqMG8uhXRPdVqrqMk/fX4
smeKwit/4iGK93Sgn1wTnQGY+wt1H/tSmyATQF0aq5Ja11lUNn7vF7X4NPQTJV0rBEqaTD6R/F/W
Sr2dHMtYu4glfJ8sI7D9Uk9CTApRSWL2eHRxF0/okyeOTKS1/UK+qXCdZQFJ5iTJS6MXEMk/qNOS
7SWoxhYZI/TCotQQpkVbBWxrky5Or9G6815d1Hx20XpU/6v5nr/p+suFV53dBgiaqPsKaj51wP5X
i7mGPZCWMlEy7UEbZeaAxDfobNZ2uukdPRwgwTtdI8d+Hr23q3Gx90QRIUrbjxgz8QS5qA1bjgnu
Ad9rC/a/aKXMdF5EmOwwIl9kmmhVD6zUj3Zrvmd5PFTtEeya/hB0ofZUIgblTOz/TpeNMwXoGs/H
LXkTEa99dWzSknTYXjoLKiWfNx38uQp3D0QY28Y1rV8EWhTob9/iOq2NnB3PA1bezAYkWK1QaKEq
lq4ch07djmo3lxelUEDo3EPNaVsEIBos+PVTMnW/j1Doz1yT5axQRUzZScNVfNppyv//+p3mfpm6
lYPBkfZK1pDpq8fgyosl2WueUyY2JE/v8RW8f1lKwJxAz/Kvt5jX8s3oEiFzOpPE9ki477M+uBEO
ej+jVW3JDLmmWPFXx/1Uxg8wuHEdAeyInIGza+p0hkOAjP5oehdQWWDfMvYkbK6U0wR/V0DWcpec
HPu7ZISTfbu83fupGfD6Kqfscn2snD5ZZxgoG+c4e2kQydyobhYW0F924cxu6xo+qdAcWlyo+Zck
trCbrpGKK5/vqKEux6haGJgpLL+3DY1bzaR3QPDerML621InZ4675VamjYAypKMw4g470Q9E/iLJ
rVSpwg/Osiua6aVm9bldXJ1cdg4NPIo92h/fpEbY8B9jcEMZsWNYr7pZTfE2qCHPjBBvyhb9pElm
x2rmFElWDd1PbIQgk35RLtH3goiHNxoe2Tx2EGexhNAiFKp7riO9sBL96APn6vZxofTWn2gR5iL3
1D99OHsBf3QyWQxIqI4txJr0dI9UHX22nyIquuXMEQ9hdA4UDKh4is5pb0kBd94hkXC1BAieYHcQ
uDPogKrbQF6lQTCpmBZNic/QH0HTYfnvS+bEfCoy6BDFXQHhOGqyCnC9Q0OZGqf/v1OZ3zyswwOY
H0q/LdRL/eSr7wpzpL2qjI8w2ZgQZ/n+1GdGNTS1cOmHrBGjqn6TvzAmKJTkHJFLQeMFH+cnsek5
+ulFfX7x5TI6gM8ZCobafa2oiMS0cYve8vbS/A4Ejmdawpqg4sAuzICQuUlyYT9DqWN+qDrSmFwq
1vdBez95/JHzg8noXriGVzgsL3CeNH1lT7QoaLX6xMqd9sGrZWCra8LJS77+kRU8fBGP6vNXdEsc
5U+wJodw/7pyEansih6S8gGw1cZUNkeP7/PfY2Gi4aDjjCAFbqYwOL9nVO+ikU8kXcKdjM9odMZD
pGEorfgXIEpfaXmwIrxqMD3DCZJfOn7YCY/uhxUpFoCBy/ykdYb5ybAxbVwKO/pFf6K/HiOlZE9x
B2PQSW7opLjbFiiYpsplYO/yR9KsBu4zZbTucxBAvsl1JK6asugQly1XP+dvJ+9qEYgJG8J/QCIL
KPBPen4XHcFiFZhAnqEoAuHiWKiig3kHKj7D3HkL3RCVZjnZcNivvVZHZPsnlWCsgZ8Jq05G/xel
RD9g/r1osVYWdMGVB5SN61VQyndoJJUCAhbGJQNOzVSwe2QIWuKLYz8d0DqCV4LqAyeRXyUH/wUm
Y4cSfTYSQpdXe+eHEY61gg6ABtDdbQC8oi7j9wovuCnCwtzn0l+iBPfhl9U2SP8LWzlpeoOxnQ21
Wvv/NSI2NUDiUZ0En0wr493qHxg4MMHfvG+iPbdPhdwv8AD3GGU2u4LAFVDgLMkHQYrLncoBRANG
6j2Bdvv3gbI9A5ZhPCJ243RyklB+TmKFTIhGL9TAiZzsXFW4TVW8kgLoBxMfXBzUlesnr+s/XNA0
KhifR9pzlBf6JCUPYliqsnqIIvQs4nWQxG5ZaDcNDUq7tmIJlzK9U3Yy8gm2P/RvYz84TKi32h45
suL+EzdQT/K0Hkds+d5HkuqpIoCjHq8CQYbGEhTv4ikt87xzT1MqpiQ2Mzw8CTO/aYbGiUvEtQFp
NiOXcvAy5Wgx0At8qQgZxzPvWKqIbnVQnkrUuwPzbDVvWOF0kOmhaZGbM/xR0wpDfts4CGt0RmMs
SB/0u6zzKbzGonPd/YP/sRI19xZSezipgIpxyxAQNirmOjlBx5IqiPi0DBk8arv+RmdncOg+OWiJ
6zLCO0MkiO227J3zpe5wHCyva5sxpmSBu2YKVUc7hurmKZI5KqrBYJ9QDYl3ynCqfrCPclTrRr6R
fAMgZTursaIsNkCaHke6bLmyEt6b9YPFojTefsP+Z7Kqrh8dbl2Bo3J3RB8XP/WqzBRsuT6cWIQS
fXQmGIfD4ZmPum/pNBvZ82Al8oN0DUdSl1K4dhIb6uePeet6bje5UQdRACwIx3vsSdnnUoRRynuE
0jPviQ2OcXc5pCkPiOGeFOWQr3ehFwbJ+Vel5EjcW6NLM1kD3xz2YziJlj8PK4zh2Lt2KSOEUzqk
p8iOEZrN+2LOgb7rhUguIsqLe4y3rqtJaT92lfD63w6JMy6etu2MTecAcdMaraDoCNe361n0cdYK
t+zE5VfrCD+zJOTB8jId8UvKVgq4dltz+l1YoqJyKogsjgiYi7NHSAbtFw0AQIefYuXsEidvWoF3
lP7GjBRxzgxEnDQ6gQggJSjPjgfHXwhv+O0EYnQ3iXH54vBp66Mm48Ex1xLtQvxyz4gCZMYA0BGQ
PlRSKMNFMTWfiI+IafDquDbBKU9LEIoVAPhjnpS6+y+coH7S6O8Y5GghzDFrURtJCoSpGG/TpZcO
ghUESLJQCJ+X4ykPlDOQERvU3/GsuoaHuFQzgq+CtfuSeu1cgOdyROBInejJHNrOXm//+T/29xVu
aHt9kXqHnuZloAsykTV1wOpvh+gF0L4yYoZP1V2B1hxwYIsrcGdpi/gDUTL58kAAizmUv4HUM17R
7m1cH/LgpY8MajHnOwSi/a0UCBrR6NY442nugAnp5h4Urkwy2vhgs5wWhMw9njYAyfCgypxRsDpe
/DD468kDEo+Se6fCyQws0Z2W1yw1mGqYBarIiZjaJTcGWnHz8l8cB4kz9XBCSFNrQofvUm0JrYUG
oIE0cW8jhjOnU2Y8kpdLFeOTBbGBUrEmB3G64Lut9d9JVvESfTA8gx7aXSaVIfS16WAO4Vrsq/wx
Yv/QYcHgYCcsWbw95dul1BUY+Luglr1uBDUbbXMPaNiqhq/YEca65rXWPbv/vJAeNNMxZ8v+Aw7S
liT8MDZjyksDpHh3+tzws8e9jHUFRZswG4KI+nhOsAfCQ47La09ym7QOPCn5pleYT5nqIOUTG8YK
1yCW6tcIn9qGVVcE2yGST9kEl8Xo1NhG66iz3YW8ZAVC1VismYKzX/N+s4Vk7f+AKnD325TnodhV
eBQn2CVdHgseAGuifa49gokvJCO0wRFGoe2rRVYM2IGPpj4c00p7jQaazn8Q8ArfYx5hsZsq7Egt
4V4HNh4J1t/O8gA41qEpe7a3yNHdus3KpZGjnDG7HupKkNC/0iUcwTHfwFeSzUo1WblXD2QjQdcZ
tiyVbt279iOCl/7xkxnba9M0BAC+fCXqOLps43IXFmXwiZ1xc6A+2BsIIeH/r2Ga4xWILhicPbCn
oDKc+2SpqSk/G74WfdPgrY3cThR/LtNL05AMD0DAFSc08r0aTQznTLOf1HTa8B+EjUJxln8qHSQE
ZrqWpf5A1nSVx68rpEc3AXGQmiw5UiwBTpw8A7EcQuO8b+S7XiuZp3SnMtCnISTgIfL8oy2Z1UCn
j/N+uJ526j/4YyyIxrf63bUO89oXI5th3aPcrESKYuPqqzPfmMiD7QR0N+gCGKE3PKkqhNA507NS
vPH5GIxwMfrh9sFCvAZGHp0HqZxpv4s1GP6fMcv4sauiWehOOvQ/2XQOV5TiS6POYjf5Bqi0hkjN
V5n5iu4YpeAv6xsH/g6I9S8iOtKMbi2ZNE6FRjUCI1oZAFfUqn2Am4pixXKSEmnyZyf4ZUnGnMic
HIRSJBIHUr4S2eYFvbirjfwSSzwBS5SQ15i1Z4DirYQ9qaqvFqGEUOKN5s5Nx96htDHssjkUTYSQ
JuOwxTWg0Ts/v3eKHhqEb/Pdvg1i4LIgO1pFt5nHJ1xSl0NcYpUx3JwwM9iRd8PLEx2bcYFS6O8k
rp5+Aod8HkNrHU4cLu0E822K+KikZzCT4MDTweREz1OF0HkKETCQ9Fgx6NkUdauo3zsy9KKw9rEy
G7cd3GbNQyfm01Mx0W65bULijzLAlAVkm3Ymudo2g3zoNIe+jrsztUlTEQ6fU3EyMBLOXUFBIc4s
oPxkM2ITXx5zCZFaulCrbe9r30kYFswhFo+ECUMuMkZrxmkmUs2Q+i2D7uSjqdPEI1nRP8vGEvHL
qtscPnsjdoVMGp5rGHF/vcCpvCZS1O8mUQC6VMhJNBQpfOt2YUiTArgofwskUTBuYjFIx28i7dbq
PHOrimH/picoAI0sIWp1UO1wYD/Pa8qjPpDJ2YQWI1vWX2FZ3SQIyqwpo4BiIwnhvU37e8U8S0L3
0VmxD3NUUSkBd5zPucq+m7BxCQzwYoNeBGvCSbhkAT6G4bBtIRp8oe2l2bwZ+Mv/a+bcDp0UgyUM
Qm0B1Q0XiYmqpdxtVgWD4c8N4Yl99Vx9Kzck5MfOEb1UBpaz20kF7nLTglZL7M5eI1WlFFFQplx2
q1fWqaO+4iGXSevM1u8pqPiknQUPXEQ+Sk9c7GxhL1OrXesIvNTvOtk9h0r99ERa6b7n6B7odQ4g
xIkClFmAf/Fwx6LoEf7rJ1eSZ3uk3kisL+ZEs4ZvTEMlbF585HclYwL+uJh9aAyZ5edP/3g8NjDx
4rtF76+1MZxOdKP9EhQhpI8cD3JVoeC4zdIvF7LNNFbJTgTScPvDMGF5UyanDF0Zf5cVdXbcy+Mc
4zMvg/sW84CLzuX1LFmR3mRt+rN+xmZXrmN2vS9M7/jhFPuNom79RIkSVkWdw0yma3xMabm1qyd2
e98eU4Wrv1D7IMjWep5eKycTEj0jKqaxnnVnqdeWhhhSFMA48OBwuYuAhYQq6v7Usw8fF+a8YuGz
L/9FmK02ez6ATQlCoz0kVUz/giVcyhMPHQHZH3nqXus3njP7TLIL/vMa7I9w1vbTJU8resYWWxnd
o66LID2HEhBLDiiPrceuzr3l/hui1zkWBNWDpD8OTbdkreUJAa2Igsvj9ugbEPwuYe+Bz2RhlIab
K8WlH/kQw0hlGLyMkFVhuKXbsyapBCePBlDA+RCqZs7xTYUID2F+SGhFTVNyyN8xWxQf1KGDOVRs
fyzmnmXXv9llkK2j2IKmpiKLqDdR89jS9E0UaRGQpKDmHsgymz9TTjqDX61lDOJz7417nV0p6n6z
lOQH0qwokqwMkjKp7M1HAsJRmY35Cq0egxfK3y74r5d8FOVEy4TJ7+Y6sen6W2Epeh86rf0YIfAx
Tk/NKYi6TZIEMZTN+PRtdRDFO7AUhh5iyEuUF0tCKV67RtxgVnZaMVEL6dLhihg+mIFindZrM6PF
ydI2xRUdDlP+mbKWwTOjF/+xxDpQrQKpbWYj6GgZBxo+RQcD5nzY/rnlCi8CbT9eVIcdU7Wig1oB
+bPzl5ylhThURteLCOFcNydicqs/eh2SxX+vOy4bSfoWhiOwKwA6NgUCV9qjXrOlcJn/74NyWLPs
WsXllouOTA1wDIRKpbtlbYfiL9N2jy+8XUMnamlr1NMzh27gfkrCFfrzLNqj7jGA/1E7ms5XNMvZ
WDYWd9KQk2TS4jcQDscy2OyRl4BXvTu+Txgs2zjtOC92/sogLglsDI3PUo8BpaqP2JiE5oeLSEEV
+anURXPDu+prdi86oOJ5iRhufp8+v+fPiViCBDKCwVALqgnz27rq8LEWsohVEGwKS4cXDl0CzsUE
TFtNtFqzlWG9NDagh81t8V4SPeQX5HCbGUf6rWpUsTGA2rxAMDpvx1/EmLXmt7MsNwkYuyJHQ0w2
lnBhsA+5S5pyMsIRslnbGytWARjPf3ntb8V1oMgzBI42UA5KOZMknP0JrFUv/7Y5iT+nvCKoGNrx
W4yO4yfyd+rg+ODHwNxsY6cwho06UZB0lB0H4mVcG34qf2jx5VRoe9me7hj7KFe+S4qKTABC+tRD
X+sfvsdR4rdr7PlO4bpssbR6ECd3Zj2UYhKGe6hFJLmeoANCGzZHjEE0AoS6fgaxlbyBm3r+GNpM
EfNC+sPpGSoxH7JRu4IdJkiYEFb09IUURyeoxQqkbD0kvUS6DeJkXCZ1u33EUbxQY4SsT4f5BfPw
CQNwLO2gaK6z9NWr9W0Jz0KZwMBiLdXmxSyoQDm5eQ13dbhvX0z7w+NaJZ0NIdEsr2ON6uVEQwQZ
wEmq6MaVDyz2SUWdC0l+R2NqLKRYya9mrYY81G/d7DBri85VSgUW9IDFxDcr9Kd1D+k/ylKqETbC
Mew0EQrgDn4EjGwmLV7bGgNY0JOQvv/yVl3d+zXSoqK82ceSzmo97kUPaEphoteSMnOuBjxgnsKc
BTCdL9J/VOByGI8Iww/KlOVrbwVfpzMfleh1JcpP9LEILSlgUhwS+VdG+GIXK8XPS0r1m9taLWgh
nTaRitExWE921nb6+VaPQP68Kt7HAtzm7TIdzsFqjCKccWWECNZgr+cww+Z+ywUIIR+skg5ujWiA
7NFTudQfaK8O13UXfTwp20bOeKHrAAbVjALeZWfiB0t4NYo2G+1ftF6CGzuY58ofNQ02ctyJFtie
S3WTR0u6u6o52O7hJ9orlSE5CuXurP00lpbBBWZcfKQrIlRkdsIM0dLEK8Tgnmq6zjco/J+dxT2h
R0Tx/5pUqJF2t3e1W9ENoA/lMJCLgihXLEfeOOeET3tManNQKAGizIXW4UyW6612PudJCEUVSC2H
+8S6J0N4JZbX7WTbD4tRroMu96JHx/Se50PqtP2YceIsj5ez5CcG5jhpYl24n1P+CKc0sIEQtiTU
GkuaeQdpG64lY0wLWtQvcgdagSEgIer9ADBVxvr0wfCgXAUoSn70TVhX4DE1fmy7wFkI5OVGeLBb
N0bYinzMmP7Xq/pf99jDefqDfvXiGhW6m789iAt+j55vgPBm50brX6MXVVLlo2h+A1KuFIbsoyqF
ta/f3xkLq7n8fGdsufl9OsjeV7zEik1o3bclqnOP3wbc+xC/BD4aKeBro2+z0ZBhbUx9beu+/6o5
T4DvRgJJfNti5qj2LtKjJNmR+1py0hneyMgM4OMcYRJWV4hO3rfUkehZJWWoj4MOyKwFFmwwTtPy
aSW3zTeDze/Eta0NxBbrybQ3XTKBTZP3V5TANnj8oeFLxcRNDJPYW6FGwPnQC91FRoNU1HOUSd8N
rv+nFOvWgTisYCtThBKT4AdWzoTwim7/g9zvud3up0/l3o3navYO2I//9prIf1DCbP/inNx8rTNU
swMOZ8DVrPU6uoVxCJ8nxZCUdLEY5WCDD4RdwGRLccN8r/VZFM86qiGurPZUF80jQVLU12d3YYLD
KW7+RNZQA2Ja0rOH/wPLf8IJtAfKEDOMjuC4XnQOVusqQrjRRfTyGMgp2r014L5Gj+9B1Ham+OPk
ofWgvQd/ZumUX1xuBvh7uPYdmAwXCElLM2PLhwsR880l28sm15Xh0uCjHvkuxbhGUE/1aZJltejH
dduw0iceU5KbPcy2stj0Rg00/akYymGVHMz/4nuCTAGC/4l87+f7stqO6orLu7yhW2ERvn+9iG8R
eY/ogwTQvu1Zd/m1VgQ+tVSkYiBEGWvLkTcLewQ8rdTqz9Lsajpwas80lPtCIFHRQFXk8AYVsCRb
XWcXBCAFjAQWJTa/3U3C6u3ZuYXgdaM2ESixrRyNWkhczHI7jROrCDBUESe+y9UKr6eq+SOHF0Y0
yh+AtX/CpcckmTnM0jNJtwSrGJDorB4lg264yLcTHO1XH6mYSayw7rsA3lfoajftwry1thf4A5K9
3NGOrHB3Evs2rgYxFJtUlwM+dwdmwfOZRo7PR5Gh/LCnyA30V8w5oRR8jX9DgESwH0Os8XajW4ud
DUxqGjEQqMYrGpx/jwGpf1UurAR+/8ShiOx/jbNvpz0Mk+F9QuVHNVlcsSBc7g0m1pv57SVxrkxw
9YMlV2zRe9xTfQz0pKKskQlpcrLzfk9qjfkyFAsp2NqjssTdARuwIt6Na2gCulPHeafKGXQABnw9
kKcYS6jy1/BuAD+vLnpl+JuPyLW7546OziMoXxB2Bl5g7uwLC6znBfUuke4U64Kcf7fqzGhLwW04
Pq/ekzzAIYE1WtG6R/swhsaIFr0orRnAmblMMkUw0A5doywVfbHeLqccue7H5jL/BgylteDlBFZT
AgA+/iOd3u7P+4SodMadO57FOaRDBe7JiWKvGtDOAsG2YLjcAZhR7TQPW3NaK0WB3275uJXRiapS
62QJgHZ6nL7UJ1HhEHU/ON68zlrpY7ixmMtN1qmDCm5g501+GZne0rnfilCU+y5iSJihP4Zipyli
qwEcftzP2t56+FXVw+Pncsze0jS5D7r6IAj0TWQ4VxlxqBolp7MgjPFox/zx79k4tI5+A4Gm0mqr
nRniaGKk/T9Dg35AEkeIpTLAC9jQ9GJe0PsBJanbMSL7jHWrIi6CTFfEN2Lq5gRwiGXqU9ow6qSv
WytsJz245Ygrm9BjLF0jhdpqYKPEnycF4ajbj68uN8HTiKLm2g9DtDWaiV6E+j5nm8D9kPNx/DKu
YusS2bb1ZHuk/TAfysJ2mmELFBvnntegzLoYCQ70eSywvSHvLuBu6z1smNCzR0WWvRjEkf6+x93F
i5J/DnzGP1WPmzuVyi0ktuqwlcoQ/qisvGYW5DKUX5tj/lrYAptCJQIVyTFDot/lBIG/Yp+juoWl
E8K/qSV7IrfVHU3K3IJGg57ZZYXZlBmq8H0F9BffB5tEtN9yMsG2QxtA8LsptBE6K+pAszxI5frb
PgBabwhO8CEvvuhlvODNqOKmqph7YSyTyiH/9Qr+SAAb4BKKA+nJ/6YUkTAEzqMaXZL1UPCBPBJl
nKFNoKemQIxnMb0nFyIfGWsMJzz9FWNhXrYxD0Mp3n3f4a+y1t/BYwu3tbiLMPL06XdIzls+XwqN
oJnbNALu5i8Kcn4rVy3ie1EXwpBaWv6HSKzWZ1B+ArLAZAMpmp7EEQbMhdYX1bUWiIuSrAfbLGO9
YK2eYv++jW3Tv+JlSmQ4IdiGS3k4jp493G/h0VDGWjWgibeCPqpvsj4DSf9m+hEE3jVqKGHgshXs
96ZoPgxeFt8C7xfbNkqrtM47VbWPE7MLmkoZX46RujIgEvlWLnXlB2EpCR5dWvhDt9k2r9nNjhZF
jBPVt+hbCwUz6Tgg/ATF5bqTIGV+OAGu9XIrmDVti3L1cpL6F+hOHvT0aWMr4uuA1lL3Rs6VXEMH
alEe/+9IG6sZCAIOn4ufOVtX77mFk4QChttye+oOmzr/ZkxYA0nOinviHgzfOwyZv6y8ueqks0bz
eCZ5WbUsq6ujAxaUN2BuaeC1ap1jpO7p4xjF6euG9Y2//8X1L2S2A96FMTuNk/NPgBaw/zBBcP33
N8HHDvmVDvW03GmuaaB7yE7DGpj9mreJcKJqJYIGpOUAxeGAm02qXRXYAd2pr39dap7SydiLj73r
KrtEppnW+NindOW4192RBdrC/yHWNCAkTvmBMZrJ3gfN2DL2PydrjM5HyZMcWjQIfvswIZ2p9Uru
KSac3FvpbOvTP77EcIfVKYWUswE0a7gWY9TDfNx3yBQTpuTy5GW6VqOlEsk+Cz/3wHhLRGL8xzlq
IwRHRO1AKo1R/zKlUeeoEg0/eT8T1BI+6Ue5K/IAINikQ4lNvT0Un/m1p8GGUYSsDyIFEJ3y3Ops
2MKy1ffIL53Ic2d9dF2n7OkCkFIzoaGrmPDDIpnBhqYxPGykGP49as0SWgNdo7juY7YD1HHfq6Mh
4OXpYkVrcTvijDWg3sh5OIsxY0n9LfLJWLF9CMmMGqOiUuorc7rV1XQ4R3C6GwbRLq5rAP1uwYCG
4OhqFCbfZdRi9CCMH6HYuPxm1flJfWJ4u8cB2wqzs5twJZb+xF/Lr0G/12LBPFotzcBHO7RL/LyD
P1lLavj5wMEzJReiXm/bpOk25EKycYfwMXE2pFhCjTOdXZaHY8JVTOxWGbTjV/Cs9AaQWXd+1MUf
/P6ut9/X1xr44r1ShboHeG0QVXR5hBTVvc69OydwKf859Z01vdxdz+ugrw/KWsUkMghGG3KQtPFD
Yncdfbkv4OI8PY28S6uw/MvNKOOOuuxl2zNm9NiCLSMIPN5UG3+GcG1hh1yoUFOb37mU6bBNuqLU
8f5R191zNOLW2YxeKSvmrletJQvdjS42MCnvc462hLG2r8czqavWNwHu80gb3x8hQn3fFNPYx0cd
qnLWpNIKapRtzOiH9B8kwB5aZiVLObWZBF16DMFLtjXu/er54yGr6k8C+ubmObGNzVJqYNJ3075A
v3Z83rSe/lvQggYpI/Edb0brrJpSsHFg3Ozbd6+pbRu7pCzBWgjmFi/kovosEWhP5zrwc0s9QcWy
caarQfvS2PBkOzoRu8kRNhGVwI77Lnl6NG7pgjVqvpUx//F5lowP3PtZcUFF9O2+XpUWiK9r2kPF
aTVUbxfR8mLTlBNYNokha33PSPLYgrsZ54CwtFljLjL5LifSN4gNVtZuLcxmU0Cj0yxVqxLX7mxJ
7zsu+VrSUyehoH1uTas/BkVjkF4mYJSBvt9+UH3ApwPE6h/y3BuJtpQnAADGPnww9W7/68pJjVbB
rRb3zAoxNV6AeBFhuBBzT6VEVd0nCA4G4/e+0D9I4S+rv8lvLGWII8/konPcHkwMB3Z4LJQ2OZfI
tC9M1jUG7wMfbS+z4KFd7wRN9+DCfjBmefDKGU40jl8MUlvH6JflZKIhCAr2aSuq7ZEx3EupVbsB
VYFTgAcm8ATManseVj4y0xgly8SJ+aSSkVXjjfjSysfOpEd5e3tAc9jZffoKrw1Hs4k7XsybjOtK
WKGQrJEMTHY45FpRUWXZ+NERZArqhqINeBKKXkPbnAY6Xz5GrpkHdq7Rqb2SZnbuNpU9kRwNdiTh
VGX+zpQOFLfqyq2ku2zXZEytRgWspI207ZcwHjeB2dnI3ErfPfM/jamCSBHPaE6AyDbeuX2HeGL7
2v3kmB4vEOD7HAnwjWiIVFSPYCvJn9fmtb+TUr6CAi4NZTJkyu7+2/6E4PZ7ljmVIL4PAPgvyZ+8
ewRxVpahcVJ/dmipGnZBmOco5iN9qSLfvjeMN2s+n/dlJ7KTIV3PqhllweyUvGgGh3igKPB5Xc2N
1HS9vw3b2AtbZoTN6WD54CUj/ibKwkghgYjYp4gTkDdFDoFOxge6fmKBhwdte9VUJeJHAv+Cy/Sd
3PxhGyRuzrWXxhEBo/9WBKZe4Q18YhSZFWW0KZu1U1abeKlBZqAiFOAwnJI95o7+x/S/blGC+tI/
EzvXjjTRZ9h3QoEjLPyGSi9DJmcojnMSAYpLQLxUgEYF+ojBlE3Ykk2PBqPdZMiGxoxNehYIA92+
Es4GdwW45VYeDSykvwL6/VdVqzPxnGEpGBowI6N4QVNDMV//Tj7NYgvUuyQfHnCARNd3B4p9gld4
NmliL6sh6E0+H+fTxXYIifDgWpFv7SbnK/PMrz3m9qux5pPictrD6chdb0+knjzn64iRXvj+Jrx+
Sv8Lgi7/iEcI4V+VOLithd0ocTnhk/X7KTchq3RafqFwsfg+ePpC9nekLeTUk6nfS+nkjqP4s/u1
iMTvDHka5FFLl6Z6EaJ8+g6oFz88qRme4kFrowGvfnURypQXj35RC5LU/T8jlAsaIA3OcUHONrPy
a1uXhRu/piJ3UWCAZ+JTGMG0j0qG07B0Yu4=
`protect end_protected
