`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CLCBHAuc+dbUh2KYCY67nZ5R3MDfXtDmN8o6zwcJ+k/MzWKT9Mu7pPqRGBzjjBPYGxBIygSXMapd
oM5roEOQsA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
akeU+KrNRdfNTy4kHUzMZNOeQ2/eOfTIGdgYitSLoRnC9uGN+knsi/FaHDaKIewKj20dGo0fkTCx
iX4MCK/weHz2384VjrOampwhnof537TfGD9S7847QxV8RLY6V2dfcdXkX3WZ5pXT6YpkIkI0S6UB
HFl6E7669iXKKjSFoyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
npaVwhKFqiavxpGlw8qFymh/PlHxrfqyj3Axe9+juyTtVHtz04uvO9OinYWbumwdsVI3DBOu6/d0
AvUN/4ABCKcNTaS01pgzwapIzmoeeXHoK5EuKfEDKGT7/tKMh8+vl2kvLlcJawrUuSc4Z9OPaoUG
/pQF94K2EPXHSXU5x92OkqOV6U5o+LsW6YXD8VVzdX/kdRziPVEp63PgnFQk4aeOd/MT2a3/j+E2
OpDPcztTlhYQJfMdP6UTD/+aJr/6EOlenZikw5AmKdG9O1q5WB723CRVjzHj8CweWmnxnkWeJF0d
ZcWspJg2RM/rfw5NKe9Mdo8TM59Zv7armLzqLw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4aiAC6lb7G71A6+/PbJHXYFCRTKQe6Z9vQkNLZYUKQqDv1wYzNqtMOCsOOzXZFwaCEKT2j+21P4o
+SVoZ17kmG5dLCN9KrXT4XExOFRFJsD7TsbxYhGbE2RsIAV4Wj6IP8Q/XvRjji1u8tqLDfgo0t4k
c6hvPuqBVcwwq5llf3U=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
s9uQue/YFFudGFIKvsfAu4Ky1VZBhkOGha354nzdkwgpbtkk21V4FAGja02MhKduuPzCYj1F+xA3
g75IsuYSNvSuzfijUIORg1kX7M1m2tUdqjkff5FKQ8ZCvvddpXEiBGTvWgT5L/OD1gfq+/ThJzx2
NCsFYGCgrecOKjgCXQypvBIi9EykWmsbiTedUh0Iqf8KUrdr8W6svBjmgEogo9AVRwLtlqIK9GFP
1xKdjJBy+iUbQqojoTtjjCF0LS1EXLUF29iDCA4wjs1XXvZO3rRKoZdEbwFlbLL+EnabCrUgGbp4
fnrUGTemqESB/hStRpCt2ZoL+FUNokf+pGjP6g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 89616)
`protect data_block
3F/F2HAP3OFI8Ex4YwnAz7h7m/AmJpAVwP9PiICioKEcUaXIqZ7Z2yUZY5QeWaEqoLeLfYiTQ1BI
dRo/+Fq8uiXaKYQrtSSEKRC6l1+TuWM8w8n5zLh07WngpHmjYHAJ384udCirfCmCI+4f6BQjMTSo
y2ZnF2g4aLLKqtoFqytc32/bCt8TgBezHA/PstWmOKY4D5Jvrb1qMvkaYsRF7nK2C6XY95ngzA2E
uUVjKLHIF8rnfBqtku/x7WQ38AYm6AVax84coOmc8ntxf02hSr4U1LWxDx7ktH1PaUsE0ZfKglDi
qOGHiv5gIa/nDoZMvVkzgCQc4s57MiaXG+ZAUrNBLfYqlnTcI0vKtcSv+MuYKZ/PLhsqCOV2171o
JjOcL3gKHbDcwGbU8YdJ7dLHFCIv5ja5Aze2qfy4HR9Ds4asFyPgDGTpe62Fh3fGg7DJH3ltLr19
OWUxVbzt3/8K1lL0aDCdBaNoMFNblNqO6OmUaNY1yu1jvnW/BDIN7r+uhXm0qIzO282H+so5iW9H
mEPmoD1pTJmloBdEQsO1jZkiOyDQAErCTnCGxDgO46t/OQEKAAhI/9+fjoQED7ynF+RvZ2hr314g
Vs1Nurr23TdGaPnmHDABSJu4plv+Q4OV9KxXMYJLskak9EpQ+RWnidkeZCJ78+ETIBmKpmWshf74
bExmadzv2dUz2EqIwPM+As7hWJcddT6s1g70e4GHdKCfRGzs9ETeAXBJqYx1Oz6sQuh0eNCj2FNG
uDIT8Z0OhV5bhtlSrMRZ/Wd2hpBCi+fraOrtwNkm5AfBiGalyk3fxrl+ajVEjJrn6EI1r+/OTexn
WfPyMshcyDbNd0aaWAzVi0Ty8uv/+itfqTSDcCZwppNs1TE3pz8rcnPpTW+RM8q+0AUqSdW691JR
p5GRtx7cjra+DP5HVUFpTaBEis77XZGnGQVmUsPRVN1+1EshteXTbmpAv6JHJoyV2Yl3KPVIR6IF
+umrNgKGCg9XQuD1OMsSJnqqj2Tw9xOyC1cbP/lbKxrlEK+PdeBahkAETQZJ8w7JrdGfVqn/pgY7
ECp8ZeW/hhB5g9zm5X2UHmD8FyIMdFjY8BeK5+tMlJRN1b4WAsFLGml4zcgUIZBf7jGJjBTDwoXd
vu2WhbYm8oPouxwRDoLd+3VHgl3Qy7jw2fYeJF+Q7ov+nihernBwlHVpRHNvQQ01UU7T+Hi5L7gm
Po+2+6+/nfSytbzzFmhQN51TnFBm67GPm7Cuf8RuxQ+eBWlCQq4yLqzBqxZLflU9ca8ResCCBumt
IJB/7KZuD/kiKuZROkXQgKuBVaES2XSHV0SkxhzCspRgc+GadLTEWdErSnL86qyjJoFpJego/I6u
6cdAh/XAX8fGKOWbjuRefqCroA9EJnPjRpRp1YUy3kNVyBraIzf2PJlgtugzpS6h837HJ2hr9DO9
vuKO7aA6tyvA7IilIN9JK3EsMFgpUA3GFYfZEieqcY+/3bmbpfYBdxlt/3UWLhVd/jFYRU6i87Np
cwI/cRPIpe1hkClN2a7e0hfaopDPvFrXoPpIRvimr64r/PQw9XpixfCBc17fve1tYGNqiRx9MuC7
eyCrSEaDOH90bbfX+1t7ZyydZGYnaM1jris7nX6dX/FfrTojcAmbvkCt8LY6HOOb5/FZJHbxblCM
kJ15mDi9ehv/nrgmZSOfms0EjHcm7px9dXJK/1y3btEdyS//9fovAOsqgFQbmStP/oDJLo7i7vGU
kKeT81PHcbOAE+B4dUqJ3eC1uvobAOUoVJ6LXS6Z/seFmH2XTfUIgHsP38PuRB207Ih0aG6woLEP
PFWMoH8V9KLk7HodOG+S3fE0eRiMMjCrJG/Ghi1tCRVqmNYWwWTbvjzzncmu+B7dhrREMTvxozjS
Dy3W0JWnH5doQ/FpXtIIlcB869i9DgRIJ2hDGlCUzGT98B6KXSl+3w8nkGcVMtW2QZwKTJOocUme
ofP6OYk1W8b2kFXXixaRH30PZ7xV1lFye9T47l8XzngB2i+Bgx5FAQuoy4nI9uWClUN6dccGz4zy
BG68wGoSfONvxaDZfU2XZDYCDMMl/MH8Gf0PMUnySguu71JPm6i/EZYqKwNCfMc8eP/gObrHHKsP
WEB2MdaOubRYJZaMY+6sYZyZc9CihZFF65949rmS5WkssJqykgCx0kaGFgKjSMa3X0zOFiFCJihN
W/N1LTlucInB24KCkv4SJW6osw7Q8JYtOyAavjFGabsKUgZvX8NjgyYkwxTkKd3xcTJq0Gm+i5eS
GKaW+I468YyyqGRB9HQrtRyS/QDmmutozkY927KCmlnlqLBf8+2tduTsPqfX+A+PK0F3swpf6xAW
4D/yT1rm8yE0zYd8E3vB3Zy/mcMbIba2XqKUVVtZjjt4Pl5nOZvBA8EtzXx6N0lJy3nWr8PisgPY
o+PTuEbJr+gNaVMkXLry4DlW2V37fseK/ZE0bTFJ/eo8KKz9eGmavRuffRtINSjSBWqcCXv/Dfhd
Y33Q+VSofEjDeReoSk50L/dTDQtr4qQEE9SwYA5skb4WW3Bl1MKtI7RraXDsLxyBli32jN7O0T9j
V68haIofzLyj2T3LbSHnowVXuCZ9KYThS0dQneTfrMnXQpjGmpmpOG0X8iQT3NSlMeHL3+tQHRvR
nkhuY/0Yne7N3Z1Yc3Xj0DbzDvPhADjT0vFDGMNm8vCPza6t6l4++uCKUwakCMzkznNJ+VJIAXvd
I7v0BbLnzBipbLA2qXSwuKwZkswHHUmcCTVSgTJsyjzQX4DbTxRtzn0BZwdI5BAosTqq36GW94K1
a3gIK5A7gEIIIO4E3gPvC0II3mOwDxRidnsW4YP1d19kW0iTh5AsJQzqzO08NEvd/NBVoBj71zzj
LCxadFthoGfXxg9fodSrvITixES+OvK0bjQ+GInflP9TlNLk+Kcd/OGgqINhl/69LJI+O0xuQa5j
4jXJXQ9yBbMEL2V7ArCsGGlDbfEvWFfWcRYSq6AGp98aZNT5QHiWrJDlLfeqf8DBZVkgwLKmiIl7
0jVjY/Qma6eG6Q34tPYXm2wpxpUGXJAgToMbum+qIGEUOZvvZAnhPOViorP2dwHq6H8dbRRXbRhd
HX7iQFljFy/SnNLf2CQSdBVpL2iBMb2hk7QTkxE+BUt6YjgrxWgXcvHJVCeAzZfL8RIi6gFFd4+1
PYullEX40zfo9qxAHVFauj54xwxa0188O2nVnDYKQzQ/KbjPqigoRO7z+dY81MEhgSe3MRXAiav8
fy9noKcGddMfsrA7COicVC2/AfZPcZr0T5DtieC7HLc62Wzph6/QD0JkeR3avCLDEH7jKB0zSSII
Fs0pKVrQJCdHgrlYdslH2qPtamPU4gg+dDxFqyW3pYHGaERuLlj2EOHYggMMFql5nNonuVsAVqjT
A16ofvswXH0yq7eJELV8d951QgCe3Z2+DofgdssgMv9w0CWxHwaMgla4iUaqDvQltNLu6GEDTVbv
PQRMnNrkgxIKBPjsKmbkkSlu7Mi0LwJjnuEyKzBd+HlOjMfOA9n3ivV6eQpo2ur/NAAhvQwzUIGn
zHLxWrJaDnmzUyMsIEnGj4JTzk26uK+CZdyU3Pf+o/MLWChxzKA1t2adiyb2Cc7JKkSmHAJHRiz1
NDo+QDfuQ0jBOQFDcU+cPvRucVmdoHgI80JnUF6If2ppa1EY48ld2D7B9FAT23zcpK+yD5tbse0+
x61WhGwH1/gNEolJ7264Y9XEuPusUy4SlPypSeLlM1mVs56HzhiILhd8hHRYgR/5pqt5kDR8DCpJ
nkOAd4meXQJQwCObJ2nwoBHABa2kYuU33K66VFZ9fA3X5oQ92OFKNt8uJhTkqr0+1V4mA+KiY6kO
A4bDn01vPgcOlbo121Db8X4bWfE6cvDnRzP6XR9APi9heMw7Oz62jWS8ElRvpW6z39a58ZfePfJ1
re8sfVTL42LChuITyNgXGpkAHM7woEdYqooUnAku1bvBNWU2p2gl6+A3qaIVrzaGWWDi8+TxEwdw
ypBlLeNMDw0oF1rB/G+7LTU3zb1JZFl37lsABMtKJydf+wlUaerhO+LkLJsKxO6MX62NPX/XR730
9QHTpqYSscG2PeD1xPXF/M/ES5zKfmeZoydw+bTqvye2S2iLRwxVGTChd7VpyrrRO2QUyky99cTk
bwbu1hP8JVVj8AN9P3ExVeH0lFPJ+pbF3whD/L8mfKHk5qwDktG1Oy0ybCOIPd6RUTAR6gVfs9zT
IRYI0f4S9Dbtm+BWVIcMZJ3b6AZr77rXUZxWkJp8/cZqg3GfM04dPFcYfrqAL+x+q7s0Sue1KFWB
/3RmQv7k3dV+AKUQjOAHjkq8+VCu2NVakj6BpbnMJTCLvvWgBceY7Lq9HCQHNXVKqIECGoOWTH4S
8pCIkW2AzHkKwGhxV+qmcO3HY9/q51BbE3D+siVz8jBc0XRmMO3A57icrjQYtf1pLDr4yA3394At
J1+CrbfwOsr238X6Q6F0KVOosPk46wtqNc87D3CjgbqvgUvYXjjT8r7FkCEu5m+hwuV/4jD1VOS+
iX7AzERGrG3q7JssAPyDe4XbKTIBROdSHcJ4TcVeyMandsMklbKdM0U76XJVuBNlAsBrNxjr3VkJ
wkaNH825R8efa6tXhzs4boplxabRriT1qBikkArhn8PJ/HWN+DjaOWwmSBa7cEjIWlcWKXSt7udO
HVzmTMLA2vdfSpdLAQevp7ohPuWFPYe1hXTL0N1MK3a4cYNUFSTqTMr18IjwibIVdKoK7WG5Xtdg
Xynr2qPj5nHvqklA+dgGr5pKadyYu/LwyTZENp0JO/CCRQFWyzpiOyR1t0OO46UqUSe19XCrsMqk
WU8mZ0i/l0pBdJ6Dhklp6aScc7f8kl3Xq2HOmmTUQrNUu9Q4fFQobnhzTFvxR6AR+EjjE3K+AnbU
404G/5FxtSaq0rXCID/7gk8gZrCAth/g/67Cfsb0tuAVQRbwkzzVrb1P3s747ufi3xF4DrVAtNhv
+9l5zwkZ/0PdzcJsSpKwfshY0j2FKFqDBaeRjBpw6QavZrHyUH3IfdT4/1Ztm6yqQAELZCPxjxTZ
BlY/153+gPD2rGvSnWXFEUEQaY8gFvvqMz7TXlin+543PpK++ANco6Ia/gDkqj4DUymUcJcL9gv1
YX79SEe0p9TjaDGutf+1AwO321unb4prSkxxpFApnQ7xp13qnGuY5XaMoJg80iRtGUeziDTicJvX
UTxUsm84+IdmvwQtsg1bKb6X3p/mO90qcW+sH7QS9tVWSa4n869PMfXOr/B+15kBmeoJD4DfOoHz
FjdN+T03NMx+14EETYKgQCopSfzvyWk9+O/yvF+Q5Hgh8w0N5c/1yKzyZeFaEdJSg7GaIEpGCx0q
3T+V5X2Ny9j8xH+VLUDqcTHH6LR4cHG2v7U0WMp8XRoMAdhasiSzHIvQ6TZa6GPKLQGqJtkwpgcT
Y99iKo4IKWAwSfl/xVmAb79BHIIZNmgxfwcxCdp8sXZu0o5muq0d8iNOD7U40V13iCVgnwy3RG6u
cyk2M9yu1v1koPyWqECmQ5M+bTblc4hJC5D/amHiHMF52GuvTGlN/NOi6F/GGdJxlm2hqtZBsS0l
yLb0b9sTzMKdh9iB/F3HVRA4VduOSlOwl35sNkr3/yKnepK62aW0ZyhPNcfjg3aIvvEBDIhxV2W7
cDZ4P1AtNKde1bUcPUiI6cmgabsQ1YMX3EdHp2+2PQ5N0HWPnZRwmlNDcEcYBntEB/B2hWC3+9jp
xZZTzUjPOvRMtmw3Qami3RE12D2FvLt0X+A2zkKFCZtzz1UAYl2B1EwkoTj2/nOTtiZrVPzHXhqk
kZ7dUad5JO0k9sd1jmO/X4g4OZFO+78SprVdK5dJmXVtg9InCTyROv1BG0Z720cCmPceydzVikCy
PpZ4SJYStshhXxFY7bWUgToBMnJv26pqrctbFsrPbakzKSgmed1fICZ2U7JMOHf96geVcIUKZ+py
w3nijD2O12MVuDJYwXOrg1cODXMo3pqxLoEl4QKapVdoNvXDnIQW9uxxotHESEaBTBotL7rFJCes
RQR5pCysH14N8OVbR9bigOXh/1X7IvctoNwSZ/iXkHRBABGJlFuwSO9o/g9MQB7JjymCshEh1YMP
kDFiyzY4Zv5yR6r0n9Nby3ABwSLPsD/Qy8ezboJTYzgEY2FvWPtAsY8E/fQrK/uteBDr/boW5xZy
mazO9IZsbVhHXS5jlwbWwPncToNvVlO6ai51DxQTgZxQPNZ/0KK+cUQMb985U8o8Lg3yo2CHTY4q
kkTj62bpI5KNqEf2H7se8LODGSvcvPtWlg+PIn2WBRUEKwYfw38plqkURtH/4IYGAZnS82j/Txuf
FdBFx4lVbBeKJWmeDaYE1rScVJTXWQWEUocFDhRYzMUfRVGyhVX/yFbWRFSIGomQ8ZQJx1Hna88l
ijpip/0oIXOwJ1yHutpooqMiw0TRSEk2+2hDwOsyO2HtCP+G9jYh7lgVFmjFub620Pj+Zki4eq+j
bdjVovulTPmq2Jdi+Hsae7Qt26dZM/snR950J2bpz5MnL9Mgx2lbdVEYx1wXrQ+L2wypDiV+omBL
iPiOBE1+mkgCJMUIaJdf5D5zvLSpDt4mcEX7ebFWt9H8z2PSZJX2hpPW3i1zyW69ArqVyGKDt8y9
gHnDfa2SpeaxNDBQE/zIA/HUZZ7MzP+q0OTrpqJ5YQ2IO/9Z75A/nT3TAeI9NO+aFyv0DXm2b/NI
ZRPxQ2u4yd/vXZEMzw2ENYzBOM1QzKeo31a9zuko4NdKB+j41+FPfDZhiSWkNCtMEFu6ymiOIIR7
3dPVHiy9niUPvrlXGJOc9ovRbBEmDlfWGHPPIrWSPL0yYH1aZjJUHG/9Gf0pgbjl+8ytPyb4gRMS
x1Qkzo0vvNqhQc0hTi1rNp5iB5uRByUm+SJDvC45MQifqBxoEzx2+Mo+eoiJvjFQsEES/QyCXH1u
iKAY3+bbwJ+iSSWPJ6BsE8DU36vKtkMc/w6Sr33tvI0L9qne1FOhnG53oZzvTHt/kBeH2LqDUZag
QE13HPi0q04mfuz692AEN/NdWYgwvciNfbjr91F4ZzTsAU0ZdYalPpG9KxcGII3m9NuYs9m7MIE0
lHlh2tEQc5sQwTgnZMnj8yya1GA+90hQJG9RDIotL7Tmb2RyeQnLfg9OCRsYDuDRgZEy2WcXCWUb
vDTkg6jyNn1YaLgxvcQ1UazWisle+OhlIV5x2whDiqHjYUE+vNyJFZNa5VKZAYzbykB8pP9fd31g
9QVgbxWEYAT1x2pB07jk6RcGL0ajMLMUFYU03okB45w+264j++XdPBSJgHNaUxoUaQvQwl77/1P0
tZrUbCq/Z9zY6eK64iX2vtwDw+zILPl+HZW+77N/5nAHQvt+xM5VTvqe8O0/POVfXUrasbXG9OKw
SqoGIjjLoyUStTzulBDDTAGyXRDVCf4xxVmO8hzO5Y74H4TIEhZDrt21gUNjXcz7SYbGcXqB60mh
yl3pWVpU4TaIZWXfpgQs8yZrRPcTYQb95FbCe00KKasgP8EquIiOsA6Zhi4lPaFnnnf0v4bG0YOq
m31pJKYPunKaic6aFBK7ehZAjKjhYWVtjsSYx2aeqQ0wdfm4wzy2YV2qbytJ/LA+69xpyhtsAWUb
s71wYYN5ag48M1v8fuJtRpzvX1C58p2ucrdhf/s4CVGS8ghKxDROTdkBjOB1tN3D2FY4u0iV8N6H
nsnE9c5Lz/MYsNn9BEJYH1zQyCMcnnzrsNU2cz5q98y3isnVlRt8cWbaEneAOf79I71DMJV0/NuA
D2HKkgP4oSvXXnlTcc5zvw6WilqFBmndSfI9Sy7E/ei+KFrOxaHDKQORruBZCpwaTLFpZBVVtC5C
1v7wo63p9saM2o/WiTQTzU1kvK4VBExYYH5yOc1Oyk7cfIiKMiOURa6AylckjaSnBvkmZG02GKtP
fR4B+lRQTA3TrrVrCIK6qMFoTS5nxinRMxX8zn0P+94eLQLHqZRXS57FbPRrI10mNbM6owknbBiT
iMjJcAD2uNSqPQaPt1O6z23MJw0Myt7uVIf7PxJu3BLs85352JpwzS0xhNdD9ewLbnC4nlhIh9FH
kXKm+Z+rXfUMe90W2ANommdEuyRacPWIwiIFxFXxwj1aXUFZ1/boM/ysDb0ted2c9Ixp5LxqXEJb
4kEhA7P4dp0PnumpIMtYL/U/gf+URpL18HditIGfYz37ex3prbV7Z2WKvR4xY5hJ3JOTt2tInElr
KxoIwZZtzZ4F5TVscP3AHxuGE8LA5YldBP6eHRWoIRJ9u4KXB+MJGWBkmfeYWHpqC8hAtpQZAlZU
oUYb34Pv/JTWFAtCz58BsJa5OXmbSP9g9ARsqLqWpOA1SPgJre9KxpeNrg1fOEBc+ufNkilx/m7R
mgbhDgFkYEWgaiXQiNKrFqIEc+pH7QJjosw4Ix/P9Z2ttO1nCMd+C91DzAao627I3wjl5oWpDGlP
MWmnQCqMue75fhkXIPkq16pZOsmWs+ZW7goytzZyDnsl8jTJcpPsJExH1DgpzY3j77ZKPIgVhjhj
+doLO+vYie1ckH0dHg+iZKV0uOR4DR8jeBRGt1ZwjqlS1+a7VGK9dgc1jqEx0l4tlyLIt8H9UWS+
Fwe377S+9XpqbTb7ekOnWONVI7L0yfryxlbKqFk+cOXbiNVYJNiZmbeqOF7T1pPLC2xebDbhU9Z7
O0bJt13TKTc/E8JUaOwIStIbNcc8h3/ITfAWuTUH6yT4Kdbi6N+6PYLgZzVf/3ZmSWTajXNuTVNx
r0KGv9XtNRPu9IqjYS4jO41JWzST/J+Xed2BPw9cYXTafEUDSnUpxUiLHA5p6IgsKQDTmYX6/FVc
F8BIbLO9aE9X1K4plNMairiixUzWsAV/BbkiLEAyP0TLX4ltZejic9tNDmnOTBk1tz/6HyauVwjy
aCB4L9+eby75kiXeIaLoiYwrJLjF7uIn5tTAslbnLKFiK7SMhI2YkulqlLqIXGS07wU9l/dv8Vj8
OzWJzAuKkGgM/+OaU8TreOO+CUVu9QKqjDnKBSDH5FBvyV3uq7qfBtrIdVmmxJBB99DbI6tTB7+c
pzZEYtvLXZvHu9iOxRzD/kYYS7aS4+U8L7N7Zu67uayTAJPLdpPj1PFuCBXfQtFABlp7jDoFUAtg
RZnhH2JFp0sGTkvstUyFGTV7IwAlUe1xsmWWeQ6L4CjylydlUknbLmhHZanWum8vh4S+tgGRjlhw
/257MKBkTmNvyeKABnc5LzlPyrDfJ8tdAg+feplCm5zexE3OJ50I0yHETRCgvtjkgspgh2Kv5HzC
apjP0EbQRDgqwh/ta9/IvuTwvzHp6QQppGPnyeMnfBDgyRXwXsfs5iFjHiOMnJrbxUKzdDz1+rG7
2r0h3yKDWrS4sRF6ukMlzmdlh45EeGFAp+dY0wHD3iLoSC1qlVu8aZDCpiSWbvMC5PFiisFrlTPJ
S1wZSvK560ahMTnH0aaGY2NHom2iWQfoYOwV88InBObXsP1jJsuonP87P7YgdaLHzZa0WawzrRd9
7n/BvDOUSwt8QPEXBfTuBtrGnGM4X6iKspyTHCgFa7zVGaMRWGV3KayS5y8oPWDApES0wWJqN4wN
LxyUbzPdyelhKdc2WGmCJu8/MDEc3U2mTOux3iJ46m3KyWGWI8mrLnNB2vJjeU5lOabt5gtYT55K
F2QmbG/ljkZ7FF80K+Tz6eOjSS9Rgb8vIzmjEUp/Ai2HalayB8fOLnMfwz11cxnvyHndSyJq7N98
XTIPOq3itnOlDvjRTO7LrnxP81iYKLmTVr49KG00ufQ/iYuK9pkmXMF7oy73djiTXKXXiGu3SVRJ
tzAPKsDmovnDB7sOAPO8yIOIrDC7wnM7ck9Pbyr2jtj6CiDfLSUr46EWAKQXJWG6oP5gdvIwLCP/
jfWy+lEHtXwjNhLprkSARVz9wDfjXoMZb5PwzceKcfitZVBjbKqpODep8bk05Uy7gGjy753ND5ye
VA+bSm4nYdNRofcRi27exp68b0RmOqJIzuAxt0bRUVncZUXTDzvrBsYD+X4c9iiniSKkv6aNfYzE
TphC9WntNLXF3FAt1rnYQRVOWPUY7e5zK6rFpCRc5/6N6GBrMT6Hktlm5N1l2PF69c5VV+wtsi1v
SAmqI1s7jLeeWVLrW/37+7zeqfpfP/LyYY9XerMtqXDwbUpwFMaVi5eFQyBh4hnNKhWVHX/dJ269
4wzzh6nvoAtlrvvM7waSTAg36kpXOKOTbfSEM7wxeSiCrDKj7ISMVN6Y3jXyhrnoCLnT8yrnLysV
tYszfmIMJeG4Q/A7c0fy1D/43M4NzhAB+XNCSR7buyikbxFLdKWJue2ksMy7jOAZbn8CpfgghWIl
6Ek7ROuADVzDUgQLHqxbR10/yqThX4gBH6IRZjLlTmXUe+NhpFlA5JGu1JIjgrsCygdN9p2FMuLi
ViXhgzWxAmkseg94DFuq81qd7lEDce7w8kmiBNgoNqR2kmWtwufmXanxX6qz/ZBufW7LpUMIWnDH
kqTgpan0/M1MpQtwnwIUDlBbOxb4fl19CVlPCXgpEzq698/42802CIp29f7c00fjHAJdGZdNUNd5
VZ3wB2DU0Da+E4wxcIEUSsCV9C+oXDLmxM1pYYvMSMsVX9yDNC2rq81PhkORuVNdLSadFJW+JX+c
XHpLx4QHxWyLD5JOC6v5Qd02XMWIfnaz+7K2cg8Y/A1BxIzqT+TcSTTS+hwyQiUHeZiVei1MVHdx
cTgf9gbSh4y0dVm9/we7883PCurBPdUS3Bsm9yEtmyT88whXEc3FsggUoqN5l4796cGZ/K2yf+nl
G+W2fJGyh397w5QI+YiXUCjLCLHZcK4Y8w1mlNZ7HFKWlES+vH0ZEKjIeToE2kMPRmpoGcQ0PE/V
3Napo7LXfbb5P5ahScqXnC8EHBDNrEDM/bi1rFw5yXVWDu5lWn12En6Ecf9+8EW3ZowjoYfLtG1F
aq+j9uC9Fug9mbegbOGIqMMKwkbiilF+KSxN0tFf+5re0N6Ri1tUJHpA/0ViK+RC3OTpKJJgvds3
9zsphU1hufq9C28Eyz6w+YkLTK2WYZLzohZ5etkY/Z1aI1E8Pb2UKMc2vYkTZuvXRSwEv563LPAK
CZyELLARn4fcm7Wxf/t1yuYwldSnYkT5gxIMz18cq24muTlYKbDtbkK6mdMSN0bTDRiG2jJlZUPi
ENvry1TRAFM5/t0KW23CFgVANLTkgEeNoBBWEPivx5zOEBZRqJIIeWEG6xNCG+UMTlcBv5Q27959
/CIfANbahBspWkA8+XjihCabKmOm5m4oOym3qrAQxHtoEm/25yHNgY+Rb5kDo5nRrSu3r5QNjcGi
qWbKi+ipxDnKT1mFSCAmcUrmSM0NnnE2GGDwZ6ySEjvCaEWfLXgThxnWrl78kp142qoSKSfQsOEE
K5B1zznR+PhB+jRBZBbgNQcxOh2oRGFfKZCNRdbHB2Q/Kn5IPsyCgYRP2toq9KNByCYU3rUyzkoY
uSoJGB8L4EVr29Dr2b4+KrrY4707Atbn42V20YpKO9DaPdqwef3gmRVIDianTiRXUp/Uf5FOnn3P
FSzqNcQkhy3BlBFgsvlTpTwRR5YnaGazCjcV70b2g9rumEZsUXd+OJKBs0w654nwNZCPEeUl9JpA
a18dMkUmhOGoH4DPTLf6rtU9yZz+K7qwbPM9NHHYEG7+5B6Mf3iVPFqRZYmWtVr5r4Ed4vNCabjV
AAxt5FHUbhjyB0PWeVrt9kiuOtk/jmH0OjW/AlQ67GtR/z5d9VHAqK5vRFXwsKs54m5JPsKS6ie2
PZG50A1cKWbRwGN8EUTXEAlCfKPg5zJ2XSFu3Z5UROsNpg9esvH4VexJ53lrZf669Rm4tiN2w691
/JiZn93Veckfs1W01rU8OayQA0cRdg0eobRKuZ2WWvhFWfru/Qml1zyFQ3alj2jjEtvXjnAA8DG5
TdjNsNaV2nCbiIj0uwQJVveCjOckMBm7KtWPnmEzHOaJQEXLYcGmEjGebsuJXx3SUjygeMRTf1U+
J8ieSZJwxALNjyXZjrzEYU52DuRkZAkwwczFi9ubiLQCFjh/JNgVDDPyo30mYpcCxzkg4mhciGCh
rub7WWjJfF/PNn4PY9TpTUOwNgEdl0gB4EJAPVGeK0/BrH445UVU5ImcRf3y4gDb8zXlpd0E1MsH
qODjkT7BPdnhWTHGmWHpHB2IbrkNRK/Gt2HaQRKk3H30gnksi6ztRUz947KpjP2pGNLOnqeO1TDw
UiUZ9SCp2A6VUeCcGZa3gA0bRRpyJ35SVuCJdzVPdQUSl7RtVIgVTHbQJ66p5uKkOWpwlX17sZgp
tOE4QYQRE6m3kVbMXC9AFg1abV8zeJn3/tIPq7IAvn9pwlhhzOi9bUnBjEzXeXl+ETy0hkvf9eCm
Itbm8gXfNX5p7m6saBHidWY0qnrMSkpjFCkq5Rm+TmaF3AKUznmMIamQnQZYCTtKA7D2mW+hlfoJ
PHZBueWpGuhuM8l+owushw7ruydkchLH+jeGIu8inI467tAhFPz8wQV7uKFdrczU/S02X0Lcie82
xSD3UaTwLPu60yGBPiJouLnuW37wiFz9dvwAbhZ+7JcP1goGjZ6MOlfjD8pwTQ0gJOILlB04Ux0r
kjChIHz4bx1GhAJ5sRMofVbDgj3HxX0r2Y05pCFJQK9huydHJZ6j0qYffjECApKY8H3PN0kQHB1L
YOnpi2Gn7l+yg1LVXgSarFbNJ/MuwDo5cRPmyB7OSrCiWDfDYPNlqU3n1kUru0SHjz4qSTlTliDL
RE+ZeowrbZsX2sqomuefkGzdZw7QuycF2y9oPCFJu4C/lzMegyqIRN4UhfikbmRdO/ox8kvN8gan
f7fOGW9PhHJ33+37/PMGKqA8aGU1jpdHR5tPMDMoxkjCpE0CIgb1pmPsq6yhpn6VusBn6Cep6QVP
t+lE61LF/SuMrWVpJADUJ3EieSVD4xfEL5e4U6AjcdBxXe/YQOG06dNyNsJGnrMEfsTPUODcJhuP
9MCey3kbdqC57nuvv+wFxw9JJiZQF6iQWcwqgaRRd1oNHQaj77EtZahIBARqiEacZBKmuSUmDl8c
txs0av5kJIEh/kafAIe6Ao35ln943m9t6FxPkc5OWBFfkFkHrYKjwQv0gz5GnXkm5OqvojitbRx7
aWjTFKvk50zIBQubwCMLngyDlu4T6r4ZGY1YMAozwq/XG1nurI9Hy7PTyVrGksMNW/NKkkNmYFOj
CsEW0PNfKEMDjWeI6q0IHjP0oaZaCaI1VoJoYO+1ctgqhNMf6/dcI6nbnifsen2DKAz1xG2TIuEj
EGGUMJdwGBsMD7KIJbFET8exkzIR4AtFoNyx8EWUdd7/KQqdLlyiKMMURBCsHGac5J+mqYsglIVv
IGWsX41bDhpoAIbNm1T0fOH6KehPW4GnrA9QEcY3ha1yHttRd3CZuZtPH+m9qY08O2fFLnYeWNGs
GO8Z5uKGqgD/CySxfWk9tX0RgQa7x1FiGiSo9drogzRhZ1xB4frT64RDnHbLVpOg95oPcffQPWlG
QBPBu5Ky30VhNnKFQdXarsJOI8jiPG0Ofn9eRk1wk99Eajcw8vBAXya8wUOUAITZsQuPapNeqvBv
mM51Xr8oHSKKyALHXJ8912PE2k6qYG2ZsqiZ171h5ZcCHkaR45MvQYl+BHLXQypjP1Qy2VmTEIXi
LPWfijSYWwjzThyJxbnGB5yAHN+I2qxMRnAa41SJ45tQ8uIlVeMb6VvusrNQLPkJvhlG/3CmZFlC
KVkD9EirItFOIyV0ylDWSzYNCt8VuBHokX4jv9rMB+lDacdQsLRyz0hOpXh910/uJlc8jbze9YT0
wiqYhq08kI51Tsa/0rosqvoE7zgD4pY1B/1mgH7DxS8wBY8adg9jeP3wfnu9SmCUtwbW6LmWggEk
jE41tbMC2HX8qw7cbf68+pkLNIiJL6bKd2HavVrnn9dfQftNFVxZ9bAogx+SeN2uEx8sx3DBaU2w
um8BzRSn3KEbRoOBPD3AoxWJ9RCE9jTuUuE/x1Rz+px2/fi8Pv6qtBpRZaCDWhICmk2FioF606q9
21ky/UqcSokVgiDpmEpSPmoSu8d4s3qJ7Yr5Y93VdGU0UeWGMyhyU3OOXTxSYQ647rZ26yEHvj3Y
eIDIyx06hMs3SEGpd+OvcTuiBX0uCereKgDYULEEc5uicY/uCxCvo3e5WFFj78GvN5Qz+Ub8wfAm
3gKsNgFhcwcD9OaqwPSWr3HZVVPBPrf9738TKmwqsWJiAJtls7j9JPBSUHV4WM59hQT58hUx8d2+
ImyF4BQ8pwlz2U8bm3IqN+O0HNQS/ZpRTnD6bM528FDspaUOJKgrmK86YXsPosvDZpN84criVVE6
Py2aohGpxA6mbzgXCDhsgK3twxnEvq0o3VeU5BVGS9wfN15Wt+Uxv5fspQT8NSK/9bjjFUSKFduI
J9qFDX6PuHWgake/9g9iPrsuqNwxYyGFwp4eOm5xZLraDUKT5weDxGt+cotyfnncPNaZTazvoDt7
4YILPlcNxy4apD5xelSNblU6jAvd+P8u9eEu6uCnHyRJSR0q0aF1mq1N4Fj+StpaZ5elqwLcJ83x
Wgf1OvKA8VvhdQxABpOZoEg/J5V14Huowc1CMbvz6GJSti+Y/NF+nu8oFG6E6lZlAOrC8L1i+iQ+
gtwQf7svIXHUZMpKeCiWZBbLC8J8CA3s9ItbGW9jJl4RVl0vmnfY+PMdBCs9SwKSH1f6LwgNY0Zp
qBIL/toNoSZdRVc1xMTLb7RZnuAuRuCZY1Ud4PwRBCjqkz0FrlpPMaM5iNwDE1ZzPXYSRVZOcVMv
ASJnUqH+HBSpFdP9rfJMYLofGYNMmNzJeR8QCARkR7D66EfVtC91mYIH8fkz8nspaMVohFUiVO1/
B+b9/6B2rJHwOl/38G3s1QDhieiez/P7SjDUNt7ZfFUfRNa/m8ebLWOk792+d74ueef+6W9DMubx
uQlNeMzj4EF/2gwSy9ilLXBQVb4AQgAvnPLqEAK+YFEKpTt6MpLhZHavbM8KyxddPOvbZwO3DdiM
VruWOlQLhE1nEr4FKVdGrGYWGV6sOwprN8CIdykxqucjz41KHVJo6FwCRSzyhjLJdvSI9XEkNPzB
8qDR9Ion7gRvxT6krumPnz+Q6GF89fVAcamI3GuMGsthENNFb6tYXoK3JUfUCUvkhLKQJWUSUgam
nouNSj2uv35JwlwjZP8fCtu3I4DionmKxPrwCnsalFCQ6lu1ll+tSATLrEKgypOT2uvL6fZ5/V+x
JK4oYmrov7ypHWp7HlzaBkJMwIaNBUIiG6JkzkC/m0NA+rzbqRS3LCK+ZBt4QpvRq/TD+1tukHTd
b/JVpwuHEfZ2RtOow+xXbCrdNR0zBxvT7ilYfcSfYqCDXt63G/f1O+hq0jRE6hOwLw+JafvhIBbO
P8hY7eHnlpVUzOQz605fbhLgyjuvT5FqZrH/PO25fOrI+7+xiiJieP04cjmlORx7WfdZ2CCuhIqy
bDtFfwv/u42gA2ofOift34kaKmcq3YYqL5jFgrkPuOFFatlSMdxZwc/UuSTzx9mYFjWfexoInXE+
a3mJ9e0UFqVYd3jsT8xja49ITZier1SQM+g+xaYqlQP3/JjMpweeionackSszveHOhquZHBw2/kI
M1EmeWua9Yo7IXHJL/vvWPX9uo+3VVf9NEwNx1Sgy4P4S7pIjFvo63mqI9xxZJ1p/crJYyduzXj3
9nqIAl76/dxZs2S0HfWmsa1HmE2HybQP/xuZy4NIrocr7RbyXM4zjm21a2btCrdtdGQdekuo2WUX
FsPcEz3XmUwnWhJ00k8+gQ4IOyv/S3Uoq1uTrr3wvQZBBw3wW5H26Ayv8rjkL8k7RMZ/I65vGelJ
xgDNTRFrtL1WQwVyumsnOGcpADkt/bAXhm1tnJVOJv7n6eFlp2186JRiIzUffCkeZF8xIeXr/AtT
GnFlpmvUGTnpMs0imUD3nCrsfyYaHDIt1qD2Je1LxSZV6uI/CFjVYBZh5jGYDo++jKVQWE+wNVsw
LScmaQtTNZEEsKaFws5qLGjC8dUfXUy2q8v56pAAnCxgvgOGuq/SQOtkikz6FXElLDatE2KLhEiL
uFzgZXyctr6xMNz8m/ZbbvfV3p2/0USpYf9ORTdOq3L+uGXt8AE8mcxMsDLapssL/G96HSgfxVrB
0I3pcnUVz3Q8vvt3cCsKAEH5ztrL4y3by1wo5Rb2zWR+GBAU0suTO1tKEzC+gphLgBxppbBzKYoq
wX0mAmyFqchnWeLVj8BeRD34he0K4QGlGu3RL5R0qLHQYT+BX30qIhTkv8ZtYR8u4jKKkwHJXJzK
KCzXFVGw4HS0Al6y9UvloWw7QdmqzTWu9GqAlE42IDCLBHRjQ4EAPF/0kTrW9RJsXHCD5fRzRA1P
yDw/xD7xQQG/EKmNoO99iva2jlhIJV5IE5taaQpV/z3/PQ4pLfnAJMCtNNEaXpKlMhxT7/MLyKYD
cxhPoLH8dxm8/dNRBof4Ip9jIF8sH5OPCk8m/bh0VKKRzY/l6mst7rSKIYa2crrhFcINWWX7DUw3
LkOWxMVl3tyFzfv6e3nVvUDix/XNfNPNWXenZEY2R5PV8D2dmKi0544S3pK0WQ4goToiOc86nvFK
gtkrZK7+HXiwhYjyFYRjW/TyAvNVLNeuFBxFqMR9M99kutR1cQPw4qAlPv8+24eXdORjSH2tYita
asSMXLimE4Waxz6G/oJQACNAbSrTeWojfVqImk3rvqPomhoVUFcFBqY5L8S17O3hLbIx//LPAST4
kKCC2VgtOmGVKUfK7DvsyaIte93UhHQ89yKfFsiaUNBeu6AW63rbAj1lcavAUvIQzoADZ86+ai4s
6flimZpb+3ZSY5KwYrd8cSBy46eX/xFN3jHNgi3gfKvZfWXfKuvrVtatXfgCH/UBLRj0eHvzaLvq
ZJNgNi6camMzKIpvsN2rWH7WR5uMtJ9/6ylHReduEzILBwtyflWM0bz7XTNmgWKbrglJDYR1usnC
q/t0C5O9T/jnLPkMmSVQUenv/Hw7CcmVl+QHzbhb5ZP8WPFdxrO7OVJkiuFxeJE4c1/953FbUdcq
EwsGhTChTSACRgeSs2Q+nwhWa1dmlXS6XzC2QZFoNcq0ztZFGVe1aPcNHNtjvxDnaYXMcy1NycsI
m54LEx2DiPulCJjyEPxE4Stp9s2lhRSQf0Ow10VvFQePMVN1giy7/oq/Y93hONQ3qjMkoDn1h+g8
vDcqyRH9heUazEX8gEiN/4ur98HFKcbKu6H7eKP/+OZe/K8xYkGyLFnbceJY/fBhvbKDqngiHTdP
whueO4Za5Rn3wope7Rtr6/W1/5B+tCk+K99/Z9OsRtnPeovX/A5Pa9HQavd+GovJYlEaEIQ+7n5v
Y1YmjDHI+hahw/WRG70KF1QCgWuvMNsU6BVzQqywC/enYUHBpaBH1+6Q/oNhsiJmA8cxLdo3WVPU
OPHHTM3rmNJzHijKkQ6FbcbH15rQC4CnjHO08AMIv36G9HQPuUyRcRM5hXAiHmHAyhHEPVxN/1ov
Fhd6ku3SgA0lEc9FPbSe3EG/wHmk8PotqIZRMH5JLpLQMeI/lsYATl8c5xjKdfDuOSV/UETXCoiO
mfcUilSNnAgKdVRIccRqHjXoz43zsYRxuwRUenJ0uO56fwwhG2vZxdfW+OmkU0geL7Kxp93QFgwR
XQqhQJ0VXJjUfZFIbWV9ZjRAfXWT0Matt4GKdg1TE9s4npuzM8yB6w3BwJapUbK0vLEI7GCHB3q1
dIOMmoHsBjR0fGlZ3pqC6RKhfPrwPzUEavn6SwPj5bVXbtMItzBvCgrJzLXcKZ7Fxh4sblax1D1E
SnHx9Gb/Cxevu/xuca/GxKPSdYnVjv2ItfKVM1vKguEQBDEIujrmOt/uHeyGg8x4AzpIz5/d1Xra
mWeGGzjoOrQoM1EBjJrpBoX4ePqHeL6e6hgsU6fgbDLAjfbHxvhQ2oz1rTYpPETVj0bVcUhx0c2n
vubt+SnnpXzectqTSdznic7TLT7gPu1W+xLx5Ao3/UX/Ry14kPm8NmDNwSIZt5OJJ8jyWvrTl3JU
tLonhrXi6eFJzv3BIESKPBsjJueokHKzBYGoGJ74aoFlS9SSJLr4CRItGwmm9p1aYTT2x3qjJ8gX
zIlQP415Yv/CJESvq6nCUPquVXjb3bgk7sbkBkR5LFnB1m397SNUq1pDiokivHSWR3CmXAiv3lOZ
YVunfBjpjlItyn5lEQMeVYgtDHMAAiP/fMn9fz+rSwBPn/Mrom+ZnzE2FgbcHUiJzfu0ie+fk4YT
oLAHXRYSTZSrMJKTFknqaINj73gC9b6OomoXJA60hbPy8+5+ntfEfMjHnSXu/oHskPjq4Zyq3uYP
HQOBtanraQVN75JMcQSHkWLdL3bE/7GGw0lONGPOBjTNJWIzegee7LK0GijvjcmA0biaDH85BVzM
40nCogi+e37RyKqyjsbPpREwiE+VSvcCSZt6TJSQGCq98iPW17HJhiOxFOhOBejcca8h2KpPlMSx
C1H6xOAeFyU/Ouv0ErxkMe3HFu3XUEIX/ad2auqfhPhSdBuXixkIhXiufEehLD3VPaRkRRuZEywI
LYt89xAXi3i0C07SEyePq8w6y05hIIf7qz5/bFFlT8rwYurjtbGcTfMa07dep0BnurowRrzqRNju
//ua1mea7YKvb20OslOul8OQqoRnCIxGH2ds7Sr8kMK/XWvkXrbQOPRzdFGCqo0pd/sVkDTbF2zA
N18Sf+Z1E8OA5dT82jVpMkUI4ejxbVdYYL5u2LfzNA+MVR2pcPLrQ9C2zRC43gQDV8lMdetIWzlc
I1QqEdDgr2weTUqDFPai/NKAgs98zOKkvCrJ7iV+2rWe9AhiM3YM2Mj27K2UliA/3DQ/h+NCK8hx
mqFL/vx6T0M8Gn3uXXigvKU935IaF97hI/D3fsLK8/hKFt94LJQfBCIoXDJLKuZX9sIHzkVFcf3l
qPMvK2Zo5EW/cFRMcvHSm69RELqp+h7Js9GA7aY6Qz6Ti2fAy8e09HmQvQRsad6sDdyJg9nnqMoS
imlFPTQIQdd7cknyLAfp3/g9E87Vn7CI9yDvQ/4d6cWJqzFJNEWGnF93UAITaxhO93VVlEb5Y8Ny
H3+AiguP4ULGaTl6WNN4r+/6kZsn4GOdgOdf/J8A6fgep1bt2KjbpR0qWp46Agp+k9+JWX7TH/UP
cra+AMzUOMudmswieJkzs4/u/pG0f2/9Sz2Kbs8n+1PyD8FyoQ2K3X4QeRDT7UA4b+2hZQA0xpiy
LRwTS6R4/2bpfdTpqQLIinD6Ukx7HX/LxiLrsL9AJnT5VAia66eaIbjqq17g79xYARDRMEC/Twga
KfO36uZH64rMepuhd5NxoE48IOO4K9NDNppLo9Mnd9ytAo0uP6H8h+IhTdIKyumbl3D0kwH57ehX
EC1S+sICgoeXhFq/e7BjbQ3RYZmhNZZMFaUxACIvrlKhKWSQ09Nr9sXcJJ5uiCIN/4CzS5Nn4aSh
xYNbojVXJC3xZwuYDGFs010niFryIUObUJJqDWF6NHYBCdsKgCp0S5tVHv01OGFUTsJ3lo508sFa
oSV6mn3O0WFduSUWW9+gVuI5OffNdDIA0fnMvex1wQssODfTe0o/ZYYeFzju+kzB1kUmMSgCE0SH
Igc+lQU78MVV8Gnh+9uooGk6ynpFgZM3PJx79U2deP4jPYjOOmy3+nioGaTnsTFBqhwaxAsGJjEK
N5hzyHq0kglTsHERxzVflED30r+UgcCHwdoEtQzeknauwBU5d7BnNpxuKLqPnBnhrvRS6ojWq1Sv
o2EtqOFQ9zWBR7knUDg+BJ7Sjrg78EK5CnFWGMWM2O5jxP+qCaZnDNdaSrti43tcCLI9RY/Rs6FI
HuMtO4udBybJjFUuTFJoape83BMFVTitdAMzFYjPCIbw2w7SkBLSFMLAe9vAeZ/7dg/Uusj0FQg1
M6GT0SofByLFMIGsPg0AwDIMn4jgoyxWmAWzPMIfQaBPJ5RYk9mj1OYaYLZ0gqOY6NfCn/rvdRJ3
u8pAzLVZaEqCqPIZE72WVB5LTVasN4wxn3q0s4MBHN+PtksK/ln1WJ4qmNBOVTalVE2E+NTqEdil
XkpzddFB6IOj1EIQcRAjKSOAoT+2ovCkD0WKvTzoLCeQnOdyJINjSGZE4c82DoWLLgeLyjgXLxhD
SmdLHs+KITuEWAq2RCgTdx3VYzpDgk9UYPKOL1LJrtxgVhKahPOoknxg58mrZcx9ELcRdHcZQ/Eg
lZ5551MKeb0JmYQTEjKP6iXZXhwCV4hX+/8G0UEywS1fzPyj7oskV9YOEdeLcuLpQIcOj0CycDbO
Ve9Y5RIUoiyUOfycOqElz/PLzsxSyuQ8TxraYqKDFiVgkjSdfvAfx/+K5upLkS648kCA/k2BJ5dc
4GH7OftqXeOcWfECyib3QBa7YeTgrGOdSCesbJr6xNOh3kx1dA0g8ZBjP1yK45xt98VCzv26yo3v
VI0zctvFI280Euwj8F0donxnaxvQjrgBgwu/ahgXfiSdCNOnWUoQQmGbfuvMcQulqwuStWibK+pg
jos6Nt2LzlJnj/CLyur8zD/ZhQY223O9ETj0Ef6ezlRr727WlcdnsvHBKrBtTeBbJZH7ZAqzRJeF
raaIr1eVfujKSMw/7fAn/XdRNwxNj+Zcfh8g7gQmZsW1Xh6+o/MvuNRK+0JmqI7aZtyvf53x/APi
SPqs3+XbJkABS2cOkaqO0j6dT5EK7cxfx3kWxo9lYHqFFB06kLmMUd/vvfbVwp8qy3ov6gtYzVg6
PWyRPt2wM+FeUj0aAlRt+/yrudk5tC+mlWu25J3FNyU7bgQwwX/aYb9EtoIjtCnrj2gAYFkqlakH
5OLTlSrShLf1uPvbGD2k25j2Gp7aCW6WjsEdlTCTA4/VYpmef2fK7xtihPCWCuTSHlhVAbI4aore
cisy8jQY37vl5Mw13j64LwhIZyG/mdj6fB9xJh3kw5YWTWXkBMw6Kr3Cl2eDzBOhKNKRTpjqiVNB
xf9m+6+Fufx/jlXlI876c6PI8dC3rNu9v0t9H4QTAiftlKUUdX4l19GfG5RRQt19GZA8A29Bb93B
IWj3UQTAULWfWiX7cApuaxwWzHL5LspxAxaiAmx2zOvXjh3XOjm1bqlty4YUSfMmKk8cnOZpMPix
1Wx41X/JATndk0TiQlYNf0UOcp1b+ir4A3u4TWcLTV4rEW3LioJ8tTSIGUoMK/B55u3c67tWmu6G
1lbkfLIrvWRZ8Ol1qWbOJututQ6v/c66zyka6re5CBeXipUfzjOnVTfWLx/vZvS1/bweO2ZLOXre
CyF5AdF6+eswlwXzgy7wWbMEtNkOB6hKPEjkhusLi+KHssLqTr7R6J50vJjk+a3UxZumE3Q7zLjG
a0wahVtk4R+4vMcmnl9zNNt+a06YJo4O2bLF1BTAq79f882sa1JX5wg9VS24xZ9j4AJBO2IIZ1eM
lHKZHmSXy3Go5tlZOWqAGR/nLmmo4JCwktMhDeMwAL8nJVT97RIqMfoGr60xe1Fs49X0N+yWgC84
XaYczEH2JrMWzqMZV6eZ6EXM5LLnOfM68zJJ00GHd5B1nzIbbyzvij6Rupoo6kxuAMAQSE829peW
ItfoLqspu2Wquh/NKyaKHVpzxZalzWOC5TBBZXikMCgvoj/6KgUvW1+UUJOsoSQVLKeaMadcS0TC
JlQ3NNnPDOPrcKZWZzp3xrYw3P8TeOESIb92ZXitzkspzFi9CeMA6vWCrzw/VY4M5F0S2L2MPV/K
v7qc6JHxr5qeiXQzB3Yt5y0nMTVRDXAcTS9KEWl2DAvKN4y7KzepkaRktVsqBhXnzxX+0S39eHe6
rL/BoIhfpn29bKXvtzohffUytJrUha6CbYZ0s3Y3EgI89Fhb3arue18mTAOhQ/GR2dO4MXFKQTPe
Aqe4SPWTmX1skeYmXOLsgOsyTKzWuK7ur4X4WsMJuN7JM2EfkgSvHRzE/D/0EeZ6Bi7fIqvAHVeV
It99g6sqDnoKErBHND2Q0CvhYzi0/N1rXx2KUTFQM1s7h164qGG1HjM7rBlUrcL+Gy1anITtCNnt
tNmlPHSEmxD5ZjMvWyXQtUf3TtqUbaLddwJgvPayjpJumUVzZjAjqjdnDylydcgQBh4t7MPgq5gU
o80hb6WyEt4AkuylcEcoK0/WFLXDJxcs3K/0z09I7oD2y/KqpTjtd7KV4Qm0Tsa195piAgjnHUlZ
DhL43I7og48kZC9RNNmyEuFHWaAfQGK9cy5ZxK0bRkfYgyksB7t24NdLQSq2oIY85d53CVUjhr9W
yJEiw/Kokvf7VXkukTAlkFNCyCBqTjWRT/XkkcjVTigNWzAqdwqYhqUXiagsbYIPqtUJu9hHwmC7
iJShWQg33gfyGGgrlzKq9sRfyLQptx2AAC/XS1mI5puQM7kJ1Xmi5JcmKWSK4PKSVCkg78hDEbNA
ye0H0LmGXHqXUKP0kX8YxhNacDCCUKexRp4izT5mPhzKfC2RFSR5th7JgzQlTp5yV9F9TpKIQmbd
Miqamn/xEtuazzPPdU9VwMxCya0YLCvK5RvR3fe3bLmbSTXfryBKSFYGHrRpYbxfkCl7/tOLTaol
psOBHZSmVoAnLUfPW9hASnPGx3sRMNqn03YMs9dEud8GRZDJHoTuGjjnfazm2StPdxXEQIGyNGLR
D7hQDnH6d7hejbWORgUVJA5bte3Un43Rvc5Y9sfNSwM02u9K6MDOoB7EWjb7dIVa1z8iP01y4qoy
SH1RJCYwlOiVez1ApKPx5+vMnHEE51bLgo1YN2FhoGPSWnW40JH5bDhvbCJXGcgWpVU76jIGZQ1z
/GUxyrms+nLLVqrQoqD7h9CLVAivaMLD+/J2pHwXWhHepf9tl27HweLyNs2iFofCG0n0L2YPIto+
fKmS4ypqakmW0nFrhpxAiFebQoq4VDhXpRiRCTjjeGV2HafMao9WaVUx/0qC+k0Wvy9PBw34xwKi
cMxLDPQhDiwVuRvFA32UAYTvz5LRMaEXUO3HFk5nBWzjlwCU/ZLcYgqAxeaNen7HsxY/2siNvjN8
SAYSJ014fgjuEUBiHLe9xrV4x2Mg2kUaWU/lfPSpXOZJKHFnkdfpUPCanXr6bl/a574UgXNVAVF0
ShFewOP+VobZu8EyoYmVlKE1PIwCgIdiGo27FZfnpXTVd/X1G+0g+J6MEgFNRzc9akeb0K4KTOY5
0MVNrWzJvNTvPuUHVUCsrlPS+c3aaaqlU3RLJ0UPBFIyC8GjcHHDc5ZHsSAqLVWdUz6MSIUkoSqM
3YmfDcNIvzF4WWnbDsN7VOYCDVpSK7or86HI1hVkwKVcI5PCcv4dZvfzRW8EZgdGn/DXcA8qaZZ3
QeoG9MjP4aFPVEWbVg1KNiqMiBbYV6lv+IQmqtwLMJr+xGOzOYSAyD1NgxWa1ls7EH9bVhiC9kTP
rgNzREa42i+eHAXbTG4HmNxSc5a9Wd3MdP3gXaN+oH+denFa26/+nKh0dhzA9WAJxWbJiGty1A/5
ty5XSgintPC1tLyjOFJVB5n+ACJ9QX7x42Uv3bnPjkv2LoYo4cBHt+QjjVJVxRKWNRXlypgYh+E2
IZurvpSd30Iy7w8+w3JXBZC44n77EokTf7ukWKeqZxHrhbFv51PdHOqKMQss33IPXD2tM43GeDIM
MAvpQMm9EjZbKUuKOmziUPF2vHbsYO+CXl+5dIqw3bDcFp+LCQicLHu7VD2OS7u902drhOll7uqK
Z0ZEVzJliVilHLYrphrVKtMJk8sTkyGZoIwIuCoBq36hjYR0UVALX/vTMOkDgUAeimxMpZg3nnBd
AG0qGgOxA/x01T7PQJu9Hgdl5kEloY0t+L/3pDDHgYUMfxlhVag7862s9RZ+YBKe4JaZoJMbEkNY
rdsl7K8BYQAgCkll5wg1utRi1G1lurETeY68LTG3deYlnOVvlOptg0Xb/GN0ISkN8DHKPiUcHuN/
/JWphzxS5osZ4EwMZDyv5IM4mMhbJ7aHTlJTFSu5qhnQgeIytXLEIhctNslHmAaEZJaCKTNJ296m
d/GqaXIx3TRx/h9v+4YoilJQY6ZF5BX3iQNWx7jOfXdu2fmL6qBJqfAsP7ucpOIjvJQFHrJPYv8j
ij2urcBwt42IsEha1Xw3BWkOl08eCCbpD+Fxf6woO6MU3SrtPS03n+JC3+kVbAhROcgQ/KHEwPc/
9D4iMo5/SdgRbU+iDu9l3wE/IngO1yuQkarWp+ZGWt8Xphn3srbV56FRn/oJpuiG4GMlf0QULoq8
jktWNgpeZQd6E/EyfbAtmtk0CsDMk/eU6WYIW3HRSK8dY/suaYYECegZO2EUs+qDTRXjBklJBMiY
qh92Wc2fRT5fqk04gwzgP3InFoqmiCRy6JYUPNYuvSKE1H5BDQ3YC3omdW4LCdeC0FzhCQ6qnLBm
Y9nhr2hhP8QG2lQ2hMzo2Egd/8piArPoUVFBDCqCZCaS1z5so5aO6rVSNjIPCPdZnXDcru+yGK4j
+km5qsYFx0x61UvEax1vzbN8sfgLUP0CtbvO1AN7i8dkQwz2T4Kt+HOhdvtT8nPjarmTe4V9PSpH
LA2/j7E9RmGZqBMtC73Y1kViu/NAoTiejB6eaDr6q+wP3e8iOwpNOayWDVH7xfYST0ka0wpsusud
AEjUH8b2HpWOYaJvAll1e3JOdj8dt8C5ucIrC0Wkqs+hAnANI/XvvEoN1JQ3UbXBo0NqcRj9/MEL
hL+7El9WYTBFdEJYEXz1tl/v7FI3ZuMkqjaF75fyV7/LASdBuEkPiTXZYwNkIU9AhDuZK6KJhHsE
L6V00MYeKD8OkVwXSFLHftGPnAc9iZd+qP88NNnADAEUn+GMVlg23CJtOLjmnLEcCvAaKei7XIHs
nzY0HaLcLs3eHocarbb/SqIIs1rnqrdELrUpauvasbPIBiK+4A6SlZHYKJwjXr075LxqfKoyuP79
hMtNcpkasZMK67+Y6Njvn6DC2H3LSatzxgn9kEpz2KmeyEu0ehqJ7xYFiHiZIe0kwenFRE1hN+NF
BRynTuia5e1+MmtDoFuDLhRWfwIGe50AqcPB6tSp9SddVHYQx5BNd4JDlCNDw+0kxprmXZGbVISR
gBCNMqPH2co0XjjjWrKmWAkEuiFt/8lWSif562VIWbEsgC6CXLs2bWgmnp2GYEt0AN0Iyscd8YpA
uqBsGqBuYDteD8JALGtbpj00Ujt8TqZDxn0Z34W66wvyU9LvgfSmkaWAX9CV7o++T372sMyZQvdx
zMHJSjSitFC5HIK6cUEVEHklE4nyyvWU3lCtTrE2/2WMhnvZQqhFogO92gvpNXmUdBNaxeDj6eZ3
DZIMlviH0vcEhYDUvYmjfKCR0bRFKOOzX+Gm1Tg6O7iU3N0xGpe6LhuIg/ckobNfYq9j79d6YK35
faiG2I/2dYsHGKzPF9tl/kJAeTrWoGxCUxgJ9bz6e4zlt/UYJabKW1s9NvqpeAfQn5Prz5pGjza6
1K2qe5eollY0TqdbOfksg9saY5cauTDF+NFNWMaFb/poMpVzO7HHgq9pG5MJrknvqM3pJ5rCUB6m
2QImDiIrJaKkfXKd9KrgnagPj18SHLD/JhuIxvFwSteJM+vkGtWS+YnmYoDPTCVkFpe5ht/V1I2Y
yTja5J4qOLLyNp8dXv70AbGAI7b+u9UhrAihOcGA/NcLYxIcu97RIbQYvkg6Lk/uRMp0G/Oo2ZAN
EJEI6T7xwg/FDdqjRKnahRF+HrJy7uWDPn9p0dvP1lxwaOKuMXoipYDyZjuxePCmG/djLFwQMTMm
cgpEMZx+hx0EddxKO45yK5gocetJkT2XP7ZeGmneXwybml4+h8fJ85NGYwT+U5r3fXQ9F2GxQK5A
BkFQRsYIrpBfO0CE10LqlQUb40fC/cPgGCusY92hel0ISI3NzWm0UMOA+h6xR9sKgW0lj6HnLH8c
NSQshgnFM8kz+NbyPdSA5EfYAGX9vBXZXtjBBCNM/w4PxNjOvN/5JND7UA8EGeT9c0V0Fj8cL/sL
EoV/V9aAxAYyWlNpXfMEoMq3ne34ZTbpDVsqDXsjnamLdApXyRTsHTLRhbVqGBwjRL2mJ5HwwVd7
4ntqbNx0VPL6O7FIVvk+AmVbKQDV8w27ZIvF2QFiUWFHomje91utUYNjxoMCYlYy53VczrQOpfzq
Hx+pNxA5LPos7OSTYyxaRRcx+jMTIWGZH7OD+5am+urfPb2KeSR1hAsUXrBJ9FTzwQ0PuCxvOniq
KqPffiGVt3lo+c8pvQJgAeQrvX6OunrLaDfjuPQnNuw+lG+ovssZO2vz3sZMZvPaJgOh4KiDfCt/
0+5lzonxCTaKSQnvfnQWsGreEaPzPklTFa7JfcHHdD+ERsyjFQLtNY1CtzRSEfq5AkBmM5jD4oKP
HKsh6D0sCoh8PcFkfqDZldBfoW7gIlAZAWxO0oYPNeYS9ccZDnOK1LSBJmakP4aiIUKokRC/xQGu
iq6b06sygeLFuAqeT0xP0rWpbaMXpQSajzYv65zljG3PAZEGhbm9CbyNfIEjYhlr7598HISABZ9K
RKNnbWUKc41FOPjc1sNYWZjVBoRrVvkLQL0ctg+pU061AMBIt1stFGhVFXHXV1QBmRHW6dSJJ1ZW
FofacpTq9/1d1uIE2LXPM26GeNxKZfNN9aG80CNYmTXxDdzld0sSgNsIRzEgG/64ASXN3OndXKnR
9AW3bv8/E4QxbMMut++8Xy76Q5IuNMNgUKn7xWlpGS0kQD7jQb8RnhRU10K4i2sS+cfOF30gFUlZ
n/HIwcsS4/v2t5FsipstyIbJTH32AJSdlj+4+v8Uy0vQ3d6JGWQqBfbQz6EHXM3m7pnt2kmBm0wt
wrgz/2aKLV/8ER0XGUMx52+0GRGa+reHh7yJLvDv9IBZE/9rXIezWZRSdJ7hlYzeW4K8LnflL2qi
V6QDFa52/TpozRKIVqfbLoz8V8EBtBmmgT7WJPosU1j3jwuwltwccP7ZmK8AfpcNy2ItBvECKAvY
g0o2Z1axjQtuzqCKmUoLH7GN3K/Mmk7VHdvOFc75AQxFyxbTVudUFyhjGfN9jk4u8BSz1BEd/ojg
ov/uTlSW49gicTAqnYcJvIytU8K/t4KmAk40VduyOQ5SNify2fa2E91O5exDtUe+PndezkFGOwUg
lTFgxaHA1BGgjOHZ/EtAdv08C6QuUxwKxtiT0S80wRiG34jfoYUUkxJXRorMvDbZK2Bkspg0hWcg
SPrKEw+cHbffG1jDd+R0IXrS5GFO6RGLtKMbba0ZGBV7PsxGxEilWNSfABLf1LtdFNNcT+KlIiJh
1P9SEdYfz2HvzAlGp7Vi99yd8cr59MFrJuOSdLBGjbzZE4EpuWJo+BoN0aB7r3k/gFgHW7xC6VGU
CEzUnSujfZBhrfQvCd6QtnkRp96hYDnYQwZoAxJO8qjbNS1iWP/iFavPrmvXBdMVje8zKHTlQ73j
QCT6vMt7gb/TMVA6RogkooEoJhvm5j66IVdcDIkg7XRfT5wdaXIBJWe1GHr/evmcXZ+pugQdavKl
0UXduSgcsWhaujTooUdmMr6kGpzt+eoMwPql6KJ2ZH0R6/SVemqFNf7B/kIByP4sk/6Je0N44qtx
Pv7p3Xe6ZG1DJe2AGOzmAlw/To4/ptQgducJBwncH9aK7O+slABL9m4px0hkPzanBBpj/3SzAluD
u8DqxMa5vSn8zId+kXpJhJ2BbRRK5FZdMazv8O8/IrvwJMB5Fs5lCSqKXFCu2x8eExcN0jHo+RV/
dHU0Z2eer3lo7V3EaP2uT4aGwmo2JEm5Fjj5nqRXEzDzuN8/RGwPOc1swZ9iuemdN5LkI/KIPvEy
fhJbaSwp7SZRI4/EiKLBEvtzrr5rUrSczqENF6BM8oDbvqGUZbOLap4iN5JrB6df94ojdamj9otc
fzmoum4tTM3M5VEqygOFoXgyNv11lBk2ZWeemJfWBp1BVDnUX585DL/IhEhuR56CCUEi7cfE1kO0
65L4qxkSww/tCHPGlouTHx7jBNk3RVCqk3b1NDXbEC7Xes5/P4y/s0rCtWI1zRWdeBvo5FccUdRP
8lqWdt1i3Lc8KbuMo6sOJKE4Blr0q6/frVZ3ltHc/j+sW3P9gk6LyQzyP7Eo+lZthFyGbGswtaFn
zu4alRzYcTCGniWlxKlHShYj1bN5HEStegUP3j6QxZ4G9TJnh1T/S6gehB7qHSVhOHTcgvATMop3
ZvYpmiUXh53ML0fljv0eQxVbjdd1lzgAWsCf7uZ0cwMRVNwPHZCwUig4AFMMXAFPyqVxChR/mff9
evxMGuwcF8+Ncy6TnuPfkhYlbfU/UMzl4bw3Xythabvy1eZPm9C1zOu2LgaN6WzdETieHORI63P/
iiCh6iXDLT2bXl4M5NTwrA8CmZaUzOr7Bqhuvy80l62b2uGA+ev3kC35G65akPy2rood0ljMcRd8
WyRpafY6iKTm03fMG3vmVXgpwa2ixx9dJhbiXRym9Lw/vEKlpZs/b0HrYSsd2zdXLhne5zow6SAs
6XxbIJYjJalWjUaS80N4Z2Eg+FPKOb1WoxRw+F1wj9aULy6Bf7UyitYOzbbOltyEhPgfT1hiPwR8
IS9bqFb9x9SmTH0fJx/frv1c3sVCjmNkfR5UrUp40vytkRBOB1WLetkZccWvIUOoC5IjB6qDAa3e
+DkLJETonKMGogRUIg0RPpE7bMSQ/qoWUe7M1i6SaPfzmbRaxj09gIuJaa1hBeELYiKIPOxv1TzU
LGyBMEe334oqc91RS9JMEOZfHx384JdcHEl/lVcZ11/zeJunPhZH+CYY0iBCFmBQUmXdpfcyEp3R
quVrCnOWI6U/R26HUI7ID+OSXP9D+JXsOWafECjcQ+KKxrnKhq1nu8AQzldvcvjjc9rtbayqHe+G
k+6x2qvF7L/jJkaOYwHPry3VSOHRLHeV5dB9B480fepflnBbM1Envx4sqjkXCXZNnhbU6S9tAgyg
994/+7PA9uS9fKpLZ421dN3Ozb9GcSSZsGh9+i7Cgvf7QxEEySlDKzgDuRpwHk2vuyS/Gx6KkdQb
EazxBK9XK1mYU1MGbi3CjI5tpgacMfD9Sz0sxLsj0fTLtNQv0QFbnl9SL3CxHFVSZqqUdZlHF3It
3u31+hSaXNr9S0X0Sk3xcjlyOwzq/F/odOvf5KuItadFhiWChNDW3KLGbk/Z7J6Xio9tK4msN0CY
rqnRWa2mn/APGkXJLHc4AcwZjPwPDVweRD8OBdq9zQor7E5iaT1Kd0pTmoI9mksMpPGLQ8JgRcYv
JC8NP0UxZOQARG7/PoBqTjkOAw9bet/Nr0ZdXOa+hyHmUStB9CiOhJUAcVdHVSia5Q7C6xFbkR93
YQmnTB6oTFt+ytYTYfzoyA0oe2XuVhs6Kjo7o0XxAHnrhcOdxdKO2MnZG2/byg2vdQXBj12MmuCj
dugKtGoCOlEFfbyNGAmHwSJfAozrZqzgI3lv5dQf3kz8ZQS+3OLZjMkeFKwKo+xC5dlI8OkBUI2J
hz3KWyrPPNWXwhWqdb67JNMVSOJDlu0Dt0T1vabJIWuxgbnzKYhTizBbLBwwmz5ek6BaPbS78fpI
2oFAeG48neKvHbcNecnf4T1bhhuGPQJordlQDJmNGC2J8459BSilLcV1Im7XM7tp4uMjFtuJvGV+
wKR0JjFNRjmMHFxribXS2qjnbke9wjXuHP5r3PYPZHaoxKhwfJghz8vVJE5o/m2Zg2TlZ/Wdrykq
1WpKz7MydscUlmXZYPKhhnxGm0ubHxJkaDrf6W5h5CWzH3U/NMUoCTDV4qjT+i0LLm7SnMcMgC9A
cTsH1xoz7yi2HEHISHeMWsKEbQtHTpbCqHGs/xMBIkkCDUvnSDOxtIisqH18YwatUNYveKaVgdOE
yHCjcI0oud0KQG0n2OSUOjgeGajrRTKfLBtxp23Yx0g/YVcpkODoOlOeTckxy7LfEXqaDsMu3cE8
WhnD8PesfQknBUzr8H5rBaonj+oSBKpCGhzfrbluGhTWOqWQGDWyokDm1wucylBlBAOoM1u0/w1C
4S8Y/WvQB9ZCPgW16fHo7jU6AdgMUUXUJ5vDk+CthlkMFLCl/0P/c9YZrbAI6uC/n8W90Z2gKUI4
yrw3eRm1RLKO6gItEooHPvWeTj4jc6FNYhiimpPpuvQ87ESJEzxDWdOfoLudK3coOiBI9UfewHAE
8NHx4Anqzz2zPEYV4DFQ73mTMjusregxyqIhv9u9BtKnqA7wSub38sfonXzUH2e7Z7Viao075/WH
jHYeyfOT7ycr83HJXoC1sqtDnUPEKzOZ3KMFBKOunNVT4XYkpU4J57Wr4yhHkloXDFCzwouxIQJu
tE7HVLS3NZ93x/4rowbngq7Y/UOWqSIQQ0ATD2RvjpfJWuzmumo9BR2h5KHwxCUhS1I+ei7YKLVa
LK7GU1+R7CtTLLovK5QVUcOpNrD2qMktyMBRSkrcSmKxGMkIRjY3AwkAVZXIMWB6+1XOITik5zrc
vhKJfGvwEf6k2isSHJcFLI4ekPjd1gi+z7OrjZ5IWSDKUBRTpr/4ymzdp+mNWT6UtLOsymlFuAhs
SFYz3HicRq0n/LQzZSt0jMEZN4kY13wkNCTGvZPk1WWr2SZYiBKcWE4BAvqY8prUTw8pSjdVGfu2
U4Qzynoyvo6XRMgrpy7jVqzjB8tJTA1uBT+qq0mtOpzfuzY86MCY2i0EqHp38yZl1AAUg7fyqyhQ
FSHfgdg8QikXZw8ld+qmWCIMpqcAz/NPgtqsEMNywq6tR/4Bmg/G/w7nH74NFpTsoqTqqy/108Yt
FARqFybZ/khLI5EtNYqrEOawLP6BI0xoUuxsxryF7o9BlmFqSlcAHS+nI1dwSdDXZBZ8ZczQD04t
6cwqFczjX12G4lR/3kXap2BVdzDnzmDmNU7oliJaVXaLLFWYGWnIjOw74q1VsIFHn+wmYk9d+QId
t9jeTbAsB/USOTThYPH7FpNB6ocS3EXEdVu6v2GYFy9uneuqzSTdSjv/5IJyYAoKzD4pcRx/YWmi
ILZkkp6yeMUP1rrNxljX03jjH/jsXmeVryxU7oOdV71SWFeZcLxsQr2pV6yULr01ziS+mipWtB6c
3cdAu05FD8BjFVnpCZEsgHwuuya8HR2dkZCduKYmqRtVcCVD50S9jrRw6otazKufdGUmuSRhx6op
EB3d7xP5CxLBkwppiHH2Ofdf/uMRwwlNbLVf2YBNBcyacbVZ0Tc1E/Svi+LW+ZbkJGQTB4iHoU7P
a3kaRTpUfTTzaxH0h5k34qazDMNRtxGVDqjoY/mKa3yC1JBpyrMGNCIx4/WL4snSg3Q0XUqEair6
hx6kIFqkA5Ss1fhfuwVgoe9nkqb80vsuoXAFgsPbihEqZDsENPVMQp74IP3qVHWZDzGPSHiMuYu8
BRXZRByxLc9oG9c3QhRakBcKg0mpw+z3vMv2RGooWHEtToWnq3FjwbJDFrmIzjeQ54kdCy/7zBQB
UOXquUHRAydUsGP1cVoffM8yCX+mK98vFJe41Mc79EdNsX/M+HCnIys/1VMbUHMP6zDRuTiMjDo7
jxg/EvtkeAOvTUeKDSZVW4jqwBCRW61+lvBIlGeluSFnyiiMAIXTpv+DRtr5jLd/YMX9X3LOvsyt
rrg1SM8TMU2rL53pzZpDCP/DTyLQphYe5xhhhbVowdU3ls79fovdIE4xXZ4vd2YP6/jyiDEjtIYO
5sNGZuxSKO9sFnmApmcixiyxJhW9vdF+2ADRPfeKyILOV6hu69oX9KyySjMLgSYd0wULhAJJQCnS
LX/Qsrgx97tVfKA6Zu5CFhtnsng/CUzKlQiMgdh8GXZMH+sHckRKp2rhpdIYFfC09QofxQvk90ur
QhqJ0NWcOtDgT95vBnIn88xWw63uH0T9oM/2o3ZqRmTtV+/QceGhq1ntapFH+bEMO9lGR+c1hRAw
KO5hn/f/vAKfi5Xa2x7i6bCgUOZMgObVNY2ey1jRrWbzk5puTJWyRkbmnq6XF2tTxdV3xvNIkgXv
GDSWVPiLnJdOiRjabw1wyz8/ME5w1rpjEAEC7PX5l3B1jpWpaZ5PjSWA/gB/GLh8Oo9DEnWL/4aH
627qY+Yl3tj5amIvuXIjjDPleEwWuZqVJj4m32TZ4p664UZAq1i5dbj/Qa/IPEweMqvdEmgB4Aan
1XL/FwBrooL99s0gLkBDqK+ejd1zvbg0JuJXMDHWnFF144LW9hg2nIqSdmT9TGDKUEWIBjiJaYGB
4jqiEeI/MI0BGTGVqY6HGPaTmr68m3Pe9ZpHWkUk7CZxqlfMVn9Q/d6sBlpzdTD0xIpY5yD8Fmq4
UBRKK6j0WrpwbjTb9JmZLOi0R6OPsm8t6cnO0SiZWd5gn3IdNbZa9+vwGt7ril80327n5q8CiT54
vl1yr2tI3Cooj9oKo2iuFKrKh6PmW21CYSEgzLOcyY27iYABhI+HbL6RDbfgtvdiGpGhAxyEe8fp
Jx+KU8jlgwjJkR1pkk0w6RSYmLAfotKzdLeZ0ioXSa3LVXVflGEw1bNvsfnHcVFC8DClG5TwYJnY
SiaxgYmT+alsVySo3U7S/sWbuRub3DK0Se8k9hy7tdWtvmzLYnuDqZaDxtPuiC1nu9QJoWqnneKC
S+ps6FF3yP6bcDmvlg/E6eIAevD8K9/Pl6kvgvZ0NWSJKGGuXoyuYBwe1W6I9YEm0eaOwN9ULpsS
Sv60TbfMyw8SiBvVqKcAMuV0UPy4QmOcuKM6Dl12WAdfxjtjauNG49U8eNbDJ7Djqg2sDQz8BHD1
U1UrJXq/quPM/ByhomxhFv4j2u4Va6rbbjDezrhabbpRDirlHU35/0wmUBnLEamF5+sld9Sz3jrG
ZQL/jJw8xPRm0hVjsoQOczfLKV/QVz6amBkcaqg+uLv+UKLQC0wZ7IlYt1S87OGRAJAGj1cK07ah
xHLB/M5B6tDNNjqvehR++38qzqgDDCTHA7vLm9q5uhLh6PZd4/ZzmWAL5o+2QZe/oVbowrUZMNQV
O6q3I7JpASJ6o0KkSxnucW7y8dAtQUphttzystoGaXj8E08u8vTu73wn13omU5qz70afU9PgIw+t
wcrH5sUbaUMfB6/ekTwok3/ibueXVH7tqlgp8n2W4X4hnXdix0MCmIxM/rktj0aCXzCbFx9QkkdC
XSePNYKAJkNv7ba9FYDLr5p7ZDxKJEiPoplZ6FCYPjxYiBk/aZC6YhG87xZRlZ6Hpwbr+flTwNPk
bHkvn1gSd5zrYWLUaYfVGmXmafGM2CFpJK3bp6+JLcMyb8sEmFl8MVTca7s/r06aVhkK5Gp/xZRw
1+lAiVuTF+cqRIoTt3Tio3jMzQcoDF1v+zciHbZIcHOd1fCYOs0ck8iYLWgO5uMOBshPb2lNJQXP
br1dzE6p4+C0EoljldP/Y5LCQgmGogSeOPDwrtQNdR4/Pt3/p/g/WyVz6EIKw+LZN/y6PAPGLIeF
lcS+v702gu4hwwFHQe7HQa8Rn51OWvfXavX1z5p5b7mChcFRtkC5zcoSz31pgN2NbZ9x4bUn6Ezv
IcRMBHDUU1Ovaf0AU2y5o1YmIPiGZORlKdIVdlJyXmrtvGoOE5nZGBs7waqPTfZyv+UB95hRyeKx
DX1CXhnJ2VfT6qFKfsiYuNLqwifJSUoHegaB4+ITjrfMNBz9TBnU5jjUNCL/0mXYz7qIMvS+FaFG
FE4noKZAWdfhtaXI59Y1ZvdHxjvfq4bXbW/1+kxbh3wlv8KtpjiLBjDTQwi8hGb7NItdi6/wi/Kp
h5+vGg1DgKxPrZd7m6SaYjhCNRtdxEyHJvJbPMfNgMfelsiKSsjFIL8yPIv/iy0vvbA5urq3yiKS
zF0W3Lil6TMKUYF9i+CfBMhghIJVKh7k/NEYz7XQTJ7ZCzjmwMNN2EDRKh8au79utd9rrpJsCGEx
f+m2iNEB14d07/q7t0qvRHMzJd8oLP1xgyopx7dpp5Ih1WdJ7Df8TjHMSGB9LAzmy5GLVVARHcAz
62cIDGMFiIfq2oOxnpdUSVOfsFDkKmeozJAbQt9qCMXe8k8kBR7KlKeCSBzRWbWGjxxakbdAcHGF
RThEeruip6UVUMFUdRX4y4TdpEtQmizJq5cG8ShWI1jC7+QycBouvxJDm64ZZGgo7ZE5uVybdjnj
QvDqkr4KNYd0bJRyySevubL0oKliIt2akb/8iWSMwI3+7EJ5QaIL8gOW7cOOe+uqUK1JjJ5cf1S2
ZBCxjjteqz1KeVVC3nppWt9nkKFApq3S+C5lgF9PEqUcVdK5EtwF9gqbXnv3o//nesQaTFy3jatE
24ByL7RFTQ7hQurqCpmypIeRk6uK+c4Da+mKNfb6LsYAVGWTLGrxOkWVOB0Mtdomk53TvoXcDodR
XeRxsiMoOgQTIUSNSztVAfuHzOCNEC/tbL7dFKqlf/eCWQdxJgOHoRaX1v7eUxPi3/Efk7uYgolT
jBM/hMphG2w2rbBk8h+s4bGIJ8KEONEReZmn01Le2WRXBL1zJKAOXUXTvaKURdMxCjDg7+h60jEw
KV15zlIscfZOMYWGR5CRqdV3O48FskQ9Lmx/DhSIjclqIwc9C9KeV84P7Vd6rq33yi9W8Sl5hctT
kZLwC8oXPzQ9kbI+G1/+eIpTu9vLY5si5Pn/ZDWIS0jhNj8UmdDVepr38upS++pskkbWkul9a/s5
zlNQmytOUA9zxmlIzt+aSO8dA4gTBXbC1m2s3D3FWui+zPhxG/ZLVq0jmJgMM0ZXfWKoNkvaIaH6
uUa3jS+ym+Y6L6YGNctEF42UeW4Efmu8X55ro9Jb+JUC23m0qMnbsduA8d4IEpsfxUz7RfROxOjy
pfmuKdBwAtFgtFxolsMYQe07rXV0zuisc1J2TblIHAHWxe0LVu2L4O9ULAQpTs5+oKrZFK8KD5TH
hoOyOuwCb9HzbOvcw/zAzpbMBDNgLk39J3mihXSws3K8GqKZMdsK/Ss1CP5opHjfTRUErBznzuFh
vCuPvd6K4pIYcLCqG73+HviQ4fq5HNspWM7EKHVFLau1MyguHZ41fST13Xtlv4v2uUtNcDQap46R
ruM+UxKzauWPRIwDQBOrxSc//iv/MV3aiykQmY9YbmmbZewIGgVpWgjOyVAk24hQFoMZQkv/JdO1
gbFnd0hPA1JG/jKON3pNLgf5iHdqi+mIzqz2Huexqb5DlrCNnY5onWqlg8LlmakryQee8ut+vA6Z
wDFzkvYDZWZdTxFl271gmBctNrrNq0wLgeI36VjjP+nQ2XhRVY085YOxIefNFbNQm5HlZT9uIr4q
vvyhkxtzmcFVQBRTu86ovdqYSGs5g1owjxVo1UySPGWoWYFmlpqSxb9bm9KYAROBLod0kgeYiqbj
KJ22r8cGBmY7ehdW4ii/W+Dmwp8pTTBE/fNNcGzLWe9KfZeNuNaiXBRGg4v2Ca1ok45dg55h+U7R
SkkNUVkn+eYAX1tVCiTwK9KBwB3NuOpLDgkL7kSDQGXMQ6b3oQC5YZuoKn5h/YNKBq3CoMS6nMPH
Pyd3teUCBjQ3BJnmj+ZudBJssWH/nOm1vB9Pdb32sVr3GYnumUTJ4qyEPwynDiDFgsLvOmqZtwlm
2ONwH2Ujn3priQBjswzSpJrrKa+O9G73DHGrYfmytDDgJVum1AZMu5AdRCPafYqlFutlFK+5wLR5
zwX/aatzHpVvAT9Qyen9Prs4hoJ2SCTalgl6o37nuupn1/nYnvqWlEyMuIPe+RBNjPpzOIYkmhgG
jemaWaFAIHWuOr9yOmPYDxH762bH1JmIB9ZaUCOnxWojBYeLS9nWy2Qw/Udtd/0E7ntZ9WgVRCNP
n1hjizRLO9Zpsqw15QKg+gdbhQ2nIGU/z0afHmlFHlKLumPl3V7K/tNFZHzYs+n+0/Qm8OFFzsbc
xcd7ShPG9gcjyoOYg/0vI7vUiCuT24/3gVKRzctnXUARsZdIk7mGNRyKjz4LOEyM5erjQ0hToux8
iMQiLT2pSErzKZADn4MIwxm1FycTwtCD2oelU3KqJPzSZu4YoMgA0MSx/sQck5xbpoeMMRUwhHYK
I7MLjRgBWe/0wW4mAbwVeX/Eae/Dab0Pq+rzsA0UFOLBDIKJUTiV+nr2lEI5arJQRKdmdFAa6GYs
FYfJ1EusER+1q7Gz0tdgDODYTDG1fKw8lL32IjZDz6NQIwhR9GsBZEO2MvvqCCXx3fkzg4OG3Nr+
SgEsKN3kCxsXP11SprcCY2v6TWsBSAXCuU7B+aYHg9h0Qo3aM7gk1hUrdUZkIUpllHjqI5OkH+81
+gHWZAFmrwzWtX7A8wVa/pB2evsXf0HwJCJ9X09FCqehKItNGsNsyR1UMMNT0Os9ZkTR0arV40gz
OkdpdY8exQCXositvEICJTEwyCw++BhX/HpeCexQ4kudp14P2CqAFXJtXYqhHJ8bMDCYuygiwdjX
FIbLJBuIbyH9I42/C7eS/uxCv1byqlw/JX1KNnNdDkbKJ7TXe37RFr/o3dkxNIxsb79rBnQGqLIY
pSf5Nf4wImUIhSbJbsxUvfB6ASvtl+xQTYW+6G39vVlej74+PtKmTGTIta0QUKwTkPV4kkRfgQSv
vubOKCVeUeuxHnI3oKYBFVncSRwTRR1AYDHSeYv9m6fTf1ELC6jBWGeU78WoVz07ApTA3h8Nt7ng
YtyWMx1+v9ArNuMfTB4w0Xl4tw7cF8bkz8q3iNnLZwNhufxgMtJ93Q5SG0edOaT89unEjE1ECMqm
kTTQNdKwgA1sciXc8z1VMYsejtyIpEr5qMehFpvfJfUfKiiZcTb1n77ydK4rMorFcd0yWINholYp
67cdY1QiGhncSN+ldg+mKFbdS5mcosIwRmsGU7WN9hqa6C4YmYgspAZ7CA3NSgOdb+WQtC7d4J+9
ZzNIlaWQsZmH5AAfyc7WuwXrFdkjymAMbuoTIATLOPrq4UrFqwpN9nFkVi+udd/44gZRAyxyXDdL
0FYuA80L1FxJ5wGRC0VfbjeKg++8WEXvCF6+SbGwsTBl7z50weutRoel5fLYChh1byMDHHLHvpjD
dSamYXQcHstHlkdBQVHAGyOMv3MDZJZ3IPr3+sjF/mTQnYnVyrycBQIbELuezlZZKSN8uOD0Y6u1
fMhB7nsBvuClJgl9nUEidNDUPZlIRq1uyAEv1zWna1bJ5wdfZrDna8Cj3iOVXIugc7/92PSSuxWf
HPSvUFHGJeqdTPFhR0ZtcZqxGz8wkX33Gyq/Z+xm5SpoCiK7fW6/SjNHdLFRwZ1u/clzu8sUMng8
4DeOq7EmBm66bCPw84PxtyRUPGdfrNVvslZQbZp7sUA0R1CyYjn3pSW6sGkhnk4jm067UwMB5tqY
flR72Dfif/AvYNxOMSg+H3CRDgFfoyk/WGman9hCEBTDwx4r/6T2oyKiS2TlnPozS1bl3ABMuq8W
lfd5ooJPwOtE6NcTUdjJ4FyLS0gAQ4DV010lIqhDMtDOOAVwd66tjwLK7ZWi6cTWywczb3FZdnPq
aQjmv5YiXWcPmDU/QD+NhE1eb5ctWkSoR1ZlC3RekpzZk6pjWEpDhyGe+1Ni80zVPbUBBOZ6jYn9
uICDG64wO+0loFqcrstD2+WDx/mLEnllocSUHfIaTukBrp6KAsz0d6u2lcIbSE/aMyCinRW8nPPN
MMEpaI3auLRB72bqM0zCfHyK45eDlVXfoAg9ijex25aVEtRshDQGSsX31Xanao27AtSJgQBV/Fft
oUUgF8TECP7pcZZ98jvFmouXv6w7RmIVsB32uTWmQt5mDauhxH3hrI6rL/56Du7OLHHy3GmlrYFz
lMoLQZnk/g2rEFKPnh0bQndDyfJpCZWY/cJWbrxOYuXhPy8vQd+Atrt0BbNaacpdp87X7PBV+AcM
BpDB+qMQXvAEc570u/1iA//DLLCNZH6s0IFxf7km6tRdlFUh45bqdXAFDv7EVEN1IJjeZvd9fY6k
X8mIuo5aBBQoOVZf5s+9AkQHbUMeOX7TbiLujK8tJ8vj5zsy/rH+JqXSzN2drjXj2uG6dXbAFyQp
gsGvBbNftWJdWGqdnlR2POsz8ZZw1iyf5JO7VfnIAtwyrjEVJPFgol6sw14oFlOKXxEW8ZzkgMgO
JwSB4BMlrF3/RCjqz3TZH6radigRAAj/YPJ5fz2XuD9rl+5Kbfli7RxcLWhp1XjTSOhsD8QGUnpB
AwNpe7PJUnL61ymkRq9evorIldU0wTr4PjS4jfzp8+ViIN00n9v7665iRDZIDYruLbXEOLAao6QM
Bnq0oJS84ZHPzZ6LlxZ/AOuxlmj9qn2dm86X75jUiVJAzJ4Mk9hRuQfdpeLP9SocxyvAIxOzzpuG
g2NCeV779D6ZdZ0BtTw8DvcxIyuYx8kREMamr5kJD9yBODnCMgcLiT0GMmCX64xAv11bhkEwonY7
oMqcg7eexG8tnOCcmiK8HGzeSAAjx9byD93u5MgwFG8fY3jYsm65BlABN7cIV02FgF8Vrpy5X7WV
1lzIAcR9MUe8rv84WUlz8zN6qs0uREVEIbcR/nv9LFnGRejTzi86xqVSSzatz72zJcAKaQulRXvY
lH6EoyAfehhP1U5zoW3uSWbe/7L9mLj68t9qF53XBdGJFC9SoMliWXJVnjB0OZlYwNIRJQEp8G/u
XTUvpMKwvbCiKDg7bLxW06zJyhu+w8qAQDq94sYC+/MgBSkslGnJ6DdzgeDm+VE7K3j6FNsCgthN
ji9i6Cz0LM6kQ488RLaDBuC8qWl5Ffgki8e7RPnYlvhPD7FnRemTWIS47FvJB76vF3/7gpyW+T7j
iB8hoP0TwDec/yRCxH9dUDK/e1Txkbxbe8Q+1ZmuD0rHiRlQwsRzjQhf3VfvkA8TqFVZNbUiRhkW
JYwS8RkokmsT6fqBtbRN76GbE2T1NWddVgpBd2iaT2Cw1kV9Z9n40pOaKMMKsAFqg9llKkxvfRaJ
mP3jK4U59CHLJMhH9GQ3XzHKAKpSzx6CMbV9kzo0w7JnmdD6hwpRqBUeCtVGzSF5W2/UoWizT1uV
JXE2C/p791Xhhn1jh9oNAFDnj7ftpPLyODP8HotravbG+DKlBcBgqCs3RB1SW2hKUYaGnLKwtdpm
euUR8tBTqVs8qoM0NrmRi1gtxnHv97YAd+JrzZ50VmeHt8OHIOM/8ErYw0t/vgfsCBfekbqUOhah
8HkSuyKy9KHIf/EqUZQyPSj40JxZKV1vEWnx1gsxddb35ew3bygTXVYis+69BSkOgQkyXTqv2dw0
Pblnw2x3v1/pk1L8yqB3kOHhLfqkUlZJBSdqF6N13LSwkL+kai78hJe31Jjod+uy2kbUICMXJlNA
0hYcK//9tQ5HgIksazL63awKVl9nCuALEtvIwYQbqbFmL9BRAx7gxNd5t7pVwnLAMCpFkZ9wCvKC
R0vK/sdVq3nTEjntmYs7iSeG+anOyynmE4+cHnLae7sm24LgunwHjLcldMSZqmydn7koAbcYw6wp
xIVMmQwfEXXCCdVBQbDQuaVcr9TjvHljA7vhY+OXfT8pHAIoaDjMkDcccouUB0pxm/N6iEBs+rBu
nmUW1YHQw3OkWhMc91iMFYvOxPSlTbX+s+Qv2ndYEHZ8vKYsrN8iWuTyuA0Sqi7dyMGOaqsFtrbI
efY0Y1Ue6BL7tJVv1lwfvaO5b2/faIUEk/DL7R+xbAfTpJeM2bTphnzR0AuBPrNbhaM2KrECLPDF
/s+3jYCsTH5s64HDxsW+rFq449M0F4UxSh9TpjVZ/Wy1LcB0db6yikFv8O/6uPFKKUro+3nQMjIr
45qqXojcYomWvqPoqqSEzpd2dG0LoZyaefBabwnUmP1gHreT2r92CH4WjcZj4eqyQLjeUs3GWm8Y
xWVJl1e4KoCxtAztQqyhQZhPznli+Ik9TD/8efUIO+aqPoJEHKvV9YI2dptW6lsTto+9ZwY0bVfL
34I6/W08gAPgy/eXJ4DsK8WKsVADc4upCd8r510agy7SW0hDHuMuxQdXfjMCbdp5wfbWNt3M6LJX
Dphy09f59zuKQZ6zD4vfxLC9ZN/EOCXVTU+rLfZW9Mdkiw5e0HDCLza2sPIDkeAdvE8pZBhw9O2x
DM+iC1c5S8GY/hINwBOrxNMCkahvT7RghetiyvhxIwUtTeGa15qmg+SBclN58L9gMi0bSdff3RC+
wQw6c0gROzhLYBzq1lZ+nAHJNLT9sUIrlQVsRIYuI3NVk4nk+IKt9fUwtywF8B/iRDRwDw2q4vXX
HBr76Cl97g3pKYgtI0cQdDh1fw0tUE7sePXmGPmqmXpaKVm83ZxUV2yZo497P6aC/RQ2mId/xZOC
VKcY9MFSWjtkeIKkSa5shjdfBEyy91RK74jdDOb1VtEt1c9eRwCSIsfEPtoGL3I7d4f97imyA8cR
ojHk+8uMEkYMBFbjUqXljoAcf0pwY0sE/OvuJ7s/W9kEzxNUR0eJF/22SkMxcqpZuMwm7C/k0Bs0
CN9gdE403ZVY0nciE8mIM+q7wN88y6rXVUT9RAZTj3Mzth7lLLXWBnsf+06IAKt1e2ScnG5vYtif
bCPxLNEQvVr9GjFe+LyHzVjwIaEQIDPc9Qg2Hp6FI2wh/Ppn1nq16E/ZpFfyuXiC6JGGJBDDMZoh
OIa0RME1WHl9nUAGY3DwwbeUtSvv2ISSyTOX4PFmotIBGbQmt8s/ca2ANQ4/hAevlezVEVELNXIA
yXN94ukMy6BNsuBEejd4Gtu5AQ36lkVM8c3t9MCTIMR9nyI0Dqjt0JY97EGfF0gKgaIoHeTHp6IU
UHcMd+jyaB5teQZqhszoGhPis4jMTaDNHT+R09oM/9IUZ6N89bJ50syEkiX0fnVR6HqLw2p6UfHU
gNmcnI6gz7dQ8jwBfuCx9D6IJj47YwD5o4lfMETh1ko8A98lLmyL/mi0D95VvOtZnSC0BDygtG1W
lvz1H5aYy9kKkBDjZ6e13drrmG0ySTIkUWQkM54T6gvi6JZAvNk2YdNG59XrnIabggGZCeOzEzdL
TZ/QFt0S5efhlcL+QgLtoOS9zUqvk1vOCne1gSfV38KVcEZSImTvxl3ARS6i0aSYvGNrz3x0QlHu
q1kw+X1kCj5gtKqrwgDKtlVWTnSw3d3jR9wETZwSdQtTwoN4UnFx/RGtk+aOef9R7SkIZqpQkLoW
nz6L1dkPVnx1O7QzIHhldQ93XaYgV0AAPb2jCxQoK/E34+VDm/Xsan1m46pSJ40f6Kgfx52rwluw
yNfR/MJrW//OOGdRiRyYg09G7d4TeNuRJpd4y+rlkCzgiRbbQNhSAmi+uEi/C466botPdwIjh8Ul
81nkgDfRmA2VFqeCxugm4i3HSYOiAkuY/XvMAQIFCRSXlRj5RNRq0ygAmA9Pf4LUpPCeakJvBqvA
i9WziRgZTNaZ8nNB79rvHZUsWDwTlu8cDXFdNodo6QVDXLAu5CuXi07L6+QML1TIIoLCQIpO40W1
cO/5CwD0AUvu9JyvB+l7ivQX4mXe0G7llJ9B6T8QyBrGytWhoZBqo+G9jyJeUzt/oCY94cS1uzI8
q33WrUH+Y0qr9cjjhA1mbCJDPCVn++pdUGJnnL2vz6SG2K/qtLsIu9GhoqGuurwXA58UjXZRMCrz
C4w3eyW9ClT2+MO9cdLi/fPRlqI0pi6G9IdrW5IoeohVkUw1yZgsHn/XIv3KMG8shLiZqxHw/TPA
c50895fV7T7YiwThHcnRBLI2TcDkyx2Zd0lWhZt2MnjoYpEOKJL74lGKA6VaLeRbQuqkXdfRbdLU
Jh9NR74uemwAp2QPTFeqWqCNsIzKRpqeihc9iUg9IizLg57drPg+7WSpglNIAv4ykS0sF1MKIwdI
HUxaauhMieT8HT+4mOcLBERnThnwG7cpT+x6mzc/nvr15g6meGK4pphzG14cssL+gAja+pocQ5RT
BzrrUf3+VEi1TYjstFhIza6gJ1uTKOmHTJHRWSOd2xLsTpKG92l3kki6NkpHEsGwnaf9YTPo1RDC
yK7Skh0ToAKQCu+GnWraJA/7dvSMO8gAr/WqZW1UtAYRWqvIbZQpT0YPBLmtDlLYD99MN+E16J68
UXiNxPDdS5Uo24T6Olkjff03Asy6YNE5iM0elnMdsao4YGOWXQyhzxeT/xOd6mCjtZXt8YaXPGAm
Wl0+1DWeex+WO0ErMfF07ydAAx0VSV3vN/zJ24/fyciOb8jWRus/5ZkehPZ+Dg8AwrsTTCRb37HM
3BmUEyv2hAaraK6dDADxlA/PCkrwGJx+oejFXUueWVPbhNoaCYQGza2JYquz5V2he8+VghTHdSlC
8NdkntCyrAx3cFRl25V8AiFmhfCmVf+cp1XYTPF6RhnIpgyNsKuY5S45vH9qSK2HmZWeA3rrF6ue
IuR2W5o/p90k9Rmno15pbQrhRAocW79yVUN/4RF6JDlAxwWRbjU9R93F4OozTvRdhdmAmJVPB7bP
GoHj8UuIev4TsA9vUxx0O3qobqg+7jzhtYDmr76U4/GaecRarPQGPIOvk87mmWcq16xGDfB0MFYv
HbY1gcpUUISf1pnRskPxa7B18i9qmg8EV9Q9D/kdTxTlxLqqootsHxzQjyfxzO5ZYKAy0KnrlkJg
wkOf3uqreD4fmdteV5LxvoaMy3xPA9EM/8A2TF71p/bAnbHjr1sc26oNuTqpu6WRwQMOxriqIh0C
GhAjHr+uiDaeZG+lFlRI+TiUt2w06b6iivf7TJuW1WDSqOmb8f71ZIVmhMdMh5jDmAdukt9Radsn
4JwV0fkrH4o6K2MANYE1PRTDygYsOHrqneG2awbMuIWtVYH1wa9e0bhjI6LhqLptXo+Y+LNPcgtj
TU31DZlTHKLZGU9+RZ8FWf8P4ayNT5p0LAm/zqs4TXK8eFbMeL5VZUqCF/pK53iaKfQHxGDa/PWP
iNb9O8N76PQQS6Yd4qDOV6jhbg2a3wz8RSqkqAdtQsq3aqjdaEvlBeqjmW5WiqqV+sSFNkDnKU0L
CxGOT8Te9wJR6dAlDN4NivXekWWglsbd43Xa6PjDIekyUj7uwm8HHAv7L0iggbv0vfXMjVIBzCEX
6ChlFxT4iNtjRbMT9xRjOQ0fEdoC/8l19Oz0+gS0rwXkqZgrQJ62cOrtozC/CJEQ4UhKrWK8uGzQ
tdHak+KBbtRvQ7Qep8385o9LE8vjAt719dgLjHoDfzE2X9dEjidMXAlm7LuDmEWP3v/07IhtbK2W
eoPylMMGU1WvHtp0ZUqL04kkPwgab+zb/dFSfMfEu+sxyjh+SE1CRZAQs1RGbujajYycccbVyupq
5of3chCn+rExElv+q3Hu2NZG1zSZ5sT5eUY6Bb2ZPx7Q5Uew0luYhwHDnfh+nr/vGGFJUK9aXqDG
AKSszgeKPCjlJRFUaDZ1nEw4GHxxypa7N220hKJ9gdfNgUkM24iMC19Tb0+5dn+VvYCLgXkMECcB
rStbWUojEUas6bGf0SJI1zjZMEzsrFN8MZOc6EOp24a+luV70ClZGPY8Mzuuu7V4Lx9yCKsWpAzL
+T/ZhDcv6JVilOw+ZAeaubKxQmEijGdY7GdzWBrxdLGS0dsmAKK20rDVKOIBtMlr4a5y55mN15bd
OyCIl0CXhiuvA5AS9RqWXPwDeolhmHvZHabHhpVtW2O5AtyAPiFD2J9zXsMy6bZG+/pdAZn5YGxS
Co3jSsYprJyPG2jO4PhTaknkrpiw2OPc68SHKV+RClaBwsVoTpGZ9aAhV9LdS6cA9GXoOJfX30KA
L9vWZ61N9Vk7fEJNTq9ZYVIWwCiDJYfiK14CO/mG7zLjyM6uOf93NWqLWuXZVOE+4eQ4cpWA6H5s
OG9+D7yWypXTFfeCdb92KZ/Ev0x3yWbNlpHOdMoTQIQ9e0O7kz8EMiITgHYi4E7K3+3nLyTpYLbz
z1Lun9lC0a7ZGgRNZmGfOZpApsx9HI6EIEtO8r4FFZtEbZ4IxAHHQrS+5qg1bVmrhp+QHpHmTNVA
9FpaFFTCLogs32GIoL6cIA9Vqa5SwyysVC21wXYM/MmZJrJwTro0wO0IgzIr1+M+litswuj8H3zi
FiYCH2ywEhrZVYM0DPKSOdUtf7JnqYuPlAPiGnC8yUWEq25b/YHjhu/EqbYqDztLO3P8y41VkUxo
lp4HxZZPman+bTr0olUYCRjNdgI7kIexn9ZD39hNoaUQ3PJwtReiXP5x7Swb0iqRPw2/mEXDkepS
37GbYA2hg5njT6WBfdkha/E01Sck+7sma5eJWaYh1pnA/aJYypqVyVRAed12TWFQLumcOJ7PqaiS
ez3J1nH89lPUMnAfj+f/gOM2HzMMF5FBMwiQ0Iqcg5hQhMySmWldlFFNWBB2/CYJGxR7t5wvaMtB
OYMLlEOGNRCdoxDCezr8HK9oP2sVZQyKCenV7BcAT+N0P6SOMqWC2Ivb4J1kuoqGByQyGUwHFziM
dfuDFpGDKOn40yk1703nByND+xOvH7sve2UIfqCI7De777h5UIt/KeXTvIcTVvCGsMlR/jWVUkMP
9Qr4Ncqw9eUMO/ezUz1uOlmh1iCUnCh2XnL0jZAPLx5wdG7wbjG+UJ0K2gWMzFzOpvwnKs3Cr+DJ
Tm+LOOSi9H4QZ6wlNoF43oR2/TjGdM0P5YCJfpMOhrhX6jcKyb0zUpNxc7tXAx80eRkMh9mSPYpF
l+Qd4TOuBgRtcV16qk7CN7m4L0CEAgMZu/ACpnktIZy9YDiA+SsMTPI/LL0ubiUkssI+luYlBir5
Pce+KmGDbTkjP76oPo1uDM3SscAVTjOmsvXb/yatKpVCWhZ65XCocXxT4BOI5y5yuI1aUEIJWwye
+6TRNQXPcA6WXVI1Uy7qs3v2Rs05wPv16blb/OyoKG92tAIIyCXk4P4dqz0kWIQFPvgMYcZVk6KS
avtY9gYMgzFQzCGV071SRumzWKxGEeeHR2chWoQDV//KdmgWrWzCE6ejPxTWhlCEYSB7nTOO8mWm
22Kel9y8QMEkFHOD/MNfrnOVeCR/+oTd122se6/e73EDOnLRJhjs0LXFYKi8QROuhluTDEE+BhU6
GFZl51mebsi91SGWftGnfE0a4S/RaWK2q3SC2VzpqI7ZI5DCrwsgIixnA78rGv0Cr69cXjzl2TMB
X9ff+nfyomMB5Z/ZaMbXyNfYKQOKM/uqMfTqgTv8WnIj/4q+PLFotoaOIAsVHB4WusZVP5MXigqe
RNG9Z1mC0IG7eFATgko1Zy1/RZXnHyzCLSYRfuAPOhRyyo6uygDd1ifC+p0okyF3LBW9sWlNeasL
jzKruWjBcBek83hZ5sdXKAbrI20EKFN581S/vzNsyWEBtxN0LJjJIdYLH5Nosoniwvn2VNnzDtyk
2IC5g621VZhEgUdhKJoUlEgUTtsL8IupA2bbJy6TCn1HDHTDyyVdI90FeNmHOdoszmXEsEv28YID
O24JxtS2KEtfn/ZLnKsf8tODVOG90K0P8s5Dpnd1oimvPClmS96DXVYLf1ukGfNxgigBmMuYsx7C
EkaKjaBr8MMiBnseeiKKEMEwzkJOc4bLju+uqBe2/Faw4qWUXtxaYAyh3kLxQS95t1QG9LJb8BhU
0jOzGS/z2A65hj29AAAwHYC9+oqZngtRFq3Fz13WCpLmj9C0G2w29mojul+mE3x5O1Qobolcu8Cq
rmw539QtMP5f9LhlqVztZZlUbQmd69TSEpSbDDomytyFrpl52R4EASdePyN/0s/wGe7z/EyTiHrE
QhEw0tjBhNG6fHL4IQqkJcU2bdwPmTRVslcalvtP6EhP5pwgBASEpEV4uarHYHRSPLmQ6G7qnXIc
yMzwTlXid/uosIte/aviQFeqiI7Ik2i13cElIEd3NIIXWkSpeZAtDzlHS4daFq46XX4V/hjT6304
l/gdu7Lku5tvqXZNBAVZC6T9gIEPigMCXSpkbvldbaj8hTBXlGbcWz9BSgsx46gjR8n5NZbwbDH+
yauamfrO1KvDCkLWrIZy6GukmfCphRRvw4PcAmWsDjwfE21F3qck7egvNbqGmgVUehlE4edrI+PV
V/4u2gXU1aFmbAh4eVcQ3QMAWT+HTxbU+J0SaBDV9wTZlaudK9Ieqv5nc1BgFy+4GIwpuUDlnHxr
8pdwHHkWWD79vYxlA5iubjCXiyDJIwSRNyP1QCciJ2/haOS6YEjjMf9wMWWb8Dbr/fDARq2g545Q
QJpyZPLbBH8Jtq+JLDzyStRMZEDLCZeUtBGlhmb1xLfrc2qDMsswWchQDwYossfZ9h4G50rIeSWU
ftc0erRgoXtaOGBEVGbnIBZ7gE2HE+i4UiLdLvnAxpK0PV7NTlZnDa0R7OOGHAnH3y2h6cNDNJqS
RgphOMoDTa0O5IV8GuK5iavjfGAzaUSxnUW6LneFsYOmTK/00q1R3M7zeYT9/FgHDSIQtCgdYBLR
6DTZ/rPphAMRc6gHk5kaI0674/mBr0wIwH03AooPzTFxLfDWol2G/TPGUvd8g7hEtGCWs2KB2+5I
5NBkQ+NKkMmYxvezotuCsDRzx7piv8TCQ/eh9qdlu3N1G3kPZuXk1y/xPW0NW0/yBHNWfSArKR/v
CPTm9vqpe+q96w4JHonxN7ekX+n1JRTOEI702NjGHqC3O+N7o5XLpeySQcejnDzV/iGzXQZB4Dxj
5/SfTnvpqQOQ3a2W6MfVUEaCK/EACZ1eOPXW97LUmEuY7CrlWoSj1iAi3r2MM5xCfsnZaJ0a9LvR
U+hpD/CkrMwcFQ6FUTJMnUoOKnpmXY4I9YXAmjP+kG52leImWlB/SzP6ReSX6LUVpWFnWQG4P9IS
E7gMpxdKMGqILjuBjs0h9MSut/dO1ZdWD2pkxdPW/fXr66DEKAmyHQZUpzZqZT/dr9EKD4/qwHCC
JuowaP9gZUURiYNmFYKXwT7tjuLgxlckTGBZncnICY56aK0GBcFeLvlfxrr+zc6f4uGOnaFNVioH
1r92zLDD/v+ZWxp3UvjzxjOI6A8nFf8q6y535FV24iqv5OdMnbY4SNrz70v6rW60WMLmVew/cqUU
Pi0x3HM9gFsU6I+KYNpN3dn5k6/PZZzvlsGF9y8aB60w4AoQ5F2PePzvxK+vEr+66DKPfSTwJtde
lqJPHUdjKB1HuAi9qRvyq2qtKsOlQVmOt1SmbFeUnvYfLv6wg7FnkQcr7nzLzQ0Bs0Mpm/oo4THb
V0hD0RSGwX2Z9P69gbuOkGP2GWPD3VguBxRPaXXBkcya3EiP10QD5KZ+HascC2ZEVICrhS9GWl8Z
IChMLMFK73q7Vtl7DviKi3Wb1s+8xPel5MfzqxC35gNOctePK3Z16viUr/mx5IX4Ajad2+Z1w5cQ
juY4gVAXWYDYQoP4EuthFQndydq3xQq3Bz2FunrootpI2dzRzwfOZzbFCCxAkTon49N2QxDk55Lh
u0g1Aap+mewTOwYmXJ1cTO5HjIujakmnefyceEiVGlsxDrKFKDi44HI3K48lUS6AnbIuFDJLF/7+
KoOCMDlXUu5Qpnyse2KnQ7wz+sj+tiHQRh3RlK/q+kj1g9jtnm/6CbuB72JLW5UibJntek3eYQ10
UAmzrSunLN/wO2itxEsVNhXRDbsdhHSQ3XoD/i1QvdJQbwi9NhEdFjRXGY61o6HlzH+Mhmt72BNr
/fcYuev2Q5dIkU0b4h3vkM5QCIe/Z4k2bvx8NUwOTNgtafUZZxInm9gOYqPCZtyCaBTg/o2y0zAg
UxxLUbdj8rFhF2Dj0FakiVJB2nUnw0T/Uyjbahx1HN+65WYSXfNlCrKDDbjW9teoBgKmuCx7L2EV
RpxTD+JhBFP9a23sOByIragw6vE5G0l+iPZTiXyTbjsNA1xiZdutIYrBnBr4yLE+f+XD3qGszZSB
6uue9BACAPBVYrLwLM+RApsMYWv3VRwQ7sRGN2DYskRC6rJ3iNuoyaPGHs4cBc9x92xK0UWY2Fti
3YLS3pHJ3tywwHM/WiIbTKjKoV1mMYZwYLkcv5xgn6tQ7qUFz84DWGYde/iB6d4Z8Sdtcovs8ve0
+XONYf3t678Fr8DAcEO7YN+K8SIvNc0QC9RmZ1zish2XmwH09mjZ/tS02WwHiEhgHU1ssiegzevX
NWk91JmzNGjt4f0rR1irP3D1UYgapT4xENITJ3O0QB21rurXUDnqPybUVt1id8GbsKqvTj7M+O8v
db1ihneW4LHaHfxQJMbMHPtmT5Qh+No4BfpjS7jnS+CxJumEbO/GZeEwAipQC3xmaiBHreMTdxpc
vs3t48eAff+K14a5nxRiYCbnIL5KWws8nSKLCd/6RJVgJi26/5yBmvWCppDGpX8zXXKWSpxVwNG1
Zgd7RCAgTKl+9V8tltPQ7iTR20au5z9HSrNT2f+hsbJFX/QXyJhNrCUrXDVKaugH6i6l1qApwc0j
Y+1yj6lPtrPfM5kF2T0VQ5oiK8B5P0BDxWG37XJGKR9IQymPeQxVcuah0FJPy74UXKo4pnrgj+qd
zzaVzbj+mrIWXS0CVl7KdXf7mmlKLCpdpRj3TOrpTCdOZJQS9I/IFn/HgzyNDOb+pyEQEU7iDMeH
eRn7L+CiNWdeNuY7dkzuuKYDlRNFzIxN8vIZtY55NtzZe2WdO/x6jysq9xGBYe6oe1JZbB83ltkW
ogNhFSH/La20XBs9yzIOGTeSda/XYMQis7EuEGiOqujLYwOX+9BmQyhEQKmUETjnhw2CZaKgAwc5
uuuAuH3Z+dKEplUgwfLIwSOA22b+fQEcBDGLPC6fax02GL1wI6LjZ8hz2UyZ2ojcZ8sJUny8rTF+
fE9dvhjuLxXQi4fJASH4DlPSlLcPxir+8ebFfLDVpQVPtn6E5AazBThZ2sam+fqGOVI639de1MYX
gkyho2RsuLzuEtQGDrNlNW96RqrQEccSU8+Z2hlo+kCsaSArSMZ+HmHLpNHdsJ5axlwMkaGMykNX
iAhst4MNIZbC/+yenoJeaJCXC3OMSkAbmeXYo/A3UsYyIjoGgIM/imintVZ4xLwMndKB90PVvES4
IvaU33b0QIHafpqDZHBr+el1tZ6mibUwUaIW/FjgoRktsTbGjVMHjWFuvjaYIjWR3LFwmQRJhpYb
UnN/KXhJ5HkQBMeoREQ+fZAVhOqJSXUlIb7ZFTkKevOk/PWT37nZLVO/k7EDWCrSOcPrdhfIhdhC
sinmIYRqptR4a10ERyn49E+Lp69tfmWUCdfdrAsqMOU4TUyUAGTPEl++gtyBoSd9Pe5PWjSGIqn1
o26iatG9sMNPMeSU9x7hUucco69DtZtVyFBhVCOp4mI7pJxzB0mmXfW0qYM10m4DtU75zS56CYM/
3XSnwf7HfbkgTS/33NYhR1VKhxppPNJrbkeEAVjbtI4HkhhBxHg2nZuf7wJ5p2pCK0ngvITZZwua
waB95s25X2lQ/N+3yTbvtT1tnfWJEvLihc30+Mc9E4nKrCAYv8/NKkE/UfRUYTNKQC0gM2W8uhnX
eQuy23sksoWJbPgOSrVek33QozSCHI+RDWkSa2svS9bnt8jYAJJQ/86YWp0xjNPDhja4aYtO54TC
e27UxewMlJy3KVEEdN5dVo+C14PUaYkBRXviPU/F5kDIZ9/xYM3MgYOrpztmpamV7fpFsTFveZR2
q8LWLE9tV0Zt2gpQB7qqNk3aqkaxJt/S3B5p07CVqV5LqmqhXRGMEpmtZsj4HdXLvMvVl1+wtsSU
YHs521DoI8X9rt4eQVn86nz50glJRrJkgekRFpkGsiZcaoGn2KikVaY5ZEOz8r0bEENQDZP8ohTn
NMNY+8ehwKNODBbK9FHi4VpqlooDMiazolYxRiqhdR3J7DKER89OjyPs3MKdW8tzeH7ZVkpn/4C4
FoazilZhSBgRIxbc4a53KP/NIDyEu7eft3lqlLjnbaS2n/0HvLKSScF8rhYUuiGrkngYpRnO5Iyh
wIbdJI5Jhdtt3KmMk4jMEO2gIwDjCuu9FJSnvmwcXghtoxqlNEti6qt36Sx0dIYfXq+pmjDqbdjt
BWK/ff4vq5iE/0miel4RFHFrk3IugQuGIu0Ty09SO2n5Sw5I9CTcNi8pNznGaAsNE0apJUr4crII
Jf+/EC3HMok3M0e81sDN/9lEcxS88UZld/lStmejBkj3hpY5nhTCmi35n6MUwhSRYmCM//hQzIE6
GIjyJZTdGWm3SGzhJFSW7R6dQwLfXLLynTFK4RqqL5fWACvscXP+8e6ItbH9FJOzVbQAdxByTKXv
BvrDzdy0UzgFGgRkyNOlKpAL4/IshHgmNJbawMqSFK/NA7Px1jprFSy1pcJOsy3pFYCuaTXawGQu
UHFhVUe7PlBPeyVnoQrlx4ZS8vA7r+axhMayiDMCO+wkX3ruGrdxz9CTpXL6wUBIiZCa8UipdJRa
fEM2zEss+0/HbhQl2L2Nd7f7/FtREhMyWC7u+eiawksyEcrE2zCX91uCyA/KaE6n+673r1EcNM8B
+GUKH5lnlY1vzSoX+6x/CjIEKRHUYVhIDCGUISgLoI7IsRepXuN3ywqTLcZd2ysLqZ2q+vVZGDGp
CyoD/yThLRe97a0cLq7Fmn3q8DEaRBb8yOiDbq1apRQ1Usv18d2U5AGqy7W0JzUX+YONcS5asqBp
YQXA/89KTuaMZ5ULo9KwWe+i4KkNKBwgd898jx8SV9zlMjko99EdYc5ax/YjI5NPSjydfVP+qK/2
eP1c39QEysSWtBcsLj/wz7qx1D9iKnuEgmwh3Y82GI5O8YzmiJrqVbD0uIpjwalLcyMeJsHv0Uw7
+Db5Q0XoCZxOwPQZuLHKIl4kv6aIVNpFDBsuusOp+xVcmlONWOGHWlMRMswlb7Irt0VBpu2hbKlV
BouDopjEFemJtq6P8isAjgQyfFVReNW8emBPOltgjFmpsg7nRsYyjxhzhQGjpAvCuJKP2yP1cxqF
GkbB7dSsuyiXa5EimFOw/7yUOHgY5tT8i3RFzGxY9R8BDOX74X7BiWJY7nDzhF2EjSjH/4I70g9O
aXmko8U913xMV19BNj5BWosaHSylPuwbJSGVXKQlftpffQPCUPdeC3RPwXfJXRpl7s7Wa8qHKyEy
xD6l1Am35fyz1mipO9Q+BLjnOPX8RIdkoc2v2yW3rpJ6s/zXvLyapndz2mJTQpPGXldquknFh+CJ
Ivzx7VKMnaBe9OSbdlqdC9NhJJXfrFb7lJ+EPN43QoDkYIDIU19nyFNN7ZvtJd1i05Hw9U+a5YgW
B9DabuBwUlkCnIWzZI9mQKaJB4Af9zbzWKTTbKYSON5rQrwJ2znJqDl7TCF2rPAZNeVw8EKhwDzQ
AHTXe63EbrjwMnQ9cILYh+dbgKT8mfDBGCkZndQp500ywIYVk3G6cnZlyvF4XGF9tbZvItiJ5vHK
4rnktzElPO3Tgz5EYj0RIzGTOCGRdrmp+Y/B7/51t9uTjOSDLQXJu5pOR5fr7kxLNrhDLcVncVm+
Sf7ppkXc7op2/0poDSunVyRo4SgihfZKXuc4vevUUnBamRzYKUxlI8xQvYyYOIGcP0XfrqA0MWt8
mUZlk6IfY45kILobbr935Awp44LY7hKHD9t+SrCSxYrgIca6xPKxA/TxPH5OGdFvwKm5KQlwgVA/
kObvO47bUV1mXO+rQAdIf46nZQVgLdu6HguPYe1RSH4fyhLRiJb0pUkv4wYueD/4u6Iyfs2Iz+A3
DF0ni8VBBZvfH20+V4SDr2LZIit6b3avnyj6LucmWFLaDW6j8Q7rP9x0Ibr9t70KtQT53h+/e2se
e4uYX1yHtKIBrv4XxwB9KfppY+ZcFH2J4qPr1txVyz8TWxrqo4Gglgv8J2BRDqCvA1MZHecsbWOq
Fv4GGWJdzW/Y+eH2vdqexLa487SM87YIMOOhA3aegCV640HsfcoQeeuEkpT+sNmWlHP1uhdqzZuR
uCGmRcORVlZbZ1aGyTr7b6SQkakeT83hSSNlPSEqFqOrwlpPBJpIrXEi6gIGbZ5Nv6zswXyTmEId
Kg9syaYKbxi1N8+bzGfRxfGMGjk8WQfkKYGJieDOiK8mX9eiYuJ8M9gaMYc/hhIZkPvmMmD0Q0Y9
/wJEVzenLGGcDHnKDXyiiYrnrDlNKLSLpi8NFelA4qkPoCKUfstZkdhc5X7zTxQX73hYpAbDWRLr
EFLxvkSKWPbfsCYT9so4epzerHhs34ZYROyyJkyFK4q/WTE7MICx7hbqtGEjc5rzD37F3UDCNCyH
D19B1CdcbSDG6KY+5e3u/I0Fq63p0RKwnC4vU8IBTYfvhXPlthqmSrFLfX8km1sGQHu7A2x4kmAY
zBG4+yykQVJCs7KBcWWuXbHL16h+U3hRYdnJ6SW3hCpiQd+MCYEpYqOQflknrxzo3LM01zBAPkCF
Zrh4BPNx4CWQiI/M75Yg200nWmhJqDsvunclB+fDLR89i86TnC2pFXjgM7EkzVna1/N/BstOrzO2
tHo+6pwZ5W5RiULE+M+jopzRgZyGkMAlTDo/i7cPrF35VL0bzM+CvJfh+xmMsGlZfl5jePe/OPIx
vPTbE9Dx7veGJkvFiZ1LYD4QZM8ivg5IrTcnweWGCWc4Rkz/zA/Uq8sk9oyIJSwXtRnu73f44PEW
f5oPBCzim+notwc8ThqM2d1/PR/dlxFL4Jr5ezwXPK2v2d0Q/ZWpJXVbpw2ekNNwhrFq8jePXLBt
wBywtxo1nIezqGTTgVaOGZNaSibnlRO2qOELnuikrvjmfxxptSa73ICbHJzjMgm/cf5s227yD79P
oQAZe7InNP2nnG61xAQ5yEujqkDmJ1oAbM+mx24ybx8vZzZw1BrKsOK+W8h1b6qfgXG5q3sJle3e
EJDEVLAwXScDNc9d9IeYsy+3u0PW4+Qp9VCcmIALBVtVcyacpnJh8uMlfnbFVNRW/cSvtep68sIV
tXQ4Ej62Ebrq57mJTkNtCL1jTVk+fRTh0JzXkdCWO3F1PMyLsaui2qggEO+HH7iM4ncdo7M2sxdG
99Ss8KGd6uj5NF2xddQoe2ZodvkaQmV+2fjsVClOGUvLD2eDgXG+dFdQ5WzUzVsi5yAckP1/ORWb
MixDYkDZWHW4Y/wR2riaP0TP6dgMrwh6mvT0I/GVF7GzlZEPgWTi+IxKVoyv+grr7T/Czk9Du3k1
oVlc9tvM3Q/dlzXdO2kEiY14LqnoshbHjwi9GP6jvhtdvNxvQ7v3kdHVwc27/kTSLyvsvDZno9+r
fvT5u3TCYAO9bGAK/jD3IldmyvX+skmL5uTGxi+R6ieNV1AbRQREWOZ8LKTSAaU3EHiem/aSXruP
ElJ87xhKWXxzIcyYXJJQeRniVnsJm9+259DtbjJxAu3VCEamORjZ0Bd5Bx4HAta9Ms045MX9MJXM
AnG4GRCB0CXDSnPB9GOBTQ8SiySX8IlGXr44zMbbwjgNGXyCFw/2ZY8GBaxNg5bqj5szD5X+uyD/
FU4oGai+JATwpBm+Iv0UxnJTl8KQQr8F5WgFffsgIRJTXJVYLvuj9RELA6ZNt2+qtxmnw/vsmHIF
cngTJUMlEsSID/ZtB9WyPj/qFQeeQHqHdAsbFhsPxII2hZWhk+DHvuHW+NQrsCNQRU4iPYad3PaH
EnXeVW8jLR6LMW4sTEcsrGdFAIv1NYCaLb/Z6tYgyXbThsyA+hRZQ/qe1fT5KRm4Rz0FEILMLa8c
RCzsO+QUK2JGUCWsO6f0RIZgLLKwbbbhHmbqJkG4LRV52eztXvZUmmLSWHdvLGiN/RgaauMJW00u
xrMjBxbq1IISmMqk2UmOVkOYdG1/rcr/mSfQ8xX/OwmzQZTMU8nOfMFTu19K9huP6oV83It4u/oE
9X837BxjBSE9awy5cI8+1/kAz+GyHLuoXRt6u4Jk8cpaWDAUVfBFXgF0kDi7NUOLT9iS1OQ530pT
uaMnn9HmYffL4QMEqjVx+saM54pI2kuhLo8gqBCkn8bFRBNLGHqPc3Nv/UUSMgDxIW83VddFUq8z
NSHkoJWkdRxXoV6rCJrDOf2gLDfjxJC0tJIWGAAAgBv/8f+tjb1MJCkHozxmDTGV1mz4e7DpwtqY
+PdHEPWaZVQB3XcjWe4vp8gcZl4itFmbS1GQ6esZcnuarljlf6H0f5fq2xZdCsw9BTqj06nnFhkc
jEKFcNHduGMO5K8iBhZtCTHz6rxtpFXdaW+F+gV5eGZNHwbWVmmiLhZBHEx2ex6YuH84aw/yq60Z
QQtddYCc7e+SyVws9RuPhFyFHzFAMss19gJXAjoic/UpmLN22WTxW/2CV8afAzX+B9viUPUJUlIW
ezpi4IIkqbkK2ECw4MGq7JT/1wpqfszAw5d20vJRLvAk4yg5AGumlAFESiosrt7STqOi+9QD/Das
hx09mfCQP3FE+rw+DlGUecDYbzxrXZqTtxa6DCGnttVQE9JFxVHdWlFs6nMJ+2lHsO5V5lvsAA4j
p9eeQ/NuV/mkHrRCahdmsZ4l4i3dpWbCgqFNKdv4AzCX+dt6XP6y9JvH1Ut00+Ei8ZsEC4efcgQz
GnfCdSHobabeEGR00YhHbqUFbzw2Gvhb5wE991EowoXTcCxwLx6lVN6uYWYlY9FcqBent7HYGmaz
CZLBtexC+bUTVrr/c05Hsvi4v462tlSUP0psPv4Op/6PD7szRbOBZI/r3JltLU5ZgB0QhWmlCDc0
MzU+Vw8c2NxOSA/DYj+JhJij1a0ox6/Kyu2IEBZceLUjYHY38tqI8c65iC0PRzgMcMjD85QtfDqj
ldS87hdDIbkUlESHfJtz7CsFt5+uoLgGiznvm+QOpVIQz6SlD9QHqgOgkL8g6rrrZ9nWvrSvlCY7
fASOPE5u71kdQc15xZfiuqa0RmX15f4zkXKm0pKuu4RUVe/sJ/o7Na1F6PjhqtKZ6erh8+CgAX4X
xKzqFlouGA3MFZHal9R/moLe3zX+Fj0HkNBGSiL238tnz860x/J+vHuzf/FUBwsq4kHpWA7VFuDK
i2JZb3iHU+BtTrNYpMi7+Ele72ztNBcI3q6Qyy/apKJqKUY/8XFKB0ovIY36As7P/HpW/qzQxEKt
YrhW3p6nKIjwvV6mFJq1lIySc4tqQqL6pAV+osnoAGj9zyhpSs31F9SVonEFgilzPyUsuRoGBSsH
KvsiTWg3oKyq3NQ6JR0F6JLlrI+wXyAoG7Q5MCyoyNYa9INLKqwYLr61/w9mhJn14kyZfYeX0KEw
mvNeRcv7g1f+/oWImVNOdbsgWwGBf9hXmX52YKxCJqjexFNKfRdppsTZ1zWtye69it6s6GBo4NGf
SuViWr/iiQUlyhQrSN9YyVOIYEPB3rIZaVDyYFOYGq/VU6vSqnjNp0dqjRFQ4hCeMDIvk2xm3Pze
qH+STp71oqprmH0pG61x2M6r5FxJzAx6NUAKfdNTiT0knqoBJD9mecFG8ZOE+Pem/qhtZFSyYaWr
pFP8UVei0xJnrm1pxOwfJFqHDD1lquFT6UKG9glEj0VmGg0k34c25vbwRirQqfIUgSUxSVNEsMTt
d/OBmGZRYzt73HnZSl1kHly44vHNusmIoxjv0H68PfEFagiXXE4pvkABq+O400eTO4/xdMUV8BjQ
nH/wUPdGge+bwD8kBhPuX5YVJvFLbqHB/XqvKqIGkHiOGQIUxndHClNejaeD4ZEvOp+SBKwklq9T
W00PTQSmLHXO+pFMYoe0jjjlKmbwHOGHpHunyCZTfNYrVr/tkjcIkElXq57gwSJarMy49KTT1gIe
1MWlW4ZtntktOJQQCa8uwU5emxBpKj3yo8bBdTmKIhW8HVNHvGKXDIEE19lc6ssWVOlPy/yBkQ2s
TrKDkie5tpLH6GGLP/MFX7epY8Sy9a1OptnB6fewRQ70cQjjLndq8Kk5gJZqsu1/vmvI0sB1T4mr
FMxqyAaEOtmCrO8drrxtfmypkclWLwkSPqiYGLycxJhMabfZivM09db0Y+hxX3fI9lYlKGffTJYe
bYXXD9XlS4ue7SjjnMopjBN8pDq2O5HkrumWADBMQjqJBZc2hpse1OJqkTzIf3uAIFuOVPidDu8V
rdskud0BqCn4AOgt1Q0JaZMD7uj6SQjzyMMYHmz1ottn5RFR+R3xd/obKy1LwguNCOgBbADv4D/N
vCEn1AwN+0iRhnZvXEsClKBP+xCSuqlifVMxm080ln8rbrsKlbSBbYGbazelkPqwcwZ52ygIduQd
OVz7RXk9BhYlBKRXjsYcHumSr2+TEftRPbn32Jnuw/artR5eE31v/VLW49C4MPjFW/1XLKNtOxkN
wTyV0sArRhowokA4r+KHvCxhXdgYGGIMjhS3mH1JrddrS5ymxHNH4ci0RFD3xCqQekCCO8Zo9H3o
P2VCsBbYsy5rUj6N7/EPcXeKnhLyD/4I/9SbTgvOtkKINqasugy6UDkmfBMdV60TUAeDi/zl5Zdw
HLWQXV4k1GBLDeMzTlbsk7Z3TxU0dEi1z+FASMx/pN/zmjL32aQvQi/IDjgydoiYcug1PUBKqOPw
jjPmKIGw4hMpx7SV4JXFk6y5HNj5hgOR3q/sj/o0qIMBRALFn0PTWr8YqySb7EF7vy3c6A/CcFre
jEWpHrTZ/jQVpeiECtPlHZD1EzkfMCe9DOyc8JaZvpWmf1dcN9dTtmmMKUijXj+Be+bDWmtoSonc
amlh/tQMzph7uGOkc8rcu5gKQ2ChZUftlaBY2kL9S+cpTImX6G5WWldVXvZYkL5GTeT9efkV/IQ8
gcG2yYL8D1BUphncV0c2JupoN3aNZz0k9WzYRgqx/R8vvUKpiux1RYsOVnTeze3U9i9JX7i0gl1t
8HK5f+Zmmzlxah7LSXP5EkMbOwjSUZ+GBZdQlqx0xF4S2A6nDt1sDR1V8paqoYWXNB4H41Vvlhtz
4WY7PLLTLn5+BcvP/8FGg78X51dMgKoZsxhbVLX3fcMeXqXOydipr3fg+gPOawBLFPtkH/zYTOWb
uSwBWa326vyfwjIGXO26V+hIg824I2uqlgP2f7IAs7cA74QikMkiFnT61b/+8HR3Y3wOTRVCv9nm
m2Yija/B6f6B27ofnGWEy5mpAwfzbW8DuLUbRORIXuGrzLg5jaBjaZkGqyD3AP1ZGmczDJrK6EnX
1Vrl8ftziNfuGPEGaGmBYTSYB1z2wfkMHT/23vGI4dWAWaoyASDi/n9LbixkKInwrgfMqDlU9fq4
RRbcvX53nkS4gMDKi6xcyth/0K7lTZx6BzhAFz2qXpjl5BID44/c1Bn1fTV8Xi2+ueGt4MOvXexj
fqeECMYGxqrdFomEWFI90VEovvm2d8PwHCwoYh45UJEKrpgjZYhc+wBqbJkROQTd9BH9A5dCDt/v
oXmBK+LIzV1F6Ffe0GSCiEnWRfLavDrKpr5keYYEe9FJyLxY6lvr3ktXLfi0A3yR2Z1Ueru8B9qU
4AwqVHno+mwKb29Dj9GurY3JjKyYUcYz37h1x3eHuYxfiM7OFe0ygAy4h2lImhZDvZMO1ToI1WHj
rSI0x7DkZZNdUpyH6y1/SMKwlxh9juoEBqC+MadMvMsVtyRFE9lLQBfSw4BmDu/EKbGrGtdkhzpx
qbVY4PeB/+zTDtLJbWtutgQ4qx+PQzcExlVOk6VCwEnqIQjWDXOiUHakc3BfgJyfg1RqdS4uIm1J
nFCw2CwV2kVLMjj4I3hoepTpOZaax19XOn7TmlTRuKKoteRTlrA4CjsEYLKd5HeRDekZH4TlkO36
/yHpwPGAKNG0qIr7XrutYRYiS1IrO+i08fNg3OorICPjQHXZpjenvpiHa+XbWMgfgTCBO2+i0pPB
RuYmfsECVrd58yA6oPU7TF2W0XiF9X0t2Z+eJ3mpeOBBURgA0sCuAgEkDnGSf05HBAy7STrRJaF7
ahcSqAwVl7CQZCsXSHTUOyKb/GomfuQXVIpivIIwRHdI9bPDalUN8GbiTtNb2b9Kzo0xAWfc77y3
Ihk4GrVesuP1LfncWm+5Eio8gNyntrqgtxjTrErR3jc7tYPmiqUYDeyyLdicRR3t6CfzufwDpfIV
E5AV+27bN8Ws7qOu+rnkQ1dTrVyG6CvFlMeRVC6nvLLlGSNEsxb4mH5pK3cYA7/ZQXugG/diJs6S
Xg3R6l6/d5dw9VzgtLBiqeOnmvhiZSLe4+GzDm97yYJAf7tc/Eo7i95soWSYYcuNC6eP8wMRz+iX
tv9I+vskRPur2j4d/SW42v29uk5o1C2ve02NfvhHc0xAeTC9TPSpGhOby/P+lkvK47l/4G1phETP
ExCEGovDTV4C14tsmlLyAHmFKMjHoW4A7bsxeejgAJWAgUH/pfmL64bhVGRjNvxMPBB1Tz//IxbF
wXHLYhoRlq/m3lqLbe3xp8eWYiUbV7x7EYC5xTS1ywsPJvj18mj8TdwIewjUKnaoPA55VK6qtLY0
SNiwEnwSeCSO49rfVxXuOD5w4tq81JkeUxr+HeOLocXYuFvQMgd7xBRaJm3bC5ODuMW6lbdv6t/N
g4RXP4TF4Ft5HryuaQGuxnZMWKknwduAhOTM2Pvg7DOAbYKmYUxT1iYe4gDG1xejt7ar1Ep80zaR
UUq2qgP1Z7XqHsMS5Kff9GEWmvsfQKjWUQ5RRGTabgJ09UL6w4K2TM0D5NTRX9LAOWe7I/TAxFRL
KOI6NWtrNPgFLJ+D5qs1BTPmbGNrJP3eSMWuq7ozt7UionTmZdmIoIJoFoZWXAhaNg2eZYKK78P1
hzlU3pM0dNaYmjJ+YNjWN2RK4xVKwO5Ap3g00mKP0E9dy+0wXSUv8ptWLNvn2Ac/PYRi9KWs4N1H
6MfXvcDJop2c6AOdhPWHfUfwGmSUq12LjkrFytonw5+Gwab+jPXOEgkad1jaAMq0Yj0IHmzBWcNv
k9fp6LRgb9B/C1gM/mM41G+L5ah46CPh47IozLwMyLDrFDf1TJFzxucD1qUAH5ZJK6t8Dtaronjx
lVyJQEbQ4XpfgEa7rdH8ToqWQJNw19C8VzibA4V/ziwYEgwJGuzhJo6JhDauT1uSpGPmpyYgpeEC
Rh/4SsVuVMISFKbEEX7TLFSDD3VPs0oNktMFzGUTxVkhZArX2VSZuafv6PaVSGRGmjHA2QCRMUpP
GtF8UeHI6i3kcYKtRHxEvvhTlBOyzsY5v09dLwn/dyO9r4AFIdsWlT9xOEfUyQIGxrOvtYgU8aMI
KyuHTpiEh9jWwLfsZOqnFin4uaIkY6JxmUhpTqSOBELIVlreSjLKRRMnsXM+7iw/NQsaPtXLEKfA
aJqtTSOH9K6J2bfjK744fIOHV7oAZONNCQUNH+baIQFOmVYgbFGT7pXyWIbrLnp5Qsvubyrjv871
BjU6Na/u2vdi3NLfACMm6PNpu1T9ejyIdzYdt0CKz/it68Z33VGFi3ga7Qj+y9ry0vQgvhvBZoNO
MFvVBrImrA9hbLIqYa2+Dd3TvG6lOmXfaLjjySMrgCMj5JpUp8QT+7brOFJot0L7x3CKKU4aQoz7
FMRKT8JWqE/JWFHbTwedJRGAqkGOC0a8NQ776vgxoVsbxId8B7JpDzIR6w7PtDBumZhQE8Ai39G2
5+uP1IySyqoZTCCEslo1Ab6Ni9xw+MwUlL94x3OfXKy/G5t11E3Snplk+vOFdZLSxi2OpRh2s4QN
4kuWSKUqEP+N/58T1FENhWkC/mJe/WjlYWMTLEbvj5fcAmoVB4aCdm4WbW2AE6rJNr7mAOiU9M4b
z243Uxwm7w/O+DRb4WEA1e3XH0RvOqCn4JU4HMDyo4BF/aRO0nJCJc64imHo8KkFE5RUXrvCZT+C
EPpbG2AW9fTYUl8q/AdzPuxqHRAON+y/OpNMcRvos7FBFSXJSrvUhqAIhXo/8CpzhCB0zI5x0uS3
O2CzhBz51yaX03jUsj5VyVgENd/YNq9OsLURJ7KiIU7j0+NroAjMuocrSBM5U2X6RDo0qoyjj5DG
naOzCJWhiEdL5pbG933xTHsBCKUOagZjZTFVX+qMKZ9QZ80yqBoVVg6/sQSlsSJEzOD/LZ8uBqP5
1NAnUngaXUjHcbs++gcSTtW7iTNRuj51csvKVj7t7U2n0a4/sdyLckBFg2neHOkrylR6avKkmVln
6LH68VzikfT8bwAnqtjVDOBzgH8zrCNxwL2EPc2n+CKvKJ90JCYUC59XpoEd0KpBlBF8mzOap5DV
RsCu7RJh9+pnfWJhj5BURaT4HGe2iQSPyXYymzsV1cA9Sysg/9/G045IMSKCQpWVOGaTbhIo7d1d
WzGsRUQB80lKfBLjIp8avxLIajaG0txqvZGlsADRZvZtq2vZ2Irdlwgif1SuUfXBdODNfZK1Cvm5
0FrN4zTAcWRG48wauyzWTe9fEHuvlqmbEVUvfz27/TPUkrOlO7hh+rQXHT4PsqSqPohYLxsiiJ7L
1v9hyWAlzGvOIS5BeWW7NDD3atIM4Fokx8EhiXJGIZB882bQCcUeeDNzQwz0/deo1WLWdpH8hm0r
z84UyqQvqr/rWlwlNHd1p/cfr+0TndcmHwA7M28wGD8LtGV0+doPM+Pbn+B+Qg6z36RS6hkJ3wma
UT9PGVLyo+9sAaJm/L6lnEHSk1H19KfLOb+gciFy4P7wjqIr5rLOc/mYriiL1RWUovdLHv8rJfM8
XK3pZ/ljvYNf8G2y04gT3UKYgQHTOP40W4Cq4385hmVL4/3oEBgqudBlTS1SwcmPrae4/pRZNhce
KQv/0Qm4Kz1cxEFNtwqVacQOAwLd6Ao+342C+sRZ76aoMk/tqU1RznQnDm38aP8g1yrItl110Hgp
N4ttfcmhXVYb0m+tN9DxpGWhamHlGJp0ZfVxCrViTNMMU9D8iuUlSE+IWiDZs7yzwp69OVhw8J1a
TNrYhGYasnL29q8XaV9INCCESzdOuAqZIjnZeUu3wPjppiEEojoR4e0ayldLNV2dx30+LH6G7nod
ZD/TKL3sFeimT6PRFQa6xXRRdVK1fHkmsEJ+Y85Dc3F6rvHfvCPvlUKX8ZKW6pYU/EyV/Mz9dHhf
J7jQ/IfGsAk0mIKgrgamJXwR0opyoqdVg8IaxglzZEfDZtemKcHMZbWyq9fBnPZU2iOC+uqMr30D
gphWJgynAMu6kwgRW0UgcUFJbu5LR9cIe0BIXhsMQk1h7qLBNzEvQKA2LJjH4hV6hUehWGdk9cZL
tF6zbZuKuYZOK4eIwbisTWW7mDkf1LH8HRb4SVOYoY+w7iPQxJOaL6UBL+j0Y+7AcsZFW/WpFkgA
0A42DNud746GhxObHBOhgJdBat7bF4+yKPKfBUXgDG2jineEptrEKEMqgBUsVx6ODH4ca6aTUUVC
VIzXT2m5uICoEcjK3v5yUlVTEi64eAOH3Km08ErQfbUG1kQb38Ky4yt7kkHl3eKO6Rtey0G3BYcm
60j8lsPguwvyTXZWMNHkJU2oGQ2JViO8kpRqeyM+KnJX0Sdt0AbYUvwFd/mNf2BmPFowb5FrJe1b
zhyAYe1RbCFlpsIlOIRddkDejPd82fTHs+IXFZexHAdQUBUM5MRdhKQsic2I2gqhhD3SDgP4Yugn
RzNg2ON93OKjGxBQqdbgAt0d8sICUHAtmPs/IQVC1kXe+60AR6H4QTbKqQhySaf5b4gmYcjaS4gf
o5NjqMoDYGyFl3v7YuRLoqX1yjAfM2gekwnSuX81HfQTgdCPc5eIeVvdPwV0A6jmjA6zt2Eee7Wr
N6v0o/h1YKE54unNnvO7D2V+GKyoJUb5F4+ugqWLUaSbH/rOLaSX+VNOt1zUjKAi5g4bo/BgUx5k
H2nEezKwZq5bbvGGOHwblyE8wD/tQ2+sedk+T55v/ARS0Mxzs6Tto4NN36wzTTZRLOXrPP4rkp+L
RhwkNxsph8HwBrOhHVrl6o6dbHZh2182H/4MazN27hKPL++kVhAgzQP/d+mWr+KyLrF3mBbRDX8W
emZSQ1p81WkvCTjqMIixTrZyF8p7RPnCmTRZK+oQoE407isS7EObs8TsvV2N7MzRfvn3JgabYasV
sZcfAwC1glTX7XlLKEh51SV6PdpYgUWB4PaqIXiKWgUeniyvVvWHHOsdIu0FyyHhdv3c01E44Tet
IWxlrbY1vbQHe/aqwn+BwdjYokiM+CueHL8HBketH9YHTrjQBcHvIJg7RBI/+EFZGVbWmWkqpw4k
Tt5iLeHkbXUa0LuNnWp+j5FK1PM6MFM1HboGr7uuBNO3UOHp6bu45m7rKq9CEf+Sz9StBpNPNWS/
ukxGvJx6mXB7LWYudQKvprMLSh5p28qw9y7PqtX5gRKfwwQ6kbJRAhK6nK2xgZwX0z+8rKE9pVSA
Hzmgpnb1IqPyXXq3gnBMLgs7cWxlrPkjnlBLO5zL7lbW9qy7CmAFq4p0URpydOiJDITzmsjCXWbM
nYjDRxXRKxeJVhSBG+LNakL59JzYiqbvVevBV04JSUXzJ1+Fe3E7Nn1vqPQq4gHTV35qTNbXWVij
7/FjtfF3eX9+j+Ram4N6INQp4yV/dfalEQG7Af7UgZHVaBDm9eWJhfG4a1Jw8fduiYm2PM8YLRMJ
7FB5+AasOuEA2/mlA4MMEoYIRCsNcNv8f80Ebgb5e7k+3ggoR1p9LeSMRk7LCCNhrgBe+EWSFSty
bMPGkpMxuU3JEhQKPT3lOsQd/iq5Pgg0dr8iDpzwOaUfNHIKA5hn4EIXwgHxWW3YAwfaA1WGixd8
woTblzQoBpqIrZ+EofQk5RAeGWAEjKc+4sIa32ZucWBphVqQK/bTZhPFpicQuCEj0zC9luarIG28
8CWL8XACJp3C4VAXt8gFrqqE0mRZWZ5CsaO4brlxsuXpA/yOHyeVKJC0JkA1zIgI8IC+3a4uyfYg
dB8O1lB+EwfhQgoN1/W2+MBlh7UaPHUzqgzeXwLGFw80JMIn9/qbGVVGMvwV9tOOllNfVqxTpqoS
IbN3V3jz2bECIPPNdnsNgsikchZlesTFVjsnsMz78iV0TpkBgS2TKqvQPtel5itd9xdym0XiPfJR
bveBAnicvwVtyZblf88nGWKP1jgugMY9jCWRX1+KqQU/Y7jm+tlaPrCmyB2RcySKh9KNHWxaKh/I
p7DpU4hMGDHjhsKrbxkEZOmwoD85/wIpE5tfOU2lGjiEob5oFmZfp57tsllACaEpcflDJv//cjJF
d8GhG7WJDZpSlcygWzgDITqBNuf39zmyDoVBaxUVt5iHblF+P877/F5DmOnW1wE2iwtq+S53NZmj
LGu7NHi2mYrk9X/kN8jErBc5bfjkEjrqav5UDPkTsFPHXfwF+zh802Y6BMqnnwGV4QvLdLBx734H
+OUTU0ueKJQJDv74CJUufHEbbRKibQhkowO1eutfipYW0CgoAediQz24Te1FzsfTDyD8/9Ns2cri
8fHxXauOYnwkuHYE864aRyg1KedT/JgCyiw6WzFKqSowIC27W1PHhHFi/lhIywmEFXqm89S8GwSG
QM+DDLYTzA/Jn8e6awmp1EGt83koJ5As+gplIjnpKFlDBQKXI9vgI2HW0mUx9vlZUXOCNcXkqv8I
1O52lG9Xy+cmhmmruw0KMuqn33icq84+RmldWmE0sfnHqApNRxfBuKK2RXb4pvcv2Pm30XTIjBIf
rO6gp14Lr/t0eWj0RxVaciMKuvuYOcm6b4B12EQO47Ev6PB4amPNVG5QrCGQFu35//qwcQ2jkYmM
oU9UyprnGH+Ji1j+7AgEmXBvZwZrhLGwfKeYKpxIAc8RZKV9Ja49CAk9WpFmwcEOynzwElaH2JUi
lfXUSE2SwkoI4wdchFtFejMu2HScQXTUF1yhG62sW/8pE/07amTgpaDXtoE8+hxoYonT3F6zuNlC
uLHyXoUHA66ykWSWIiS6PkyjcXLNkuENBrKisy5vThopKzWq/PWYFfEjzhiTwOhxemjhNd2AxLzr
aCvtPfikfPI5la9pe9ppUvkhqp22Cuhvvp1TBgQEadFb9YOSD8mwRT10xq9r0NInwCgmV2rKo6FA
+ilxYOu5OVcy2bqeqreJ/lTSMUiApyr4d1S1dNAO4WuOROhE1oZUAVrWdzZqRJoGH62W1VChzKO2
PgjZZSY1vxRJLt1p70Lx3fx4PIDU7G85ZkLJGm0uKI9Bk+lsfcQ2unjD90gA0CAp+y1WMZaqY/V3
BBX91Bu+v9ikmFW/g67fK8P5CuCglMyz8zGlBbSjd6mFUVhWj9nliKHdVX0557VdcH+jZv6cVRCw
vOwLSFsz8NzBO3rr9OKJ2/Kj7fDWUxI8JEgckT1nmPnrm3U5xOYdVMxbpqIN0uqpq79ruc3WcArH
94KgwXhHIZSbb+c6uItbwBNZgCe9Hjyqe3pfhGJ6H2vYVOuSJPXSO73QvUZjNiiaH/Jq2JCt2Wzd
4AjhSWkWGpv8w9PS5cV3/NqZUm7hv0HMiHVgO+zVCMlB2YSbaV0U+/YDMPG8WR+PltZoZjFWErHn
2Me0ciOdS/LbnsWHdMaSOHGZh09Vq5JmWuZLS334P3ezykdW2o1/qqFVLpKQtJGwtY8NP1bGIx5I
sUo8YNpbCLAt4YNHrbWVCYv5idegntQt+8w+PjeBNEHEC5AtI4fN1prHMlXLb0RAkCTVdwS6lvUt
U4zUlNQy7VU7d8wsf747MEK2rXRU2laavZatbrhHB+3TZKP+/CEqOGox/cMsL2P4BwHJP0dfu8Yc
5vLrxsOOHBBaq22ZouJdOSzuRG5fYLVTYhnZ5eheynPBMYGeetAIMwxfRe6K888+nDVw9Q1LOoT7
C2ySihcpRnqfYzm1/TYW+PKjkTwF85u5Z5uEIhTfkYUyywNMZe3fQxACkJilalNm0H7WH8FINeJU
kLRW63to/dBNeDj+iSjPDyTbB3i40V+Dxnj/Y+A4++7Y8mxBR534EnmzM4p45T47iZGh8/QvkmXP
+lzVAEuRpaU3nYfpGnI7NgnP8FnmfvpTAZL773EZG0Rtv+S32hSpqSorQVa/DlvgskHxThQvY3HK
NItmqCO522xUJ6DBxxvm/zVA3ZPRhA/lrKAP9MrDaDvywOQeG8qFYOz9t8/pO7h9zE+IoobUp6RT
6TCA06JJqWxUgRd8PhPEd/y3xKyXxQBYSljbpF89DOsDcUiuqR+4xzgAcBYj+AV9g9LySYrvDk2z
uk17J/xNiyVGH68v5j822SoMvKasdYb9htepeYiwfDhMkpmd2h3hfGDvq4jOFB6pB18oBrlFgG2b
+diAT0bGmAAmNfYs7IRUOMZ8+M09Er5d2mwl9aplRQvqBOCq0l7QJs/ZknVAXb8OYmsDrmThkiyW
HA3ShPGQmkwupPjY2dqt0R3QUv30SGi1sF359xF2a49iQ3K2IjFTCa27sPEz6xua+8+z4HRsQyAA
Cfn1AiVpW2CgZxELfLN8GxpingB+TUlkS7shRlOZdx62P11lZjFT+TUmdpnX1ztj45v0g+J73oJf
XurfZOFYfLfkCHAK1pF5NZiXXcQzOFWVjbXQxWgGNKfcv9qN76ARPemWBvPpHe95TTs2MCUJkDFX
0BRVGIarv4uc1YvjeLFICkBaUVTcAkuYGv9DUTUSJiqwy1QK/tI23vMRPCI6qG/5zodp9kGIlBdf
8/SjPURgG+9MYnrdraZ/dTogVQ/GY7TzavSGxEXtUiRc6NlwTQ+ewETHJkZFBJNfmHVJxJXfuvSw
UfbDyG/ljVn5GGu7hUpOedhGlFl1i55gRUWKnQEtcplmosZsfwb9fADl5udti+JtZK9H6DwQbTcE
R+hZv8t25EggP/Vdx3WWMfuWv3QrfsiFF2PzQT5Loms9oxMBBFREX/muMLhVIE6OnJQFCwbhVLRX
Oqwc3MKtfp1h6UD/bDzczzrPiYsD+w64SW65w84W2YsD5oDe3zR+EzV/DHMd882srZrUkFO5fzQf
cj16EZgGEodzMFYG/SszV252XOFiQTR6bReOGA2Lw6IaiFwG3UlPkV5vAZ2qnrl8YCnjqW3JnTu3
xYepZUP8UNJ8PfvhmmjimAzPIhfv0zeeSxqSFKdVFM1hhYRBRqiTTD0NQZ0VDQqOXRgu6IqfiUUg
jT/M/ubS8O2F3rynZS2T1aEHqSWtzkQSkKGivSV8Z2OP+4xDd+bqoDUKHeVL+2eO8s4RmKRg2+JD
Qo0WVkw813ZNQ1T8lXnsBlRvKKVLVwE8GjkdqvW1tQUxIwLi46ChU4XSA1DV3Y7JpCCtIIQFgI01
c0kK4r49GW0bTA67jzg/+bfEnXU7R4JB6fTtZr+O84z1LiybsYC0JmwMWO0EnZY8ua8ZJehyZW39
Kw7do6VgXOfwfXFHdFeL7m5DbjilmystSDt57cwhKrR0uScY8F/SKt7rGEIKiA9MbwLgZpO8aaVO
WRfwxCq9WyDoMrx4iszS/nWrXZ6iP4IQ+51jnbstMIXdO4ERs/ih6uanX0BKD9tcT6IfGSThu4No
T0YfHp86ppmby7a+VjY28nGTVPjbZTq5SPceeUh6fV7s6iCs4AIN26qt8JXOPv/Zm7Nw6GifnBXE
Zj9A5tm6LRoJJnIDWpH9cyMJzQdDFrDK0vUnhZ79ijMuXMKXFZURmHAm/RhOhTwV2yWoqX5svFj3
Fi3CeCSZM1hTWJz2GcmLkCwxFtC81QlVd2XjqIIxVPjHeoDZ/wRGLwarmaD8vyNPL8qrcvMjWdqd
LXR26fizgB99Bvqt3lBAHMnLz/EZ/RZEeI6Co/1lXnxqJfoFo9QCb9qubLGvlQMiYUTQqOaR8weP
AmIsiWkm6GcW67/+3er6V+HffL9qSkdFxDmqkypjEVmr1PXDL8suaESbuPRc/HhntJvyUtvJi+mX
FrWpjWHN2tUpQAeqECp4t3oB/xaMv2jhMyO6vN9xfW4N8VDztz8gRTx0O9ER4y0+flW+kU2h8Tp5
uaTM5rw6C/yq37gudK5ARsYK6Tl15BnmFst2pPPKDhMl7iZC6NJnnFvN13WV967jVdBKElMIFC2j
vJNbUhcDv6wo6vA0Mvhlizyp10G+++XL/AxQHP5TBQys6xNruQznMnKUdr91UKp0jjnkrXhSaVJa
qIvLMsdwMqCpuVUQDh027ZzhO4vbC5tVgPQ7nTOq72giQbgjPiDKn+K+3XpNdjQ478DlTnaD0art
1TDrad0Mrz6gKY6NJdQBji+RfmWOtJGrSCKRM0Vch8LR9WwXx1K6lS94etRCWCDiql1VLXMIBdCM
AV+sRLdTiNkCjOF2pr42NZHKrN3WpYnPmcbLivafGEXJDbyXYsaDqxp06FQ9eAsZPnv0EKJHiaLd
P/ruADegpjMgSl9pm536/rUKIKE/xv4qCPQxzWRRXoE0yYYEvOt5dcwgWi6hlePlkRv7s/sYidr7
tsuczZ647KkwEpmUTqtwFe1pwGoEEsdb+42/wn4Lp0Cy1aDKt4SYvT/QxSm5IxnMzXWVkgLhMpmj
wVFsgjfxyM312SwX2xjWnYt50Em4LiW6v7E4rYU2kaW+T6EWM18kRKk3tVRO3poH/p815YsKCSd8
k7BPJG2lVl8Dl83b8xjwf8Se/rgWqiqNZayHz/aIy7Ik99tH0sTJP9/eGRoP7KjE8llw2MiV51Ut
fUy0qmd1R1oC6JcT9QTKZbZOpWGRNJ/U797tM2UGjfXWEl5K+27KGXmWV2r6YQhhsAhesgySyx+R
1hW+3jBZP9NzwP3741J0xfFiG5YaFofG715dcuudAL942DphIESveq3vK+SfWualf2oZfZ/oVRxd
/gj4XI3+0zjWnP+25YcmxKccQGoT7lTFcW4ra34yR1ZgFnsejV1tVWBLJTiIm5IW9kHSVuq0N/7L
YGd/b4gxdXnnHwAffOE2PoaSOiMDzMkU/GwewrMKPxnAxVhtPDkrGxlYb882y9zbCrCf9TaDOh0X
A2f7HxnTOyhdjZnp7LgK9S3LlUbavOeZInc7T4P4/L5XapMEsIwOjeDNP3yCW92K+BBGINyuNF2q
JkUWP8h03lkNptJaVTPFPyb9bX72OLXcmJi990+4cOmvqB/RcAPNfQLlebDnq5vhOTqVX+TPcD7Z
zNrbxjPOiE2DwCSgaKQP53sixCgNMQmXnhzPxXSscvFaeoseFUrVFNfwpmFNLoBjQSoe8vH3XDFa
jNnZh4s0M4pfG5ZqO9MxgiCzZo1Wm5U9ur0NfvGi8I3kHqbDjVzRWMgHJi2Py2Hd8NzpXaOeI8D3
IoVyc8rgVfXVyoTqMqHE2xS9wsSITwfA1AjsOqmlwmkD09ZQfY+TiT/hPgsBwtWKEnLv9YCM70Lo
AM0DhdNrD9d9w7YJ7cOTIHErnlivFKi1nvH2NMD/P//9G4oD2/QBNpY1OYctEqwDzXvAkDMeUHGa
mimUGnKcX+D9WBERzAH568GGxi7mBLeFFEnFcKj/y3Di2RIQ+nzy6AYhKFljwXtrL2AlLQmR/p7a
fJiL6Fbhy9EdUcl+YXFgUVM/t5ecVjb2rpzXABuMraFvzSO+RFEqEZLZ3dvZNQ8LRcotNY+b8tn2
jfFDDesG6VXsBYPUnu2f2vDR0tNpe79MhJPSZmyWX/B2uDT4Gcjgh/OCBJCrnc3MZ2rO7Np0HDGO
1MGOyTDlyRE+YbeK9/9DDQjB54Cci3wKsHKDjgUSEeM1bdUpj35jbvmtQ2UnQ4wT0EHDFESw/5Vr
fe6uCfFNZEii0SOjaIxL6JJswIdL7au88kWcpeJM4O37ntYAqDnB2NtjT+KICeOcvwT1JufDkyI3
ioxUYmjC9DdiO7oWzIFdYqWoC1Tv5DEwsnzRt6Qr/K5cdhY+SGbFRiw+oKG8cGdT4LzYu6TKY3cH
vgn5+hL/v3orAQz3z9QZtqjH8N3PlZ8eWPz/YNVqigOsFDFbK7oavddYQvX4cmk2mT9TZxW6xIBn
D2rCCsJoTMh5SVb/SKjvampyGJUAQmrNlEpe2mXwKbYYObOsDy6jZfLPnNEwdZiVGW+E9wm7carn
CSca3DoaXbwdi/Qs2Y119Oz0sdollEr9+u69iD12cUG2lf05aPWRBY3gpFbuN8ddGGrLGajvIw9v
7A2cpo9O3Zsx6oybY981BTG7kcAAPUxnJhY2GTpWjhbh1kvO0V3++hmnxdOrOtWbpo7bmzgo967p
JXftxr07Yt1w9SPw/8nRU0RnXRif/2KauqjlyEB6BiSH19PgCcHnJoEwPeqRjvomX4t2CmAhizuX
+o2X/GXKYD6Muip4tBuhtNNk9+oIJDbnSOIQiKrc30i9/SazEB7lGC2fzawS8ADfSJV5tkeLtzfy
ivl1TxaKHhMrZ2BSMRtcm4iD/yCtKLmxyblFe9FH5eOjkUJP8I9fE5eJgHf7FKojyHb4PrzIfRcO
KtbJ7f2XmVuus/ETsyCDfo+8pK100+nvGMSToYJrymhkij/cX5v3Ed9Thibhb2cU8QOXNbmTmykq
X2xBl2MkJPhxzH7zsNmc8VOLC+xPRpq4aBoKcx0WfTiJez4YcFTIH0O2PAO0I+vg7t3TvMjFLH7S
QrkV+YqPhgKgVrZE0AIKgxY1BCWW9nakarur4lp0vxhYF5TnbK6tEOG5ugFZKJ8VyZzrlzJ3/SLd
uHD/+ufclIYykHrL2DLlUt4cYDUGYkPtW4VVh6v7eEckQm84/gKBeIKWLTcKIQMutmBQfIfu0UuU
gNPNuGvcmeeaDHSYC/PsGWDKDS0ssoBYY+eTEGGRDUR2dy2bz11iRgGRmCwKUJsvqbiZxb/phH4r
+sWO3mIZ+y8rjV8cuesvRYDVCi1tJyh5Wn84BtuAWBNnUQmq4VV1p13T2gEqRk3MmKG6YLZcs6rR
Lpqmp7MmimtxqDm7rNKjDFJRsUXQJXHa6eLKfFG7WrtjXliAIX/VKxtps8jjMxtzyxAQXobfRip6
ztmfVHxKS3/OUzLg3qQfM4wqoBpP1OFxB308/dGle86P3VgzW7y9AyKbyI/nNlvZeorErlHuFgbx
LO/6luqlxDEgMrpeFxlaxqcSjWrOOTtYgENY+f4GxAg6hXkkLGrcT8zK1+aX6X1XnT8wr39FIVHj
AyUDDRRbFb5eS8CZkhCxU39lm7eTdbU5LfkycFpY5uWeSoKnjHuuL5Tt3Huw7hMS7bCmAQ3in8gA
57Es3oeDMBDMeW4EKceNshk01TtyL8HyVyFVZ9/tObaC+iliT/FDmXjrollYQoL5/RqHqIAuz5gB
RIHofuklKXICOBChNlJuXZN6gwaCX978raBqFftjRwd66FEv56C9JqSNXDrxb8YmOPEsMKs1w8gn
2eMRCD2sQOBPqTMjRjDi0Pe1aruOu75u25aGsHW6ZS87j50MqAvOSXP3OT3bBBX7CsqGxQUXJqIm
yhoQ6J+PApT+uivTwfnspDr0TSoNE3uTFfW58mU0qVSzkJ2+Xsn4mmPSixChPrd+WW8jye0aEsed
kunRR4FVkwPeCgvxopFiFl7s1MmNCEB7khv2yLGbpF1YPN3WWJShibxd8VE/NknZTwYrgdW/kGB7
iTJBpt4VtcMDRvcBksHCr8D7POhuODBvqjsdtBFyTZe4RtWbXAlT+wIlOgJlopEjoyIjSbKu8G81
v7NaIXwkz/O0xbZaNqIvrlVWe3IAtMtXU7RNrPvs8QA4/zpUj89i1G9yyk5Be/VVS9o+EkdroM9+
mx0LrItcVjyGRx4fLgH0ON4EotgE+eT4l1CKySF2EsXHJzmuu3QP6syi3Y2NZTjk6jnds6h9mI+y
7pVGvspwPC+6yoDmpV0qb5TAB1McDelQTb8MA4d2bQ1QGCPdJJE6wvi6yo9CcO9ZZnDHq1oL481L
1dlMhXUimBj+q3fDGOjbroqqItSTDIvqrrjAe7SKWfRcEme8dkfVBl4izWaIzAZnNpyxEMbmuSMb
CD7+iiIGb0ki8WaEcCIBjt87gw5Aeen2lciGFfqryI9O6O5zmZ4hYJmXui3gi28Y1nCviHJr4OW0
sy7+GE3ZHp/Sww48dxq54uh/ZdfnbGZSN8iV0bSM5x+hN9Da3bSxAyTdoKYGAaTTsflwV3yDHehh
oPgJ9mD2QKP27pt6+2f9gGZDqVhsLEKcASqCS75bU/vDSEkMpxO2fVVA/T7UNcWN7rZ5tCVnhSHW
qbApO+XEPau0vbxiBtrEqHaOu7bEewuaVmFyx79MgznnvCr14My4b/9lmmzt1DfjbwLA/E/10syc
yD66aoYavji7pNWo5TripYFQ56pdigzkgspizytmMKAAj6eeN4TN0TYywETvbaVZl7Ign7azxkb+
gIfXhxXCzZE8IQ+19RB4kDFi+UF/0dIx/2VKo7DYHEzU1+xL9TA29A3BJ2RaPVI/JCLlVo2jrjH1
Ue82TzuSRhbD1GDeGpqHo1mE0pheD2F1Y6KPldcnoyop4ZmGQOKoy/yLn67IdJH4SptBppTJSjCn
ZEQFIbqGNN+E1KSUcp+3fnjYGdF6sG+QMx/k76Tkbjn1gnqiZyRL8WV1w0nl9jRPWq2L0x5QXCWs
gHKSymUwvZwUwYbOdbNjvn2JocRuiyjUyp9HUJ33QezagXL127VjVis0VG2+HhFScF6zXctB6WgB
zY7bwCk0ZTVL099dGR6OzPD8tU1A2QKeLryu0AfTzr4h6PvwacelXrTjeh2V/lyadB199Jy0xDpi
CYNIQEiYmsFXKKoKPRDtTAeju1TP3tL9HXYrhWrIA0Ig6LkjC6FXIOD1oG4VcIgHt6tCHDinDRBY
LNbPA+reyHr17brXMrysz7CATB73raLDeWH/XpJ2mS07jcS0W/Jpvkt74sE60ZmjeqajePgn38Et
CtTGW8XA9Mz8vwMZwiDrDoUmeseBd1zl4lheMoPZ4ytZoDUxx3Y76opQ6hcqnKhlpMmE9/upRtA/
t6RrhFoviPBhUD6BLsBFJyv1fLOG/gYfZohhn1H8WqneABqtuLd7+52ZG1hE4XaFonabyzs0GFUU
bwzujPQwvCKGjIqv7gS8lwCYOH0zdNkohLof1u14EZ15Rrv8U3YKPZAO9llTEMOdAoUMXkVAIcQv
9dp26ZtCMhrLsQvGqAUY1vEvNvJ0P8YrWnOS81D//dlNIiUDoJMns5rg7Qt99YBG4kxGtRTL7DG/
t7IATpJW+w+/PMZF5R7DL7vF6sfV871qjfq4c94qEtnHJPG+9bhnjDZFotGKrCeLg/iq5eUK20aY
bd4lUBWUiLO7EHzG/13ld4VXt/ruoVMWZ8DxsEftjQDW7elUti1vqRkB9jolO1baQApQEKqo/sZO
BnVYPrlclwr6b8vTBw5Zg9QdYIJae4PVdw/lgzWNQ7/DZm6qK4P5jiEX/lhBzV46sRxrBx+r8zXr
8AOtDSWpPPE2qHRo4RZQaN2jzWw/WxaQgkfbTHRu5pIhGlKyEyn6r/Fvr0M8d2OT8DU0/meN/wu1
N0STRAlaDGlggUnfuTyEu6FMmGcz/bA4oJVJdOUBieuvrZJupBkR1W2SJVsAq5Vo4fykC8/WCyaZ
oUDQBY0vjO30HOtT/lq7pxzcaMDdc52qN1IA/N5iG89q/sxUVRIQoTwYcTZF9cn4pbvFtMkia68/
6+D/pXPtWpNi4K5K6S5OuTyWfBSkKm0hpdQs9JDvS0Z7EhX7lwv6EuddI/mX0h2WTVWcEm9rHWxb
xTq1xXh4ViPCBLMZGHSrNB38i3woec9TlXZzVfeBpQzKdFgIFGYg4kTsjz/vO9FeTAb2ztZ010aZ
a5MuZjJ9xYsVk5gqQp7eNDcuN5R2RozJymaUWVJKgcqBufiWtgprElj3U7JJ7v4ha9jw2V4c4THH
wdzzP56UF0Px9k/4DJ5E79DqNWNv8H8GBXW2wvf9KUgBzgOIzCkxU0E3eRPlgKyjAgWyV4u96mFM
2okI+B/qzkeSOtCby8JilPLuh/uDjmv54s5R8f1+/0ZyGbW3oWQF9B631CCTe/jGRSMk2FvC/y+L
5OkbtEoKfvQwEtB5NVl/2z4FUIuLp7idtuTbNeX3Xh3miiKqbWArj7DLV+Tx/ZuFihIo6Ak9Rp+t
lK/ux0RlCUncH4FPfZkdPGuhV8e6mk0KqSasZgcqMQfFrfzQ+hxWCyprvqpZZ3RA35Xd1YFtiF1x
6VBtBc6QR+6wBL0VKCLwQjsT0S8FPUkY8bVZLlOVwwU/T3N4XCRvjovkuUbMIcxUOwbv+fUPyBmv
jWn8jSwgwsaG/qlWbcWfPF6J/t1QRQHhnB8nWe+k+Ml09QT+VfGQ2Huiqo54uuZww3r6nV0U1M3I
iN+tPWvmcmekZ0ZcxjeQSfShf326KbJXRphkXtqibJGl9M6d0j+HtmxEocF9yxnv9pMWnb1wEdpL
0IeBtnLCR1fviqTsBLgtlPssQV5Te1sUy3szRlMDml7eKj1+lUByDidMuzZNgjY7JfBkqgNea9zb
+wIyFI8LNdFYvipqvv18ngaOe3f7rp+FXrdynCwiqgTvhH4ykfW6+xqsAJg+qUcprD1yziH7ytEW
8zjoKsIREOBWold7ulvn6RHONqb5vp5zZ19rWS1kaeHOvPuYCiB2MfLrRXniJ5RaE6MQpkypmdf7
SUf9Z7/agwgCnIwWBhPOqmy18cJ8QXURjrFIMhOjooIMxi4SMwm0TM0yd1x4x6E4h5L5fb9OXyUU
/cIp+ia1mAg2k0Uadd9FmWIB8pJ77UGEtKI81Uu9SRJGwPUZeetJ7eSbaLUclURfjsQ6AVLTTuFr
PIuXZFpV/ur5a4z00UlI7b9vF96RfBaRppfCHWJXJ6BBGw0ST9IvAEP20JhLOG5iI5+teVJlj8QY
zBHsy1CmjXcLtotXT/Gzs5O6/fy0iySvgg5z7hKerP7T32lJlthJbYkjXqDTMRDDLwoIBgn920Ot
OS2slKTxoqoVYS6yuB86DZzuWwqigbXcjFnfJG+wr4o1S3/Cz0SX2Dp4uOSgrAbYvF7QUZKrDZIE
ct49MVH39/3LMPxa1g3ebWNIGasiznMufMw75zojsjsNA2E6hlbYS67bPI20KNizsj+mJeOepZgz
t2U/IGrbGcEhcip4qUnjCfBknfvXtusEe5E78hVaUbI39sJfxekzUC7qV+q20gxwLNcY3ivIP8qS
rzKtTjHx49wwZYS/L1OcN39iq7ehnY7wcY7Z659u1EMt3ZuLPSRFJdCS6N7BmUczVcVJe0KesZnK
aJGFjCiw5jUFMe6mppET7vfSc77+sMgSu2Fb+EAF8N2/rvOmZuFw0RPsHPoXYJqWbP8j1h6E1e+Z
jqpbOJVeyY7WtwCi1RFW43bQSC7+ch9t8ZwkhWbJ320VcoZgTbqEOYdHuGsmS3nkB/JJBG6Y/p1s
fzY1ZLFkL8gvrXYPAqbXcbyKVvm+yNoez+hRcw3gDNU6qp8d9N03jhSTlPVBr9oJ39vb4gpis9xY
kI1P39Rq0sa/Dc88gsUkSJy7+HfIWnSY/tnlnbhxT6cK8PcjGHx/Aa4zsC+Y7Zl6EE+O5PvnJzQG
ub21R8zv4k+/lXURPVxTCWryHf3HlV7PfaWiK8H3vKT+2obLLeECfHru2nHAE75FpiRpLDwp094o
rSsPZwupQc+cA3mAnpzNLqtomTo+wTINZuHky3DJxTmEoMFOJd/mXM5RI15KEgSG9Cggjo56hEEX
lUSHlxCLnoWHKsNVFfUqzoYKTvjZ0C3KBgXjM8w4rXT5yaP832t8XkPQFEyCO7ThYdxXfT6AKhQ0
FGe2Q8CCScrS6pEmR6Iha7LCJ/FHEdK0M6IgCAstxRu0JgkkEYLY0mQejzxrLddMgTfiS5CvXo7p
J4iiGZw9E8jgm/OoTTPfXOjR65sA6jQSgs5Z2+UYmKExOv/79Av7b6EoBUpxJn/ZH8ckpJOuFlvs
Yi7tRoU6+rIuu3cnFtl4IktvKAe/kTdcI9A3KGrsXoqKccXszczqF9gsmmA9FSfFbIsIBeSuC1GG
z/8aitNqUVwD4h3TJ2PlZhEuM3g0cBAQjB5w5pRhx4nc/PxyROYRSt5UYNkzIj3R+TXEQUKvsu/V
7xqOayR+g/gzAcYkZKW1mqqZ+Kn7igsBORcHKIXZpBFUnx9bZzKFbU9214ALT9UynWuUIoEFM2ix
pNUnliMlQb7kZFDfPaL0LeKSYgNS0a6dGegG8w5ExL0KePvyRzPOouEKBRAN5jC53hwd82EIbRI6
PbjPUhNZTktDKjCy/CRJlZaXwOdMgvtp+11qo1yjeA0ZUxcNOjETgIZA1RSJ4g+p0Lb1ob9ezOyr
98aLWx3l1QhdVHlbewscX5oiR8KONxbar3p4ta6KQ3y2lNhPnxU2rJfnSRTSph57uK8MuKqtpxhz
p6jeL1FalfQSJ5TZgbTO0MZ8CxyjMcdnrYsXYzft20i0lZ6iNgeNQ3cDMiyHUsWGZteIRXYAk16i
iIOkaEA+B1o77k+NyMKVvJP2lvgZIiUtDibtiJ4gMDUN90Yohc8Ux2SkUto63AUG0YfIPrGwFiBr
00k0+9Nt0ZCAyxxaJ7hu2zcxGfH/Ha1Qockv/A9uWxmSziFqcsQfUr8gGWMrYb4yd7A9jQcdex9l
0haz6MsH+jTiyScEUZLZGiUlsDFijhswb8629J/MDLY5OgrTo5bw39f+eummIh374Uo+QM5zdkhH
EHBrgxIXwLMd6WzlyI7Bsui7R+HUWM3mwoIL32U41hwjj5yMkcYpUAidUbFFhoIop5XAqtqfbIzF
n3YuUrT8gN65YuhEaGOa1hu7BpWFMPqfr97Iig70LnGyFN2DXzdR9h29cFJ18z4iG4R0oJMM6cEX
h7E5+/6BK8V9RPMhABxxNhJCs+zZL0BaiFbp4J+sbSWD8meHxnQV3ZlnRaofvxpahUI/GUqSPZcr
GAJePRqfW4A7/w04TgrTqIBxRkHrtgrFYKE6wVo8BNIaOZAsdaIUfrTZBFbwjB/HkkjYkdt4a8Tp
icIlNeuBXdld7Q2xqFDR8cJlXmQrRGaD81KxB5Tbwmo1xq0ATnTW/jWj6Evy9n9ioSpq0pzZrqOo
UcI1Pj4VRpfDHL6oTQwrbMx5HUpQ58N3DYLUFycSAsLFZiADY6eSR5hlk0v6B+IcHSgGT0/rsy8Y
frT6IcXcZq/yXCoTddoJSbSkccdJg1u6N+W70RPhQYdgJ+j+mmH6Az/a0dV9gMoNTiuxHYBh7/LS
T7LKm67cWwsd3iYFZ8U5EMznv8aM2he5PaDfCbo8Dj2nDz+n+htz6fYRYXbiBkC8bI32vO393UUf
PrHfXZYqpaMcGSZQPZdltmT6OzPt2CepnDybq6BKlCMkkIVhQZP+c7A2FoJJoQ74na1iQ/x7IDwD
YIany8lSsk0HuAhM2ny7f2UCvvqYUvqMD2gH2+r1w/c5u2rP49AMMNbj91X1wIUXGseBKeq8XUqF
WVeTrp8JWc6mGlA79PBpA9ZIInG+D6699IlQhxO6S/kUOHwShPLafnYayFumsJLbxXTd9+CcJUp7
aW+jjSuMU/RaldvPyaHnmdK96BaL73uOqj3nuDI7P4PbaxXn1zOiYY7zzGZqw/YaNGlw5lYfXTIq
FgG5MfQrLQuGbAu/Otke1QrBdI+HiuSfLT+Q9h14VLRJWBxwXKS3cVe4LfMgj3vGwyJ/lG2zS82v
M/rUBcYoCDpaRkqsuxUT+liOTqIcJV2bavPpTFG4TyHageQkfi0P630WYctjgLtizyDbwC+PI7iB
jgLpdsroXiAshqfPxmRxEYaqyAgGnDvqojAPF4ElnE0FiS8Lf9HlQ5rU2A6QDMZv38p3SYihWwvg
i792HRJQGWTXKtUn4MIJib1m4UCxN5B914VPf8iAH3Oz8WWrotSh19j9NRERKJven0l+R5tutjoa
88oS7xuH9ly+M7qr6SnlnPl5XRWZgPQn1DzzizMH1B6RzarZRCH9ZBYm4l034167OxHo2UX70l8O
Z9Cfb5ETuPo6eT5bc8/PnB7QNP1iW4pVSJBLlIX7bfukVO1JVJ1WjrqvaEWFU1cLGdFXNjyPRqKh
L6B/qx1gHJGQebuE3xVErsMBfOXe8aCZZ/1WDz/VlfmORLXFUojCyPdIqjXQDTGUIbKsIj/aUHmp
HFEPddkDR0j+Prd2Kc8jMFnOQYuil3atsND7Kk5sThi/esodXTxxO1N2++is6WoDb/CHHB02RXaN
0uqxoVztPeMqF12CzooG1QaOUOGe2nlTGZG2+p2JNrUhNB6DS5RVNdt3PN8DiI7GZZfavdDUHXXJ
HU4QoSwkIdmkgy3otU6TH6D0n59wChf5ZCKpArTX8jdOuO5PuXslpr3x/D+6sg8LO68rGEsUZvCe
+mLkOVy9UlX4IDnaRpnaAuPu3QBt+D6xglr8HFzQAl1sMk4CFjG57Q/YYpY1K0YNlpJXD8MvZx6T
aCKE0uVONPl8UdDv6xc2KSUiop/ROxK7+qAktgzrtDILd8KmI1Jw6VaW4CQgv7Tyant/jSt+lbdS
fMGFnK1r/bNMLo+QlHXWLGYprv1nO0yzBgV4+oUK4HsOhMIVMTqie7xvkhHtLv6rfVO/jM9mWMvA
vl3KRCWGF1FPKBtJptjmFkO7YK61gpFB5V95uIkh9VwxfMUCA9nIwblGQCuB4VvJTzXW2yBnDRCX
EDmmDq5DrMQSQHxZlHs7j/IGjXhB9vUvODlQW0peME7Z80T7sO1uxrOIx99HVg5k9JH2IQMtdHQk
W7GGjIYQVFjtosU3343NLU3Yb2yb+Qwddp5Qqpd7QPZHgfzl0Ja5QJMXQM0gvCjvZV8tpm9QDedZ
TQFJN8YhvUlh63JxDrAnplcZAdDliTemNhEfPVkm0uHFSdcYs0PzcD3mfJhHfIK/gpqBmu7Gfz/e
tmtOv4y+LIYogax8Ch5XlA5piHYuqTDYgU2xGId/7DwrLh4KVBBzRT4GTgVupwKUk5k4ogNJVs05
K423UPKuiP/0g2zVlzo2OXTnMjCGd0rSYm45sSsd4U/oS72g23IHE6gUIUCz6jHRSnnJyjpcz1fL
QCw+0rdRB1y3ClN6WCdW45Y5K+ecKz4ayBKIuiMCUI2uv1x56vmk7RXU3V99hBDpRkWaNPEgjvHr
XFYF0mlShism+6CiSVeHCm1S4o381Re9LS7vbzwGVyjExzBDXhOfaJCs6CZTA9dAHjNIbrDzla2O
gGNdCpCcB1o0GsB4sqjVhjcudFyR7/wSt5+IJicIOYfRzvhwue8nTvKuFu7td0ImgcqGY4PXbmt4
d5pPWxW1rR8q7NLeeYa5D7lwnb0ELQ9xOlomo5bZ/24hCQCerpvx5Z6cpaQ+iCTRS8pHrcD0JfC+
aMAvvTGKpWufBRkgpcCxRyfIXvxfOrFbsTYyQ13gY9D/37dK2M6ymG/o5ZeihMCvj9IMrK3YQPAx
mvBedF4KkFnMnGG7ogrVQizqOBE+1dK01qYBez8x7uJJqP/PAM5aDUBml0GrrQQQcxhLIpDmbyVT
8ZqkWPfHa1yikZmhPpG7qAOF4YMk7XkNpgMf8rA6o8pwY7wT3z/CRXYYrG+LiCil70cghzIUclUl
wN4Y2y7LFToUww+Am3hbS+Ul6PcGEA/KHFp4a3cUKf5HSLRrIl0X7v3MyvQT+exNR0duqOUnRweE
kxbnaELSC6GI+VMOmosRg2naVx2R+i67j4ylG8x8hEXlibBicQNBr7fYho7itouT2S9ShYSR9+jK
JOAccns9GVtXJ8au1xyRLvapFFTTk5CvZcVk8X5ZQoA55b0lQu4VsqIPt9Jt8BbC/yagOa0m6+Do
oaiay9ZetwsiLpJIlHDt6WC2DC4GRUIm29+V0jWj4pKWSxNBcBrlIHl/LxJeM5unQLXk3BmG2Sxv
FvESai2HQkmR2q9RsLURUpRkmu3keqopau5EoMS+GJbZtXAGKd54INadGpdGUF3gPXooUgra0FdS
h2jwibT83S60qyPwR2iWCl1Ut94IFwpvoMpYP+riB36NRAfiDgS45se5JTqRHhi7eS7bkGxuzhUX
TUhL4+UGsrFs4PWCRm5tZUmTRpsE7Oo1JdDBT0A6ra4cejIKzLljthIClMlGOCM/fWyFdW0Qzowe
905SpTF0QECmCkGjDEmuQBnq/+gxnA/18oHXN0vabL2G+I79x+XE5Bga8dAXl1h5INrPytY6of7K
ysmoZJnQu6+lgiyRvnZpKyyp8OyQALmjuOGq+L7y/w2e7Xw1DyJczhnv6i3NYP5+rGTFrzwK52nS
Pubw2TfhzwRIsEh246aYqmuviMrbjP9C5XIpEg+7E9vcllEZJZoJ5dOvmvrwWyt1BlFEx2fcjUCK
3eughGAb2ZbTB1yL2kAHOiP6LnmbLYY2tQ1BUYbPZU/oshdCG60uTMtX6nab33gKZt/+l5QDE4ln
64fRjoAuhakBVGOnJYoCL5xCO0UBPW1Y/hSHX+vgccJv0i2XQax1Ev1IauT9oql9tbwv2x0y0dAu
7IVkYnsBfqliRJGMT6/f7xqD7gLR4ipK8sOB4iJEPX8RtIufP01Xv0a5oWAxdRglyhHM8a4WwHiN
TID8kdKz0I5+/au8zHwKylgwCCEqO4RLOpHlvRNkq0rp7QZ2nHL3T6luivX/YzRyFyqFhDQjUiBp
l8UH0ugopn0FowtMGG5g7gr6NrjLCs38T/rJq8PYj9gwDzajE2kBumAmhJPPC4RdBNq8766S3Nsy
DikI/5tPGlpTc7no9CY7j4zyeKXPMN4hl0TC5iy7eBFz2Xy6IB7vOyIN0SMiWZ/RuvrGMcb5KqlV
yl7vlme1IY+21EZp+Gr0ZWosYNaslUBDCzPcXdvW+As8DVLJMvvg4WFGfmNxU4Qt2L6IDqBKJo0d
s+cqgRt4Y9pQtSYAH9+PuRu4r7/nnmY0fErv/JuxxWp2y+gIHjxLTkk/5jRSuiozVWIpmyrbHLb6
Oaaf/u4x4F9cIxCbiXHoyftOlnSjp3Ad6Fe0CMXLSqPPv2zom8xLyGddrcp4pvMBFZo8Qs4GX1qW
kGoh+6vR3WtSnaBLm/tHhxRuM4MLZct1QE9e1FBiFzfdn9BYDCVxigMbJHTtLsvZLbQDWpZqOITn
zkUxZ6wy+Oq/RSTcFdwUljNTQ68Iink4Sh2DsiekIeai6Xrpjjlo6XGMV0eGvp+rMik1VtVumTnp
HUhTEiJU/ZOiG01CxDiZn9VZKhB3N8lwL/ZOcvsmlcePER62pxdH6EWywD428pNlGLXyre6x0NPa
biefeoFVl0uyGF+EkLkmfbHjFksr3IVdOQ3PpM4uqdbYMzbNac+iYe7IQ2yTzetXQ5e/skL4hCky
KkM807SfG3fhgrfewtwUdbnXec8NmEXKtB7dliO0duFW6kBcUw/4M8z9CLFOn3rcYFySGb+d2IJT
nvSk/hAXtftz3vlIBNszRZKZsRmlEqoSmOMtjRhAwVKGE7XZ29HjqtmLleY3zyrLpSv9wHPmsm7Q
7nguHo911W9nhLJOr1BmCAMUB5RsYddyTsqvJjZgQXmJIbA8iobaGIJsz6152oKFJvLnstHgYqSe
dwnXBRxeuyTzyUMaFPygdqVgJce7hEH4SciauX6c3gtSHlHKBFITm22sdljJqStW0Jnsi1nSgFev
gGm8yUAjTcG8MvnoD9bLd/1Gm6bQ+A+tc7ofQnQhT/l0PA8rP0nzXAwFaBMNVEktJDHViUmxJ8Zv
ZCMW4PX2NELstzbSMLBvv9YSSyqU7us5K6KPzFIYziYRpPVO1CSKHqwdOojcRazrur1FTwTtdtz7
LG1eB9er0xiQ7KS+ccQ7rV6W9ss05q/oxwdEqoGKuiEWOZsTirYUW1Y/heGad5bVqddHl1F/A+Pe
tqkOT610JtxmtsYuMwdHYHnq50JNhMImeeUtiPmEb2TgElex90P5Tbpx+eWQU8gnBEqY/FGRabjY
VrYtzIWNLmhO9Pn4vJSC6RDwnjErX+LX4M8O+xpvwLW++lk/mur8PXAv9S31qnuI9JOQgogQHe9s
3AX0dzBP+Z/FRLGr2csIUy/xv1oRYh7B1CBQ3L3hm/3I5J93mPT7sTG7iVJFajKbgB4LkVb2X4D+
yA8NNImFK7MrN+Ia6KdwhiBFSZqngKhdT8dDvVsR36hswXvHhx8j+KsV2C8ukB2M+TrFyET3YPFI
IUr1HsPSMmCT80gA1DOSUafx5pzA9ovt5LD0qGvtTImG/Bkhm8BketSyUthbLjPPvRcigfUYD5LZ
WCeafqwEbSSfBH/KpN/mIu9CfijvP61zsacrFBTRGQ70gYdnqhQs7yp4/HpSTyWpwEyZwcHyrThh
YgsT5BGUTbQLombQkYxWRvcyLzpGpgwcgFBJO/9SMj3MiVhp6NF+c55vtk7CKbu7LY3TniHRGGTW
81f2E4y/L818NBZsok0aZAIvOCGKWD88tak+XoOaIXGogZu3lxFC7xtZqOBTArr+dHXVtBR7LBxq
teD+HQtlX4b09C6KUwlnp1adSUca9ManODuz8L/2gj1esmPbqDwhL6FeRn1rMpE5hST2hs6rbW0H
M7t//2S0twG+libGRLr7o61hXMyYUJu8e91XEZeNpDQXn6391Z49UDqlCT75QGwABtT1cviP8FOT
QisG8wtg2P1kHUmZNCTcJsQdVQ5aDdNoQ4KZwCQqfQDE18tobdbfnJyVuk0nDk6xy2TvkNLVlfc8
MLXiJ4r77Lf/GNir7I9rPJ42U512DKzH0EP2XpyTMk4tSIgAxCUhxYUUo38PvQTRUhmh2AGWbx1h
ZNBu2i4HoCgIBz6LGpb+fdNh+W7tBPiVjq7tUkXvJey+ExnMjiEydOsQ+UX09hAiU3Ts0amh+hJp
ntw90GB3W27fxyagbEvAJ2qBM+l3qH1n3aJC2DoOa+Zgt3Zar8uSTeqpuGUwLkcBHbgDouyHw+Fz
gxcCb6DpRYcpUL4WsKNw9A1oaGcTSaFjmI8PV/+uZyfdlu+3RYm+uoZm0/ne6YY1y292HPW/xidX
X20oOYKedUDa5n09QcW2HrnLxLsJetWPV1y7VbjkIzm/omneCyN/MdNuXYpgJ46aFHgdOmaxjNxj
H/huzQIb5U3kTt6+t9EO+1b7m7Jm/Suth4czIOhJVSGoi/ofZD4byzVhfFGk0+n2TVYeTCA/E2wN
iW4f39e+zpbY9JjQY/UPQoTfTPFexxExPdsMYUmi2krOGQ915yHKZCBfWgznRpwByFsdzNY9IUNZ
pXmopd/ObwxICQO+dSA18ljq4ho/fK0GD+3yfbDWjnuK+pNZvZCmI8Y3mk2F2eCeCujGgCdeup0d
P37Pj8e7emO8BdjgUATQZgP1dqNS6XRZwlAPyCDlsxs3NU4kPIPNtmceF8jmJXF7q7By1nzRbLqw
E/U3qW+0GBreRIlleidBK0wiZ/HerdVP3H810V6DIxZXbp15+NRJVFWUsyfC874nQHBQAzR36PRu
y8xkS2p5Yw87d5eyguW8KGpxJy11mGAt+09ouWTSuyGH5N2EEmn/iDRxZh6/MvsaG0lSDM1+AHeU
LlL49E9trRy9ZW7QEpXkE/M8jdVfWJFD9+SwdbQpJkk8CVFps2eW3jQjbpK+TcMQ0T2K0mClMC1T
PEdLWzvhDkBVXhv+kADdOCZbpEBLr2vJA0Wz/sXQKs07bxBo8scw2DIye7IEvWcz4embuZ9FIvI/
PSWiATK7nwmkrvOK0OLyQPid+xP7j/gdIzpKIycDAH5+xq/TAMY6BsUBcJX20uKl0IKqJcxN+FYb
vh/xxU4AI92i7bGb42XelYgegje6oTkFjVvE1qaFRJS/U7Q1L2I45RSbBMRQAxv/r3N7jovuw1sS
JX8g+t3UPhh2d9pw2+d8xbsp/F2lW7gbLQJGeQcXMj1nv1KGE+jnAHUCzgmcgLV9vv1uHxm3QRBV
jWZ6y8QS7eVW8rRu5DyUIPHz7EOZMG7J5lieyjLkHjkVXTqTf4WOOFkcSnk5fXUfuPLxO1WB8d8I
7wSDmjWDPILzaJA0YE3R65QKPG7zR7YuH7bHL8CRzG4uj2eOKRLuM1mfxFks9/Be3wdSHhxEcAij
Ejif820HlTAEe5zWGOgGo1bCqbiCwm/wzYRBqLa1JcUOokRjYAysQkzE4SDOZbWz6QQgSQDBpv7Z
xV5cf3GLmBrisydeqlw0DyUiPEBOgcZOLudjg7AZABHrn7WefWFBLD6ar7w72h6jfHzxVrHum04/
cQgKKRw84wb0SKEBhTjswdUOGUGXM7UE/PCrTZ6/trIRFYulS/9Pyd9wJo+6XcJkQS+sEFcptsK7
s47OuRa7So57KAVsji9eDVW+dUKl4ViZ8yG2HFZGpxl5AWBLsQidWcdc42ZysWnjiNsdBHgOb1aX
dgAzq6HNZsUSbhWThKR406F3hZOPYJG3V9AyU7vJsnruCycnzu+QLqqMxObpHGjltK+ZLkB0SNXN
dGHR6t3tGFk8U7IxszU0P94kHwbakV4YRUha7WAUfslD28yVvN/cWgAz2TUlnB+I24sN5oiDmgFW
bJaK9i+4wvOnyjCie3GmRybFj/9LPuNAS8jOh+0mDG6URmrA4bTujYi7r24G/mBkuq+GDFmVrMqD
l9pso0F/ySvggoSRaxJ1IJQ+P770RLIaoCy2al6QgvUlUnLUXkpH3MXG0GBSOvOEccmYyMNUbdm6
zVQ2IrMvYuc0y7Z4KhGBx66il++MututFyQEmc/kd79vwBhG8Yah2rdZPDDNJqBqDJq4VTBL5a4J
dC4yp8By8g3D104rrLYLokMohQPhu0Rh56O3UaWcH8QuE6Kr4mCCTb8LyjYI1KPQinXIichy3Yh5
ikRIydGDUOilIFOKLl/bfLp9IgaMvMGWIpN2S1KHkB48fJ0sCSsBccZcRNdOSvwD6IOmxmVrSsqD
ww+PI71KaNG2slk84yZLsEbOikqO+vT2QraJpO6j09Hn32fSb9J+I4j3yYW6xCjrYtwrWsv56A1e
Ztbp6A+b4uZg1oDOCIz+a9gJa5o8W8L2THX9xwD7MTlNj2DLosCnVueof+Td3Zhst8DaPpwx4/Gt
SAJohp4WZE38ggM6IYn1I58Xwc/M1yDlNYZbNOd5wDE2RcfhmYokguotfBcYbGf38bETMSuPZZVZ
xNoAyTTNGi444+UKdz02XfWgAT+810D9ZLhYJ8G2OckzIGj/6QhRdPNSzCXDmEiJIq+erDeMAjNo
W6esl8sKahPfyICfKRrz0AX74XgB1jZkikEpW1C+2tW/xpHdD4N1mpUnGPWWrHIjai26+Asxw3qI
rMlF7PI4sLbMJSwPNZOOnZS84xsgptMhbjdgkPp9oxPZkp/kLQPQXGCv+0uyZbGvfKjnV+EuNx8r
CJ9dOEnQsC8c2JvB5dFDjQCCWawN+EvH2fjg0w/j8KulgTcXlfKyR7koMeVPw/+5LJW0KgJ8MhMN
K6xGphfVu8F06FSnBGxClLgozgwow7db2YHU9RkUtJeLWUmfbL9sqA7qZwCw2XCzpOmBgbnFKdwJ
zLSVqvfi2W/576hdIVC4+95A/rbFJ4Eg1XpmdO4ZW2KPGKfo+fGGN5KU0teeDT2lhwn0k7wS0Wtc
1t3cpyiH7RXG1/nvj1zYk+iB9sSTNjdIkTjScfDtDhpHL9VJ/Sf+Cz785QA5DAkU8EeqJ5UE0cwI
lHCfJN2mVg+bHgCNRCWZp9d8Oe3v2NhHy44wQ5x694tjlHU4090Jlno+z4LheG+iagrUooSxYRaq
rb4g18LIeG1nDRGQfVcBLSY+QPsIWxmz8D8grH7jAoDgBebt7i2+LcNeOFyxuFANWp8tIfTztYmi
Duls8YMuRDuDkCJcz9KM143GhJ+xPP+4Vzz+jO5djt8nLObFr+TMKg/CXQGIVt3knlPUXxeQUvjw
Xldoodf5uBQV5Fl64DCdM6F+Ph2KP5The+ol+2wjv+qEZKPguOcNf0hbTmtAaI8ISjNrZyHy0/Uz
UiLrQx2LA6o5OxD3zTxoBSW28KJcCczUgCwuWK0YMEUyS7/M4xU3Y1/Vk4nRrBPkYGeJPwGups0/
GopMnjJ2X+L2kyPqiLKfbLY+jKBdloAekK+rpWpvkZe1Ae2nUPlyPjC6IKi6K+Ykty+1brdhc6Sz
3zicNW4Y6//FWmLb7Gj9zwSjwPi2/nLi2oosYNEaHDciYRJSFutO8rp5vZs9vvnixOIROkVA9rwM
5sBW83onDEbfoVwOZZCyo0EKX3zOAqMGei/IK1JwPmsYcCHFYk5UnToCxn0x+948XTnUYqsHdz0y
wuT7Iux3hiY3pH54JfYDgNqCqKk7jve386T4Ld1WQNAwUeEgAAsRo0+ImJPUZCeU1KgIBdcQavwQ
Vxws5yZ5CASZiIYdKXwCX9ctTTZe0oKl0g3AQzGJ87IpcoC+TTzv3d0Vk1BCyKgNvQBKScukLv5O
H4I0V/4G+tcF2Bk/F78ZMH7p3LKGMydLLwi9oer2JOMxryazJCtor23mWO1FkbQBIqCE3zu0qYHr
CW/8xybAW3k/PuGHg08lnbz6cFVLmRE13cM9OUL19tzZEI7xNpxWT2IogJ+I/+IEE2qCBqouLuRL
dW7JeJFy5n5WG9wXY8hv/5V6TpPOmXn4rvdyZ1mNbqBLb0pCLA2LpHFpp/gSLZ8Ffpddf9rA7jWk
u5+Lq3pUkdsd07qD4g/L9HQAiyVlGoqqo+IZFW7ms2a6dHEfUU5LVxg9xoIlTqf2Aq3LzhWbV1FT
m6+zIiyEge3tGByE+K8D48wOAnvVUYLeLXca0+FwNODxdb1VPKlTklqGeLbgSeLPodPifz7es5vS
hj05HaPVuusHbyBcZTR3zWtKY49roYDx29p7Ar9/KNyZIFB3GXxzb3wZLs1huEeFmoI6a9min6Sf
S1nvnH219xX4/NqS33A06OlIv5IzodNry4vCoF3FM5X6LSUghzGDrGIFZ0BibMxebaYEzB6gcGac
78UTsnDtVDi9L5MVLmLNZmThiBje0tw14oK/KLp8pA6DlgYrk3FeGZMwV6yRcu3KAIxhgJV4xs2a
RijIRbJg5kYW9/0HyvwMmimDdTepEgWp8BwQbD/UP5YjwRfUytcjZUhEqmCDCn1rCYN85G9oThjn
Pt5bR+Ebk4x2cStqWXeaaWNd6VQjoqtCdU0cTQtHQnsGPl7l/zNCzT+azQRN4ehkLLE7YCXJkXH8
5wME+HjV5cqMm8CpO+YagLSVwQcfNQKK3GiVw7QpsQx0kfWwCgeEGkLeIngUla6PFLmE7yAWlKz5
kEZUVrpO9GNnyGkPX2NlhgvpNnnZ99/Ibw8O3yl0JbYsiMOihymXqfOh98HiGQa9gKdmvNhwWkvQ
TUL1kXvHVX2dpK10mErWJaThro4XFeXj1Uj8+NMA9jsGFHPviSq9xjVdQkyCXIauPrYoEX2wp0eD
bD/NUiWX82ZNmiUCPUBEliYzPXtf8KbnpDM0mQTRQxGm6WnzFtheeqK/kCM7o+ueen5dgIPg8VcS
rhzIgMYYQXBBajVwJsk07jsNmFeNtlIXu6caisYLv4jkKJPn2oIprBfTRD8s9+V7hDDqNWzma+xI
UWTyqPt0weRZInJVGNcf1+d8+ot5RkEew9Dl1/UKs887bAEFb8jV7jPxWvbqvslSAwFhTRC7vRDf
SYB8HA3V6e6NRWQdsMEOSDPa4Y8ePiF9AZZVR3WFURGkGCEC9+Z5LQ2Mb7PagYBmx7EGxLHaMkJO
2eE483AjKF8qHLZXpQucYjrYby2Shqc/3gwyahVeb1wt1vQLeeSQKl/n55jCFw+DyX6UAsO+eiEL
bCq40HJxo6BGVLMBlxLQc4kjTTbBZfAKzf7KBiI6UHF5mdMEb7dxmJjR83pLHFdgNCExf1NNDM1w
FtX0GfXm6xoCeIvH2AVWsnNNw9vTNueV8jox5NVkPH2ZgUmmZgA47yPmkabGc5FzgUD1ni3VhlRL
HFySLGdLKbZjVrs7lwrC+8j3wW2txflXzFbst7jpRXJbbD5C5JinUufxBkNilD0nUFNYSjO+wIOP
U0BMK3cNYoF/TKaSIQLFdhUOgfgow6kW1q6b0Bst4mUpiGckwKVSsmvjNUoXO0mTGqdP1hkPtSqy
u78sUPhFvr6CmjDFo43N2krxZA0pQd4djyRbF24FeFyq8poOH/pd2GZCXTb+AmYXxLP04DADuvvV
DFF0Zv4YLsidcyjr8OHPvoil38SJ2Kymzq9c74ZBmZ/42W5+LcTHlOLD0OJ1CtuZIxMihxYxo6EM
NVpYIu4mblsUp9SeT41rv5At1+XbYQwEDF9Dq50QxaGYK5PP5bKNR7+1/6AJ7zLLtjNyZ1q7d1av
tL/c9xy/SHc+JSYZblyoz8MW2jGnGeAAa6ySfBKALpWtXtztX0qDxr5DDEnhckZ4wEXBXOQDBh1a
jJgpwHg1vy5e+JjqDKRyTj65CHE0m9Tp65k36rWWXNhIeLol9/eFrEZBzUnQG4Yed+74m1Gnl5Mf
gclSSJborKDnTIqQYhoQWb3QePC+iDjbCqm/s02Pj7pOiQfXD6Oc14AlVUzFlG7KmdR+I1nrbzhF
kDgbooWjLmAcp/FsqSR0YxUZYUJjXpKnsMsG2xJSxNJJdJQr5kMjpWTMx2TfSncSppUnc3VGkdE5
cn7RD1Mvl/kxb2/LxVN4MPTPOCTEscmKC1RGSj8j3C6O5U/sxU5nUEFN2FR4/9jxMOsviuGSnK5s
+FNY45tVrstHxRqsa/sWqR77D4aUXMKb5O47dYnEjW4w3VIVB6ZPX+OTdH6NquDBWLGAgjYLUDEf
ZJ2JgBDDJKDhmnmKx4OFOIzpvZdzmb+rwjc1kBouLDb13C3XaBz9HB2FtdFykRxp3gkntFqDbVlQ
rzYuAG/IRxes5A6j3oqIxRgEgj1JlUMNqrv6dh+piloqKrjt5Gr4y42hoTthBOZimU6g9vuSr8Hh
DhONN29C/5zgXEFu5pyOmXtipuTSksXIlfegBOrXiaDkYyvftyAXo5/5etvA52AZb2OfPkjk73za
akvFtebD+8jI9IcJh2dO9TN8bK9ReejpBWncGnwheXI6iiQNtZTH4K91PqPAIIPDCEUoLsWGljHA
a/PPG1DoKthbKwWE4CmD2ysrhsjfHw838joQr2vzk4df+Gox14jwY7tCGj75WK5J05Ria1KXuB8a
x501HXg7uQszYcKGr11LsIcCxsq2pn0lpne4nosVhBBpdKNA1VmUvfnRbxxYpMLV4z56jkNwbhkW
68PcqcCbekugk9Y1b0IVeuXdQ70JDoZBmjMR90nxiq5PY6i1Vh3yUCgeyvn4YDSR3SeNa80BW4sE
TS7l4GWFicL/a2lRi5phkIuxmJfcnNf9vgT/EuSJEu9Bw4OS+YdW1/nyfW6Ele+eclHJ/Sd5VIEy
BT4DddkslPJ9N2VTMpp8YhHuI+wCrBAS7TbbSYvRMvESgPVBEnT72E52XUzeEWYbtl1COWLf0k8Q
t+U7w8HJeYIJBOH5zNh72GVAIKCPHKZXArmGq6+hhl47cST/RBfSpPA+pd+MpiFrmmlfqv0ysI1s
Y610VkUz27Gl3Tx4N1m+gNlwBF5Ldqgd8O8R3ufAL+Pzci+SHvH1dIDjTHXhEyY/7uTgE/iisIn/
EK7VgHBSoS7XzVE84jGhWIJPJ60QFwgjzl2Fm2Fjx4wngWFTiBPfXDtseLHRrPLLitacj9UDuiyX
322aNEzNS1pTwTXCdx76nSSV5cGyq711XoUrFIa0cvSFyEcDyFTFHbjmE3dG8uJolsajtnlBHI2I
HmT6butYZg117+B/ocul0gCzMZtNdDAadt5+JXxIac9k6XFF2fWcyatvoL4jqkLawqzGG9gmR6jX
IFGv8UIBjEnMuXr2+7VZop2QJtik26fnO6j0rovkw7wU6NhW7rDajf+uscfI0GmcaaJx/fgAYAw2
QNnbcR9sGJxnsRXX3DkLe+plH1jqIcFD/K95z6CxpqZfW4xZT+58cL0xxZvB8tEHtjmfAIOzpiub
lJ9sbv75Of7ZhtVSKk0jg/lgLLz20WiVeGoUJim57WTsybwA8JUy59JXuW51ruWuy7fGquKNPtzq
BVJnAtcbN/n0p0WNIsk8zYjAK6yFW1AjEoMK06gyO9VIozB5ZVk7OL/jmdItenuen00aZNm2nRTs
2ZsCkd7YJJwW8Nh4SuJGr3ZQERbp6XuSZ4roYte+swN1eNMCaHFfvtlLkfPsP2J3c1RsktFiwfut
3kkaaGShvsStRTIMyToiShUfzC2G0OlTCGylWjd/39B6ozOX2kG3GIZOwCLSA7l2WR6mlMLdxRY2
gK1R6S3Tj75nRi4SLSCMr/7DeiIaudS+ucfXDDTDZpLBsr8/hJsdyKDQQHc5hSWybKOgFg3Vqw7r
X+qc4hzMKO64NacCV9Dpi9/ArsenkP5QFHPBk7vtTbra/uaSGxz/KOGa9FKRw1gJloE1yk2orJ2Q
cO5nJna1EnUDAORXy19cBtMBNq2dLA1Ateo2tEEw/64UDYK7m3kfXFIMacvTT4c/tI/yI/TQp5th
AFMBaCawFwh5dfkCeBwThHrUbtNb4ROpl0R4tWlmOuuSHiljK9TkkYBodKtIsS+2xICeqalE15e0
+llnXepZ4GJ5URwXH6IoV82J1gAgdaQNgKX48poxaJjiTp7F1OmXqdiz9eopDmWQlnfESe//etEy
a0+svoEM7v3zWdnTnw4j1aPhC4urZVMhZG4EOj2W+Mirs10v5iZIxLxBvA9DvAXp9O/6MHmgZqnh
4VCYT+khWrI511enwpzOcBHpbz2opTgx3ocPgMZ/r5VNzCQAleoBgJUQgBM9fxe7BfJHKFu+a31c
BmmkhFOKzI++mz7FpdY/BH4Tp7B8EW0gA82nO/2m9+hAZlLHHPTvYWcRGnP/BvdIS6fseT6BuWCF
8OymKJtmXWBIOFK5bK5BL2xNMGbuDxk3B8YnuLhxgTML7C5gewrzXd/QDaqDd3ImRcLZE++MjvJ5
xVCCkMH4MQj7GmsH5laQCQ+3QyTlzT/dNIaszgtHYSkXQtJ/d+7axZbUnsqoTmB9hGsUQRRXovqF
+YqsqLywuNvF1iLkbRpTFR3vgRzE+DA7AxA5j/W83kGAlbRLJiTcaNzb+i5yBbA0RXs4ourq0KQo
a/uNsjb2PdEGMzwOVpnAtrms8liZKSellGd3wYlVa/KPJj6e+7pPZ9L6EgqTvmUBRXgolYI9Xwjr
RltpdpP1uonf5oz+hufiKoxrtWHEuP8flqyIojL3jprP+hQk9GDP+p86HQQ5Xy7D0KwSfE/1RZpO
Ndj7j/rCeEzSUS+BLZRt8qOF/LeHwQs1r7Y7n9YD2+RWdgGWE59yFo47Te9UAY2bQNvUaixc0olg
kvf7VgVkfXhf1WLWNYzLMhZtvYxS/yMJxdgTg1zuVLsO1nNrd0TKtw3szybv0jgdYBo8B3qDtvou
21eTzmmhXyxmZlFUGp62EM1Y060P0pqnxexEQ2TU9O8tnXAGAxbbvUpro9piijY1NX0nb7nXk4dR
GR0o9qDMy1dtBIACYB+jNLSRHKnFXpxqjfFXfS2345+6QkI7iyNojWGvR2u/n1drxvvA6ITGt7mz
qvtAuH2LZQjBt7ILBGjZHBvkfzrpdTGFtmRQEl944g1KHhJtR/ztpHSTTVrrRQvhW1i/n9FEX4M2
5ex7TKz50UBEhqvMZP6ceW+JjgaV3GBWZ7ihZQHoxsOyM8FRn0Mz3gwY65wVx2xQuoFxtN4P9btz
Ykrk1N/NjIeSZrsWhFH+3+iurJ/xcZj7JrfQBVaWk+7rWv7f0MdFcERMz50liAEgQFlgwEnMTAD/
x1gCmFtpD+g8Vh1mnGxH9p2y8/85PvxxuW6JqTSVdQ9pHTHYJPMIKDHOk0O1RtW5ofyPvua1HAWF
/iun5wYZq9ed+qFAqSAXh7BUAgzGZGTKdxZW4Rxfn6MNtMKr8xdhzmdLI/dL5Dt+Bx1ou5OQf8c9
scszhXMe7mkqICrGV+cXTSEDCyHgNU9gmkLyjTCYjXk0gHEF6Wy6EoDXxsL8253hWIUHj9OVqiEQ
ADzyldiHgtz14jjjJF0TwLD1L7qTiDpErfnCRz0y+tZXssZXar5ZgXsT8MsQhn9tCSYMb4BMLToJ
9xFLXLtg0eIJzIFq+11k5Tpp+Gg9W+ALdklOzSqsCu/4tE3Ns7ruhBVa3bFBM3APd0BSkyJgOJ9Y
7tcjwNNrf5kvjWQ3uxVEzbMAIkz4Ql+yQbBXLtUtSkowcQNuImazVymRxh7gLyoQMWBX3AGT3gJD
E9AxfApeYkypEWBFybGoveL6DMS5QDmj2qa3PEKqpbEa48SBqkhhClqOaMv1CMEWhV9iDXo5J2xd
BFHT+QQJgBrHYqR4gRs/nzVwzrZFhgsAPxQVGAIXeKl5ujoBVTZQaC73xWiusaA5ysyLPdTpB9ek
kN0fW+3ce8w/UfF1DX3B9KjtWrZym3LZ+S+Qhxd1RB2o4Q81JZcbkhnuID947uN7xlY38K5jPHkO
X8PEjCw97qnclYDsUC0+bvaL+CUe9Ak6fJIhfHvriin9FcbjqU97SZ8QOyuQFQZYOXsTEodyUunD
YqQ/g4ClYw94wvUGOaf73X8J+x2pIbDwUBhATHhYM4puFWlU+uVaFBhlOZ7AiaDOnXSeU5cKM8fC
N1VWLjV+shxJyWAOGoAdm0aAV9dtfGdYzFLpIZJpU8hu2bj//dnQ9KfeQ9ZBH2csLppmkFucm/br
3hM8nkpSmgyLLpVL1RKJpTOmaU6TJbsz2gpLzEdfggdAMWbq8D43hKTKsQevvZPIYAf1mjHzWvhW
qmvqZUpKGTVdAsruVykx8Ge7rT9dgCmr+JNDumw+j+INFBerNeyKiX1LexzsfLaX73tz6F3bs8YA
5CMu6BAmh3VuLfMM2VrElAi8KgVukVmeqNWPODsSdIHvUcXDZc4/YjQ30ceC0yKxuje1w0ICjiqX
xZ7DW8Kden8cTJ76beKaSI5lP1nAQnhGvojlpmbADrxWjfVE46jYBvN9aNaXPkGs2XMC157NNvZl
AtdKWdbg00B6BUdrD0YkP3vGnVDLIyTA2VXVqG9iuusIGDFjzGkDNpzl3DrhSvfE/KXUbaDdncO6
qdO2hwW2B29FO4eBWohO7o4RVRiDPYlaQkMQFH1JdPufqfjSwR0In+EhA43GmysBnG9+Jy58+2h2
QrjBDbnIdsn946Uhiiy59m+HZ89jiyOs/5F+PAm9NVIrbobnWAK7jGMmTQDi7hNn85PFIpWZF517
peiGXXxa2q+DlU7IPvLF1RiQO+SuIeszxw8S6DScU53XktID+1l6+kEjwtIPi1qFYkEvAvUXBivi
V9xJ+OuwMqU8NSvmIBidRAWvHj569wri94TUUFc50Pc2aCKqh90QVxWdBq6E2BJkpBvwzDijKYon
+gPt1WRK3sM6x5LauJpublrL3jl+SH11uCbBGWRoIkPZnfIrx9BnchFoDgIsO3WzRRz+BTHxTgj0
htUNtiX8GA2uJRXdGiZ7r6z/t9WGQ2F43z9cY/+dQoLqkMO9t8enrCU4mSXPBxdJ/b+2Iqo6OopC
3Ar1LpfUWlldUg1NO5iOVNqB2S0CnR2QtlCumLWI3t+eL348L0oN1wU0KGvmlQ9Kv9IU3hgKkahx
Bu4hj2v/J9wx9uWHlrsU1bBHjTNQz7R30EQVA93QZbACi3m7mUxinfY0YrWiKh5yEUClc3lnW1IP
3vqpCR0Pey9l0c9yWsYYkqVmSMWSd/rKjnyXzhGc6p1ZBHf98GOJRvFQ+NZVFTD0gNpDl4OeyDGg
PczTeSjJ+UZjr5sJT+ZW1ZakQ13HpAM67cBfnJWIQPdr6EGGTzARtKVnRmDfzUr2yESflImQ1Buy
RA/y0UbabRL58b03ElDkh8K8LSTKTokWAE0D+s53rlQ6zkyjb7MgmneHX2X+jyXIbT+yk0bD+rpb
qykXbMu4JMaTWdbkURbteomNLCpnnPPna0fLMjuCoMThlkugU809cgdvy4pbYhG+3DMBI6LWP5cp
5BSHFnDGHL/7p9tAProvlJxslyRGiPRmZoNMITRZS1A6dfW/QmuMKSq+QjSbtuGNacuEqA4m4bSk
RbRHrfMAUa5h/uo0Df4F/YvxfRcb5m9Uw09MCgk50QbmuGGPXTQzpCRFtD8mC6mGLWOd7+YC2FQr
Yi9wMkGoDx2WpklD+k8J/b7JOFqRdIN4ZJbOmT0gYGGqwjwdKVo25LvI1hziTgeKGM+Gmn3DqXn4
120PiIzP4TomLOWdb6gNYfOYFYoaQDbOiXOuBPrbiNirOvluXsLFu21brgXFcAa9HdS1jUOQRklq
WGPDG2Z4PSAPc9YTXf4Cp1bkVhjMabfJ/yBM+7qpwPAujpf/HQODvx6CO5NpImtawt8Eo3s1ejWt
NEcHePUPJimjj/0mE3MepLiEcLuEFysqRyZdP1t1ceYnP26vTB6H9I8w3y7lcqFXhEbzCOGSUldx
N+mhBVCx4PZp1WMRYMK/bLTG2M66UeiQeL975tVHvIVzCCd7UvMOD2QnvKhT4VRtdS5SZG15ax1s
0JelBshWOtz9aamPQzoEHfglFsqTwa0NsHvu7yFi4QuJBwuZ2BwHG4CB6Btt9Sok0buCLQo1qs3C
GVuVUChc6WvWskzqyqrI5xmGc4jJdUi+OVpyN4u3ScmQEz3yIzR94Q5Icz+Gj7eSczaKdLY2zy0w
bl6ANx5SaGya8GzH+ZyYxtVApofzJxIi4lz6N/kLBzUmIYtslbcHhKkjQP4IGP2S9SYGy17Xca+U
oE4of07vfIgaIg5/Bm2D+ejulwazybzCRst5XR3IMLMq86aphTGfyD428LtDNej32yALvJfKGj44
2fFeAOdPXCeKjkr1acgeLvj2EYanE0NflomOkZrlahbEgv1x1fezKGlrfwb0BkinZENJZWLcy1gb
siJtBQzX1nDr3L8J/aiQ6VMHkWNbCdSgdaIcqa72Q2wl1UdmD/owmrv+xo1EEBpBcJjSldPMfc0h
3WY7dZgmao+AeoEIhizGnNPcZ6vXmdyfGed1Bku0ekx6OIB3Zihyd55o0O25w5npz2NHAOfj+A5j
Z81QEcXToVQ/SiqnTI/jSoMxvgdddwEnikjNanyRNL2I2gyJPXTKewIUk7K3A7LQsKtHyO6gF5Ht
0OXh5lUOFC1n0u22xrXYJQT2K6Nte/Qk3oTC5aMD9I7JcwAyhmZo32znOR2yHWcSP/W8oUzyH7g1
KtiKIQ4aePsH/tq9B7b+q6TXJ5SsUu1559nRq3k9D/I1q/m3aqqOu93BUZkld1cb8kYZWKeJf0GN
63Dfe1zfNrhyptitOco3FMe0Vv1cMkhSsdk4DhWl833PWD51jHMqQyhBlGIiDaJTqoksLU5Lsm5J
TwB563h878KGZSq2WdmnsgqOK5y4/3GRy7FL6ChYND0cH2CfBZNzsC5dG9XgWfnS8ztoaKm5Sc3U
ojsns00XmFtJpb+4mJlV2lF9nK6Z4H7dGM40v+HR/EJ+wJO2BKMhYUq33uWRNHaEkzou2eebCOAU
SNSIxRRSi/ZXuOowDQi5jW2jels0rv09erym+wsybY8SoZnRj3Mi0B5S6p9e4Z1D4qIol0lrwwAG
H0RK49B7+2CJdsYaIgGA2nBDeZe+QPTQOBWj1DYHJ18MITtwTSyutazPNgQ0OEGkZOK7XQnh71Tj
zfpT2AsothzrUtNhusysu/vYfgfLO8ZMuIOKBRM7+lz2n0sgu4wX0Z+4kki85o64bo80lRfMJm+X
hughxVkhblPo33lyfB1TnnEROpIdmB3Is1MsnFPx9YBMffz+QY5fLv6/5RMIkjtTpb/IaTjaALEC
QyjSGiG+iA/9YL204p63MMVDs1QOLFuqW2a94yYSpCO5LrmaecRVWDgr/6itPjbo3l9l1VqhP9FI
yZPIlk0jQKTWLq6aV8PFYtVtOpW7EMIm1VKiOhIRDJd9Cuu3099oT+cZtNorU7Sxtd3FaJszJrwT
eFx8d8PIOaHr0mZS4ZUueHEdsxcUViPmKXIKb3bZWoyAJWbfUm/Jyz25iyGLK0EerhuEUgt5K5N/
B01svugK+tyA0tcxfNqyzA3IHXXLvx6HhooKKO06UZP3eHC2LsvCC5pVvnNw+35PgW2NsBF/nUgI
0Xh/YZU76lybmm5ri+xcSTVvINhL/5wQTPqTMRnbRrN35Yk2fzhOdxFymHWOD+tBdaK6LUBgJCV3
rutC54aLKmeLayVLcW0Ti7qH6WQD2Ppi+WoZJjUTXb/5OG/8K7nOSoXPxlgte7+hH8FPlMRRQ1H/
CboCSoRoVQyv0pgdV1IwlBBJNCCACIgTXkAc+a7aALY4ENcSUoseIGsiiwGyC0C0SZLQqmN4Aeso
eDCtTCZWrsg7QM8cYI+vowzQs30bdEY+KGoaCskAYVSzrRcKTJG2wdfMBiejEOKVXGVo4LPa7aVz
SCAva1GYBCRPUQqT4jtdG4spJHPSwRLe5dkckyyTvTkF07FX8gXI5oJzRgvG3PUFpfVARx4B8ouv
cii5YtaGQepRfPFLcHuwzEzPqEPI2eHQv0UAKzrSlCP/Kl/U31kTNOH8l3iLkTTI4uhJf4D+W/9G
0t2kkSVT8IVJnzFiTfVWbR+XVRp8kB2b8a4YLXhEp/EWYT5in3IR3yceL50u0KfxVV7KmgL8d9if
+lmhALd9L478wTf12gWd/v+mrA4uVXLSOy8WQ/qw4uPaslWkCbMl/q6I9eZSbYJXwkTqYia+cuoN
+gTZ7mRwyssHC9Q19mH0DFbRIamyX1tJHgUJ0+HoCtvBqRWBpUHxucoeMLNbqAPW+UYknBTbX91u
EWT+AEHD+flj7CBcd18/ahAk7Ge2gHpsaBIcz3Q/064nR/nR3LwiCt3PfiV+nRYLjZyOJaUNEO/w
LwPWc2H3JueIG6LlPY/q0xr2+CcTQuAASVdMDJjPaIDlY4HNz+KlaMmqFA6hzjI7Hp/gsuxydUWo
D/1MSEh/CUMHFVCDUX2kOcYmzDB+xRw515IrBniWzy0Vjx/x9S7qNpVXn2I2LtpM3M4zemCflVhh
mWI8nJF7RZMqLzv+sIdHe2F/9X4KPopLsuhet35sM5nNZyuFOsg5WuFa0FHFQSf/QHXX4RGGGxqm
m7wHIqGXvRiZIQjUAIMBSTdkJ4FP27IWDQZjvxSjPIF+QJPG6kFo5wRF5ZJiogCR7XkqrmXCmpE/
0o5w8DGnHoC1sVutK74K2m7SNNUC5WTaDX1oyfSTwszOCecbXJP0G6ROBgcn3yQseJD9v7w0R4On
T8uGavbSPVkNYqsbLaUJqwc8gebYCfcM2NECb4t13f4OttV8ZdlXOIa3fIYaFf8J0ZgL37ySmJF3
B9BiBgK5Nk3LvD52FFjzvW9GDWD/sf1rvjXI2V89L3qqDvOnuaAyi7C7eOeWOX1gFHEiop+dSo2f
Bd9FLytDIeZjK9W1T40HO9kRZSnD4TTI9qUPiA+gk/rdg9VfkaIs+Z8Gn8mxklenijtjYaetJ6Lj
WqMYsKfcGPmiHLh4j/hAzU91n+L35ZWudMMVgRC8bohOrCufukzpwRcppnycVoXE+N6uE1xTp/8t
/50uVj5hQzsOddUVa8ZSCyfaJqKJAtoYk95GLjYbfT++uEpfOGrWBwJCUIvzPPG2K9PDzbY0yu8U
mwlleMOYA3o0xUejv/SdQzSngLydQWOVfKgjsxQAjBgf0dzXhJe9EbQml7ejYa3L9MHBR8XeGQx1
sDrqMRpMHOSZ6S6upQ+kSkse7+d/BU8T23pdMg9FcOxHN3L5IgrTU+IKEuSHDJpVzmd1DVbs+kpz
Je6r/VLMzFQb0xspDUyAfywaIC3uPAVizuSSFt2Qyi9tYNwGuYxqIoCeEjvJ+XbLr3qqRzr2+YV3
cIl0jSGoqicjPJAQgkQrbVl7w/I5TmDxqoyEDvTx5yYhPxMSm17ISYFTzaZbye5ZbyTcezy4m+DW
iAKbbZN6rh02RdZc3QIhgAie/02V9BkBKUsHCd0tgXma1PWPvwBDmd0r+4K7X8GXTAvU3ONBK+IC
k3LhvnGobPq6dfQkceipM4OliRpO9ydzBJTQINY8sBOypwht7Ov+ImFmwB+6E/3TVPjOFP6K1uDF
JKBUTjV9cfvsjSqUZ8qME4APDeHlYFOn/JvvMR4TbExjfceN2U17S1dtWF97hgjjzUiWDF50OPla
gROUPCd6Cns/FjKVjuAdHbqFQ0BKUnvJTQkpDORZJjkEeW0QjXlFXek0IyJtvt/lOz5O40r6xsK0
cUBn0R2zCjaT4J7ijda9DILhFd2NkATy4/hf0hor4Ppke1Ku3YFgxZczC4Uxz+uYmqZNZjzhYVtR
KCTfb4F7UBt1J16dPTIItgfdjikkZicaKvFBquVX22GUm69Z86hRONaEMSVtWV55CpNQR5f331e0
ecAkAorAxH4dPu6qovaIRKfPeVH7SDSlhZI2mhkRWLlQWw6IPdcNDldZoWNl5JGLY7huiOVCH6Vo
LlrndHu5KjcmaYJWr+hKmtLFXWJ1VGY5B9J2OiBeht53y7IPylF9+822tepxiGuEYrE+LBBPqBgx
Ck2j+/Gioe28iFEVFLJbwbdbJtCvC1nMJ45cEvXs9qpLvRsPcs0lgLxMmyGfDq9X2Qn5cY+VCEcm
EPuhGRSkw7qlHYb2af6fvlcntRZIYjXSs1RXqxY3vnm6E5cAWT6w1Y6wWrvVja4v9BMBhaHilmDj
aa0mI/3ReKQ0PK5oaKwFHmNarULRqFMybypeRTl9DiowvAl3WGiw2pDVUC4uSiX+4ZHojR1necam
MJvjFYsMy/Yj535cx6PSPS28QmZp6y1FhN+SuTp8g5vyW69sqH/ge1f08hD358/rFXE1WUS6A9d0
FiLfl9b0Y+3BKL4cQ7ZycCX9NnfXfnhhGwySMEZTB5rWbRhJShX2abx552MuZDdKB1egai7Vh7BB
icaX4o8DbHNSA6rfC3qG+eG6xk2AJi2Ctrz8INCvqrh6L8KJVx7iqsDuMt2gvs7SlBz+hyZuxvIS
L09YNSBU7UvPcxDT2o8Ef5SuMjOLkv8gBO+ylWtN/vGL/OpdENL7lC+K/KJU2sMobOHgmKpLO/Pe
kSs3GOQ1JLuQOh2GStdTNtTkjSiCgKRrWKRj0r1bxTj1/0sSpsGz0kbIrvZ9T3lNTAMTYX7erOfh
ClcKIAd0ZWn1tLFHjEg66jhRlgB46DhTNhWKgH3mHxy9VxEqoFZ1kB3xIcb7D1JZORHM52lvD/7F
XVCl/Wp8UVc769BiK0Ec/tNyKQmlRC9oAYZ1kvXVlI21DnwOSMshlOMarr+1AJzNQWSQd8ot3gQx
tHzICFHptnyy/O+c5JuZCd6ljllaH3lHlcdBJu4A7k8j4/YRNvpTHQmjB3BIAaEfUlahGxJFTru/
Dppm08SqGfjVurW7DQzGS5y186LChNT0o4VeLrC477KBPbqhyVP0D41jeZPdyF8EkGR6X4+HmUpR
dLj00KxInMgOGXMDQr5GLiilyzVxd+voG9511E2RgPBza+Z1QQUArPyWghj/SQv+D2ydT2Q8G84A
Z3JGCU1LU/i0OfvFP06QMOoP+xKfythTN+hyAKaLezFbA8JE/0zknnLerSapPYHATtMjBakZiySt
gD6Xp6y/uzGiSm4HJNnoiSiCeI2vizta6S4b9HkbhiaQPXk6e3e0VsUVttTuud84nF6DpHOO2xFC
twnmPuSqBidG0Kmf9XfgYJ9F1RFGWGlKTTGNcH0qrikXTJW4PxAToGczXBdnxgUx5Atzl5zDpPsv
M419ePyHgf+LsdlYPq4XyUOliI+sA7u/fdxpv7+WAWqHbH5milP7oyUuEcZXKA55ax2ieEL1qOcr
RqkEHbsyN2S0zDJhwxf7R1ix9UQf0Z1RPcXBHLmwZ7NHDSXMj7nS6hHC+/Ta5lEZpVGsC29jTklm
ygMA1tAVJ73pZIniYmaCpcNMbpVHes0S6kslpnJexNaUxxWj4VCdY8boCnMr/GJ70VGdc6htXCWl
QEaWDubHr5R/wQTgACLiiyP04/V4U/vaT1wKpLnFstE+vmmWdxAd8V1lD0tnxOo+IEgEE/PuX2IA
LhJaYh4ITJ28PqVnY+3Y74AgT3EMxYjSESFctot3lFDpzkWn0sm4e+fZ+1ZrBwwDmgffMYAfBjCx
yOiG2nKxQoPAsjuJzn/GfQPty1l1pDah1qxU3V7gWk/IcYEHP3FCGfLSkfZ3ZUJ73iUQNIca0Ig4
WCkiUR0cyPx1iVAIWo83lGzV4tEzmKkYPoBFGj1Z/QzJ+ABej+F7l9iAA1QZkUmcqBiHaTZFM+6R
2mA1OACsqdyQQbPobNw/8qoc0G+fooJh4BzNn6nkWSg/Lx45NCJKmUUxRRa6R+sbLIs5wguKNpC1
MoIZP/Hb1A/HeK1d8BDUUzWVFZLYVzlxK3Vmdhazw1YQG/GLAt/o4brxk8X/z0etXlO2m5mfYiSe
R0iepgeE8qdRwDOxVYhU8V1yHZ3KtgcKD65Vtnq2+5Dbugv65Ex0R0M/UOQkxKxOY4lzVrBbcxHQ
yUQb5Cn+uK0JFHzQm0WIg7k/jlcdmOaSiGPa2hRHEyDI33hqxEa7U6bSyFDe+KSN1CMN4eM9czQr
1QD6KEVV/kcOEEuJK47s39KYeMJoZmLUtkU62AkXjNicjGFLw9YfCG+s8cowRrEd+NAbXOIkz2R8
5e6FwgTMaFUh43bcCAXcGFsIq5wHerokKVrs0GP1gJL8VOcqod82Dxthy9yX51xtzVsglazP5pl2
eAVtzLkeQNe/6qB6y2ngRvoZLbTvlR64XF9Pr7hqC/A1piTYCUbgRhdhYH9EDGp37hNcCddxCi4v
qQkNCVHr6pzzQ2JRGPMH43O2gt7CpCMbeFMXjL46iQC3li8xZBKrHbStBXxnTEDAMRXuHtkuqz9I
Ek8gcn1OzRaO9yX+1+wP/0INLqbHtEPePGK9waUtyIWRN/MsLGNOHcL7gcn3JZAkUHcWgvXxf6hZ
mY02XzrbtqB6U1PX2N3or6AQQeiKWEioIOHy7xOQbhKJOevYoABEhx8wazSkkylyBPvrKN17DTa8
8rfatoiq2EUwqTHlMm99d9mgMwfXYC1tX7jeJjAVcD9z45j1mjWzecMgraEykLtJ6VfhUtaStQy4
WnlfS4KqhSNQgkJe0y3gD3gEZfKQEdyshPUXJmB9yYLElFrPtugNz5gMnq8Djb4lanWLqu5Z8BSs
rB/YCVaP0rQqTCjuV2YxLEpYxCNtffH9y8XwZP/6pRzVA/74nieQjgJVujjRRMQGx29eKbsaB0p8
jj2Pu59rjZRnRee797UyITRSJUQsbLgfhPkG/BpflQJJlEsIWXK8/UeWrNFIUreH/P3auvSFeYfS
crrcysIibTC8uVfL1HlZbsprq5mbMk+EGxj9S4X3sOBwU9QIrxndhx4MLpP0n7H7PB1ePY+gKgYR
klBEEhTxC7twgCXKHVZt6NjtbaAM5gvHbj6BoK63kImCFt3edxeSbf1EzFc6GbdI58t4xwDeOOpY
umRcb7GAXfcqflYlRPPOv3zwt3hLLA/lV2Gw6xY2vUaGi+ZWOwi5w+B2FvnCp/ilsFjax+nCjY1u
grGt8QgzKDJ4dpFL9qCBW5pHYP/CBTLCYHm2uEmA80gudKDW9lk45d6Z8oUbLnKxB/fOY+/It4jT
FXd/aGuK3tqDisMqMNUwBgyFEU08GHFj1+aWdpQPnQKB8/lfLmgnqnB9XPq/IGlk7SUeWsM7R9Pa
3bol/aldmvQeZ5DLzQLzn/bLVoDC4o9G3+w8IMjj6u4QE842KbD/uVzmvpFGYvL1EcvxhTnAK4tw
MGnZ39chkrRUjen+QDBz+X1AJyCkXKx8YsN5iuJRA0QNLPTkjqIa8IuqNq1DdzJXhFMmfWQPUCMs
9VYVIQ62iVYkgGOQL5cnOoPUsfnKCrfts/mdskGcR1yTScY5XarC3eTY32aZrI5mk94hCPyN4i4C
uSkuCqO97Ce2JLfMOKYINzC4o/1c4vDiugPZlL0vO+pkPIQMre47psEK1z4ExnYI2QJdVPElAR+D
M912S95D5PF5qfR1YaP9Gt0r6wlfkBWBA9G2W0R9OaIOirULOy5zKEXuTtlCkueQsnXUcu3AySpy
0lvmikQkWpAOrpFsggcCVf9ZK+6vLc4qjJmSztAZmQsJsXVPOQCKlGdr369JCmlIBnsAnH5bi9tK
FB03TdHxgIKBQDxM6BXZxVewCuZCjPAh363U2kQ1o9pMu2Wsdr8AfvDHEzC5eAO+SZVmsKValq9F
PRsA8OzN98I5sHnsHp8tA7FLjxff9MUup76KclNJRy8ZGKJ/8KTDBQz7aiGkbXzhjQVnCLXcOciS
PumM9Aan9GBghMF5yvMTA+7diO6CJ4248DYtiF4B3B4Fa85nU9GSO4PBzVZ6rOX4a91PB1DIipsz
Vnf813c8f7jfi8e0Apg1YktL0EnVurLoXEb6IXmML1mk1HaU+8MTecAvKs/7MwwDuR8BXpD/fno6
sZUckG4I6iqsFJyilzoF/g1ZWBl5Ym09iDgOSxLIf5AzijyVleF1CxvsrBwzEE16bFgmmfoQzXKy
FTcoH8g2dSwzzePO5mJDAs0B00sV7MVkWP9TGV54ejXGceo+VorrsiBe+U5s/sFnzTPCECtZpw1v
2xBG3/aRtE3zDvOuEvijy7kNXXr1krj4aYne+AWTZmmG8f81z5e+B3Nsn6dIGT6z2MCNbCZCRSgu
V8pqSEbeANLIg2q0pvaMoT6NqNvOOqfnPcudzwLY3GKSUBclaYqrAckd7fawTLGdT9Z09vZT/SGx
cD2qHb/hmTsX3J3fNpiINQct70cmjtPZC1+ub6uE4mzrx8yOQr7JuXbhDOt3OJ4uw/WKiF8VM2Na
aGVeypeiiHoPiQWdmRiJrotpH2vxolPKWSjS3nWeLhb+tiiqOQ0IC65oOiXSqvDhHrSr+bM3iJPo
QhjV7hfyPfmIGYwmK5jV2Or5eGyPPw4ZcUJdVSGzL+Z3EgHgvDxJZNYngRliHZjZ0at/x2zV5JsR
TOcky9u6shUXG6AmparMhnrWr2aZNPHwTNJ4KADMRxGakoSeNqymE1Al7xXjAO3xvt3gNCusNeBa
ySC6faQy3ziM/0C6VBdZrv0fj7KdLhazgxbJm1X3zuVXG0dc9vZdP9Gb/z6Hps6WeMUkRX+MsPZW
7drCu0tqTqgT8rFF3vgMo3DWFpVqYuZdlG1xOuQd6rm6zbInZ2NWZT6symQR1z+sowO2KasZh5Qf
0GssNp9Hu/VL94b/2pdUeQqJsNhMKHfeABFsMtBmFVt9qjQ8ZZ70BBc3wXoTzhN9zuOGv8Wi8odD
G/9eSEzisKYwOrRXrfMgLDImO0WHdWxfaC9JnvBgwqDdM0XoKebGW7JbHYgNKBf+B7gs+AG2XJAW
1vy8WXLDb55PsEh9VPyNts4bq+WAj11BQk1NxoeVqJVzIvTTZGErQQ0ItNdGINQjmtghWBqXl1Ys
z3xx70UBSfql6QhkFcAQY4WWIgR2URrIRg3XpM2ljIWAYXin9lD/tLF9as5wcf3a55RqIHJTTrgg
xn5jWPOt3WmLCjf//nGMPYKdG50nPgMnLuAJ7MlQZ9YOJzWutDHSn+hSDIU8ZGG2taN87L3ifbYY
rm0iIh/SgHI6krfvyfuP9ekScIKE0URZZXwXw1iLFQ6rwRxYLhjtpOWZxCkIqDzO7AlHxkJjyRfF
2NRPAiUkIKKPLozD1o19neZIfR1ia64Vogqx4KF1h7HdWJ//k2jKZS5aDBZmi+UG1Tcy2vAa0vOD
arXptmESdHFeMB27pYSTXjeUKxxObtwdQxyjfCFFF4Zvt8CnaIYnJaUc7Lid0Mfly6gCnRZxcrfZ
ftZ3RggkC4lszsSaxosUbP9AIS3NrU90OGw7DVHlnlesuMSyNEcD6pmMQ4iYX1HYOsz0vrbXVqnu
4KSw9aWHlrZQ88vDUzH1b8ivu/DZAW52CbkrVuhVJyVjSW6Ran5vycqLq6u8FNnYPVhzBQDest9S
rHY7eSJTL6qLZVsbwsrTcAR25bBLakVfYR6vScS4JTf24ep4ymlZ6QSINaJbuoWatYnJrClWcu2o
SFKLcGTryvlFHIx3lPwKUDEnScaw6yPJdq7Zbv/DZnWQbA21J0T/VZe8N/ymKxfeJRsXfRlw8D0P
h0zp/iLtOGDLh8wbC5heajaVn6asZbV7vew33wYlFZES/vjBxY0S3Y3r+GQRiavpTXoAOv8kgkGH
Shet4xQFgelUFRnErX1RuxKIW2FuUr70b343R5JtKc4jIfRK8wistzlvgxDC7nZpmhFEpHDbTx6f
Y4cSFDg0eIh2O9tvSOCx3D/ZUZO6JBmaQf0SbEnGdLBiFc6cDZo4t0yGD+pHvh1eBH6LKA7QibFY
gopKsR8aGzkPJhxWbcKIDbS0UXxK43CpS7L10doLKeGaUyhczRuPSioiN55CsaE5wNojiXY/hghX
Y1IkqdIqN/PQu+67Bqxy9eegEOypsI9PS77WZSzjsvCu7qaJ8eW/Ze9z36IS2NFoEW7Y7NHl5cSx
dY2Fp6VWWPYMXlXa3WJumcNjpJeQVIVJjaFDnll5mHma6mbomoYl7cp7MkYBytXvsLdA8npgoeah
4YfnjTbcKsQShIjSicCiRzy/TfpHLrltEiw7D6WHswoEM3CWs1D1VL+/FeVzK0JkELueUNzuv0/4
M00H10pJea9rSAIwCYLX4Vu3FZrxlF8SJdo6Kle0wsvMqwEO25+Y6ro2Ii9EJDM3xs1fvgch46Cu
388KEP4g4o5Pucebec/bGzLdt3GIDZ4w63iAoFm2ImZZ0sapINXg1LFXbm8i1NG/O0dBohhmxFTE
oSKc/liPXHfK5JVHgkBUxsdCvw6hp76qC01HLE57X8iDR8wuXteD5Qw6j52VIegcQTRmKReLTo7Z
DWRzjyUnzejKO8r8MCXB/m3w/AeYt/QaPpLpnc+6/BswHwGU0nOFKMLbcPzyZl+rI8+tbEUeRZFe
LsHGOUkEFrCt6fOeYiBlvX+lND4gfe5NE5dlJS8vNjj4zaYrD8KwImekFvB1pAXA5NChjbdYYHx6
dezKqDclfdapJpG3MIjIOOQFZe9mb060HASuyYcF4RVrJ7hDb+UnmIDvNIN7AJKXGFmiuK2qC9//
3oukqRH4L05AfrboF/RLASMc3D5L48L7QxdRlXnMk6WA7odCLVdsKhcYXqpHrf232LHHVO1ETebS
qwvnupb7+MtYouR09J4flL+QzLMh4LE7zTgUowZSjRFDVZX5ppglNG+FHtunDfUO2gfx1lcVQM7t
XWn5g3NLQu6SYHmhK0A3Xl0XwEMsRKGgnLsIj8n/vGvbXGwaJ7cgos82MSqpmrGlvpqPLNTHmKNs
LWVVE+ZXgBvudPtdXVoa980k4qNf45tJjZMJmFIQhtNMKN/oAxPZPA5GIPV9HqauKsU17Swvwsb3
MXhYEylGx4oQIxXx5Z2p5KH7YlEiTnsPsMSgO5J7J72ryy0yvf0FRCk+EpjAXPNlbnwLiwWjg+vp
sFAjIqUm9DiAb8o0/fM2yFp9nbYLVMfofTukdZYxNNkzuB+DPCm4YIybGwq38G1f7KpMuMS0LvBY
t6ExRvDFa2g4oVsr26OI2BGhvIxdD+wfZJ5cM85hgv/EajhMvdPWuJVDTFqzTU4mFYAlRXv33ftT
KImNLJVk3v/n5K8FQ7FJL2M6bSdDxmtw4AAAHc1uu2zVs5cL+81DrIWLvoOZuu5b+hsvlpD1O01e
cAz/N9TlSYkCyTut8DPGqzT4bC12k+QxSmRPXZF650xM0ZhQ2SfAZj9zOdjIo5VkqHlRyeMjJ+Bi
QB5ZKj4dR3XIc6kBN9TD39PGpOETDmXG4qc1XUrnzyHkxm4nRy94mkGv9ZMmIOpBUvhrxppHCOgX
KFDxDSpv6rOJvTDBY/6MbS3ISbsk5HtFWjRqncwd56RyBko3LlF9Hhurfu5GH7KNqYoS2zrXVQkJ
HEIdEVxDbyQmwmDQVyfAUwD4ylkPasr3bXwzuqOTzaz7VhAZ241w4FeYmTSdA0EEq4QtpJtxeuWG
qNJ1GEeITncwnx8XWsdq1XlULXSQeex3qGCZV0nQPvX+dLPIPgU+Wg+tUaE7wIb5qkPH7k04IGkz
65ZBMePrgYbtbnb+N4pZbOV242pQ6g+52xb4vwHJreXqvVQ5xR99CwzCCngTVTyE+EdkDc2H6qQ7
Eq8DPIYnnmXkIXZ0uXzuCdK8cUQOmFpK3Kk3+V8W2xBNaYwcsFlN3mis7F/RfUOH/y4GwQRIHu9z
ytOMoUIpKRACT+mxJ7+DkVr9adhbMiJbybOsWnTP0VaM8lf7OXCNqp/0po8LjdXJmemEigP8QQIw
UjLX9t9Jb9WaGrAMqf3gsY80PWWYoCypWIEQREERTckPk16x8R8JlHNFrCK74nr+M4prXgIgtaiG
VkmnIqEmPIqpmTt5EkXbDdOgihFvQNUv8WF05S4+ebrnPspznU5fXdZIla3jOGkdnsjkVDshqEx3
e5TbfNiP9rg3NNuiPirPydlW9AZJSyXgsxzJK7/dfVrffdXmz/7seVAktLp76WDblWODdUJr4/LX
jq3gHXtbeVhzFAUF2O/bHjQnBmLAgoeaeObv7BCyovkfgx5/Qieny2xAjyb/7W1em/nbyaDIXR3l
NzFzZkt+kuLXnqKCsxKPlDrHp80f0ka7NGCePygt+bGn+bzJg16P429qWam4dVfS99IjADbsRbfF
HDte2vIgy5wP3i48PSvtsol7q9lYLXA4Eef8tAyRA4csyT9HMr3KBhEf5172md++aEoxR04eC2ak
lhD8q9jke9V6wloGJqLAdzMnFnxQUltE649ZQSddvvLqcKjPnRYiFCx3sZUJjIC8c/ppqfveXC5X
KmLMKYopOGFkmplw34G+huFejx+BGARXUgJn78FQB9Qe+BKtTXAAzOMqY+BWXv1zbeuJxrI4bv0G
rtj8u9Z5a5UcjPf8OV1bTv0+Gaa+X9zmE6wJNrjIHmwvkjlmyEmESAQiTYnPU83Eh1UhGMvKFCBK
/IB21IS90B0jX3gUCt9Jaj5qFsX1Y9MQXSt7RX7AvSeYTb5B3DDporIrUomZk+VFfip7F1SSkO01
wSOpGZoOdLojM/8KFMnuV27/RQfZXJkNidoozx2P4uGqEF6uNAKAsjUmNPKJiS5gtsho9jTCelAA
rPL1p+QBkLeIpMPc25pFk9QOJG2A+360f+7bHHdy6Ce4pv+CF1/DULB00AnqXRcHBKWj+wnM45NC
cZEwTs9usEqohTIc3CvcdIPn6zCbcaTfB3Xwg8oNkfzZsDSshDenMw1VfwfFzoJe4dQL/2/JZKVc
ETZUg57QhzjFb377F4+4HmX2GQMGKCRmh/sebQvb2AABspFd05jOriwtI1/D7y0kPx6km7+ZgLLg
2Beq/4CoJLzZ0icMBUeWcXBnDGvrcY6AnvHm6aOQe9K/5+vLfOL3yG9VClb45FYvlFhlBOH/+ajI
UqcP4xruPh9J6iW8EOJ0MLJQn+09PdE8cIrjSmYf4B/O4mRoEptun0gQLBvcCSFL8qiytdHum0uS
UfBuoPpuoO2Y94SQRi636KJZGeT9dLNHR6TGDSaDUVKUhZE695tCdQtJgYPj3UJ58+SRlzwbbFto
b7Voc3koxGflMeNeIc2LYEP+LjMupGFdQGnTBMiYPoAoHGFAbTyknezQxSSrOvaVvAP+/9lwMN/7
9i1bgBQ/OKDuW6kgLIkA5wCxq4ZoGT3UXYCWPTWfrFqqzKkC2k7TSEe+sGiF0kRGwI+uEbsMLM5o
jWZJK8plZsEKh9MERhQEfTuSYS8v0MqPBuqAJM4KZ5w2RMS2sCGFXpjPcfrwSy4zTcipdqpA5YrS
9gI7w6NyS1g2t7HJaDSnuQmSjiB4WhbYn+ofvE8tRZBMIpGxE4eAwUC4oSV4Ycw7A6n4PwSHKysg
NBfTkJzjT/Lk9ASpNQqqBxV2Bt06M+G8TLCrG+d/TRyjRAeMyRznSnjYtt8vj273F1+L9+Ppf2oG
p5NRBaNig/sTgPNaqKM5cFvIqIB9JLDVKc9TZ5jCn5wszIdqYuQs8osKkhH4fsW9UU4OcCDEAtvq
E8laHWQL569SB0C1iW2BKQkX2L16840J05iXZjATswWX5omW8P2f+fx6NQrmyWkF6UY/oqMNYEO8
+4EsHlH5ZJoRNX5b5fWCBypf+8AsqUERuOF6AvvS+TWkrKIqW6fHoVF+sFhYnPwu1Fhzv0ULJYZU
jSDLNcqZ8+GahsKbNDdLnKOAMq52T0SzQKHlFhi5JbNlJivNHU90H5V7chefeGAhlfHLbcwCRgPO
4vZWRJX3Gg3+n3GUzUfC0jZt3UBMY/3SRuMVmSdvXxkp3IByo2Aw2ZMTchii1QFOY84Nv9a6K8Et
Ue2cKCyt1CPTEYcBgccAk/Y7SS4ceftfGKzTQPvKUbAnbHbeGuHi5TKLV7WVjWMA4R1tVUZVzw5Z
BWbOSNwyxYDoHXZY9iPWOZDTEBl39mEGoN/weLiiI3A6lSINVr8fIJ8o3lNul9V1/oxHzIl/q6E4
eumigQIdN+Zn8fCp8P7xxcDEUSPRaSU/W8s+nk9RILz0/WBhtBSG+P4HocBZtwvrrPJ61Lxjto3R
UXmlmEACBhvuJNFadBHOz/7zEp5NWkwAukGtuHLW9tfNa1TJONh3X/rLCMXLLrhodgTjtm8QR0Xv
D44DChaqBufUnRxg97rEu+KfqYIRTOXaHehtseygtLnCRn5QK+AEq585SQcN3bq5plSzrdDEJCzr
P0Za8rR0mge1gdvuMYKMdCaGoSimwX63i5icJ7lRctvDAc7lsgQVWA7ozkgAwLyrVRiaeXksD1Qv
VXHfdCwW5MyyPhPTN3xmF3HaAqi/rkyYS0n6wIeLSHKAWwbdjdGNeFXPQBP57mFkJ6LIGDoarHYV
nQfUgiXustQU7Bu1PgInPFPQQ1+FF7VIUl5ksagziEyEOkYIkE8wnpUce+dBMuV9kBSbNhH/8MIE
E/gDDGqt/CprfmovyyJql8rB43/cChZ62go3dN5vAY/uLMcMlA8qQpom8RRlBt57kiERq3fMwiPf
bGZmMI4s1RDIOrjGcogMfneBaVc3/6QjLZxi9VnkRL/Mhyf3nqnIfhkkwfPgzmpo9fb/FwfZdn21
cadS+gr1vx2xI5uaoba6b7Z4i4hvc/clAB4kiaJAU36k/KdQHNrnw2Wr0XMYQNf1QYWmXrP5dJGy
Thc25f6ydQMTnNq/Eqyfsuo+5LPZR0uOAXxRX5mBsRkzaHIdBcH2ehD09bQySGoGnDSpy5i2BFBE
p81eo3My83unDG1X0D7+kubHnTNC1ucgytpI5FluVQ9IRxZlGFd54qTKgH62RJ6sbOfrBQ24KC1q
6syDe85ybQYnCm5RHOxg+uFdp8BU3H+XOG9DhO4QmixIYNEOLQUVN20bw5UCLsLne6i6umXHgBdl
vtgouw8xZkXCC5wUswRWhiIekABY3PehE0UDC47SowGrzyxIjhXRgmLm4lX2xWin+tjUjQXKZKlq
vHMi1oo5sCtpzTVhR6AH3SzX+6JicU6/ZawKu8Sc8YWtW7AThmuqsv02AchEUq/5F++5cypgwCb3
FpbaMVHlagP8jhGRb/Hbc0npbgSXYYVaj+KHlLXYe2Nvsd6dfkSrRM/lFbLd/rr4X4DPmUohJ7Z+
FgFcLsqrTiborHgufkF/fqow0hleTIHEntdOfMSqT5rd8/P/19jwuMhaSaagf+eG0cr+UWC+ahQz
9Ce1+Z+DMjA0txgh1Gtwfk42hxZ6nKMA6hHC6T9SzoEeogYOZzyC3OBPMo/qJIBs4+SOU/gJWgzL
M7hqc07IcRo8tNG+bFHMlB4kp1pOfbCrybjgXnjRYQK8k3UIhpLKNt5kCWvCsiANjY8Jx3RdM/wZ
7ukMa72kozCS70B4gUizfGa9hfshqPdSHtAe+s+AU49aQAT8E4BHad6Y0vpnnT1m2M0UfG47mC6m
NUq9GekXE4dzcjo0dyrDEMTY0CP1+x+LawxZnAt9tFEyo0/QKTFivDtPKgUQlIJB97Ja+eGhnUZl
KA/63vc3fbNYz2W5/vL27euAOfGuCLLF/ojLKr1TYY9LvLPU9kEehClrkJYNDsATOSr940Tk07AY
ngn83w95r5PttTA0Ey1Jpj+5QxG0dojTdnn96wMo9nacG7FDBSxtuNzSF9cmwCBI6Yo7xKEcvRym
nfMULy/0OVYI//vtP8cz6ayC5O5z0CB7hJz7dpq1UNPciwGBHastk/eOym9K9K9pfznBgjJK4WuY
FE54w7lAHk8WOX0Sgl0em39moj46DiKtUZwGR70cFLuStOPw5pUZx7g4EJm2Aet3PmUrBs2Wvujf
WYxQJRfypE313Nf2Y1UjZ6PkAiBdJ7icCAa3KRxOGB4Gyb/dHwzXb55bLCNQDEpjeV1/VwP+p198
d5/TLuFQCsjEmziYLW9tBce9x9x8giGPomAy3i0SbAP67TL34+IX8vas94P1htAXKUsYy19jrm59
adwM59M11coyjUxy3fKjs4Ulef5pFzY+7dqLy77sK/zNvSh1373/IL2lDJh30jZX9R7tga/EWXwh
Q/78Dg048HvJKqAQgs5r08/QquZSb70UMDdzTXmRjStkEa1zH78lyzirqCp5FsVqjwEAsaXVHnvo
kw6wM31NG0EON+u0cFvAQ7KDJMKdoU3Bg8aLBk8PdYh7eu47MTf2OcyPgrpwDsNa4WbaKxGC2O43
uROtU+zjRf+zP/aSB1m3Ajr/AefmsTcT41U4O2cqJcQOiGCx0WqvnW6e0zyb6pkGLObVEM4rSmk+
zjY2EoaOnSSvULnSL2QYqzahwRQoBnIKAeOFOJzJpcV5qUah9bpAMzhzz2Az2kI9rkre9aWNhg+2
AVKgZqn2ysHZViK2T+UOg2GxiOjGtJwjJe2cXb/Ok9MASzuyzUZVQHeOxyaDvqhqbvO7V6+TKWBU
oTzPws4MYgthQRgpWTF8UvRPzDqL/m1N8nEiNoIaduomF98EuRpGELvqLeN4lpmFKhlGUTp4Yj9N
Z685UOLgmZJkgSCDsRyyAluQZPpi8UOqcxKzGoUCt2zDHAOtdV56uneJSE0/xZ67BPtOQPcLq0gr
jDHsEEeSbdG7i3ZlzsbmTWVp/uRig6Zu0WxPQ1VLRfbnt+bp/EdpVPR9jBlGZh2k2II9u30GmnDp
pLwseWz1VgNzHblMr9YJ+WJwGuG+pmiP5ed08mwvFM4zB2Grrv+LUktwleb69bMB2w0tSdD5JsTZ
ZjCyd6CrHu7Vp1JdkLEqk7ZVQAsaROdkhigh4lEZThg2Z7Fp1BDxMEZejIi25pXMW7sN8BOtgdvp
v0UZF3mM49VPEkCpkvWPm/aN6ActAwlLYaiKcSK+Jj4X/WJc4hVq5QJwf0RyUfHGcla1YMqVm11c
+AV+jUxPAEU2DdSZxb8pDcEOLdMiFsZNRHeyPyUW3DvsqeTL6xz1zWqr3wl54TQnfFb1I8BBFO6x
DZZoEhwWJ8OatNydvXzx4WF2DmhgewvjbLXNw81WlOvcLhR0ShVDIJ59XXaSotBcIK+dnjPkpiHu
ZV0efgMXaoneY1piKlTK0+nG+UAMxtUZUJCNoTjTpDYSLzxie7Exp7mGSICGdT3Dra/8sX2UfblF
//x2hil29nM5ZEq6G9cNEZxgr/vueFva2IOVp+GnFwMMqwDoMiIXC4AjMqASUUqD6zN3m7mH1KBf
xYB+CnAuxb9+A5VDkO/vjro4CsWolpouPFYb5PmjsweEX8x5JnAYF715IFHFyI1ithdJIWqwY0xz
V8XB4H50qpeGroSvuVewnmjjniwNU3ZSXVyN+3WQ2icc1ojt9O0SvGouwyWptzeLzcRTiakCufNj
zHddO89uYTpu1NvIkbWaHNyCNINmQJ4pdZQfl5JtabjyaPUqVhDzDgGmVysHzirSakaA69cMv0H0
KheaPL3boPLoByw3U7i2IP8ypBecB7XWzmqzXrYZbtbDKZAyi1sz+WX8kKlnhyvY0eFVKgkTlPuB
0WqiqYwHylaWq4Epvf4pgejCP2oxCZ6B/7YIyM8CwHAfxjBAII7i2um2azSB9E2Y5EWlpi0CXssK
f39U99zsDeGVJiAAjHvqrVyCtH/ELXXDmsr6FGCOTWEsBF+SwNO14S7/W7K+00+QjdfY0XWvzW30
m108M47hjuTPiuzHSZNZAwrVVio3W8x/iKrIrjWtfj3TsNw0wPLA3mLrFw9y2ZWrB3IFN5KMbV0l
5hsn4sKp/X7xSuYCVgScOYcvve3uxHP8wwhC/3SN2YDT+DH876n60BUImdOomMsqqg5M7INupOIS
KnsXYHIJIYuOnNaclw0JYu3hHQJYE6KJvmb0cXRqlBESAmqj8cG5mP2pYkIHtKze6u3GCllvQQsD
LAgNV8UEay6ueH21VHMB39rlA9GNLjvo4Y2GNaSPDWqsX2Y9a6Damx9PBEc8tgDuGBpLcs93SybA
Y1K+skQ90Hxx3GQeHw88+AQjEWTgPSu/WPkcVqxeYaG8oHYrSBs3ndCf5sQ9t94SvhdekbvFRgCS
OnC+/09QutwNBtxjl1uTwL62It1dztrHm2oE2bfXr96rwKmYOiv1LkFB8bPxw06TCx2aC4C87LW1
dnaUViLql9MgSSf3LRi3ACFtplo69KoGDsyu0k2oYPhJHov+Gi457jBbUy6cpM2/5ykYoqhs+wI3
F0ApDmjwum16r5jFi7phKJKWrMKTT9dK8dBcK4i7U+K1I7nBk4tmFY1f+NaB6kUJsc1sn5wydh7f
uIQrqF2/W540sGntO5SJqdag1nedI2jxF+9LjG9nhUwyNkGKf8rDLYiyrrCVockiom7fEoG7m4df
ELJz5YXK8ldcDp9MAqpLmg1hRt7XZOp5nqoTJfmpWYW4GV6ixCg52jNLJgwjzXE2LIk04qTI3kEY
22s1z2i7IYeSAYc8/FtFRYmu35/tv+A9RA7ql2ReM/JJCeJK1Kp+Y461XeRUEmg+QYkb78P3jyKe
y5AVYSXRdcNVEfDOPci9MJ8hVPdddbEDbU6aVhIPV/HYlqJY5odstGv/uIBcpUghL8f2g010I+eP
BcEHXuvo7j6x5V1QPwUVAIf2kdNNneZUkJLvTzbB/gy1gqtQAlm83xwYurzydSDeJcD2knWiB2tR
zREkUb+ampXjaRQW8kzC+R2NVVbCVu5/duGGSmthZuMh8HTyD+pguaQaX/bnCB2y40swmIwPq5OC
nNFYikfArGFgfq/IqpGow8tfLweSZv0nbEIhLKUV0f2J7fDPD1ouOrAliAcE4K67Nq7fFoDS5Dts
R2i3asZL5cswLouawSe/CyB2X8SyIhTPduUAu/XwGMpZ8mSzHoA1iNFiusnxJvYQAxkI4OxGc/ci
AtmpQidY761feZZXvr4pCOWPzulPl8RSORL5zz8JbYMTl0tT8q2LcWUSB18A1IAm+DIeQGegtaSS
tme4/8dknHK7cwLTisogVQT9WrrOEHenECZFxi+vHoXcv+xykJvCBUP9JCQUjkoI3TPU/VLb18v2
u60z1uL8xgP/Rr0x+iBxM88Zx9zeV5fuGXFHgH4csWSI6dGEv1bzIR6EWxNIOLrMefL4D0dJaEX5
YESSujJFUTnxFr+6KUX562FKhiOICYpBd1W6yhzO5XFCmhOgYUQDYtvoH/A81KvWfNbxADzHbQz1
JMEA0NMT/1WLqXgYowo6x6qaa+dclXfBLz615OAYtlP5EG035jCqNPPGIEm/r0wRF7gY4OK0/M0Y
lNdHUPw9yJVRb5hmB6wu8lTHEQJl38GqwFLJbXaeYTS9cmlsKYgGWUgqRpvPJmDjxKFSae3TYCs3
yxIIDuP3byQBcarikxSKxpTE8URua5bWo4i05uX0UspAzP0IhWmV6AqQnO6yjgJJ1cmQvhhAbWE4
QbRy9KN62FAUcmwFzVHf7Axti7GL85c6DeVBZNHqij03/WvguhOkINPbGYp+kW2ilMJUdpFgVVZ8
Bw8AZEg3QHlU6S8MfIrYkGbdd4co12UiogSMLVKFp/SxkPkiaHcCRzFwHjaEP43gNuZ+vOCvmmZN
AZbi1J9RDDIa0f2ORhfBEzaycbmMF+chff8z+vsVm9tJd6QSMk6mhD3Byd4XvS6zAt73a0L5Qio2
rfSy2O83UjtVWYHPg+dUrfItAIksdVLARgA+eotBL1j1YUpzB8XrFQEQnW+AvjbpuCmqstPbuDPW
smch+WrKumMoaoQBUdQhd5WsdjleXLu95ESLzI4fqJZnZ+O8vZq1P/Q2PNoWndnS3a3/tCkYVKUb
L0JJcjqOP0oIXlGW8+0L/itvA7/zN/9FIhXbBjIwsA+3PL7/Nc17gsYHhTYYtAbpfAhmdYNsb9sV
YgKRH7M6YLCv2V9SJW98M6/hfgq77aU1SxK55WX6ei/ova9dHuWkh6DRtXnOrxAOT97i14WH0SuB
HBmD2cZha0mV3KAEk+bYX6URA4gaQ01h53L7Aicbo5RF9W6LmxeQDSmZRY+dGqERhxATj/niEeKB
lcYXwylNL75sycQLCFCFIylhtlUg62eikJqKaFiO934QLbOV3mYAH7Y7pB1gE667GAPIcLCFdyVO
4/aC451h6Ne4k5vyqPZh0YlnAJn+jCXA+z5ZwDlT6QYDiEIGm2naSy1NV2pjhFWdKzrH5MUQpYVR
HP3nd/SOd1zuJo2tY6HmblD7ZQCoLdjWDMMzk4EbKql5jBSbR0uxVG2k0zPJpTcY33ce03N05hmU
EV7UfL4xEj1K3rmNKtEJw/OvRwQ4/L0s4Nlqyc4OSXl9TLSnfAgQvE7BC0euysOrLL8wJm3EB/Wv
bl8alKWrfkEJ6VNfYtcob8FEw4bQwhaTMBhkOMQqhv1ctj+cOEG32Q67ACy2ARcHUkxrkbgtdtjK
c4x0CEvItz80lnJA/5piE2UmYfAaWrVUZafYDyXpXwmHG7Envg8N9mSUr58YLqq24/zxSmmr+VXx
NOYoI4bnHoI5iu/PIjZu5WEpmRHby0+FTVmvSCBGcaeR1XS13yMfWyWfMWF/k1UESPgyznlwSw7j
sj0pJ7w5AeAPliZCppYe7ObhBZr9tD0g30JYHUQhSSrsy8sqn/p/IoFaFBMwxo+sZg7JJKWrxHTe
+nM7blAygY4GCB9eUDMd8oSWQKOlSJUHoxNPktlHRiR2Q2oeAgmGbbhxkXCGlqdnPLoUZOX1972m
wXbBXYxB5QDbGnEuASZzITTiK+ylyf42owfY2OCqvi9ebhZhd3PWuJoYeznXx4M2tNU2u3Ry5Ruy
+It47OBjl+9F6T1xkGoSfgOJeOW/kb03yZpsL344DkfGvdRMGqjHTl8E3t8qUvuJJAc3TLAYqtng
a60cz8H5mdy/qfbwJ8cKjoTY3ToHQfedTgDR85MR1SRQAV8cgZCybl860UaqMmjg1I4XYlzaTIFC
3JLbi+CqV/3sUgbLsTcJ/LS9C2C7EXuGrQ3CWX2RIjPzjHHoKMn+GAnLCfBEEpolX7ICEZBEs1oC
YnMyfZTUgIExOnuisyyjYl27rlYTMGJ8OjlrVDjp6qVncqslm8ThjwwnA+ZwHqDVEQ61KLHBuTHq
7IxZQ666p1QQOw5m0zJh207Qp6rplBqK/J+0Z/sUvPzkhwBkfzVPW+oGq0MGhzIk7wBA3frnkg0E
GG1H5CzI+5uq2bhPj3VRj2C0IB4SMM/yxJZ/xADLozps32DrUXmJz8uNG3ZCjPFGjMczT5c3DVlm
hWwKCmBsUvXwyAx2NnmGjuOW/xIlEGwSX5u9ceWt+p42+wT6vNRCIM7A+FTgyj8pkXMMXFBmqWRU
pxXZGLB4OwYkAQEqbC+4kBDSvhi1xI2SZTJyCH3E9eG53a0Xfhyabm0+XSQ96gvRcZdrEJAmJcll
nk2wRaGlP3KRbhVC/QjciLnx3ST+jIz5u9+vYtXPn2x+ym3O6ZP/6L3xiYz4J3dB7NkWzUzg241j
6PxqPD2Ot538eoH+l6vu+TE0mgHDLwB8pl9UCcFJb1RlsodZcgFXKui0nbEw08hot2T3eEk7KyNP
aWlq6F16ab+/YpKQKcSjFmyCEVKMorL1odiOxZD33CH/gfwMWwtoZdWRNv5vZCLpgZ5L1RVlWVPf
iiAyEW+RLLuCX69R89d7TyetPqr/J1Pdwd31sJqRR4x8oPOO/ZYaICXbbdBoOIY6WYeHlMJw1pv0
PzuSfQIfZkSl90icD3hvyZzMj+GvDHSKV3hOC5LoBLvNs7x3ahbVo9E94MpFn+bUK61HPstARzXc
ErqvCCNZ5CBHKWnzVqhS2Z13PMMpP86XYp92kUb18Q4WwtLLQTd7PoyH8BqU797gpLtzb1Of+25L
EV/wFbZOtq6gBvD+mRH8aMGSkAAo7Q7+sscBOMJe1BBbdAqVZt1qGNffg+xWjMwTGobz1KO3x/cR
8J9Wgen3wVhLZMF3tFiYyDtvTlC7G8KdOYQ8/wNeQATR9CW+OHuhdI2sjZ41U6gAG66+XexB2abK
gfN6NQVmEKE5jVcqDjLsHBJ2n4KRgfUWw0ukAhs8nszfuSiKWNGk0HRbL1Rp26aG9OTod4r/u+SS
3rWmq4E8NqXZls21rfX9lpdtSJ2ttfI8iLyqwa8hZ1aoxluVhbhZVQoJ4lZi5PKrM+1ZcNqVQXKA
zS1DQCckHknAtWkUlRU/wWLl7VNn354NB/k+aPEkY9sHsZ13ZsvBQD0Hojd1IcThOkWjicm3bXzU
xvSXmFtI6fN+c9Eaun5GQcOYshdse/j6I9Ax4yjwClnkGoNVUdIOh9vTfTKgsPpOyWXCZDAp/jDd
u3vt8+h8ri9NnHwizHflk6umBY2FTKbYjCYfosmeRSJAFqj8ABmlhdlYbIpNtbFWDjhT/QdpC0MQ
nB7/6TLGnz/dOfpYqK+a9iqqmAJrNmjOSGL0+bakh6gOQ6aQZb0DFKDqo2zgB2SL5po8/JIptxuj
znHmt0zHnLt2UjUSEzcwBIOChtvsGrO3AL5RLXhyNWnzHG3Xw9LIkRfWTKjaG4KHRyVuhYwg7DPE
5wrMQYLaKL90jcMoF6D53FTlbMTf9mrCN9kPrhHL07j+O8btCUSq5OOVLR2doIdiZr8EBfnTY5lx
+fWE8sPdPSU9K1gI2qTHNdbFiNuIIFs4tOFAwGYXLmSpilXURRTCio9sXuzLnDpF3KD6QzOxk8kB
au7b4K85uJYi9mZKWiAaY10RegmImcHpSyN0KgQHPWSgN5vzDUaPogN2SOOj21gjLU1M94qBLqtu
aUJDsfU5t6YBf87Mtu++TGm0ysLLP+ohfIzT8UtgP8MMGgFqCjfMptFcgGHSl4tsWOXnOSjN8Z0z
r2dmeXmu9a1dzrXngB25rL+SpCLZEW0oli8DHddWsFdYC4TMUxhEAzQK/Vx2zxGeOxypEd8QeeyD
g1BfqR0vIIXdVoFLH7NlZAxEJoPmCf3uRkzZHhJCcv7qmT6fImSPKcyg9uxLxxOA32HanPcr8Ysy
r62uKPRRlihYktUojEVJqdBhOmIAaFafehooaxSd0oHo+NWBCNyNejRhv/F8qAdA9QlrSpDcyD9a
sWJcjItmrCGJBQ7ennrD67hksc99i+dAJY+EXKp+CQ7on36zOGPjV0osGHJqxr1zg04fIHG+fj5k
bTUuvgHRGdnY9uER8n0FlDl3j3iKDLSKpjuk1DEF5mhPvR5/Ls4tpEoDhyKneB2jr5Znq3FX4pey
QnfMst2TtvGZ9AYMcUFlfhq/nADNJds3vaGqY0TTdGFdaXfwXr47wYrsZHXzJ3KNHNKHXME55foD
zlurr1AxxrZXxgkHJt54ufgrHJ98UTxh8ABEVb1dj95f7FM8S+9MwTVHb7f4RZcgS5LdokP8wpqw
TmeP6jR93gBCJTIJJWxyxzHKvIyxkrBSQW0InGCw0kITB5LlPOglvvojIqnZnWIrRP2/wunZmvr6
w3driDjWki4nVbfoWcFh5HyogU1Xtt8uUqs5z1MKLUTtVGjYifLZTq4t6q94b1s4UvrqhtzP8m/2
pfEFpAMi/N0UrFPh3ifASEu1sGHF7eedlImLodmGLC44lTuuByys8fbooUuRYQdNGQrp1blsLhmK
Dcy7ZDLKvkyCT1hJbXyGt0PRU4m9QtU5oF4CXOm6rhfjS4fi2pjixqUXgFZStLQ0pvbMhuj70+2y
A5SSdJnaf/YHZWhwdfNQdPplZ0llM8941xGua3Jx7L2xtDpf+L4SnKh0rUTC+rwVz1vzMN/FCaJt
gi4Cf0qJdaKyZbcflP7Xu/kishFYTRh7bC0Beym7HRcVrupaLG6kwHS2Qai2PY3VhZNUTnG/+CES
JzqEdHKaLTy2Y2V/GWBEzA+Dmr72WYuVOdd991NXc7IWW8t0LFFxa5UvFt91Zy1G5trzF+xVFEvi
4gPM0aHy9rm4IZnD7WbGVK8kY/1lBPVMW09aeWmB1NmdSdb5Tl4QWW8oqJl0q+r3LawcC7yQHaQk
8fJub+t69EJwqG4SWGxbhjPU6kgksEGKsXf2BTdN3reI5P8DtXZGbpfrt7nYyLskCXHY+FXI7cdQ
RO0PHCKecre7MAN4sZvmzlqrv/BoaaIseH2EsWXs9ZZedyGmvd0FtvzbYhmno/gPGvkdwTjcXwBq
4P8JHzOe4LSHiondSxtDOtm+Rk1jmncZu5UAUhYde7YvesIzFhw0A5o50b97Ja1/6g2LRrslDYlR
19w0OoxigLw8pEehtXgrexKx1E2lFRJSxTZUSbcjHoHdyMtU0aEcv7Fjh5eWN/ZrKemhKp+1YUmf
pP00Ao2Ru6x7iWffFkrpZ0JLpPSrYia1cCVj40nTv+/SAwa/54V+q5ZIYPKo7d/UfKabk+0feYEO
k8KWeFf7vt4HHG9HbMAH1j6QjbkNZBP+I9T/FElc/xkcDCrbBGFg0lPw6cGAopPnwzQDVEmGlesc
NhyUhdQ0WE/WhqzTUOUBCLJQL/IRrsEik7gMlV8wL5V0tBFUX0QjpediEsPzZL5pHidp1WhZSjzw
sE4olbagqkLbmum8FRuNK8YTya1bAHtivyvDUBA5S5QQ04Pergq4XeogLe9KwkoVexxmwwGJW5Rb
YHYCdG4mMVgUPVS8uOt+BnAp+P3Z/IB/LCwLygNsHdRsw/WxY8J9Mhbz5Qphb/geanAcqmOvIEYL
fYjyy0ieJ11C1K+pkTIwJzRnsEiPbQLrL6cxMbVlT6o8KUwi2IVFU9qNXeGfxtTSVuCqT4bXS+bE
8r/yrHtQA8R7sWO3eWNosbyLeBRq6j5z7wjM4/LBAhSLFD4cA0GOAwNgVCX+ZyZUIgtHIji8inhW
IdPyZZoDWtta9alPoVJezcgYU5nnSmelG2CNwQ89Bu6kcYOY4+ZKnapK4OhZCO6OC+XtBo8rxTck
hIfKZERNmlp8yL+kxio+fBLYamLB62M/9WMSsEB2L/CcaDTMMRuspIZYb+X/wT0WoGbsSUqxLPQi
peSF2PcErw2FbDZHr1ZF6tLCEGq2f+ycEo+o+2NdjhzceLxu9unAKoe2q9rTvpeCv+XXeL3dVKcM
Qo0RhEUq5ZU5o89ELldVO3Uc8NeYSEUEjqwqBV32W9zOYmaCiJfKvkVaXAd6yDVCZQct4aqTHvmm
iPMHj24qA8banFF1gYMxjNF5c4sbeBKJyWbJndSRddcwtiC1vmUfPzEyplkN0rGsWxU9xQVrDHPz
uuKX1k1sU8/VqcSSLSFrikfuzhAHvs7Y+xbAZ5iShWRV9jJQxzI7a3gbXUDnzvukhaV/Oz7wsqZO
GWIKqm7xI8/ClFZMiez60Hy6sZeYjkZ48mcPbxWIjoxo14J3ttFOs96luW26Y3tM3v420ps7VanJ
ZzUmpz9hALvScQtJdd9tdVfibFuDelBmxI691iqytCpCJfWgtlpsdZnTBjJe6OM3ClghlQrI2LA/
wOAwB8F8LCKOHmwvXiR7e9+RB7ZuVg+y8rrSG848nNFYn6W0L7LMSAbGAQPrboEtnFkh5cbiqd4k
S4snm/siCtT4MXgyeIFxqSQ6O8vUKYedDc1VbO0x4R81N1352VBRzXnaWFn4tET6hxsN4lNfDbwh
2qTIfmVUxQQPr3S6s56XXF5qY9d86q7HqDHLzHnA5kN1H39bnufZnDRVkn1EebexrpbP19rfmeKM
kmGMeFNrBMkDKU5ruiAdmvMS407vtU9107BomDvKUDzgIfbs7K0fWXixxoo9pf1QZzpnp/zFdfAz
NnP5YdqaQxmompWQ+3b34cSTstj2c8GoJ3peJZWIHmRBQhoIk4xAZkAE1f0AVG6ppQjHOjXhkyoH
zBzKPjvGxjMPJpm7sgFwMRf0TCMIokuAS/RQAvyfW+AKo6V3PHvkb38CQpBUnQSPeJtg/GzzXwdI
jHtoZWiBeclEzxRn5Lqb8l0yh/YyXJ3U1Paf7MHQ3+JV3VLskxRL1+o95QsvzmnIbZO85XBIjT2C
N6Epd412+KSGCgc4RXTIw1avqKaOp+c9HryHdo1zdLLkq/WF1TV842z8eJjHWo2v9zd297NCj+Sv
6rzJSaT1hMmNkmN+
`protect end_protected
