`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
iZtBW5FvD+4JM9NWb7AAsPG7Ur2AvDEa0sOBEqmI71Nf2Y7aohqedIsWI05qANQTl34mU9yxk6OG
qlDX7gvq/w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fAmdTJMPvBnk/xvwLGeup9Pz9NRCvuaRALYwkwyUKNqqNgResqzFedzJNzHMaALl8WpbKyVD7taH
CckykZew3mfRZfULjbQnhTDzJ6MRQT3KKGC2NdHm3vX5gUHkm1QhKcdkj7nK8yivtYGb5SX+2g4P
slHL/+DD75Kx/dZfwe8=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
p+tDy6u8xSoeOP/KeRtmSf3d0Msz2jghPigcEDjvuu43VJeyik7toGsoBzepVpGvn1H3WJ0qL76r
8v4tdu2hTRdNLc30DYNw9g7w5rRbxzR/58n44bgTnuhIqzzyiddOyjcMoU9GyMJTfBADmHK+UCnu
2DKXXVsoTxafPdrYgV6Mh4c+QbQXlykSnXUcXfEuNd6jQ4xKGyzqopd7czZRR6j7R/3G3ORIxfQW
kTnTOzEDZzUIB1Wwe4mbc4i2CSpFvtUN62ghLfAc+UShCtsoNoAG+Pe6z/pCE85rj31J72v9EIru
czteqopuj5KFtRQM3PzS4f+GNC/mQUqkdYR5TQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHuu09X6tzd6vlhX3Z0CnNSScJxY4ZnX3CGeszc8a5/b+jLfuiOvdkSA0ytCc6AVDvovDRRkNtfb
3pvdA0H5deV0mTU7cQGoZSkWj5ueoBT79iS66vKORUmwhJpE5hfWMKYO4ozKcD2tKeM+47+osmyf
bd0BbWMvxTH+f0DpnOw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nk+A0ocFaLzK7gYnI2FIBIgo766hl0ULcw9dqEDZtS4WJkUjVhxzMCm2KHbX4u9jbpzn+G0lq1xW
fUtgSyVwAtCV6KzluqhaLJ67icijtByXeLC7uG7KTMC8FFpAMAYYmLI0mfiRIqcXMmFOuRyERJSY
x4xOews+Tf3N0blRovYNtUoG8+Of6eqSYyJoo+bp2kzbH4p3VBysMlpFqUHFDZH043wrXj4AJOZE
GOAJlz9WvC5umtMLoFbcWbJDXldQyjp7uMv3T1jNiUHfPi33Rb8ppbBgeMAxQRlePlKVfAiwV3M4
Jn2dtp/9kzdokK5bYkUOhY/MPlhUB46+NSfaMg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 50560)
`protect data_block
q0mAoNhrsgPelstEwcjfW2x2YMgyIsS9ms1RJTg37RXdM+8rejJtokv44pZrhHCv1/AoEWHca9nt
zeHBqImGnZLFXTafXrfLN94PfFvlo1hb6wIlBz1nnxm46SRhXisPCYSgXzL0XKDrje7LasOGokrx
jhDmfv8Fr1qh9mOCDRaUz09kr5BYibeFbxGAy/zXp2FUHqwwf6/oNKmswKNKTOiIVwnjSVRgIDRV
4RxlZVH8XzPR6Jdg1vlfX1qP2SvNvwxmOpbf1eNBjmA2+a05ku12J9dTEpxdyhUKq3zFA0T6/qst
EejrHhSTHheXtfyXHnnALYaDzsiAM6kLZyN69gI4Eybn6Oe263kW3sPDkIUzhM++lbOQX0pRQrDh
jsYPsisP2F5+72rr45D2tNqsoyrmu+UxxNeaXZyiR8dtuoSu3RX6bz1EdtNVhWpJFgJsY0h7ADpG
zZyNlEeV5SYuPF3fh3afrTWMDRt2sFo8p6p/hj3ZSAGYCwDHKgzO/uWSiotEB34Z+NRD/O0w1GCz
Dv/Oehu/Si7n9nrKgW+6Lyj1C13dUD+PfyaryrNkcNaOqPMvofzN3ESoDnuY9dDYB8OfP6cviqri
7mTc5mglhb9ktrgHZeCGgArhilxKb+IyOr5sknhkBFV0FW1dpdAqnmHxSJNBgrs9pGG7U55QbbyP
13dzoMq5Zcox7bKNADkXiznCix9OSTQtIuLQfJNfbpyZU/kiJXXlf98GN5jejCcGF9tNykBQsfyW
VSC22zRu7313DPj2Q8PgW4sHry/lsI1z8ufSmyFhcWFxPLb+DWHvYH70N5IGfXdScY6F1oJXKfKp
bMQVwIXB94zli//9LR+4kc4JkXLvqat3C5VGy6fDhHCUv6kg3y+TA3N1x9dtuzZJxiwmyCsS27Fh
Nio9bbQAXWZHXbC/nL4iQm6xlV6LzsYpvVlQEYtUYWDxdCUYr9xMclcbpZuw0ruq6/TNUYMy3PpH
vJni7RH1i3N/74WvDD6uZ88ZDYn7qA68Thr+wor3Om19Fzli2b0binJRcutsI5+dpSndRYpBQBAe
5DwcqJUJwiOknUkuj2v2DCqNl61yrDHJIhCsaxqUzORPq7BpKl/J4o1dLhAAV7NaQ1xe9wH7ddfV
iTp+qJjnXALGP9cQa/Qivfr3UleIsZLbrV4HIf6MSiV3mVAawd85SmTKpRPzhMj+kpknL9fE5aCJ
7hZqb8faa3EWGtlc2EsiRABjWHyXtQmDSbDljT/QDS1JYmmbTpV+vN2QQspNzVv4SmKMtX2IAGKl
tiLszMj3lQ8o56DT741M1EoJh0FhNrHK7GMwDID4/8saLnVDIwfxqRQEilFf41THUxqZFLteozQ/
NY4osrziU3tRdnegDU09m5oRg6KnPUTCHQsAsUMEW6JqbjOqRKHU7ZiDlJPrdYiHJiDjn+brp6MW
cIQvkVArLGBWeaClSDrSjtJhevia0HIz9U5c9dtRuuB3tbPXQ++zxduqr8yOsQ3ZK047aShrSXdu
FSfmv1c2QH3L4XGYCN1/9/KwzioQtW5M7cmzTGeuS2otv6wqB6eKgqZPfei6pApDko1VkRBru8kk
Qi6Nowva6KewAFsewl+Lt8uvEnojbPQ+++wQ1HMJ+8ToJCw+ps2A+qxUsQckt+y9bAw+q6LmCy5f
c2mkKrNrygM7ymcFG7ppPsZhoak80QbDRIwZvYvrfGUOMzIeck9y2lfmW9Tp9Kb/1EfwJM9S+jdp
NeEGkCVwmkVw6nml8MoTGKboYlyt2jvjdvf2M4pRNbAcPMGbLDHp3TALEHM1dGyZHCIvnRRUhM5d
hHFxfVTdSEwjHNK9fPRFNUBwpBbOTdKrr/8ltM5FrARABn9CMsSHNT5cZXwOgm6p+maV+VfpbAhk
qpMchMFEulp+B+D+WefQdEvBjv6zR3ZTtNMvR5pq+auN315+kFwCw0stdV2bJb9gtWAUGNpjifeM
LGYmAC6Crm7NQ2c0gIGTkFlWXkIK835pTaohIg/1Svjw58j3CvGovtcumhRRmCozqHR4w7ogu782
4j3v9WgSTslFjlMkPuC0Hm9q9mrPqQXkJ4zxJHpOv9MMFcQxAfvLHmpQva96LIOF60q2ITcGAhN7
uSmjJAFrBkIx33z5ClHm/fbbyoM5QZTOu8VMSbeGQeI8nbcJ/3pJmO6P3Ujpd0Ly6HMpUYvKbwAF
vT/+04IExUNjN11MAFJ7OdIab5y4rB+jfvsBKo2Z7Al9Kllp0PZE9d0kGSC0doPQx3fNB8+ukgWo
gLlkOAzxvmy6np0wCb4ajRivqyLwtu0hikQ7KiGVaXhuCpTWeIYuXxQaOkqZvu3azl+eLRkjPCc7
XH208LpsBNo13S9Uc3B7BxQM7TvQsoxA0D7yjJ0ZCOC4gyN+LmOTnzhtmd3K4qwsXh2sgvLiMKz+
8t8CLkkHZXkyxWmNb5YZC1GKKWn0WM19znslu7b8AoR0nGw9yddP6S8CSCjL3LsiNUibD+hvkg/p
PAKOwZ9s3W2tpg15ou8d9ews0AUpM4P9EbhPd0zvRt6MhQx0vGAO/wcO0d0CsxtybMEmx1FfR5EQ
mmGbkrGiyiQdKDLXiu5PorQWVKzfc+FSWcJdHbFMNIbDPIToiFGKY9iZsmzikWZk+runC0l9GKKY
H0X7s9iyj3FH7ZfR4ubjrCUnH1Ji9y3p2Pq/i+BYDGeF35B9QwjkRoRQ5IDTRXy9l1cUrHFV9G1p
z0wOtg0Tr66/KI6Ys3nzCKHRYy3DGwQ2lKTsdO+qZ0J0HKaXVN4GwgSjoVDYdThdSf9pmWtO4VYw
pFXMvuzA68m3kcNellnx+QIGrnzaqQFwLSkBkaGsdKuath+I78JaehZl1FKY/5gfqoWrY/G9OOOi
vgG/NJ3L4KDgwVcS3B1M9BIFacby14XGW+duwev+51hg/SQSnN/n3M4gFSGvybOj5qNlbrLVy/JA
62Jv2P7YOIQEY17s6hq7S9uWLumJro5aVI2gteeTCe7/N5P2gFRSuo7lblrRIJwBdr3rOCWTKmtS
dsCPHucqZkzkObNhNs1yjBD7Z46ye5cc44fh+8RYS/PHuQnF8jxj6Xh8LiAgKfmZTw+EX1RgSA5z
zpaKKEwEPU1Pf3ZlE2TyxO+L++ToptuBRgq6VB9CrBbUHH1wRx5d+Lc5yLmNpf7k70N+2SgxGEZN
5zFGg8cUteZeUN/1UVkPLVfmOUioi0vVMYNea46C/hHoxL0UGcWG8W7HcgA3Uy84HUNCjuEqRmBS
etoAw53dCfVs2rAjycNXjiPArvapO/3WiSdSXo1s3aFrFe1PhTObTqyzPiyrj/V/PNJrxYooC9EP
UVayLXUKekvg1ymVV9ZKbNlamQcACRheymMmVVLZ6JW9AVxATU+4/bcToS5DMmVYPUJ2Pzgzbc8a
YfL1xinlwdwtM0cMYCRFgVWAFKjw/XyxB3cTjZp1x+bjwDoV5GxYgg9BPKgQKcHLgru0gCb9kpsa
ONtmMnGdGAwfmvUGdSWzYncdQXIlXfvRETi6C0TzkqPjDB5hONHmuunsiGmAKzJ/5rWgVkMKnrG2
sKLhaYMTfjwQ74xByFbG99Dmhu6qlHUtE+ilGJMFsAgaXfx7iOV87qGASaE97iGU7xm1oGd0q0YR
1bkY4TQPg4XIX2+lmryq+L8H6S9xKeFCq7JdwlmFVWsCpIc9TLSWBR1NM//3fH+kvRW3aEjuxkSZ
TYcPF0aSuAfi4J8OhfZT5XRnoY6DqfcsqLFiHzDkBTdH1g+c6sdbE0nfsVxW3QozEYg687Lp3XLr
GdfWLoftChiKJSBlc1DmpVVkIRBuWSkdl6kJvcKc1vRE3CVruWf1DW2Q2Wnk6lEfu8HXxUHDFhWf
1tChHMlLSRyIW5g6UMRw+GPpVtvbaqbnVHH+wdGAHWHisnEs0FS5Ff7Mw+pJVzZcAzA+uR4fSOAT
gVXPa2bGLBPrXq4r78Fhfj3AdaWL69OYcQ1uLa+uUKOTGtr9qAlpIKMkQ6bnFiYoGn+sNgymcnU0
T4IideQ3e9O/nBW2mUsPh8DN6Ge1o6tw1YETZfM30+3hwu6RJeXAPpAD0mOOeLSo27gq36kovVPJ
RGuB5jNGTyuljXEJA+nP9tTjGROuSn+18cPND45VdjbMFYzXBA7d85bVCFJt2jhAS9CIndAcmlmW
I7B8o91SSl2mRQq41RMAcoISSPfNwNbkpymaFZMyuPr0g9RP37uSGUzNeQaXmWqe0hOWMv/2jTpx
RZjFO1vnZHEVQ90R0Vm22TjnWlPp3DXZUBSJ4B67FZbYWYquM6qcbMlTI4jfpmjiYRa4wGZAo6Eo
FKDaSly3GlwdV6Tz0jfk20Lx52OXqX5FzcGm5YeB5eXQc+aC0hs6DH4mZgQuoCIK3VluqUApJAYp
Di4Xf1ZfXospXmtKbq1tH7AIf1Ts0/9MkqM1MfhBGjQKopsGsr6Xk3/kLPnIbhLDFaXSH397n66d
k0Gl4hnLAglvArYAkGX/IixyY1k8KODrRlgffW232mw6ofkfwRwyiVPXtN0i9kLpAd11SR5lk0GJ
CjiDgyEDJYasPYpzNFsHyEcrynOHQYTgZbzgpA0pH6IFirSESmDn5c1qdgwUHAoSUeaOSAxxkaMg
KEzYI025xDPMEgr414QTEbELQtAYGLoXuNOPI0tabQWXyHWB8yuJodS6Dcvno+Fyp1zoem5ltAyM
t5xoT9mWdBRaK6arzn5VKW4AB5/nl+DMRq4Uzp+3Q6lh2M57IjwXFGqlZY/XYEmFLWBYqGwL3CD2
SJTlm3Csri2zwvMl849/l1mQwLx//anNMn+CYVkvLbUSrenfmVxb37zSrungvn9KW6yt5BHNqbZf
F7YF+Ec2c0sax1BBecp2gSQi1NU38vsnpsP/CktwWaoLRTNuJAuKiyEvp2MfiZA1fWTKPPEPYmC5
Lcxksc2HaUJ7LbNaiggT8iGKxd0dAiBhV8+gY12zhRdYzQI0biViuryi2xFzEUlLvUNcDFwyaSvF
OLiLT+qXkgdBoAN/Uro7BwoxRqK+HaC5hhR9Y7C8QP4Pz34LGspaWkOw+aXQheMU96j2eAYewOBQ
HD6afmIp+U1HFQ7I1070Z2GiXVZZexaM8VdsaMvtUYl0cox8irxHgvMTiRrrE9h11on7qeHZ3Ge9
HQpDuG1OncHkN1lIADTnBVbm6TTr4qk92ZpOBSNd4IuOQgvXfFW3y2v4lBl4VeUCwKBQY7KO7XJj
UmeBf1O0L2nWP2W0RTEyttteKCdwSwPbBSDjjXjrBL4OEcpf6T4pkWXnA/6rCLVx7WpY9pCJEiwf
TbvBXWDsvweVTJun8G0rGT3/II9r4OoEwKWRL20ImgrHEOGn9VyPnHnx1UK4IrCW8ALxp3bOUejr
KAS4R5jtc/iFaZcaAndEUFUsHCj5sjkVaOpE4bLs4mVPIGyWKGR6H3GlgZdFeYqdYlzOW9ASTPFp
RbQpekOqSdvVV0aLi7f24iGEjTPKLrLKlL0Ht2DNKlToe2RykhTj267rasZfKX51R1vbhgF3Vpx/
zqfzdeWvKLW39lFKfKB3MhbJssF5h2IX8bh3W67cvkJCJwt0PyJRf+/oELsRjBCzhfBwGI27+eJm
tkgSGSMeC6mXKsJJCQFKAcojxYQC1bHQOXVroeQKsYyFYU7O6vcJ/RK70IVo9z8bwNEF/6ECYYxt
iA6P9b5/WRvDniikS4dcvnLzvTIznvUZv3JmjHnCozOlH7NMJcT8isppB6s04fKkXJyWMMkIjeM7
zPgpjGpQixR+Cj57UIUrzn7jjbwo4FYsb3GwyDmYDyYbQsKwRBnuhQexA9Tk7s45xIIoizk4SnNC
QmvK7S+hJag+BG5FcflTN3C+frS8G1H1WP3OKkWF1QfBic3Le/HeGu51Rz3cynKolANrGv3UB36b
Cpy/oXDuoFkfuflFYMEav2Z1ei5jIiXICLhZsdqCj/LjrDst0j1RoLJhaLje+7glRTwYgfD/vCc+
2z95XpKGJ3BAyyu6fjU2JVsMR8d09q2YoZQoSwrwWv8Ki2+tozK+51ykzc5H/bsrxqSrbe/b8HH3
TTFuYqcuRz/Vr53+Pk0O5CeUnIni1ztmhprDmW77V4gxkJeAiWpuNo28Y8LYiqqw9wjoZlBtMh40
07uY4cpMrC9Sx6hFVlGrtQB34OezvGLwbLlrOebfyQpNuEKQty+XfQ/t3ABwmpGtvM8oIKGvL9po
4+ro86E+n02HDlI54tiRJ7Hpi+15yqZnaUOseCCY082dkfjXpR/kHtvh+ilY9uw/qEOphpBEpxZ6
S4OQ+xDZdgjl7r4kbz+n3/F7APzQLEM17NCQmJPuM3AkhI/3fKXm5PMfys6rOcCFRzTjTdRMEXnf
6RGuA4hTwr1qcQxJEnnB/5UZ6Uf8B9pe5dSHrYn6vpbd3Yl2kTywnlYpYYZOmITrYEdfFdeJhLCx
VPEbk+OJEVuW4YdIytJ/Ncala06NuWdPNMv8od+u1n+Poq/3U1Kevn43MGOytbuDHYw6f3w36cz0
hpClc1JvZXNZf12jV277VPI9JgxLYRlC7GB7R0+8JqjiqNestyWSmb4S5CAMMFFfsFgkXgn4wAWQ
EgEoZnuGRPnyjIDSCHFky5DrL830/KeCoHLv97qWp0qBAg2cpVzH5QR95JON5OC5y+M3xHwjp+9i
GEM/7FTuItG/x1kC9uh/9C6fFg1CXYFYDz1kcjRd8WYyMXF9pAd2Ugn4zLluBP21HXVX4K/HmJBo
0RwyvtAA7Pu8n7KDXINNcoy+sSAOdCRcRID5P7D9CKjcYd1WDCAzlXGvXvryLLHKGf7GjJTjAZdj
se+JrFSDi1PNAAgdhnV7jTuOG1CdtlOk5FEVoNx5IlQcputHgRPsGZp/JAkfk1NVdh8XvBb+/wCL
McZyc2BX+uX/YK2KxeM1wabXZybW1dBbbtFeiBzUe8Psg32UW1TF1XAEijgvqGNXGuXYWpVehUhz
TF5eSnrYItSO2yIfGFZItSIFkUdxbubU1tW4U7geQWLjxiT9iJF3XQm/il4cYAXmXSOwuWFNd4xh
1sIZUdlY/I7wf58MvL52LYAuJbRgEB3vJvWn19lyj3ei+8/cPchdp7TAePFJJ/NIZtDZutHNhkyU
hP77oaL43rcmrnViMNbmaH/7/x2qJQnsRNgzz7wPyOPXZYBgWC6zePnZhysqaV2DwuCxDEFeLGtu
YeCoxa8jIDy+Lzteb/wMTD3L+qUaolVJR388w2KyRn+gFylfECzqLA9ZUIcTvdSv/H8NQ5nMapkj
mtZyoRygN4pUhV2uhXDp/mmi6NBzWWpNhRW0bPzdz9F2guVXJYR09vcPMAHdoXBhYabdPsBHrdCr
XXNLP/viUmE8xqvszM3ZithVeTTnaV7wuKKhUfvCoY59R3ivCsPax+azqtZKPCdw1NlIvBJRzR2r
M8JyYJv9i9M0CDl6uvpFaM8BcZ4fU0zWRxhyExtwaef3Erfd1jiZR3GxXHgKoKc651szHooQjp/Y
fy0zIPqqzAifgGMWH+GyWh4UbkCOvsz96C4UuDEprld8Js+qTBSRgGKZ46KJega5LHdMWYacfX//
PhPP1R6ZTDBi2TKCeMaZ9kkXrch3nZBk3MuEweQB1GHLYNn1g0zoUkvnOjn2Q9IgcBfhrZ+FR/pU
OlGbVwHS34Y1nmZ1NYquP16eCTEjgON2L4d5slrPJPVM1S2NCbXAHuxPzmV9Czlz2ue7nk5eLrPw
YtU/sYfU/tlSsOtHPDs0HuiQw5a25NOYThMernYFkoqZImnTfm5JMT/EZ0AUMZu9e5AzQbtCAi1G
P5AKM/GHEsFxnxEgXndto5oe0Ww62auRhOE23nZdertdMdC1Pn47v0El82bXNekjkQ627Ecz6Mdl
MyP9+dZCzvjyX4PSfMT3S7qEL4YBy6RkIrV/H+ZF0p//iEWBm6MAVp8VShbUESrmWpTNOytMyBtj
FNJqRy9jIMHd3Fw5i595U+QeHEAxRRtfB7O3Pl4/e0d9si82dKA/kJBKNCztJp11FdQuGlYLaxlp
3/nHHYJ773wpO4vtbNKIlcPk/kZHvNCaIh4BOeqJveYMsgfkvkFtrXG07gtdlAggY+3lNoUL7Zkn
KD8YVqbsi6nPy9X3oW6FsjiOM8OHGGpfP6o7Ugqk6FszoHlCFUkP5CzPNPOHqyRc32Visutjw3eB
Ch+YxtAsu8eu7A1gyEZl2gQXeDeyskPXgfk1ecL1fm/Sv075Aeac7+wpjPGA3soOHfE3EJxkMUwG
1P6W5ahO1M2U+f+Ra60c3lp4gPx74jqhgi0Lk55yn6KXrsZurQsEHjo4eEe+0ajJzl6Idk1E63Jt
MfupD5CWya2wGn6lBsOp4p0w+ielAfX2a4KM79KzAE1hbMmQFqsfHxJRA27QUsm9pK5R64i8Oa7y
BoqgD9iF/zIMCaXvbpvhXdtFizaFuQKgbT0hjyqPJXKdp76qTS5bQBLaLeeVRKSSHK4ZOjVs2+SQ
XxnGNbLLu/FpYnY99n8Q4RFMkDDgCN1ryn+BnZFJFCwZ7E/W32a5Ocd4oPEEIBGFsNOvIaS9qQnt
90Skl2tfv/vTKPoSJ29tfa5q1SW+3j3+yIu56qRHaN8EePc2UQQWgMwWIZh+lDn83ruUK/LDesCL
rG5EqM6e4wQppR9bgCD6mR+zGRVNSAjLclkZn0RieKbW62HCTMRVLxIOl32VrE9TDiG3eJijjtVp
Iw4WvPFEqbTFzJ9JnhaD5qv4qYGa0+4QmNcS9TgCPmR1hYsrjwXh1jX+MXEM0aXmTXPsTREnDGPG
Emk4y03CmPDYFNNk0nzT3knq1lL3uABKg8dI2LkHSWohqS79X1hocOXPjMd306Sk9RuMfhhSQO6l
fYlsFN/TFwqmAtncseiH1kv4du14Na6vCon9wMKtK5XFaSSCPph59pUfRCm250bv4UhuKwV+M/3U
IIymUrAu96VT3zAPV295zjsHYaqw/+9GyqFSClyyqTeC7Yp12D6cQtcIYM2LUSS/JDSvzC6R/zC9
D4HAeAJBwqhlFHMM2oyWN4dqk+z/0TWPSZwdufPxjoMO6cMLqPJGXSU8+rV40vMGL99fk84yt9iC
NV6P01aSB/Pv825gmincKLDhFeC7vfAvPvevg5JvhW8xyERzHG0f5rqj4B7oiehkeINyM2LwAKeA
9xcDx+PEY82tDu+FvF2v2uT7C6GDFaQCvK7ePRyNJfOPRcKzDcBCHSKNgeU8QeweKsXgTRm+VQwC
d0M+nxT2iR7N/xEjECspkrP45C+m4gMbQ9I772RCBgIKb3+KzQb6Ke8eJsWTMEzImuMk7+475pPC
MoV1sQfFRAo33ed+CEaYqVV1yD8/kJAJzoQM3tydq25Q+IJVxOM3hbgi7dKeEXN8krBV4cG9RlTR
tR5DoA2H2NGLIafk+xMvU98V/p1bI4cGjObBjxArrVIttQgwukvaHY5lW6Daoyku+4rrRwe/1I7E
fB6VmK/6DzNvYFds79fZh1piKPx+LTtmgjd6+hFxv9KqHSP4wTHcQWAaSizeelPoAQ8giHbyDzfJ
Llik2Kpnu76delUf/UcItzlcFFhKOi4WNeIikdsbZMkq/5xdmIqCxe8hkDQQb6bjd/YJOPT+lhyn
FyVb1XE3d05hKRD7dROYGVHOWtjibV57cr2pHPd2D3U/4E5rmlVxhhqY8kK26LWmC2u++NSNLYB6
bAoXCb631UBiRaMzSZhFVsadDCiQ8JiBTLNrLQAwNtGukfMOSgX5IMdSrQ43LGtcaXQStm3HosH3
uZ6Gxa8eqe1+bicKT42f8nHgQBhfWVgnm1+ye/S8oqPxFZm+f2gRCwz1lvllv/5AZCJJL/LQlv0q
gk3dOQbX9Q1CLlR9+Jtc0rP2E0hlTC3meRbWA+nfG0rOxxkTMPb/9ko/ZQVW14JqXhkJtxamhdjb
7+sS8/6dRT6IAIcN+C2W7DmhB/1VZnppH4tQl0YVjarm1ctWjq4sYNjGXqu+Nb0tE0c/1Y3EpoTs
p/4ASna7KZD3B56neMlaXZ2VjfCm6Vp/W5bQ37ZEGVu9nr3MMCYVfQ/Wc9Xe5wJg9XjrAKcnrzqc
YJ8YTwCq7Go+8HlxKIZuvZcQsXDQskC5z57SKuQLGh7uqC+osdzPX/+qWf+SjVxi+JeDjtwP+dFq
kns1f8mfVJOsn8/7gW0jOdfKnRSKWZvdH7vtVtj8Gh8bMKqqIoodHrIjzoPxHGJBF+yS8RSFORqc
ltD6uMgDwBjc4+EKA0p16DYZ93F/D3mpv7w4sfjlvnrDdGow9TTit2Ddxsro4DnPNchehCL9PwGr
2MT/FfPPS6/m11rQAX46wrcpA4CAP1eB7BHICvigeGHxLNqGm5km5q94Vr4Z/p7WImfhtyR8kCDe
RW4spiJbMIhzgWcD8JZwpp1aPySsLN0Yyq5sUKe8Wi6FY9NOn6/rjguZosT7QjTHfU4VPPHZZFjb
ixF93ePvoQt/YrLk4znu9X6n/NtUxzVzBfOWblNIVjz0jJUj5YemqAPKzX4P1FlNOTxUN9coMxWZ
eMKhH6Gz1vKAmu++e1fBxCjXjR6DuZuFPFuz4XTjizo+fZDLdOatUZXObvShppmiNeDqZ2yv4Ns0
3Gan+7B+8cRmXyWUyM2KV4vHheiaiCiLBEH2mgl4MLoYQxFTPDqsmBPwQ0eeqWQh9H+8jnTvj9rd
HEAE1za1scaIhtxSEily50n2PaJWkD1xwzZko1+XxPnDxptpmF35eb9XUL4HaEY6HF/nCEABkOlV
pD0UsDLKzRgKLNCHoOYfST3opXfiWvZtahnNsL3WNwROvYt0kEq5M0kKxzNIcwWnsfuZzD9zdbTM
Lam6/diot5zkZMUTiXPZbVtQW60bSfAVIeSlDKDuACLAMkBhitnueRdrmhnv4KrC42dixTie/6ya
2KPEzXLlzgZp1kbPy6jaN0VM9Fvh/7VynFqmjWRPBmF67Qa4u26ximLG0ewMoIkcnBRTlwaPCtUZ
pSH8QZxhpFjjpirpOsRX1s0LZvjWQFJQfuweyCmwAiW1JIKpxKv2TGRP1rmup8bIBz3CHN/pEoQK
WqHfV5tCoExA0DXX4UbiWivVCngao1qgjn+qG/In24M22iaCVFHGwsg35qXDtNw0g+bnMnhJpKz3
/VubMBi+6ufXI6kgSdrs3aPn9N2Z6Ii73xOUGsR4Z8VMGGb2XfMnHia2uC09epdptBXsQ/w7noqn
Yv3pXzRjhStGCuI5l/EL4NKMc7MA2YIgDPsT4eP8k2OFGeoPzbXOSzagifS6wavEw2SOneXswgQU
yAk661hbjOlPasJi60db4fPoSGnpt3PksqTC6C5SuuQTIHuXr/FaRkccyVxBtBF175w0WtuS9f30
UIBTiUVOup6qJ0P9oUgMPcfhF74mMN7fGhTgkWt/JzT3I7xzwQyx2ASM3HCah58OMO46Bei1psW2
iy8b566so4nbwgNgSTI6387nutgKlLgkDvvGFVEXt1htwzK1sLiYvhApVBtQiVOAhAkjN1fQCSSq
6/VQxoYNma7gzSjH5zKwcS3xksVwX7X7iO+bt6PahIV+Ph8Evg8qfjl8y1izBTuBiSZi9ZUot2aW
7Id1aGMdvci2KMe7Hw26gMdzS/T6PrLkEhC70A+16b68JL7nDmAX50uGOiGxMw8FbGzu74nuTgmd
0COLqjPwSz/ZqEvpqgkOr2FSvrZBC4A9rp/HFSSkW/Fld5JgAIcRFZsSPVziJCBebIy50Q9pFt+b
7UOlk6PeFazSzEPeDBIAQoBRGTK3w6g9grYuh1Mm8dSK4+4M5G4ANPfALYsMHnVgeaIdINI/fhMh
5gZbNfuZZKXXdMa7iVquANVbMVwknt+UKrxr8/NZXp3DpkE1nEfyQFWUTrXWvoUcPzpgvA0LYWY0
pbSx2Jjypq9/swzH6okhwQEkLSZux+ByB2NCrIm+gfCB2hvXvFkFdU8ClOqW0uxwFyhU6NHUOX6f
hoiBzhd8HZP4Z2I2bjzW/CiNlColEjsqYkk5Y54xsI3oW+OUgRFb0ipKngvKqDcvRep5Mn1pMZ3m
IUvpxdfoxvcpyGbI6M+ogchdGyjPDTltY3C+R6EbEonhdzUw+P4psBgikW9QIovXXr04wz7mi3kD
fsZJkPbY/3acK0fELMSYrYR0JanL32Wl4SNphAVsZoWEvhTeuXSv2WYOycAOQaWCRbStsnXZIjVa
Hj0THzLJ547sF+r1VYK/Q1ooXA5uQ2y379Vts5SOF5qczm+aRdMIT7E9pCo89C/ijuJT4X/8KVt1
inAuR6Lo2ftVxxy1pFVbkZx0xpziGWN1gNs1CZ8y9SpGQVenGr14/+TzB953+lBB2SgQhGV/kTBC
S/OmdFnzS8hn85dn105xVVfdpbGHcJxSVdkbjiXX0abj1N6v9xQL+kYx0PXbv5UT7acYinkUsByp
wQ0Iy3PZO1gIl4Uno+6Vu01YJn+gq0BnPztwha6ZKdNKOhc09rb2WAvE0LK4UfSJZDOeWa8enr4y
q9uLvSGc3Y5JHxvAdRRmqoEEqJZiqY6nYJRvjkNT0D42YH4+5e7FOUNTn/Y9r6Z8zXeOzKSuhY+L
WwVOASa18zHpMRsrHiHqkBbuiAyyfsuC1C7BlTYGGdikgMUVEwFAM8h45hZn7VWuO3pRif6UJZNP
t72BN7LAEcx7vNWlDLjCKCvYTM0E4Q+buuuaeCvzXrxQuP02yrlu3IdFF3kkp0WF02spGvso7DrZ
2kdOj56RS0TRgdP1trsr4HtpNiy5YqELEHKid+XHIruZrrW6etZpxJJZaceGuxsu/DniY3bfHQE4
6rvYZ5469PP3JNDPPJC6i19CpSo4YBD1f2DRTj/CXGSXVOkIDXaaMfxv8DbxL8t58YuLLbSbmd5J
KZV3ctBukNTbYAVZHR80zhKIQzH+vbG796W/9v5+1lsuWq8So++9ei83379wrJ2XKwNEszbHR9BY
6t9Ck90A/nW0QR9xmbby5I6ZQYxlTvTkaHb4ommWuAjJoOrmzYqSrmN7YnDxpEx6T/qdUPvTMxLb
YXN+mvvHe4T9jwDVLKtmIN5w/60qBlQEz5m+OYSWFUdYWtUjogTuW6I8xuqWMNKuxt6YLzbydE+H
2spjRVG5qY0j/yGAuqMgSMq8QCSDgQ3z/DgggQSm8O+U91cJhRseMaFIEaR3uvK1oRNmkW/zddL7
h+id/8aJ1cod/1MRE8ZMHQx8OJJD+vP2kj4FOxUSy6GKmZ4vluIfJGTLScel0SXieyhtSKZstt5F
JAC8DAMDdCQDrP63+HF9me++8LXjRpKN0PYu2XAxArvwe7e9fSf4fYvUYJNVR4iGt8GQIn6l4+ib
5t0J2yhnrrS5tCAoa/sONM5NvOFWYawLZX0eFyf85AJNx1irRJiCQ3fIa+LnqDp8iBKkWbwylA6u
nU2ZoVtlqhdAZGJI1vwZ/7ypegxpw0+aSopEE0mYS7ta7gIfQbZDLcp95iCH7gmGMZp6+5q5c45I
nuHXly3XcCUoM/cLpGdy4R/yhgfnSCeEUaywAeD4kFvPPvO7+Sc7Wd1oBbB8RNtMqLk2vy+A5ktO
g3NIYHWkQ+bv7YjD7pFmwzX9WyakIP1CnrLrxoo7bjCtDZQkMQ9Uu/SucHXMJwqssTXB93ZRna2B
aC5IL9P/+Ghx2+wuyUNY661IoYk8ELNEyArp3B8Scbi3fKoLb+mCRCB227QMH9HIMv1Scd20zmq4
NWRvReG1KUe8xsw2mlsfp8SlgpkJpKz5SPuwJEHY6IC8JhU1CQbXjhdmkUA7QwJ/YGt3FSUkdzQP
2+Am+Z+5Q0nDWBxabQkFIlXc8k7qsVID+6nr/FcfsrKGiEH7I6iF11DygvFCgeDTJIU5BdlZ+ztn
LIf7YteNy/sgflpP0s8QSe2hj7oud4t2e84C0o4pIXTHPLOHbxA7lCokbnRX3H5FFRp+icmCoPvv
xH5tq4DSRBFCBvO9b0GN/BuD1lqtwmb3ZXBQqDvDzqRMuzup6HUJ3h4I5c/mZP09sELKliYxHbmG
QsLbhMF4REoyAr735ZUl+QqlrQLN4k/O6V7EzBTa8Y4zZuMi5eXyHmlWvm/3LBtgHPwY5zyLHC6W
ydvAc3Y7JW7cCPacp+RoibLDEahi1cgCidpcdkwh547ihUvH2Epz0BQJrEk1bbvchjeOf5aG2w74
BsXxo8wON41X19GPDKxxJT1jUhb7keBpqDS7pcttOfNl3/HhDeKJoTEY6BfvvfAnqNdUInZo4X9c
jLqQCmK8zQzdr3BvlgfGPl5LYqPVYS89pFqQg0PAtE4PkskBUD7VYHAh80AjeGoRVAI5PtIVdv7V
mjkRqUrYXWUawtuAL61ps0Vcm/+c3/gHii0bXip8LG6b5OuQWrLiwm/HgYeNUDWvmaXhDibee61/
GP9xxF9gpv6uUDwKzwyaQyhURRRK90FpoWetN+p46l8YtN9YzV+2PipOVcf5x4KNdL19G05H7TiP
/GFFAZFzmhVuFjl1/GaTTGIwRuSyNYvp+HoI5KvOGngAeJDXDjSeViSM8Dd+TfA56zWcqoBFDKzC
AzTQubfmkXDOPukL2Q+pwogUqhWPsK1RIp/pC06LYW3yxkSQd3xtoewz6GIbbtPwzPVVjNQx5ffS
RBz0ap3pvhXpBFosgj7gyakKf632kAIJ1OYxkczyARrFoeoMBg9DQm+4/IdDx9yoSG2skwmaw4Ad
l9Har4k4DFMoqUhjBiTH9n/XiSvObYX6J07YWFaEOh8XzNa/vGkTx+YhPQT8vbOCFg5S/ysJvhm2
RKtzDzEK6v+28v+dEtAVnu9/6lj71Mu2ExosIWXorqAzR04HECMq5WZTMfkWJlyfUjzrSvUmOg6S
Wwe6NUINmgqjoCC/9UbNw//BeMOKHka6Fox48f1o1F8fqZdkjrABFn/aLELwcp0tAToFKK5C1b+f
deltjFNUnINnFCIToBQDiBb7TFDiHC/mcuY64K044QxYGTEOr3WrwXsmF6ugXY8hSjLKiCBrttVv
mhfj0krxqVXD9oSRa0mqwUyBWkJk3HiaBFzsMsLcKaGZhBmeqE5PB2OA/A4e7fBA+0/doV1At4A5
WqaFsZyCCK3GZ1WmZviEAsN2+da4O0OuaKNYZuyUHBCHGTVr7mAgkvxRDQSBCdmtTtL05+Z6ACo3
/w5tYEXwMDakyyWyI89uqnOx9D9u+idI+41ss0Yy0xNhYFHELUJIc272rff4tHbsBiCVfwaS3cnM
r9jCiZETqewKfvlEZ2+otMyGDV+CElNGRn9Xs4yh9J4ZUUU3dfahA8PqjRwQkDOYrlK9Jp5rOUsW
qiL7NOdS2rmA7M8wNXfbhCR7BTFaU/Otei27VXk7QXF+QUTiDGi/mYZPSyrHkRVIXmJx2AnQEaF0
G2qU0SuP2eSaRWxuL4SfPHXFkb4mPJTk3al5f1bfmF+vz/ACIUedx17Xl0zXHMPBjW5e4dUmJQ5s
7rjYikEr+V1fnVyGt2RcYkNYJIoDexkkdaQ7KQmxYiyyuJkrHCydOIn1fPZokIJggJS9LETLjZw5
vwJoROIvArDOHgLuQMKo34m/DV/4/tddy5FO8m2jnbttI8JewpaazSxxDLW1TQcjvf56OY6ahYUp
ivHCkmviIsIbkg5QzkiG9br7FaI1Bk3f9zscob/4qwChaptYLq8yuk0o+REeb8pBbT5BkLF8JO25
jzBpWaAiYxR8YYgSe7mZgtbU/MgjFzgOT4+Z/6ICfwIH18VDKG03hx2nshLfKQsRUdxHIp2GfC3a
E5NacHHrRCitD3qV3bthPH/lij9mXMO7tqdSSvOLXQP8miVM3OGklGBQlBytHfICFWCHPXEmF8+a
WPUbs/fDt0fKAgiDiIlUwwxFfwQ3fmBGlz7Of/lUkbK4/6qlpgfwO/6uAvJ6aLyWK6xPigBxo6Gi
dxD+gf+QwMP7z8oLGVU1em7nJQtv4Wo3rUSg7wk30q1G5YDzMWz4l5KouByqgKUPs2tLDdTCv7sQ
Six16plBs3WdvPpU0qwhuHL5fvxt/gz9dUGLYLSkEzHtD0Y1lvHYkX58vUgk4zAbPczaqD5X5bqW
BZWEv6BV8n0cxkMH5dIx9iNSZ8WtsAlDgzC3TqpSnmtWcc5XqeFpAjCEVM4+fdBt44W/m3rds0Pv
VbpL9+a7m0/Hp2JwTQA29HNJFglfhPws2LqyzG+DbDkPrsDDG68bCrQtz7A4HluSCQBLDRuWEult
fg3bKsMmjsHWvC0CCucCq10KnF1TAUJhUBluuuyY2eR3hLt2a3Ddn9EQ9hT9DtqA83nhtpyEtgHP
MdHtdFC86BHzGElu6rGcd2HK4DqrPWQ7SEddpq6QJu8s0yLch6nHL5d0tCBOxTVeJ0xYWS7bjNR+
qLUkzstWGxmqvcu0omRwttVcKK4ovFxOURJWeMUxblYSXO93KA1ivCvyt3k9RqqNy43ihAe25jy5
rsFCjGLZGnBE49ek3qhIIVKr3nBIQO95VEXXXylC+LGD9EldeDsD3UQzAmA70f4m/0PHT55dLsR0
tvXvTHgAFhwmtwU63urOFU22qqysCeGiJNWb/CpJvBd6Jz4bid/GKU/9v3oxHg8HzpnZsRSFL8Kk
N2TLLDlreFNRGn0J6bQsr4ErqD/JGEd5A1ro6lSRCmQpSN9bWXqogQernj/MEUPiyPdGL09AJS/S
eThD119XdFek6BXv7TCV3m+bgDwUqqoXvB34fSP1BDDluLLuHeOj0/1QcweQDSyvteOJuGfmR5oq
hRQqW/GpKGU37h16P6NQ3/oA0TcSF88nbgoFCsBPwe3mD+z75FzNWIljz/Pax3KoOiVVlt1vm+iT
8eRb9ugCu8q5MW973SGgaxOL9qWyjN9uo47fU9GTgzS8xqKUHrUhqtGMwbc/iRjsVfbkhsedFwWB
EQRevD64eFFImy7o6KSyojK21mR1CrDn/AKyVXGp6Zsa7zR/bHH0FIWgTtTAzIoqfj8IT90RKatZ
6kyq1xL1LmhAdjd5+b9Vt8m5gFppTs194DnOEAXz6FgwYe9oENKcwmaSJO16VsCjMCSlwnf9+hwx
QzKWFfZ13s9GOjLeB13x/LYBRPbb8yaAeH5sJP8AxVC2lkroJ6IEZGWn3WHnDSnLKsdD5st9f4MF
6qTLNt9jJMzIavxANXdnZHv6KPEDheWy1Fu6IZ7rNNZMIkL/GoB3Q48QANDrBQGZp7qREkgSVwB2
AKiFJPtNHsxZNtn6es/73Im1ipOzR2lVkrgYKfwXhxfTcz8Crp10re3+rvCVOmiOgLuUNPhrgne2
apTyQUf/p1HfVKed1X363q56lMRNHlTyTP0aBFukUmwD3aR54ffaHNcfdILydZ+TSIRX2xYPx1OZ
kf9uqWQJcx1tZUBdhB8DBzjWqfJXP8WgvAyXRevAwssH74Ybpv2xlKl1RWkaD3jg1nieanljL/XU
zJtQEAr1KlbSjjWRL9cLMhIq4UwsKGqOgzWiIDlHj0V2pRTkzw032QClHTBPsC7D/VpUgWpLmcVX
Q/rJ1kRYeiVcepYLv5LKdMiiNtsRL2tKpfZBnztu9Sks1baCunsMR9/LmlJkpQMfQfTt06E9/2s6
eUXYcaNoLEB+h5H3c/nRW3baSbAfVXRy/9PMsTSXQgA3YitzA3M4Z+eFTrpWJoSgdAEwOLJpIii0
/x34XM7js7PwHTOydgDagD84WTGGTtCFI8kMv39gqX9pp+hmm+r+hZQm5+yJtyIi25V5Ehfv+vUM
+qGiRR/i2ZX7ptB9fuMIkR8S/bMI+aG+OOwjuO4OToBDAsMRYEB53qW30BD4ZFFwp+Lao5iZ4tr5
WZ42S4PrmVAdZGi9q11/fVUzn8LBZxwdb24f4DsUoOk7yBe4dxcBCcvluvp3cOlzkZ6P7CbjTMBe
BNiMQZygsDaI/QDozZQrbKQAMerXuF0xcxPPSPwCJ6/WFp2rIRicZ/kH0p4lcOVTlKNdO/wzeeKs
Z8eud0wM/qPnHrDYhdER6EDEXwjw1Z0+xplzbe/3Rjg9JCIJMpGaa4X/vY1lB6GU47mmKnOXk8nF
sEFk4enuDt+iNRq+pmPNiQmWK2s7kfIp5hc/+a9DIWD09wbHn4bazUjQ4Sq7Nnh+Q/SOKdTyu1yH
4Nxp6KJpBFNh24lHQQ4BoheJaVT0JjY3ibZnoY/9s1Zy49tRVHRWWQCgOehnwcqpsPIaQOggGl8s
SVOr6UmPdjftxqN9jUhOJOOsdiIqyYME6liomNiqg0kHDhbyruhrXBLFCdkNXBtqOsiRmNm4zAof
XS9UfQboFufM4pG9SqOx3+QCMGmcGEpOSdVAQcZIDuUO4RWLLz2yKu+MDR4c6Lsfwki0yjx75NWa
WCe+mGVn4vVx6XSdV34vjFvHqPM8MFaCr8rtm+QZWF98O/Iwbft6JiUwumlrtGJevL+lYhx7tnnN
sKGJ20NqPNT1N3awEHuU2wdVXa5yEC1ubehWW26j3uPPOAaEYwSAgq4vm5LA8oXQ2Z6093Xb8u4S
Po6M3Sr7HrwRA1/5lF/00ncHMVC2cKsEzM77qJZr9XSZf38F2/TFC9wMoOrzkHIJXfALUsrhR2gi
HGWOMaC/+DMxN63YpqJ3+2NRj/WTowRGVswGB0QvmtQSfclC97Snj+zGu7XmaEH19Dwp6AbEwHSd
07YQk8o7HL7gKrvm+DJFQwWsxZUgwuQjDHBqqxOvG9Wq1HukYlcY2Oycx5NlOXHFI7RhRZrBxdEi
SVuxyjNfNe7wlY0lK8NpK6h1FntrFpRmMuOEny1Grz1jq1KO9VGEIFnAPffvx6lukLpTh7lmzZNh
FDwo2tzhaECIkFikdI1EQSaW+TdzVy7gXJSB6pE3jyD4lbRNxHfaqNJCOBDn6KC5y5pISTuAcx6H
YxeX04t5qjnwzriD2dPL6iJowLQbo5Y++Y+FkVq7RD0bAzIB3L5oSgRXH4so8y7nbfruRd2qGnTq
UkSn5eTAHXYbxzKOlCWCF5t1TCkeilkhfNpLpQxwDlNfref1R+7BIY8pcRtorf4Q902EQbfqmP6q
v3+VRGQTCHXXt20kVjZe2nHP7/C/Pc82wk4UW5crUpbutyJCGQ02+6v/1biAXDRLUoGcuX6VRJE2
3I8M/Hq/mDJp5K6YxyTntHZZLsrJWfz5mL5p5niYZwAVZkSjGScihPUNreYXtP5tYcEd3i40+gR3
jgN6z5vKvFt+y+vVJWR8IC2SbiFBaLP0s3yztdaFmra7UcLciM1fjk1p12YPVLhdoTeepxjiROR4
eQlMAJyZtUyGWfbCKeX7CjKBeVGCRBwNpfEcVn1RYJsnV+7j6NzeC8rsix7pjHd95DfCXUmbSHCs
wf74dQSeAF3Qn6f7gvgnWGvf22Phtxq9pBEeEb+4R2renoDvyz7aCHkDz3j1sJx1QCLhM69VaWGV
a3wpm71M9hs7c8tkOPLcJvlJeZ7+xE5trtiLH4BdJlgU6A9ErSBNDg0Rs3vjDZ5bkS66eB3okH6L
STod4PJRk9Z2BkLCj74BrL8plT3A1EsAAE3r9C1L1QucOLVyOAiaX9h9LPdBBVkrH/Lnh7xg65HD
di3Ok6vC/BqMfCTBJ50w9T0B7JVwHF1nem91bxeXYa+J/nue0/PskvqNeqbJvu5Rw1gDGF2HLmHh
bMIlVjfKYtgXBCRdh7R1tVCvTlr8zHrFpzkuThPXYofHbJHk+CSvVHXO0dckQv6pmcj04NSNaFX1
lFIKXGpZgdsHkdKKdDoRlCmMaFAUk2rQNOp9XLpVGquXYws4bSJR5wRrv+YZldHRJrFpZWcJqjoJ
1VVDa6jLIPgKl9PKLequ5GK4n1Dyfgcbo3hI07LIeETQGsT+egVT+EMGCLFKg3tVw1ToEsGgfzx4
9tlfHQhjvjdDkqDDRVxJWYDoxHd4XSoCuOHU3m/TrNUCwzMfhDoNrpBmeteYCOVc55rLEUUZLGC+
z3PWvFh86xcgi35ZK6MyXfa9L7z8Yl94OdGF5PvqdZLQJD/L2kZnHC0tsq+gIXc2WmzvsiclG61F
QTihzyuoMvR2tjWZztgxXN62eWWtEDUwGnnTX6GPZhNPOvPrH29QRhZm64DXK/8dYLrQtDq8FVHF
j2Ec4rasVWueBIf+NfhQHywpJtHsbX6pBvjBt2u//uiNEDBVxBY0Lap1kltYNvBCy6ral6wl+bmQ
e9nUwlXLbxmICcjXiM9qEbJPkEuW97OkddaNmHkRD7rM/paV9jOLtGYEwVETQ6dC72cipZy2LQm3
vyzZYVrKBACSJz5QaIlAY5JpApYhMn9l9ljZJFnXb+SVPYpKH2cWQvxdEboyu8kgiyKuOw6ndNnt
5l3kWGXhey3JrYVxxgWCWcLe639b1Gt9L21Q45pSfeIRJHFG9NthsWbfZRTVauvg/Gz49OCLRc4R
jWebf65uab6yv1QZews1WgaBWKIFRPyNpV+gK3MrMdssKzPmxyzWpgk5rjMaFhyF5fDGWO5zVp1s
9DJG71cAepKOudboF+YWMnA3crpY8ExuyKmdPNn9jP6IBUQX7op/XE/0K3gROx5avELM54I9urbS
QSVVpfsu8uTNXfTUr8kS6Q3mZPElI6cvUJt2Cu+RojoOM5Kjzak+cr1SHCTr0M7eHfPSa87iF3ez
QHG/7W6DfC/V4JRJk+C9nCCQR64LYYFBZVlOf/CPN3m/IYxSx0UPiO46j6p3w4NtyMGoK779e1nq
PWhyTwOdqlihCXO+i5jeqUnPvex1MHqTDup3OLVe7EiL0kSQ5fzS7/PhaC+NF/TYG/y0QGYd0zEO
/jOH2CdKSmPbMg7U+akkP/uBaDrlQEZLN5zmiIs8hheDUgiOONYJeJ60GZXld8NQJM5noiTmUK/p
8qFAz90fFXEqlieJxlSP/PUqVqOt86fJkorNavdNRBxNLVY49wmSghYR/Elp6zLDkWmPzQZy9oKm
kjNW2fIXAtRJXuAlqjjgnEIsfnYzq/Sf2PADcS2xRyiPuI9bZ48Yq9bhsWY8pCKaFV821YmMEO8n
PKU4zhs14qhpZxYkmqgyoImVhS/vOTzLd8Pm/3ENWoDQjCrp2x5ioWwrzIEU/ToBv5JjZaA0KZZF
iAIr97IJ2LVyeLeitbfz9SOc4AvpKt7kidNU9qcuN3P15W0e/xrdeinZ+mhdk9+AE7+u9wNnrVtG
s7VXNRlcQMFdRI7iS6xKWOtcgYeM5BbOVDD3BI0X1Jkco5OY0b1B2z/BQ3iEQ3mJjSyxMleOKd43
pnM/8SVrz6TgZZI6280R+svFIiqaqS4asP6rnz1Zd93le3NmSX8m9I6SI4DAj6ZSFnK7WHEYlk2u
7EMsciwJMsjZOUYSIOdl+wr/sgXoWJZUptwxv9ww0XSNJ+j+C/vDQg0xSV1246HHPhnAeTmBKVjB
DmxehoE79UtH6rDUG04UypdqEp9ePE9XcmAQiP6Rx4YTPYTcTgOYsa/kAJoPjxtizI6mjYV3YVu3
4SqA8e5JIHOl+Nl2qN0VZUm2cPQ14bqeAqH/voIcvx5aUjrjt/VG28/GgBpFafNNBGbM0sMPERmy
rLHVTcVo4nOzyV3ahOaQcZdO+ings+kL7jddlVOppdENLEkXDYXhDkXKNOGyGrdH1GJvmXmChaJl
ZqLa1D/kuzPr9k00dmo2Ylt/MxQRub/BOiYXdc0IvmkGoYyjejognIyVi5xqoBkuRAcgORVfI1ZE
r1AvrLuJJED1a6BTTfFX5Fk2FNk5+Lw7deCdU/raHHZ9vN0fE9ugf+CRGKPPntlI9S8nsxrSRGl2
ztRA+2klKlxqUo7rWJ+0cT7bLIcD8ZEUDtaZ3J7uiiwlhc/PrQTdnKNyhjlObBv3TjfW6vZR4bqB
qzP9675HbmIypLhg9jAu4dxrEHcOAGbmW3c51qK2YGmJV1PAnm3IdSBsX+8jZDzbxGHEDD5XUFdr
i8RmfFPsQSwL4MBS8q4WCdPocmkBFmn1vyeMXJ+P06uGuX6KC3UR9glp7z3EwzmODqNfsj48ZS48
YRMOsIoepKRnMFvGxD+QNEy9jfdVhLlVLLPn0k8ltexMOeSGsKO7InE17/MvSm3Ag8x+Zpj2TbT7
nid3A+6TRzwQmdaSg1sXs3N5nOrVc27+FFUtA01OmPylQSbYmvLN2R7ihck44cvpGnjG9XAQ+qvl
r7spFntrw8gKXFochv7sMXMbgY1yUfDMAh8oE7c8O849RaYXJM2/xmNhVh34S26d6X/Uim3gVSus
EO3XBsDJkk2br6UK9uNGIuhpUtpBiAaPikSYxV7uT1xPkvyMmUy58otVufYC8DBRAQKs3TGI0Ng0
FfnRCQBfqSNoORkiD26gEfwcxZNnA/lUvAbKkUlITQOJJLqLi2NIzRLLR2aFDA7gE7XzoY/ShcQ4
IgNruAITBWC0DiDrkEd2YbWUN7ASu5CRpiZ5ZAOXSoPbukEq8muuJlIPh01gMmaR4sEjMGupCNI/
RALhpoep8kEUgTc1tt6+q2EaENA6wNzYFjGZJRPv7Kivx3af8URu1CB3yxZcFHgJjArTeHxEYUao
WXnsix42LJXRrJWC2DMJ5Fg5AtG+xdcQpRxOgZxvaITbc4l4FPDGiYWHwoZcoxyN82HSmQ4QUzZo
LaBabd1FtgrJiLI6XIKod6WCGPwcE4BRfLSFYIc/189HDkPhctjqUTN6lJY+hwfRgIqZ1ZfgX/Ib
NI5EqSSP/YZctlOgB/ZZ7OPdz6r5mVGEgwXiNjK+bVJo0YtEmkSwuTzWlB+Ka3ep2rri5E89E3WS
1844vTJ0gK3lqmQ4RXZl/vqlHwn54lYbAQTkK8SY18/N3gZ1ylTZgHWezyvMPYYlP3BQihPuvCsH
DQriNcSWVmHa/2179xChwIrSlyPU8Sa1JNr3uMaSn0Y20NwNDK1rQq43tfM3kZgEab5HJn7ljv3q
0Y7FPjq54POjT6J8u1IfAiyPcBeHU6iiJHJ/qV9bO2bBQGdGgq9T5Vm9mKRXh4HVNPCZ7h6mWZQ8
q5cQ3LcYs0pkkB1/1FxKeCSpp320icckzqhFvpFiueF0l0KY8mMDkdsnQC7y2TY+bKHW1CaimET5
MDr0nCaaClIxGSiWMXn172fwCCuZp/0JnHVMbsrM7uY9+7kw1LwW63d03hn+jRXzacbruYBXQF51
B6mE5zvtQcjdQ2Jlt873JrGM8wNov4/vNEVndf5nrZoah4oxJHPVK+7ALnUlpLSMQJdcW+ge7hSw
XNj9dQsnqp2d5uie77E6bSDJYFcR49/goAf0YB8qS6sK1gtverZ3Vki6IafVWmBYeG039LTsFFOO
ic3/sfx4HjCFf30CaxP/s0XarMiCcwepaIooTskHw0xeW1pAn+cFj4UT6BgOi4747skVX9CX7MM8
F7p9s5/nEpD2uPzgACY34vfwKepE2d1FZYmwJlYqN/NAPUtQ1E2am2Twik5bUF6cJGcPlXJZFMWs
Egt6KYj3ErygWhuJzasmJL5pdzMSUx+n7DBt9j9BM8L3L+XtrQ7Ezw+YyOMTkCnh+ScZ6X7TtpNZ
RZkI5+mxe23RpD+KTggic7EeB6vrPL9GReqTFxZTSjpcEemou2z0w0sg72kDuaci7J4n8oibPTpU
DEIcqOOmoAzcV45NpzDfZTiXey9dQEuVFlEjBZVj+t/+CAVujb+QV5k8HCM4aF8ZMh1BBWpKGYNq
k7nZUpn0fx5o2vt/zfaNueIZ45Hv7rGGVXHa1rltCGDcb5s9ZfK+zoLDD5O+NNq8M/KUp5MiIC8n
NS6o4Yvtfv8MdvWxzAAK85mxDhtgsV3SX3c9BPR+Plb99WtKME6Gi9oHo5kvk879gufqiybeqZUh
Nw540D4RRBqCil6iDldFBCkMFuYjFyViode30gULWRHOLYVl3iL9nINtuAqYQ/9XWJH7HBsTPMFD
tFT6T6EmvHlOxyWRuV4pAuUXDLEkdy7oMOanQs7ijWSIruVZYDSKsrtDqOk3XDMy6ErZLZrJlyck
3IZpbvizxDcDCZUVmYhNovJKZwP+rDegAdaVnnkXn226Opd2+0i+XJLMa0unQZII/1t67Huau/Ks
+TXT28r4sxnGzxbGPLncgJN7qYM85tDL1x06xWZK2r8ROG89XxpAwCPdQeH3d57PEnU4P1DpwN2k
XjP29PGK97a7h/sFREqxttgVxirwLDqTy9/hv8JhxH/b8Vl41kLblPQpCckjRWHgKjKY8TeTKVZX
TMnv7W8vxdHibN6rFubgNeO9ubXGuRlNb+JR25zLX9pZnKXZqD0cWN/+KVLc2OBjJ7A0mXqp9QTt
2pmTo/08YjMde0BsJpoaxyVBVj0Nn6/5j4rAteRq0LQiEw/xKleo4enTaHIYXwjCGgULdai4O/y5
85U0aDBoFA0J6dL136Q/YgQSJ6Rv6u1wiPk0RPzqWdJDMQAzPNXla7X/RwjazJ4vsVRba241OFR/
OSdaTTj2MehEWqAL5j4WgEPKQTKguq8ErXj4ppfw91u2WZMzK6zQ+mi8w7bKjEG1EXiE61YsFAOs
EdYY1ZTgsmhoNVIcDId8b16A5aNOhz966b+G5PvTsDe8iw1OvGKHowlPY5zFLc4pLCdqVWYNbDMK
dEmGD8ZKsvq15GciE/UIHRzbkUad5q2Nzz8RIEd3fm1k2VXWUEuB1Fl2qiDeFgzeyHYKiXJ4XjIJ
PqwCrhJ4cXWOrYUg964T4EhsArzbfgiGBEY1cv1yGOKef9xWszYCGRc1NOBEDoxsl8RbZjZXrR96
/TwTbRNSSQmr/Um3kSnTRhXdFutbf0S5f77ei0OPHZH302uzD4kT3G99QrUfV1EaXc7zeY8sAzo2
RY/RefZrDQNusU1oTJG1VL3V8yxbExTa1c7+2rFSGXB5uydeTdbBgSLlB57rTGjpkURWNgjXoXUz
7UDKrJSaZZYj7rv0R6gaTxo2D4lC3lAlAx4iOUTPwZoXDktBzhG3HdaDgiFUOwfETnNOZ5WyTnbD
7qI/dX8z3eA0Fr8cXXKrJ76KigUP5U3ly4FsH66xJARLAOpZ3GJATu7a3mUlWhDq0cmksT1iu1ZU
61ITTx/NOBM+8l5y7iUVMhfQHtTbnMpsqmetV8HkSB+LkhOtkhypEq4c2LtniWIMMKzwtfmnTlJP
dGK+NxeiKbzTNnyEGgFmX+42VfYkhGmGrxTxI4IxjElrPnpFqJoBvRdgj6G0jbamFCot5piNu9Io
pP0D7BOPWBHYf6Vjta5VDVNuV1iGTQgb1zc7YENIJjMRboE3t/dhc+Aazz5Oapk49qi+HtgCP+vp
pNIWyr/fIMLMWKzaji91rG4+4yrpwOjHZJpq7GMXtVZUm3atA3mcI9yJkC230DV7yhgcBlfdMzBb
/Hgaw9jldEeSdr2hs1EPa5wuYutyyA9ao4tK4bS2Hbng2ywIlg2rQZkQa4mIsdt0M8VUPrtJXqCR
wagcTtvSt1p2D7XqfXHdYg2ZrNjiSZ67RIddiEyqfVSXLcZe1NbCOv8Vn4hexZxJ0MFZ8z81qFMT
EoqO1cNh9aPNyN5TtU57wyux8/7JV5TEiFNhwI4lgV7pIlr5WYmAbw2h9RxZL8VIuj8PWV211nGK
g//xXRo53dQ+g0hS9p2XE/CUnXTyZWOddZu12mOcxxnzQIZSMub9/s65tieObE25XGK2QL53AOaw
eMlFtNg7PFeWv/DcGyIYrD9kiMq2uCBLOEJtFipZ3Bi4b5DLT53TfDFA9VIsFVEvn5GsALDrrtgr
A1c3lT5TLeXmK4eYrMab2gWPpfUGftLSKnTRgaB8m+5Ym572Dw2QvZOdsEGyV0f/KdbKcJmRb7X9
VCadOphhJdBH9lpaHv/80zGCt6/znFDygeXYvKAWSe5eD5BiX0dkiF6eSS0rrW97wXZl31jWkXru
Sudx7pPRpAWfgmqI8kCyFvXrM5vzXoeDGixUm9ifhdnHey/iQzPsV8faMGvUu22vTCUDuD7HG3zq
Dx3lhyIhzpH5apEwl31bwY+WYX4I0JCOx06e9QgvPkDDzpbvXgARbitPAybImvu8drup4YIW6s+J
/8v229qKyMeyyAM99PF1nmGOvgyXN5Qj6YjW1G0zDF8azgrgAjkfmEmWtoyrMx6tPQtbXOu+6Irj
A7PqOXMJ+Jwm51OnP51uT46JQ7HoQyCv0iTuA1/u2gw2992uKkLgyOaBMZZKNJTE9K4zWuMf2zdf
heY1cLJfuxYWK2YmLsds6OUq7chsYEfDHqzzOkxRImRESeIOqrmE9KkRGs+X8Cvon8kRP0W9WSwX
HZzi8zgOzn6ipRV1SNbVNnbGrcpFg8u4FHyIU2/aEe6E9Cdsmb1u2VmHlfONWLP3Q2+ErSeG6A9T
IMDKqGKd4O9K2AwvO3KJXcMw4iwjep+3sXeOgvPMOFXBeRGz3dHj3kOHCfuIXgkORfX8rNB/amvI
bpj5cKxaGntfHugzT5gFzEU5UqUTxFhDsZUGpiN/qBgI6rGPc9D9IPTId/F2BZ8jlV26E1n4fDYP
jQWsJaOWH4xDNCmDQgPS9NDir1GC/Y/5C4oRGSevU7d+eglGFMA1bWN/n1oFenio9yBc5nC9WmDj
BqszrAVvZC6HXGXUVza8BfTlnPB+FGj/xoWXHw5LmZmx8faPElIEYilj2EyvjNXK5oDxvGO8e5UP
zCaOi/R4enpQt65/ymNF3xdK/IBaGuU/TSnrwFe/OhW4NirWi+cwBJi/mWX0FhayA5wz084A4V3O
/HQm0hilgfuROTbN2AmGgMlyqZteidu2Tr/sc/fGDekOWV+VX8+lplOlSh6YvzMw2KzVPJoebogI
kDAWXznidR8vuZmU9UsQTaYiaVkl77CZ/ovF+D10z+5IPX+PJxtlXMZFM+HsN/GwY8a71axOxjCZ
k5cvuLO0D5XT11jecU4G3L9avtOf8jGa0rqJwaODQKuUTFsKCbnRgkYNy5/LwAXW/VcRuRHZNmE0
0kxUWgYX6YZ+OTXkmhyz41JWyFc/udmiJ6ldtye39YPxqpPvqQ+P76yVl6kEWl97QbJhJDmHPFGh
gtdDPv2A+n0RibvZKGUd2XL/rCWiMI3cYBGda6dfmGwjtBLHeR3KjQzw9B1JuxywdpIb9/cRvQjc
/7HQbsRsAKiEN5nS2B7a5OppFp5bL0tW2arFbIyA7qUxRHv3RoifavouQN5PSQujnEmwOrB1NDK0
C57W6oc+gDo5bX29zD+rbU9Y8CuKiqFelgQ4L1ZjqYLxTJA7/+6b4FbrXfIccp6JXeLvbJ92TMGg
s9G+ZLwWrpJ72i1k5GlQdwVJMQYKyHqAYFasvNwE5niHQQyaIqj0Hz3etPogQ3v6FgcCWovc1V5Q
d95vmCNpNs2FXFh5wqCt9mhEVH6sKF7cZrz8hgDYLl76OlYpL2gZFs4Dzm4nKlxLsVf4CDVplqsw
Yt13uixYy0RZ1SWoAOQV1f6JyoU+K4xEkyOfj7UK/N+8tPWhrCAgLOz4SHIaY/J5Itl+vOLffYxa
peocIgv53pzLUSjjZaQxQ1zC73mNxj7DizAW+zJxjF3RmJpt5aTVyNnd6PaJNVL/HmtTUMRgxrgX
MiRqnyh+sP1eJuuPaKU+Xk5bWL7wFSnIpIc99RnItvNY4tTozy9zGOCu/+PLwKPLbmqUrdEuyqrH
/N0TjNfKPxb+NO6tQuy+3rSnjeJIItBAjcNmvboxg7yJnrubc6hMTlXFMBEi4GLMRdb4W42U/7L+
HJD/vPPvVbt9iTwGMiZlWcdcUrfvRY5p8JP1BUG/Zyp/wqDIRns4fDVJPCqxTt+yFOTED1iqJTln
qlNcKk4zKweDak0vhkCw/KxDrKlmaE0eJ9ni9z0tYMlwUMN08zRQrhf4MMc/jrvQxgh0Au0vTlv7
1Jub88m9jWAKOu+M/qVd28YZFrtn7eWadKzTyaurqUWq2eRS8Homc/lndoe1P6w7wf6Kt6JIXBH7
L8JZ4C7WE1Z4FZowv/6nOFSadJaj/UD+CSYrmlopcmc8c0+gpMVryye3dhcc5DDZZZ3bIKk1isnv
wKbsDXpYV3m2TP8YEvXHu9RwxTjDUy1rWdrmbcKdHvhMyD2M2fDe3gk546QEtd8WNVscyGkT/GDO
FEvroDQsYaZj3N/8yKy6QXnpuHoCFo4vJ4HQwK6pO8lmCDcrlEbk+cs78SCMTa31tjBw120KK+Em
p0TEa9WnoKA5yUmiogHQRgR3uxWScOABvvxAV+xfOPTD+FQwVkiEhf1OHGUAeBD+HFQnrJNiALI4
huLw26GWUqr5JuSHte4vBHciq9DqmWx4rDL2OQIL3ReeTA3OFI4AuRDr4eGsnecclPpO4OhXmc6b
fqFvCmdAkAwkY/SHNNPfLUZ4klS1McAdVp9UKWrorx87V+daa+n9ab/EFBedzbzrCfw4I5F17eA9
UNAqXguBpSpAAphGKixHekD0JKCHfMIJOd7d4pgYkDOLPbnxcjEZerSl9SdMk6yIF12lebJYiIIV
Q8dRpcMJ2KCdevAf0JP7tpsRzp7YhhiKt5QWiiSflR4ijIt6EggCd7sKN20K2pb9HGpSz4Q5IuDh
ttfXkQzhomcr2DRSaXOtknI/Hi/NFZOUMgJxRp/nD4ptbz0pbsvVi7Vb5zHn/AJVhAYaiRTPhgCt
oeWHi4Fghy9K2pf7oeDVp2rPEJoc9k8VGWbc+JE6fzNq+viIicLJC1/vg5qziOeUVJpWfGnuvXW/
HLhPyC9/JDj5RpTEGXaAU86UDVwQK064P0EUhi6Az1G4Fmrtme9y0EHD6+/3AfQaVApxEQc0Soxx
Sca4xpies290c03PxyeTejs5zmYlQTXzQFSPrjJKizRzOYAw2sVQtKfHCVMBeNSkXjdDPCQxtoqj
iRC505kocIfXWQvL0mX2Strj7MjtZWduCCLO4ZCdPZ8T/FUHqt1EmNKxhgPurm0DQUvRWV9rGmKu
RkTMkHPw5sioK4i2SfQHMCiXV3VLMY+cgrGPP9/7fl+JZm3aGLLkkOOnaaxQ1T9heov5bgbPB0UE
lzs2FGdRvMLKa255ZN1pOQba1WKl4vAYyFk3+aZ1d6nyVgdr2XELC8JfjjiZLF9s4r1dxz/qlOhr
eRr9th/eOjQycBwS9yoBiH9AseViGtEAogbxLUpEBssr+JpA6EBFv4bn7YGFdtHFBhmHJ/npAcoI
6EdqpAdPu5ySJ+8pF0ylj6zFWSuUgWIpvbwDKzLnNWQKduhhOTGnhb3DB1V1qFez0zI5CP6rr1WZ
bRmzANKnmT7+XeJ6yGJPGIRCQpLoPqHLD8TRzn43Mp6wrmA0Oj/VaTQWBBdZqx14MyQQErlhFIHt
o9I4DrVPEggzpnZJPPD8SuBkP593wGs5bvEAdEz/I5znBb3ivp5Cjyubiie9X4BrH9FtKNahsJsq
5wr2OiU4mvHO2hpegCx9oi9K43pvV/4UDO8N6UCcDi8TVyr9PEPh0DB7l5f3ItJ5p2E7eA6Adyyt
b+p4vSdzdtyNJVnfIsUmithywIuDV56g71iFlzKrkEs8CWIKZK6hkunrQVqsw75ufLIxdddB8Eg8
69K3C2GkKfv9/apVKiCMO9gXRkQL3OhdWSm07aH9F96MB3+UNEJ8LiQhE8feKZXHydh6Csgz2JAC
uu+TaGSxsYizC9NkF+bOP+bmvwSvA5Zifs2rWDaXOK1Gow7OdnLtYw1LuRBF6J3aGa95tigodc1y
Vap2w7sSEuzO3/efai0PdC2qBTyQJwYGZsCVm1TyeB/GSgl0RTmeGBQvXgnAALsEumc7x1zeJk+h
GzyBpdyYKDgDTUg1eKKxinDNno9wmYZ/AOX8HKEoELDS9pXBqMRSikvitaPqaecG3XXMMwzOXbXm
PuBwbHmYczuUDt81zjdvggN228PuGhzMQZ4ULszSeUbz5/3wCsUloKmrQHFfKcjaWz5gIwtxJy2H
L2QDqfGOI5ZdHhwXoK3wEeglcjqCdGpjmpCClJmIWpP2l2B4G0t4WxdFrFkDozmRzTFBIJZrt7N6
DFb7ouG2XMX8seMIU+aPwRVc/8r823/R7XoYR8CAq8HxePJzFRllImE0+ub/pujOTddJurhx0ePb
G64kMeGnbSXwVNsxGr2x841npR8LygXIrTEDZxAQwvITal2W37/zVnQjrwmv73QCG1HGwflclZYe
aI4eicJYkBphkfE4tuKHJ5kRUFa5MdsyXJCDzEzVHQDtWx+X/09gurZcRXXCMZjgGvdFM4JpQBpT
Y3EfOFYeWbii27ldknnwRsW8UpPKyXZitJGyqOZbqds+gY70mfmN6CqzTS7Uzmdlns0YfjtfHITi
b9XVJTzOV64mVnIg5O/Hqmh4JvuF8nY431eq0SoL92fbbQH2rQdl+BF4FGoCshKTMhvNpLc06HsI
oa9xTwUfjOMy3GiJPZ2FGtqFdma/lk0JlLOK5M3xX+KynTCoHmRbdGHiKGdrQgR1Enj66GXVIMsR
WN5Kof2VbWos+c4MGHDLCzFXyha97ZYC6gQlHhRb6f2UOXujS1ff36ri/qH1cc+eU2NXGShje2d9
c9YenfRVqgpgyc+zVr/B1JtOvH6RjtRyRxCaejbatHvXXFpkYasKomgZGO6bKJPiVqbgZ2nhWcEd
9W+gzZl8UoN9C+2ibDTmYjIe47tlkgIf7vFQlJWldbNYh4zeceNlWZQW0NgYRLaogewGnBisN+No
FaweFprZXCKvsN5rLmsBURi7JyFP4ul16/DqGdLQ/7U9THGINuBvuP3LCxeJdyuJHfO55+rgODAR
wDL7CTGAukvc8LHYB/phn2HMmpP2aF7wmNT9sKrkcBXK36Y2Y4WJOdLPAbAuj2dKEMoHr8pK6fHh
+2grqfkA2r5b4OiTSkwsOPfHM5AuoLBzcPPFJSay/P3a8tB18sT1FNDNgCyqGM+Wpa2ZyEsd6QG+
QlZ4gQj730eTEj2XWJEKvtHXdgUOpuZqsL+kOu/D8WM1UKksodFTFStAOKXZYNl7uUtQHJqDLB2H
M7I+5NgdFDuZmFcpJREjQgQENO7VbluD7F9ZvF+rcJHjG5nogXyCE2g2nvsMZ1dJavZGTcs/wQtU
UD/L2BqfaKlNaDaVTpJD/FGDc0wNzjJNW3Ar3v7n9tmm2VyFtMgFl+IS53acBd5njZZG71EiNT4z
HhmJ4RFlXaXhbMrSw7XKRId90ITcj5O4crf34y8u+ChjM8eRqLMo2wDGV0wEpsMt2YaAWyF9wAi6
+GHIaT+1AeLfW01xBuAM9b6RUc0AC75vlGtn08GzNbc7jg/i43y7phS2YtLWp9OEeVrHeZUPaSsF
NOHcJTF1gdKqwnSNO6yneWwzALtAPM9LGxxaTnR3idrmV8/bIOnjGTczyqPVSrOp73MM6UHnHrrj
OJSlcIhAOssw7+30MSgLYZXkkHd6yfOJ2JXRr6AWYzsogLudMIpSmTjiJB5laxanBa/uLab3ogoR
rymkq/OgY09GpvjSqXvd7ciWHx5JvysIq8tgUXIOCuLPCufxc8pf+IFKaN1FVaeY3I27Y9Cvg1r4
jCDhXU1G4PYXQWl4lpZN9t2ZERUMDRFZqllTjs/C8eV+YbsydIQAo4IDy8j93sExeuMF6wLPWVqm
FpwpNQQT7AzWSwPeScx3+C/dczrVkpyX314Hg1u6wxb8qeD2/Gfv3eKyozByK+4AX26a+SEbzWYr
4SmJKaCNkiGe2YF6CoQyUN2u/VUUzdY0NybPPwWgxlrrDlAvc6t9FuWA2RPCwJ7XL74qnsX9Zud3
3kzlJn9iF25YW2C/HW0cdFHZgj7CQ6MTEweX1QxxVVVTVhZdUaEi0slw9aeseyDYmujj0x6JcS/J
nuv7Ge7oPmmq4BX3P8G3iBCJ6wPx3a5FZz09y8ugAg9qfWy7/61DOyWtWv/0hhpyH3sTFTiyw2Ij
VQfnwIauVP6dlzPLUjA7prHAat4P6iCTpySvwfGOUzAGfCt8EDZXTfEk1CMU7BJdMlJ+Ky6CJvVt
2b3APR5DM9doEAZ4f7QmGtwVVpcst938SJRZy3NK4JHShDWCRtfVGtmhnKUSZTtaZwiW+YmaXrO4
PszFY9AH1AaJSRu1v7B0icb0eg6yAW/btT6PYaiy4d/jgYA3kWGAjVTfce0NsA19fMTMsdst74qE
Rk2SCstc3Ph515ECfZLHHrgApEdheuNZsFywuXF9mYl3G/rd0wLsUOqygptQB31mF4BaZjl6oFta
yRaG2ORs57+KGdXOzNws8Lh/0Fc7FG0MSfamBpXMXQlB7dOTeCLq2IAsjgtriYz+4Jw1asOfwapL
SdWUSkjLYY7K8w7uB0qO8cL2pDITJAC0bUl4Em0RIfTfY9igOoBhOVAwaL+0f+YG2uuQ9jTG0ptf
OEzG77ZTg4ghaGY6i5GcUE+gCIUR1z+wJaqxUMe3l3MbGhn70kmYSLYkk73adt8gXE5bI7RNObG5
1dVm5iKrkoeGY6tmcer58lQYxoPsiLxU2LQLa5nvK5OWmXldZNaPrYGubkHefKb6cx/6WBjAKdeB
A4/KQLKgHUG9xwWZdUmkURISOIGXk0bumzGw9zBaDHC+GifoZuhNS9C0DKo4NlRyzbGv9AsBEc9E
43yibU56alEpi7IV9gbkeSFvkphY+cQ7/2u72BSvcodN3YRbYBdlHqLA0lJv37W0fJm/ZATieyDE
QKdzJwgiLCY4CY1kh3D3NPNMpqQg2pn0s0zT5VExU08k+Kc5eGN9MufzWV5XI1ZqGSiBJ4/OlMa3
tr525UveksP37LhKDOb0IJLsYd4fmJukDQV9CchQFyP787XDxuF8hwkC5dbVBaFT2JzG/9BSNVtP
wExuEr7JTsF4hmi47j8m4XLg/ZrEfxxQzThHPVUqdzCkijKSlUVIaBaAiF6oQnpSlXSZYzk5HUdg
Dnv3FIEwxZhX/hWCKwYN/IMA1hNFWWUXa/A03DOJutiCg5zCdVWmxCr1rINgARN5t9E2oPOFLDUW
fLx4zHzHPfacgIic3f/2yh0XEtx3u8+rXfJIAGbpLK80zT2W4pjv8G79eTg846qwuLSy/W28sUWQ
Fn/WgzG2ld+t8cMO5A5r2Un0plGWszk2Yalfm6Wr1c39vKiUkR6xuMQYFgVU9uVN2rx763ZqMRqN
NwCGdsFE3fANZ9ulL72JsbsCswvr9SYZHjuEMHAFwNHqPFYfMNIKj1xpzr+g9jd3bmBTGKAVR+Jp
02Mza4AC9cySMSQQbfX6FVJPq5z4ChQaHeNwlSLrQ6G6FDZh2xVduuTymKpzHl6gXADSUsCdMrg7
OXy2uMGabagQoSe13bW71JniMGM1ncB6CzKWjHkwmeEKRsfZEv+rY8iCWJ4md64bee1crgJCJMrm
hUEhYuvF3HkWgd52n69SdGU12quhbs5JTq1itWMhb40LYqIYfyO0WvIZnIHSjN7tNsVBkxOhYhjw
o1d8WddIwU+CyHM0tm4pvyKaFIkr2OIK21c/VI6bL3c1kMPT+UJ1PsUUWVU1KT0IV2sEu2qtrNNf
xtble2voPvK9svIXOF8oon0GaNiXRWvxF8otTHz7adUqtvfBOIcl5F28RQkaD0Zm4kSfPMuVAEm7
dbRTLyco+JANSqgqWnGrVZGLTV3hU2kKzqj7C7cy2CWdwFzY2h45K0KK62lkN0WdrTAYvxhnTiB1
0xSmuVxFxaGYiZpFxk7LJ8+hMwsL2+78VuV9qyl8b+mNjIGjmYZEgDnw7C6F4+HCxMLNSqKONb3P
MKhGOTVK5aFxe6JwzVMSIgZFiojIhUsxhaNBK4MeIwwdfcGVHEpFvSrIvacPuPweIGSTbUeeA4Ve
C2/8H2MibgvePaGm8IKc8R8pYiakIlmQce0TC3LAladsBxhWpboV/Oisp3NBKntC98lT0dQxxn7H
/jvP9ffzxqHTEyQ/YDgPS0ROXx6AVtFkxIboOEICD9XjtuJzQlOEM1jcb2EFkLW0MLKIilkFdNMW
n5cuIxrX2JDIL9EmWarhTw4n7WOJx4z+FFzZi+xC/g9VE3qEZmgJD0cmcEETQRDR7XZ3fwHG9ksk
MtgXrKIEtcUunporNNPrN6/4/WM+r4T50Z26mTL06Tv8UGGuRo5bxWhsVPHq4o36NuxTx2kSy1OH
mhqlCngC6x7gO1QVXpYn2LdBROVX5yir5bEA/pPsqnn0IrJiNYpXmgR5bzP5XKTmlY8s/1ED4b93
j19YwM99QPTKCo1cSsfXjj46RVgSeRanKQElv7mbt02MF1bkY/ORfoV1Tm+aYh7xORsg8Gnk2XJp
2zyD+GJrE+NrHqwlS+WZyzZpKTwC5JjGAxsO4drw0tSyME0uu3tSJgYURWRY/YgQ74fsal5w4616
eSPwgJqPy18MbMm0pQxRt7/v8ogfAgbTxcmeNj6g8k9pqvwANWLvY/2VPiUw03kl6rYXLKun488+
IAn0x8LO2ebNxmndLVA19U72y2o/LOnLm5HyqC3V7eNg2TGUEgn0HWIO8XvkmrmUNyOucH1wfCdo
DBRGewJ4ZMBW84tgj2N4P9p99JSKHKLRtpKOWwuhBk7MnjIZeE6YfBZ/KRh2Ks8hdSQZ88vX5Nhm
ZD4x810JnibbSFoBoNoJHXh5yx9mQn62al958ORBcitAbdJTEuHOjp0bcwbQlNA5vK4YF5nvXROd
lCRqXJF37s7j32StxL4vRDXar+0qs697cyjsYC1cGMzo1mX0hAGPsknUXDjd1MVdOeETeM3gWQ3z
YTJDO6zDSCTosxW1NX57vmd6Kw4bAXFtZNWlyCkA0AjzGJBYkxDaUmJszspsLADY08TcwBZwuCZ8
OsH//h5pecuuA4OyLZIc/FStR/tWUaL4RRm8pPT5XEWkaDEGYl9ICnPshbq/1WkU9ykGm2TQ4aUx
cVV3JWCaVR/3oW1ERrcRjl40lRgTIGHKRwu+Ip8LZC46ZB8UBdpO6Nsfqoh/ARdDTiUdymvRb/wn
B27vgbnKh3F/p10cDv4cGKLtl9xq5dCZGKfeU5tGP9NApvXmU+P7Ur4DyAt0C95ZiYVYr5xdHplo
74MCxpFOcdIZb4hQsRrc/cwrpPDC/js5UXNn1DUmH9m5b+Shunoucr/E2qu7eNdwTh8T8JBOees/
nJw5B1gJaDd0bZ7C/g7+Tld4NJgLiWjKrsqj4A8vi5PMI4sKr4TV78JjbT8T+Gi4Y42BUVKcuVli
6ActfshF0kxPpCnx0S3uj6YqdK7bG3QR4pffFA5MxbgzAXJdorNLttAQidwGvCBnyvHUIZ4Dd52Y
WpePSm5achWk2waLaEYIZi/5+Hm9jbdfuEuKxrxWapR8+YINO5NYDH7hsy6vZYwxFdxrluSleG/y
oRQdolmiZKs79E8dFZDeKJ/cbwHkKm0AJlOfUhnSKZVmNNYZt6EakXnX+QH8GsFB3v9hi5mRqbvu
xg55nY1GLmpIKJyI0A2EqJRDgKJc/09O55cY+8rqsehee/0k6vw2kuQ2wNEFdvyXb2VuHxmAQC43
uo6gzBS+k2i7a2C5M1Gzq+xMkqskMftGhDvOYBNw4+dncpz2PK+A18CQr2xJd1pT0/TP5vv2nmmZ
BRQe6J2SA8DBTjWVABbxbi/qdBR/jWSxWxsO8yy+6LkJuhQU4osPJUtAfH/dxfBDAq+0ZFM6ORxr
Hl5rlOR/h729ABDtPgVWVWyw9ysRNQEhOBf71vrXxNVlFecahD+/SJdXe5Eu8PM2v58uQJ52eRvL
84CIrH2OQjPTdP7w8Z6gZYM2oXPqPBqkND6AFUbhjTyiBPkvqGWeO5ewslY6hZ6Ved+slYZXrQZK
qr7G9b3heuaejlMERRfSm2pARlt7Ti1uYqXx73twc807Vd7HzaryWKP3Px/S7dFGqEckMnNnZDoH
8KmvBTNx3AsZeKU/FgDdYReY5H3L/Uhb3BYzlhpx4hMTH2p4dYVbXvSOTEpGCfzz2KRm3S6OLeRo
amFWYMuTg3KCQ7UvcEEfWOVUUzrxEg2EwpMYkfCdnglloDem8uWZr6gIgTJKJpZJYK3niHgycO+g
lsoVgBQyKc/fNjWl8nMpcMsEfxlNdZCPDZHvtmethioACkCHaAx9dShhyrbmiEr8f9f3YYKo6Uq5
wH976fIkBeQSjGnQy7DUSebBpr3Vw8Dts9pW7327NjKTFt7EQ31AJeXa5CGM7VPchrXe9wdd1Rli
MaaluLm7Y68W6m3AGCUvMJkLyQwzBoPApdcBVWCDVVJMXIuiO0GeFN1m+Gjvae2qGEvJkVSo4Gzc
lSX0KR/krcyMztoixHPPWihZ7LTmttu7d8SM5HebKZC6cg8wiA9a4DqX2azY2T8bcoR0XHsswgus
GiHuB6QIMTfnqrZXQGFidbFtmcX2QOneIHIBotKkaQRZO10SiZ9PUYzG4zkRpEnuSc+5iYKf250d
Gfr2TawAdkFNFEm8Cy3CrxyWlRltdXsqnLv8rRz1Kf2tlTBV/wDm4Kp02cCv4svV4DewDt6RrWPj
vmr10QQC3DRHt7jrUSCTnC3zuKWCmoG9ZCSWfwbXC9zTw7nfcr/rhGqBMJpj01gSyTeqFzbRmMp5
ZljJtCxQmtyJBly7lhrE7Pmz+EEVRV1TiZU6cgjnzklm2oj5Quv7Rq7qRaX/jR2ptG4/ShQYQkD2
7jJHkLLDKohOEVR901f2jmVHVX2cjOGLJmdf43NidsojIMq4oI8PpDA/NLzbtRpz7IIf3AWc9+mQ
BgzF99JBQpCm4ZT1bgvqTZ7nUicCOchGP4JdgoAJo2TVyp0kyrE4wx9s7V+Pw9a/b2kiPRsBa6uV
3F7WldNoTQI/OrVYXlD/cxfF26QNfUlOgPeCpxvuR8yKTO1xArq/ZikA+AgcIu6KKi2cNZf6xp/9
3YzaHXOMkvIFQHcsDvThBBHmE/Aa45lQUImZFWIpqded2heVokywn0lx8IWgXNYwi/FkzAwrwwIH
qKpZTQrJ7qZ1qaYfcxOp5XxMyIZ2aHUPLuosOnr4HQIsCjDzNvmJmZiGadPJpw3KLaA6c+RvGyYa
+m+BwwsJCG98wbHmpHO/F9bB25I+ZfsorC9bbnDJON+hBvT/amhmAbQRTOcgEm1ic2EbMRfzk6HW
GLCmaspufa/LiIEGe0Z33lWI/PosVITmMWucZMU15EWCER5wJ6bEYSeVy8G+G87Ld6ZKscVWcCw4
/BdeMxZC+rTtc1U2oLXsxbg+MWIvtOkPHZeAL88v/6qPGMqxk8nK1pM+lBAVmc9cuJLk3W+m0Blo
xlCry7ptbWc6KWMptew68PFHPDqcZxdQIRYdH194BXNQ8zHI9tjzzAwcJKp9gZFV0qYaMj1l55oJ
FydoeCBDTWMNnj4PN1J9GM3hEd1HK2CXe6/qH1PdS6Vd6SoM5C4HWhwJCn5uQlOfpO/El0IluhqK
KE+YOmn/R8BOm1CG1uBxSn4uwo/e5xW9wxdBLyU5eYEvblKXqjJkeBAxHZ4b88pQMnfjxb+mrGjz
Llxqix5j0rGwi//1shV0XEfxNV6unRnVok3KRjj55hmlkcosRt1LzOnqC1KZbD7SdVOIgWFvSkoN
kHgV7ZFSFJR5c+PjV8QtYUP1zwkXjO5YIV5HrZdQfr8d/LOZNadfE4BGxIO++kcrPxtUAbVDfNPv
Dgx1SqmtjggtrE98wqSX0vqC9WLNNOKrmtcLBupO/TzkhL+4/cQbPzNH9OrLIMG5nvrnzaYPtk4e
wdpWcD4AyqWC9ER1bjDL/Tcv1DLuujDIOOOxaS6xhSpsGsBvERowBuZ1+YZv8EtX9MejN46PTRFI
nrWMbAaE+D+LcU9aFPU9fg1+iLm9Y3LMhxeL39a5i9WUfDhaukUW6SVcFD8rE2qMJD9F5jjAT/Bb
1j4XUde1Ht1eMeWVtDRme0AE4PD3ICuGbfBQuhJedDl+Fn2QfiCbIuZWyVP8Bltog4tgqhFxoSIx
BbWGYKwl/YNw1m1hAXj3KaA0ahWtQEfiXC+pJfhb/yZOduCTDgybRpXrPCpc2RjMbocsonJRnyA+
cCsiix1/kt3a6LHYueGNdEVMI1mhx/urquZY372aSXliq+gTu1ctx21PYVA6d9nFW9KsEXQKvnsV
rvtEj44BMq2JMMY1pIhNWud0rV1QUiK/KtPoDU6VulS7FXjMuTmIPRB+1Qjv+nJq0/WCei44SyDi
VD+6z7W3EGWPxSYehS4PEYklDw1ejNYEK+wT1n6m30FTMxX9bm1SrK3LrddpqNARB+crzu5kdM7T
kplFfog5VLIaN8DYU3KnJuiM6REaPbe9R/haUSwBswDnN1x9V5ocX2s/wujj5DovbOGKdNG2Jjtp
zBcR0vdGlNkHIH2VUImnoRLW1+Ll+t8dLRd9wYl5q6SGpt25ZqvUesnncJqt7kDJlQlEOA+nPleA
1U1u++wqe006rlxergDNia4Vzkp4G14GqzLXDu5y6/5q1p2yYOa32FjNewD8pv5fK/J5xF/euCEv
Icy/k1W2v80m7Y1EDoDhM95hkfb9cheI6CIrw10ZeFe9umOvNXByCGVj+KDiXKx0lnkHoMfcY0mZ
MmFFios6B5h+0AfFN3XWdnQCr3J1Qsj57yUAG7rQ5jvgH/yNqBAhcMVAWm9AF9fMwG4y6duQM/3b
Z68E2gpAsD/92zgtY00t59phU6WTp4KNJxpJ1E6m/nblbdHrUgwGqNVXAgyvFD2OTj+s3TUTVWJr
+YlZFJuY8tLURgrNg16EHkUr1O+soGcT0Fs48aDfPiGxeZRagvfQSXrKededYp/4r8q1bKpDeJPL
U+j/8YTEJU9yYxEuOLZmync4AEQCwfrKtmgvOnLl/alTBsiyfPgIiVnmyESWe350ME8W5dR2tPr7
BcIaqrjw3sMgzkze+BTZShq/MHKB820NzdNRM12itBUmZn7rRS/mzgNzGVAywmUqhYP0WtZh887D
CJAheCNT5EM0ldNcSW+mfUVAfKZZqEEkgfNef2B57IjSF3rRUAjZmtVq/zoOiNs17xz2CHTBH4Qs
B6XZsZiujxN693G8Dj9pLOmGSnvUCvWqEBSJsw/QcZ1NVLB/K0dWNJQz6n+9ONMmXSaYpwL4zvhG
V8RyxpyAs8Q4iyv9/v+cXuYwhsSDyZ7iydCB00Gk7qAoTgpvDvNB54nWvRPkWVZWEFl2vvqgNpOJ
d/uaecOPUE3sJ+bR82ikBTOzC15+PVOyOSi2yAi5KtWltcx25SGxZI3sojSaBeM4aIn1ynBZ8vBr
lJtRuCvwAL4ywcr5prtwCAW2Lpt9hW63h6mfOy2+IGBOKb7TrRI01kpsNpu6OmmU3NxdHUYO3/3q
gIomV3h/wzUhUe7Y2kwrOU0I3hSvcqqubqZuXcql2iD5nwQyTMIoDWfWPplV1u48pBWijMxR2Bqj
VwCJ409FP8JtzK9BtGNIU1HxPuVQcHNm30tFA+i7NO5X3Ao96FC/iYDMLyytjJXhNTY7amRYT+5w
bAVdDNSC98bfN08CpVo8fGxaOl7JtTv7Zxg0V0o9XV1mcPrTlWw9BAzPLuG4U9RFNGCfdo2KtpYj
hX9qIFpCJIWpWflCqceBCzFhySsNGUSKqS+vRf64UjGNeMS8Y2pKuP7jdf7F1IkZZ4n6KhX2SDxk
2LDYQ2H0lJs1Kx780Y9U28Hfk3Uctbj5bETyz8QhtQmiZgjhquRNKqmII06u031QwHgOAqFQZuiQ
cLtLsxsS9f4+yzEgv8u5TLpAj5s0V0CtNDz9wcnKrh8QmBhbWNQbxfqCQCQemkUvdtsYlka+Ptl3
XAvYVq5SIupkGrSsh6BDbtEf5IJP6J3wGnjlOW2clMNS/vKL4xmgBBIEAhQpGpYJe3b7w323/Oaf
IC/d0Ygw4qwuZxtHiBPPaGXmJECZi0S209Ne0uuPMmQWgk6QVc6169MzExnxOIRBd82waOyNco8a
7LWi8r0vrmVEeRMKnvePzV+PhUnt3TVfZR8KIRwiQ7MD4PHpPNmWM2vTMITXnJk7nars5j+mDXrP
aiidp0C24Y9YIOPdZbh3qVxVFpxPFfN1NVIINT++jzuNAbAUp04j86qhvJ9Qfz+KyHNJ8kmWVWfC
/sfKqTOb83kmdpvgfQujNbeiUWvhLfPvG0QpKXxhaItqAMmdfRvhC5nlg0mHEdpOFrezcrcrN6pr
4QNogT9waORfHVj29/dK1yLU/ZNjUKLzKgaWcbkPW8/dzavedISr7Z4+MH6wDmBAzxKRcMUsPfUk
VAfDoKit//c0VUkEJyGRheQvnummNLuXaeB95egeQe16IvZ4QyrIhQBQDAaPeHr8OO5splzhPDKh
5Fh6JIqQ4fH3uNVZzdD8Hx+VIrv9gq7VU8O39bEiaXc7iBnz2oJiZezGhp71pI+e9G5nI7zfqJc9
qSU7N9Gszggky6z7QOHwOu4N0KBGqriYW1Phb9j8MmAXK8U+cWeCOvWx1Aqq0SHZM/GUhjUBrBnw
l0qjTBf1ffHacWTUqZmWw0hpnANLIOsrzfqt/hyWMgS07yh52NYhLqEHPnxuT+iZNMl3sAYTmSW9
EeRQLZt1uMXeRkXlnRQzNer0pMFl6PQqo3YTqficN8p6eXs+9QCfgKQTfJ0vx92mR+SQ6rUSK8x8
LQwPrvYE3PsyAgsFSK0IXVYNzEJQjMT7dwPniv3FSnSk8y2k15hNhjrQII7oVDTuO2VN64Nag9JC
LMCjN/IyXJma/EJ9z9DFT0R2dFIxyU0B6t4aAF9IgF40Ac/U+MQkx3Tn14gJaYOZw/yapu/YkO9d
HDvH/P9QI/5UYHcTuLTV2eaYOhhfSeIxQ6CfqzangpwRPwcYZeWT/AO68wYlCZfhHsQw8krzed0R
mBKx/YXG/upszl62A65pyM/tOf4GGxoehbM+q8BBgDOud2aARgnLoCtipi8q6VXYjDgZPpCX1oXs
x8YQzIU8coXRJZiGrMzoRCqpqbyi8LjgCTvlJkjII/SP5A2jfl1IqYPwzxeSNUchApS6YggG75Cl
htgoZu+BBKwMyV/JEMM113tQk3auFF1GnjcQaBjl6Vtv2JxsEPUAEExx1Pn0nejKTVdQUIwzn24x
J+0LMBa7Gc14JaOFrPAv5VU81H0WRe6i9Zfydyz3w/1ASIZrLrIezQR7faF/ZoryMPN/0BwjU2ot
Wb9GHsw4OLRDMYV/qDKglqvH/IaWh/usUFXWRjaNkqNUmtY5nHAZFsOkmHV53BaW25UXGEHWspO7
5S2EWsOYaxGPWbGAB45j2Ls6PQ9LqG/E9ytOLQjoowDRiJNpWZPXuSLnMMpksBdQo7W2z89FJvje
uX5ewgEFlaeFoqt1K5UbZMvern4d6TVZvSfy1vFKIcAB2FCn1RxYNkEoMqucVXMNPTf1OZKSAe1D
BHocuebDS3igFf7L+8iP444htrlgEY8DMgflZ81+OKo2KYvm+JA5TMNYlJAYriUcVVz9/hraRmq/
mMK8mNL/yMpSNW8Zl7YYmP+KQa6itf2B5DvjMhvdP1J/7mjEvLNvyv2kEvbkvwK9ydUlUV+6P18Y
84RywOuhrMEsadK10Ei3nhVnqktc8Ql325JvA+DmE3ytWO+EK4QCVOYGH1BMmisNuXEpanVJ5DsB
K+Db67d6y8VQeoF5l/lr+iNxC407C0JZKKPq9OeTjD8VuTw7tspeAGnDm1kC3KzeDhegVgmQ9Jyb
flt/tZTYu2qMP9ehGY1LRTftxCHYcIYKrY0LGAOUxkknpiRNl8JreV4nt1HwaKbLr+tsmEYs0iZI
Eiaph+I4WirxUN55poNoBdfz8fZEOyQ5j5aOheG4onzZM65XPqx+7X5MoxSc1cMPt0NQx3lueAza
V8+m1tU4EIStIMlUirrFtuAn059T0MnErKVoZ7mtS6bLlTjB/+7x1W95b38ClrT2vylGS8yhXlBD
wSYQ/tDuEtbeTkxVp2ub8VdKC0VeBzogTjw/XwrQgP8F89trhbuSjsYe6rFhjtbz5xsybDUroWj8
zDQyXCGOkYV7ej/K6xd7v08zfwh8DfhOkbAIHr1RyU2sjBJq5o6CI6Dn9xTZSHdCWPURAtjeikoc
WErFo6Zx0x92xhBdIJSm213GveZXLguzAcOIvVxnG9/rffP7hf+0HaqUpk8OwCJpEbAQnl+P3PBS
zvws80AYxc/8dJgB3GkP9jNESjdpaomdjkWCrFOQs0rpa8YvdG507bwUVbUJ2az6zjrrka6CuhhD
RVjvm5I6krROlWmPGTd6G/qvhYyAXJoDJQFQdGxZfWQmxqJWyv83XJd5QjbEC1mrqvtckd4xSsou
s5GsSgyHKaxr1XImmU+0z37dgxWc/xOTarwXL0/KTLxSkJOz1RuzH8Qpa7UC82wohOvasKznr9T+
BpEYgo4SQvxm9YPp+UiBQ5BdA83bZlHb2aDEwmkTzQf9rWz49DxVDJTr8AhNvFTehqjOlSQEg7lE
eibHT8YbysFEbSfUmPoLDiKURztY0r7EFvtGAStEwBpNrUdAMUnfkLjnyHF1kAUtYQOuLVIud4EW
S69+On7jW3gaWfaGY6VopCUZIl0vprVGQ/Pwl501xVrI36mMWvteHD9IAkbVbrDrK3CTAcGgeKyN
UVeOoS2P9zyNRLfbHHSjpKkJEe3lBlANYWHIpLsIHLKb/8euslTpP2aTl/oiekTtfXmzge3kIrfr
0J1J14DlpTES7XW8yNv6gAXJvx6EVGv8GedqOGo9vVTBg0PDlnqw7E75jM8tTg8o9g4igasomlFl
Q9E3w7NqghMJfNSmAPM2yUGKdvPNMrCXR2BLpOnNBJAU/iNzGtMSW6VUtX6deEq9ZDAQl0GhwQ5b
r18QcHRl1WvdJU8S8t3zxrRhe6ElaTeAcCeXdeOEwNwczOg7Z0e7lTuIv4oKQKq7viSvNF5DiGsz
LROWTdAuJRt4WKYHoLzwSc5QdXDDsCzxFdSsxUffP/lF2AjnRDROy2mSetYDGDeGKi6UOzb3p23H
qDZ+huTKQ7pHY/Bbb1gNyT/mqCh+sp+4Df2Wlk4CdHPzZbPjMsqjvVErZkUnDzY7PZrtCMVgoOVe
KNyl9Pk2D1cK8PLFTFy+vnFxg3JJg1mrdzrWOIPLADHl1gtZnrh4lX23EzUcrc+RK/EHT+sx2zLb
Np1vyweU7Fll6Lsg2aK8ix6xBrnGOe+SAdrhon+BSbMyOLVKAxz/CbAW0nPpfu0RQlrP+oiiR3Mx
8AVb3lSLhAXXbsafF0YF7qUN04QffyAlqi+pKmOl9E5deCEggY6sgjwyGECIzPYIXjE8WZrY9zTI
HPRVCyK7sMba9xd/3OohmKQWmp4/3cncIOFCkj/6CnQCXmI4FzIDXiRzRLLMCeVVajEqascWth6x
H/DvW0/kRiLZ8ik55sybZ0Q33JUq5iZ69G6wPenrv1jnuWtbNZL3BqNpM7bEIMxMHjqYlO92GPAn
jPsQzCxFNTELJfSmtfOrYwSJdu6SDEZ3El1COkWgsXhci1hCbAdiHC/qQJIyjpA+hWld/7XTz/Nv
+6dSzRqUBOBsLM2PltEWkzXR8RzKanHd2u3xFe5g23Mc9yYN/8nz5T7j6JweszXmqMEl0naF9YMK
Xwx/jkBRtqVzpvqaRYGaNOpQLKPavtsRK10uGxM5l3sWQtaiONqQQVKi+DiEXCe243NDElDz97EC
xj84SfeCoR85S5BxyC71FSHQxN5L3YJdWvXlC4feHuc3UptE7Vmsx8VYWE8Lb7pVALwog/me5Mu8
9Z5m5nqoaWWgg/YbsCqTZKxK0EHVCvT8tbkoCU0o23uwNPusTf5CAZ2Rj0qAWpe01Qa9g5jBNTHR
EiZACKDg3NZ/M+ye1moa8c4Y+hYE+k23AXm9Uc4T9/yAe3lUFNRz4/QCkJqLpqL0pMEbXoAaOHpu
rcZRfqtwI0P2/21QpO0nhabvj3caP8n+NKsQOWFwBcToVJI9gejhtYfw6LLOl+WmBS987WBrfUyd
JlQwzfVB82rcBej4CsRqBZJF34AhK1Eobx0kCq5fiBazY85Yx+MuF9sJaV4CbkXYIzwT1sqLTEAU
6pFociAQp0PKwx6wWZw8RHn+TsUZI97/pD6qKtQmzLXIcz2/C2BIHGBmFE7QLq0cFU5RSb358boN
oelGqgORuQ/MVjRcS9C1GbHdE86Uxf4urCLdsL0hWbs3odJQ3QQke+53O/haYZjV1BHzvtKt+V/z
hyQX8pncFYwl7I+M0P3XIL/QxZqi0wLWMVRklIOsYR7FQj2D6AGnM4zg4HUJT6ZzpHPZy5cSib94
bdRw9Bnd+PHpj/NLRQkYMcu4GTI/xqrdihHnJbKV58LIyVkbf6x4WMIPolqBUnqaUB29cMlhlAJT
DlVpRo6Oo9UADlu6Q6/PjjBzRUuQ5wPkxzZ9HCuiYxVGET7eA4qTKrMePEZqn1S0/SWvWb7uRTr4
c+q5SDdARtJqv/tGFJvthBiXW4kECbykzvB5TFYM8xQSgs4fT2O0CasdZ8l0eNA16S8J4e/vajvW
HkMYQltIw0XdWuHV6l4T/oi8IikrwdiqXq1mMglHuKqUSoI2f0uOTBr5fURU7XDaDbUODXEuCr/X
JWL8GJrA5PPrBdeAew6Ke1Ghdbj/yagL4+Mj59F7IhL71DLrF6HhzJYXRrmMbz3v3bmwXFqs2rdW
L3p5J3FYBGuDieshCLf4jpdz/fIBM8Hn7C/LRTYKHNA9iqsIzKzOPoCk1U/IhOztovkaOfeWzgaU
Cy3LXDO2BFbQGTMI3FM5lw/x7kdbbWul74CmYHw+A6Eq38lq5bj0J15Qlk8QwS8hPEmqoOdwmEaH
3yoevkJY3laUQ0k0d1/oaEk3OTPTFcHSZTk3Zigm3jkrjLSZH7HH4x/+9CX6xyXKgXZYwiDKAY0a
mMFQcgmP1dsYQRXKtMboj7FoWQj83etJ/D3HwKzVGGuNn2+J3qHiTAeA7Na0I/ZitW3FW/bWzIYH
jhJ5IWCFmyO2SVtU+zUt3M7Clku8HQMLuQfARYyShqxAY18BGZxv60K6zvxtdFk4yxzGdUxZcFNc
Fb7HQZ3k1YZl9MidNfNpUNfH74ps+iKa16y1o0BQoyzunMgcOrsdevLVmSc9wbm8oxkX1gsRbbPw
yHYY+WxnH9pIls66cUHtj1dhm72oy4KzA3WP6v6+SKJGUWXJuNLzRU+wLS2RaBCOlgAP/RDpXlQE
3+jbLv+auOBe7umi941BxLomSCxbTRffemAZEb3uq9b26tqFvw/w3vpDSdR+R6oZ2eG4CEXsMdP3
Ehr907RkOodZeEeOVfVwew4ky8xPp9uhkGG0/xE4Dl78S81oGulMFgs+Q9dIgtG4Xopjn8MObjDs
q0CdEpWotqjjjGGeUzEZLf6dsU85hpVxp6u52q+wMlSRUrILsiz9pbvImPFNHEiG1wKn0JC8Tvfo
w5JpStRQCM5PjN+sWW1K5kquCHQBtHzuvQezKLSVsAuHMAMT6iK1tO7rFwt6GN6VXzgZYDmffUeH
IT1+bAYJa4QOvr7N54lm0Dh1Lk9D0d3rH9HfOpMwiXTUQX4gMVqfSetCY3ch70XKJvTEL3f7sO50
5sNNtKQDwNgstUfyzvDzFmhL5Eso2Vm69/RAlI0GYeSaA/s4KFRtNOSHQiX6AYnmzJ/bATNr1Ew/
8Too4vhDOnxC9kqWkDdUsalnrjH2iMbmYAj4tRgZyEHEx2I13FVBbut0XbQfLCugNX4Bq4rfRsNf
pQdzSBm6Sr6OKVnzIJwPsQjWS23UfaWb5K2TuEtbGC1B67pY1gCuZeWDiCDfOaw83r3cii7DrjCp
S4UxuLur5JQ3KjhjWJ7n4MtEHo1PkmkkQejEdBx/mSH0pCVuw9xcmT0nAf2ufuzw0COCvWGtGz9z
MIyNKtf1nu+g1+ieZPmB4iNUXW+yJTsKUTN42m001Kxszz+WZnFQs7uY9bgXoNq5ppxKJhU5y/hi
hZKkR+ILHBDYNTe7mTVBv+DsPwYYybPlCIs6MOuEwDMtesPs3KptUkhQ3UgynDq3Lyue16FWZ1sK
usd/QJyt4ckryferNb0+P9dnVIU1PlaD9OC2U4kNdPDbRYwJ1mhUjOxqC0MFzDvlaazKdsiXgu1S
k/N7YIIZdsYUyNkNg/SF04ENC7weg+0PnY1bpdULVhUzABG1+QGpGGSfmiesRE7ncRYp9uK0GuFH
SoUd61FTmiZChhrIJlh7uZqNesY0Gwd7I7bH/FOzQ3bszC4H/3PaK7AAhr77lni2sI7ywrzfdGAO
kzZWnn185jEdacLBAdYiIajaQj/TRjSQtAC+FCtZCxllwKodIIhE7TL5xEnMUpNoPt3/af1Wev0C
WI6BMBJf605nb0TB8hZmCqpSANvuEKS7Ffe2xbuYMOuGGRgE33jKEBu9Ah2FmZ0OEEO7WEDXsxHP
V2UXzdNfRNrRYLJAG6RSWPIKgBF/nLs7aJ21DYoEO9s9T/SMqh2SV+bE7tYEXrVJubT0JB5h8JfM
fnSh9c0ONzOaq8xuCP/ciJeGfKedqIxfvSzSNJm/mcvaqCAiuFxgUjozIfjFhmadvAe/k8mAZC/a
K7hTiPb7qix5OKaPlvL0Nix/bszK65jEJM7nScBAnq1TdXCbqH5x9v6QtQ3KKqC61lwoi8Oq0AP9
4LM0JIgghiO44oftHC2dR4/qbx8nkRXDJWJgPV7PF/5tuNM3ZqomllN4ncr33lLwh2iYShRJfJgO
Wrc1nzNwdVMqS6h2KCi6ONA+ddW9hZgNlcXiy9y5bpVhvtbSj6MEfcFpJeuUWcpCPeiAEYuSnmc/
wCMixN3NeJ+HRQFPrsS1fvNY/kkfMGYykoCfg3K2nplX8c26pReXG4jepzD8qcZtZLK13tlMbKHt
kuRkBPVhR8eYtA6K5zNCdaldEXF3rRRypGPZi9VCBBPyGKrSbsHoucLWjE2sA7IXcB0bLrgDBbGC
5MeDa6yELvtkLVJ0nETdN7d9ntLAxc65fKbPqArzW/TQar+2c3njrUzypSMHtn7/lnv+DvnpeUWs
VdSf2RaOBTyBWvZAGWvvhaINRKNAgFo34/P+qmJHF2G8T3Kb5vO8leWtGHMY8bL3mvZ/EwF2RzGM
qOgXk4RURJuzNB5st0oDtuUIkADkLY5QdrdFmBBlcf3+gcTLSwxBsJ4FGZyRlEj1lvm1yYbNdYSo
9DPdPbofqDW1CWOcvVv48R4v6SCsmGwbwy/MQsJj8HNR3N4sOLE7rylpGlw3onhPEU/qskMrqLgl
/MxXZvTudKB1xYP4tIKKMpNXSlQLqAwLfQZ3pbADxR3+3UQ0DzN4GvkN5bl/eLy+4cJzPpm9yefy
E3BiI31iQ0XVs21b6dSpH3yxHoYx/WE05qkvQTsnn8pc9xoTVsT4shMf0XAE+RpFqWB96wjdSt/Z
ozpuA+pg/wcEA5Zp4Svy1SBr2FEJd5JfcaVRXNOD1uttOHDi/ghKvlHNjQdeV+2tUtufEA+n3Obj
6rLE9RBr3YjAWfyGJcTvdOu9y7mc4K2O7YDWI/HkNxBE+sGcV3LUMn1WlREie+J4NpPb/UnGaDvK
JBMD+diz55TqEY93ONn0+g8zR1Tj8otzUaxcEXLJHGIIAEw3g+hRWahbO/Nc75VOsIprz/EjCHD6
CobXFaLrzqdihiCYx27p+CeK5nWsEz3o9a9fgtNFztgpAiRTUXTsS50gVgSazhVqK3bdZhv+fmPe
k5pqZ9s0VDwzAr9bFaJ/K0CizMfj0q8ITEOVZNTXyZ935HsHrnKSjB4l9dJ4Tjsz0E0iUNDtAQYe
yZgkKwQxDKcrpDSCplj1zKhq+6QvnCa2WffCQ1c2uE9aYMs3ZpJC8c7VYM2ZBaDGIYMTxm612VYY
JyQuGHgDqH778WfQHFvGujd1tjRGkpGLVkKGLpV6zY743jjQguNaoACmr2yIHAR9BVOeiIzcRj8a
oZmH4yaJ0asLS0zMd/8xTxQ5URlJqCuSGaFT1zHkhHbIzBLpGsOkl5cwU4Oull9VUOKtBv1duotI
QXDG0pHI1ODsYzoG2KIh1xL70QsS+SQ0GOo71JevYmeY7kUeYc9WtpzKoQsq8HUzsboUPf4Xyck2
e7Wr8br2rW0gCJTKeDOGJezKuxsV/NVyLVEmu+ECoMC3thHxKE6DBGzOAQ4O5RIy87ZlOsCd0xT/
hXlYb5yqcvzTJKZj+9hHsJSSGGlO9kOXafU4wVPN/4GgHd0ZfIq96Py9j1oLkl5VSyLbtrI+xS0v
152CuG71SLfKsk4xrDH5QZHJ1UBvi8Xg/019s26agUXe04DxU1HEsnvvDteSUq3u9ia4MyEDvzBJ
LjoKg5V0eRkn/Y34iTYLq1UQ4SR+hbAVNKpAk4RSpijVQeEQmUXTRgX/Wu1qhqNgKp46fgSJxFCy
e1JycF18oNoTdQpsuRzWBiSJlSw+DZ6VTfF/qaLYoouxCfC489uJdaGc24tvYZWqqLUJvm4DF2f0
Ler7gyJC43qI6xr8qSmB+UdY6FfpQdhjQzwM9OpjAz2CrfgbAZKZV3recUD6w+CP+YTGyqxWAvb9
gE/yAtEz/hOslqG9jmAh3h/wdZ5M3Spd7sd3/qrBzdnp6BcVSTTmUd+rsyzKIr7kMrk1xjk0ZkUb
KYR2ZpgHKg6pO991ygSe+rNPp+mE4qjtPyKuH5hhDvH5kymNeoVUEq4AewPMreb182v2L7agQDWx
gS8oT547nh9WRi8ZjQBf3apbB4OFD/kNaOWan/0uSy6QaO7KgXOGxiRYihrjRPUZEfUBBViIVHN3
gCFkyP1Zmo1cAu9k8BwPsg+fknmW38HRpOlsvT8d5nTHMh/bmpQsrAaaK4MdqpXMLgPu4bCl6cXI
yGnFfoYiiwccIcxrI0FAPJwFeh85G5rdx8ogwLwbS4iGIEDQ6Ze+V+o/rWYW3bPdlhxAkgkPGZLy
8im8t9FguriOariyimh/rmKMRNlHEil2+VNQersMRnDc8PXqfDpc2ZVKss3noMUdhwsWhT0veXEp
KnUDu5/ptQoHWt5KVREPT6BFGdia11Xrc5B/nwtZvqy1JraWc4ki90/jd98r9J8riDmVsGg4jezf
oOMqrfrRme9GwZrETcy8O27Yzd4YIdwhmjS/vvMpRiF3xT+X99d48tqOiw9oUrp6CI8swJG6cywR
kpBaAT0nHS6wH2MPKSka6zlTkw95Oc/6ppbljROdHF5c1EjqYXRYg8bGh3bvmvngWRV+TTpBxwuK
v4wBvEl5Q303Q1CG+5FmRRTEXX5Rrbppumzkp8gf8dPlCXsFYhgAMfkk4a53aiakPASztS8nEvfI
n7CDr0/xR63gAFdS27FMZ5b4j2/jSKm6C8ZhhlBJFliDyswY6PmaXDdBSlQt+hpmHdGF3gz0WABM
MYx2YEcasXCqpzQxOESa0aEzkwKE3/ZgVJjaaE7O5rGRpG7WTC4VUAn7sB0UM2OP3aKySVw6/WSj
jJANwef3z/prlyj+1KwpKYLv6cC884PFpdSr3rStkyJzPe4bOb1kWADH/DHuCtEwksGhcBjTVtwU
Gs8PAD6wTOo0txmXhuR1QZmXyGsxkCx3A0SSgXjsbRUiRWU2VKRxECckVZqkYyP1UrDy+jqmcDRu
7ZF25VVjaMqj2TqdpBHUVrrU2bC84DmI8jifv1pWi1AFY0N/V/tr8KavfKHOea5ZT/6yqD64Tbxu
Lc829T3hVdMCTAc77oulNMUSlpTluBRX+z3Df7mXq50+vy673y98+BvB4ztAAaj/R0h8H2gTJO1C
0uxRTEyBo/FJ96uCdnV0GiYlqCEnomPmFzNcA3apg9/XIPu24EHHs8LSWVmLPvFt/z5u82iXlWU3
SExk9bfHc332zixERAH9lNEwqzQwbKdj/OBhAY2dklmDuFfg4DA+wri4cZONhkwYfNIn73/zEcJb
M/wBS3EJJPK0hOgGhGst9Y29MBvmJzU8qNt+08h6g8oCHjbA6OdRLofJ3ISEGtPVrxlGK7m1cv3W
BqUmMVdBDJsPrCeZO95TLTG5I3HAQheYUwac28peWzoy2r3n2eiBgezWQFO+XEsVRkWqkfIemeUM
RTT79YruIX1IIumo5K2+FwyCjxmwmiXftV7PBT7NsRUpxI3I0ZMOg6OhEdshT+sC4S//aUc+Se9a
69a9aYxT1/MgTIAXStqpeYukGfUvG60wO4pCDUuVPHBxd3MBQqyfJ8XqIDMRIngbgb4ycPbLdbyK
/DAgDyoDWgJ2sCxKnQYhQGHrlRD9h4c1xsS29E9JCn179/tDFArZIl9LeYvQ7U0057scPp5q/CK2
wh9orJDAdrJgvwB/ertiT0xCUyro1j8Yw92/DCHYj6+h5aMyTfurXmPClsWp0WtZCKOjnk6o2KQv
OcDR+4iQNwklo8EqLK+9eZp2bXF25MesaWqk9Q128PCo+CAr9vBtqS1dPXi3tsmsq9gay1zeJSWE
zL6u7yxwLzUSsQQfz/ovLCsn2YLQ/wH2grYFsvRNZCMquLbrJSJI3Xc8GlZgv83YJao4h43MAdX8
5lCaiB15ZHfg55yz4B3QW6cRrjxbg+vb1UxmdZuaX1kcOfYiPWuEnJ/ZklNGb8mx7E59P2zgN39M
ryA0GZSpN9GLYa6+PpFrCFG2GjQwg/8+eqBWByBnblI3RmGgdyqVou7u6RpNeW3faPFLm/tq/Toy
3SCQAexk4w1bXnF10m5swu4pTRyCZpzk9Ptf3ST+7FCy2Pzj1+8kd048eshGTik+Erclafys5c3R
amb0+715KCSFPM5lhOu3hsumkI2N4xBJ1QAsQECHNQ3ksxFWOz7fH6J3G7Lx0qJCpSX8pHRyxBGP
DxeK9bPrplJMmhQFbw6Oluqfp6iarG+lT/kQZXxjZ020T6SWE+9tPBGnAtr5jCHXLG43HiX8xFcl
FRqIFxDoyA5+PbdbBeRROnW4q+N0QM1IxMgCBan18Rkja6mz2oVDDo3OcgTloS3CPZtz/VubaLez
wNLCowY+xgGIx73UHTCK7KdchDXc7IRPBSlv5DofjxY0keRFkXUw5/WMW0WPY9GsuD3kw2rE8qla
i7UNw98HzrK9GQ4CMcIUjt+atg0T+UsSotB8ZI1gIGDlG/QmTbZCR4cK3mS5xSARoBURnV9NxA24
3tEp9NB6HK0vQfjYW8IU1yL4VKzjIkHYwE+Ww90BxfJtOV0UvIEe220XsNaRLB9hNiscZIaeviFa
dbzHC5EalKcYXQlmmypA5cjYwAr+JLyz9t5mZOMmH6M+8d+NDHMekzR1TLCPkR7Efj3pL67Lhpx+
WTV3ubpJTuOrfyXGlt7x9bhh6sv7JWqvIPKmb/0Rt2GBK1SsOgoDu7SirRuf7l9cl5nq/jSi6RB9
Z0+lGH29wdBE5/EqQoaf4SQPE4KgYwXC43zZ2EqrROY/MwSXhvzxlS7qSxHTddnFf6ukbjJwtlaj
m9wt1PVf4hySCw7SKYdDsWXelK75v20JWxBpUANiCWHw6F+BJ1yjcvyj6DcGt/r+IxpHW03YUFGz
j2PNEWPbmp2SWnw51kvCRqr26MB0g8/gQRlFmQVJ0RcLg/c7qDdiQto2ob7pvpGyxRTQpE/oyzUl
CxICaQF2gVvK8uiIRxi+dgQvHo1D3jXPe0Clbvqkqd1rx7Xf2DYTcwDZHDZpXcnvXkQz1m9H0z0R
A4y6SDbNtTKjHEb8yqlKp/0GSwjxcf5y9M30FPHmwo9tue5atFauV4mog4wKECZH6ouE6Lampv8C
vJXenaLshgg4QclMko0Y/057kGqKj48pjdG4BQXTd2EClyodz/5curnVauVQIoCS379TJnZZPAZ1
rqFqfnpGJQG3h2EBdrPono1Q8JEBaKgPMtdGxKvfRVyXHRegFE3/ejwJQnrc7UQEoSBRcKpHtUaT
FD2vt+T7QGsl2ptSm8l7tcYSQozmaHmYPPsAbXGEHV1aCBHesqPjOJ4c7Xz4Le1zj4csK70PCeRT
xNC6/47FHkzLijus/q7Ih6O4fD+ghR/Dc1emZmJxS3cg2dmQvBCnc1hW8mj9D/x4FXSKwTzNbaIw
7O4AU8NZgOoqeTwaSxnZ2bq2QUpfSjHzMyi2meJQ11QkNIvzztzmB4ish5lSmbDfbM8q2N1jyFBw
xAXZdDStIocZcQ2iWcspn0ifWtauSzxOUdzAAgmOda3AlZ0QvEDLpOpuhiYY6Khx7/fIY1aCFYMx
vtL3qhjzwsSD6qxdx7b912D9TDXARJBfZ5Y6wL3XSqHLRavX3adfDdCzvxugIn73+pOVe+1N85LM
yG+cV0qf1bYSyy7CgObk3uVao/Zdqj7uwjOfOle6AMaoCSHPXq+lm8nKOyEc7Qn8qajQ3xme7EPB
Uul9YiLndyhGrliX0+jz8iPDIEpAgURpQslEx57YW2EttRHGvYFJephRb9/U/vItI/GhWHm4eKEp
A/E3TX3PzB7LPTlrdYSB8o65OIvRTxP11B16VUudVkqGB4mFAw4R+oza/i0RLuiT2NETmUj18m3a
QR2oSXMAHmalasa6oqnKpt2dWVJC73Tgp8pDH4pOrm7tQfQZV4CwcCcwznE9B9/6X+P1YBVGKTdo
HhDNsN6AAlTYg0MeKBedFmGAU0A3Veh4wmn6ROTligvtH/tQFUztZALxzbM88Uf2/uH3m9JpQ1u8
hsnUoCal/xs3+xyFrfl98Am2mo4hjXEhVa30a490dHiXraTMGuwXgIk32ByDUFMULVIU5ePiU5sg
oSl6sF9O4CJGDIQ1TlkM1QoigmEDyXncHbnVaZnLc5JI/PmlQL9szUgjUckz3EvJ18rXvny8FHLk
NiuSwzyttezmTFDEZu2Nw3H3/yF1e2dg0kQkjmqOsDMG2+kmtHEY/TxlwI9jRxR7GEuYEJS9rMzN
7yLQR3k+NghinIEULD9//6lWLPmXCZy8zU4dEBdogWA94Rekt161v+eoCoe/vAngpmb9JPmY6JJb
/oGu1Ggz7A0sMxov5oaajmv6ERzI8R13ef/W3LT3qMJtfYNR13QI7i4GDrB+lZymtzpFm6XLkSI2
v6tGzUrC51wiXVrpig0NBI3550hoXfMVvlQiUKuhKSCbDxDBykE9FQOKUDP9FP7znqhlIZNRRmGu
66+ysRAUs+7FywS+2zczcdIo4Bt4cSyATt/l0c6M8/KFQlsh3OFXnzreX3iDGiUg6kjhhbaO+gAl
2URwVU00Q953UWJPT1GwyrJly/+ODdVp32/tDItmYDLicotkSL/TNuXiJ5qh2YWYcqzR55n5eV+j
wzSy/vKmwOAmJdJegSdOaAzZVV002Vh9kDPaWoDa6Du3mbyxaNgaUOVDIvOKxR3Nen77FfQWWgDx
Cov8o3+k9aAoZKnGPhci93CywwzZKthWnOZ6QJ8qVZtSCEi6+o1n8VmLzed3OEis9mbrG8rJo/es
+nvaCweRL1V0lYKicEck4/UKUH0eZ3Zv9MV39FLXJB9GYvosjRJKQbD6nD0F7ggNt58mQTyoLgLO
RLf1cwRE6wCEFwnzuBfcISBs2JtD5mD9PjiSLDKUKsOtVXTKDn4V1e50Ojio6GBBgfOKvYwm+Jr9
HH99jjihCCHatgVWDrXfSEicsk0u42eNf69Y4rYx9gqd065f/F+rMa0eObefkSQ2ECA3S74Age4h
QTN9/fqMnUTeaNl56HYTAEOzG4yC9ljd3+gcz96XMuHUasv8oPREBUvokg1tJGjU/gG5wzwxa9Kg
dmt40SlrtLCnB8JkM9PVpQ1Jy1FUkeqk6t19hBVi5RKy/Fnvmaoy55pXQE8Cgzjv2TVe7hMm/uO9
QAbygnak/0cbKdu00DMknrATb2W9/fFhMiaZjOZ1dqmhyxitLwN8qVicCca3TisCZMTZ+cryXAh2
L4rmsTFFNO/l/D0/snXV4maqG7SFIwnRsM1Mg7/lrOV0lO6Ih9nlDxfTfuWQr3AZRcu2MkVOWeC5
SZSxD3mtCtPXGgRYUSjjBqh9y47qQgKyC9qK7McdhVFNH24Gf1ewE6jXl0/m7A3VM8rTfIsCYyR/
ggvUYKiQ/XgHA5DnBd0RGsYfHywTE9Po0dJBUNyJ9FhLczGoLoUWTqZlQtoC8Wli7OjWpjgvXYqp
BRISq1pguWIbS9S+nXr/eMMVlk+i7h8pn4+4w9Is62Frmu1XyjYt8FI2gmh24mKaGBksOZ2FhPC1
I7F1v4mMsQ/0/zQqJFLmhuOBCokptD6D31EPyEZBZXx0pE281pUoRupcVyCXgRcmYbzpQSzPdyxY
QGsD9+66QwLNhSbB0AOZvsa/U/yRcrsibRq5fpEbIhS0n528kVu6Akn7qQO+JNYdoZUD82zUl0gW
JCla9YJwqVPalaf54Hy2Il0O9wUSCnJJ6zkQSHprzsJgbTaM9mNXzmN+dgJelrRbQF2fHHtvkPtp
QMr7jdCl038Sq1pwv7+g3T/P5lgm2yUPKfx3h5kv04O798F6vPwmMRCxISTmqP9HEAE3nffvjlxZ
vDrlkoPxeMl6dn7OJGqj4HUHXPxK/hQOrJcf2Ki3G+Tl8kXk+T5vQlkO2vodwSK/t8keAVSoYm36
nqXeNKzIrya2mKJVj6T3rL0kOQBlnhQhV3hDt8BwQ2B2NMz4mfJ4RL95M9QTpT8yr/QMiGnr0/OX
x3Q9Unie1YfG5Z/qaftf+zFRulNRJ/wZzbszik+NkRGJcZccTEjdojn1JTIKy7O2bdhJaopZC3+5
Zi2zBZ6PTL949TCYcMEjz0KGerYh2egG32cgyhEoAsH4/dKk4SRAZvuTEAhHnMEyCLylH0Sin05m
M9JdPrBF20BUuM5kAjPPm1LscqYahwYFWXvbFLw76iJp5rKI4MUQJEy+vLIWpWK46Foqc3sXnHCU
xPf2fKeWm3xMDwRfZsx3YG2ENGwfJDuyY7NgiUdzCcCnrjQnabS4l8Xg1zcwLX7tpt+Q4gTmjU3G
msfblgTehaXB5DbQEbF70vTTm51X4D2fkSPHUWvYwh73XVCPKkyEJXd0vh4oy3bpsv9DOzedm27G
65LI/aCvPPBWrzqs2LxGR5F37tlLOzOLisCQFFACoRaeozuuJmC7Kza4WbVIW2T4q9RkKqZwXZMM
b2gNBENv8/mpFIwogP3tzA1N/CaCAXQjXR2PY8BAwX4JCbfPQfLR+b3fYWmekdSAQc+jkuXmwmPz
W7OlP5y1REqb6sW76Cr7SbONgl7r/h0fACyYwnKDcjqxe8lGSjKBK+j5zXHQLRU1VxD95tIjwxOo
9nWK349jPdS+uAw6N0hcF6AcNwzD5AIjHzBNXbA1sbZVKM93hw1R6wYDGMTGh+boj5rdKW6obPfk
SepY5TeNejLHuSv73TgNHsCjQWCftwNfP0l/uhLlvvifl+wC0ZWvig0/MBcrU5uSdaqlxFXqJgmj
9dkA3fjLxSvGz0JLvQqfUGMt4pqKNSIpZyyaH6xEbrk/0n9MgxahfljsPSzW64GDFAXiNCfkyA/K
OGrtgF3xqaQF5mEw8Iuts68gabKwicAclgDOl+r4hWAP5mcuUSIxF5BYIZq8xWQvKOv0biuH62yh
UPHmvS6fKUJC2kjeeTbdb6i0XAw728iBNEBLs9rfsTXfzvpAZ9cgEyte82mvKdkCAWskTL1IOngY
wpk3EnOzwiHUjEFqeP3t7RDzk9iDoTnP/BNimD0WQgBTiCIJQ0zr/4Mfw1BFXA12qhHtXoJiMDmu
Oyf1/QMNZK82h5xI0/C7jhFPBMCXq++BnurEBOGqOyYMQDXRjXw/tuBdnZQUQ9mmcM5T6THW8LrZ
q6lIXYdC+OCdOeFgsbKTXg1XrxslaIobkcMEqnOZfflOYySo75XG4tawtHUvwvCxt+Moui+l1ZUj
jVv+/amVaXMPSXF3Sqv9newh30RuKuyl5glg+Yzm6i1JI1qepLYoSipBWdjtdkuhkjL3EYKf+12b
FfZxt+vqzjTUjIvk32htq5EMg4ZA5l5gWUJ6taCCiLhXE1g/awHBMQrfrsx2Ft7Y2ON9TT3o0vAD
82gwUunja/DBvWhcMjfXkDc2F0V5TKY+Y4SuA1h5jI1EMLjCQX4iNmFkIxLzZSWIyXwKMPDKZnJF
qmzhfVaDggeSeocf9tO+gYPEJ+dj516uytW4eyM+L1SohdhBp+3xse761nbZFIGTMqOxz6I+aw+5
vLjCg7PV9fjWIqrzvUo64KMP2QrTl34Jem7wywDxXelwzu3iCEe5acMkc6SUfacl2i9BKAVZNSsD
+I07obneLZFl1bdZjcahUY687+LvoxJtTTxGlmVmXeOUG562EPsXiqyEpUNXNxT2CzD2y00qPeUa
OgwKelQb//PcN9FS46xeW/1hqhaPvERnTb0Xe5dxz/J3zZIbxcQMWTP3g7jUuyWQVf+QTjTnL9eH
ve9ZjD2l3hOjeHf5Lis6KZWv939bzwUxjnMT0YdWVDXSRggs51RkbkQDOAiU0TZfjYsIH8lmZq8G
5eBWVhc8nyUMQEhEBOK72LPSiQMKB+zlU5jloJ3U17xVNOY9xD/DzLGuOY/iJBld9C4TAKpPubkB
XSojlybsvJwyE+wbSVc1VIBAtwpbZb6lyWxwGQopA4+m41vDBBsb7sN+74NIn4OEQQk3LBu+G6q8
sNx3gC/2bqZ34wl1r4SmwUep4iKDMqUShVIZhDPt2MOjCpTE+H98Q8LsDcdxkIy0mYMjBXdlAHCl
02rl/36jSo6JHk0qIo7N3nd55K2HPhUdY07ebdWTDJiA/8PSWLkDZ+GgLxj6U6OdJnNakgfquETw
909IHi3ZeTw047FBEQ5zhSWTytT6CMr0fyQYxaU0Dn1gP2zSay9n4F//Tv9HL+4iEvfWUZ9kWbQ/
1sX+XDY8wr9fqnt84wDuj0rA5NuaNq5GSNQQzgFN/hRI5hv1uIr2yUR8b/6Z84SjTEiJ6r6h4Bly
sjYFzawOW/8vNtJ4O3+3Bz1jME2J9vhtzDRVqiO1/Xfa22kuqGkC/Z4Rvu+f5AhyQhfdulqzYaCP
RBnCWGCrctxY9m2zyps+NjrU9PsW0EMt4CwEEMzRPH+hGcACn1OyPwgDSRvboQXgi5nWLC1LZ0Nx
v3fdNzcD9GCTflbOyGARUUtiaZbSOg4zsKp0ii5XLGQuft0qDEv7RaLofw619QfdbO/nAhK96e9C
mIOLWhp7BdenEZp9LHj+ELn5ceENVXU69l2xX9bUxvUGaMQWIjQTKdY24bY6PJSwqXtUCwLvOehu
hnbb7ah+PtmbNge8ss9GJ1TLc128MnPiMJxZdjYeS8vOauFI00mROQwplmEGyZrXwDbILEXSD99U
F1K/5Ij8HdGpwaNJoAL8BY5T5fe0jrPnqkYZ7m1Je2zk43HuaWnqWWo5LMqwOSnIS6J0eOcEAmOk
zhtdud9HWbY2PrSwunegOto2tiZLc0CVXTMLRfwOLR4ETs+l7Kyf0Z5OVf4H/Ll1/NoNTHhbwLgT
ZE8OY2nn2UXnVm41OLStwc/KST9TfBobsisd0T/jgrqxeGC2swUHnlbE+D+ZLtkz5J++yBOHC9QO
/r/0mVN4v2r95qSJVbVX7iaWCERgFSmAjLxSs5GR9Jj4C5zviA3VbX5giys4bYA0wGi9HAQZStqF
9YVVp3219GdXJPEcEYgL0BEg8d+bdWxvveT7/O3hkQTdQvqNd9YNDsQPkqO59ckpDesuKHrRgk3j
mdWe9Pn6BY/7IkLc1N8WOc5DT3VuZ7VXKjOh0myMUJ2SwDrPId37+H/PVxOFMmW0Qb+IVXNxOlX0
slq/GBTVIuumj/ELJXkF6YZuFx9CrcvYhbqnASFPq/Hq4B/V6f/sB+eNNoROhpwwVc94Y9PC9iOz
ek8gxdTFq6IwltaUvAfR2QhAP0pG+VOxXoHP0lhXFgiNilzUh/6MbaDjNOhzf1qeziwA51lLP/0p
aQHXYC9bGUf3vq8JYDoi0ZmMGekIFSMHFsMoYVtFmpVZutgDHlElWwImiydopKZVj1DM2YjQgOnQ
ntZrVpOVI6UJfqkL0cfeRlXI3lO7oJhAjDdjCpwiVddb+th/X0Ke/plfOTqSf5yfNl57MYbFrVgO
qkP9VKBYMaOfgdzdRUe5Xs6icropV48l90AVgWUwfKhsjO1rqwxowDY0lN/Rgf33vDCj6YX3t1wE
yR2/czM5MXdjisaiW9pRdD/4ESoMArt8PbaULKl3BmHKS8ipQ5jjwJDy32YV34VwbO7suOBprSr0
gExqBU4U1zB1Ej8WMyfk48gU3jKCEHyillcPOHWo8VzZ4tFHOVFtvzItDn/EUVCSSH0bl9Oe+Kbp
bOEHaUk4ckdpMpKZmLSkOC4AsZvT3udhuv0qB/s+qZ6JY4Uo5TnqJ2ywZPvLcSuhQh4cm+6v6T9I
P9ixjhvfqKnaqWAJzc50HZ0+Ep4DW4J9+v27C466AGqDoCSudtClKy1bl8TZ90bCD+xwozn0H818
e/bNzsKowY3U06XFCVz5WkaPVoy+8EcoYc6IbOhwxiFKoamjdHcom6iLfPU3rNO+muz+zfssJWv5
gNzJ/s0F8ml2dMZ3DqmLfYIiLDZ9UCvVQ+Ab5g6Xyi2/pju1VH4tjTfQY36QulW7rK3YVA3AEIGN
085OIkLEV6Q9Hq9H2Hj5/+tdfgMdXA4Fqe34xWtAMGypvqWEgDQvOi7D1lCj22szIUoZOMqXY44d
KGazP3uEW0ARc44oP7IiMPvnYhrENIH/u3VHzxT+h2ZZrOyfyrlEnwDrzeFI1XH1osZ44a29NO6g
2mUNyAcR8qJD/vcH7ATg6rZbKbOQpRGXJwMY3Fac5pH6WNM6VI0DdtozancjB8/7lmUXWz0uIibE
5YHkqKJ6+foT4b1a5KDUt2P1vRabYHopl09/0dNYg93U5M1GTsV16qkhWTSArT/k9JxO4aa8e2xH
vk94Six6BYM4G/A6JhVFxYoDVyoUM12CevisCjnbWcafLDWMSHrjddM2syHSqz/Ltoe5uQ5LsNe/
MZEFAGdSgX+/nIGrmN8LoO0mIGw4g5MZLqL6SIcp6OjGE53AhvZgQJbxPz4mxr0HIyg5cegdq2/O
FYgNQh0KHsmIJf3lk2FhbgWYEW9xqAdmgYhg25aijWEgJW9iWWX9sEJY/BYQcMvllZ11J7PVfC0y
1D7lfOQyQRnmfwYYNauuie25SjiWY9ZMMpUreFRQe8m9I4rzHW6eOaNt5XvPC0x+vf1QnQm72WIm
G7/ABY9DIvsx02AoG86mlrMhiX0jfvTOchRKoazl59E3jPun3Yv1un2RP2LHZF7rZb6FrgvR9wmH
1/Tpb1q0P/Au2ZxOLh/3nFII+HJCrIQlfayVhrUbWqxf9rEXXzJUtCLZYBcwmeuIPRpeNE+JRJHx
haqw6OkeG+tBwDiyaBxNGQlvHk0bPTqVkASNNCIioCmtlaVw1ZitIEtDo76uohA8aMdc8DuFi0ZP
f+AW89kR8lfvsO5zSyXg3Sp/C1t6IBUChkmvcveFrj9ErDNdQngRfhWnrFh3Upw/k4N7pOVXNfVs
mUDvzGjT+SxYIw1q1gozOb4leKdAKZn6oXh++tGKxB/a3Q7CxjGpbCrkm2yRSLEQV+dIu2USjt9R
C+M1pncvF+PfFxPPstJ0kdFItLR+Ogt62coB1wKIRV+NRj+0LgiRTU9cHLMWEfeGKOLhlXFABhG4
GQaoC81ZyKuDQWa69eFSupFcM2m4w6pP3DjkR1qSiqGMDsh3H+56AQsWBFNgq5FSJhPDX77DCH2Y
Mj+F0ZIlG8i3AEt/Y/8/MgKCxeAcNSyIbxXzT1cUuf2pg2DGL9zmYOqJZFGIZAjKhF4QOc6XjwIi
BBOlpn7R/CwYuSdPvVSz3VHF9/8cRy/4NwTsde7nyoyiDRGEdw+ZcfeEC0NxWcUIHo6nL6MZGxrp
EKMQl4qoXYYD0NGGleKk9QtRlDh4CvqYrRWwu60VN+T5StOTUyJaMwDfsN0AZvg5YuvkHZlcVeO9
0eXE8ra6yOfYx+O+BXcoYub0T21e8diJlQskyztUsx5+Sald7mjrDK6MQ6bpD8IktpqvwtCmLnvO
h0Ppxl/ANzKeA36SurNtfLVerwO5qnytQGrRjpT7fce3gssdVNhyU4fqAuwZaFMLuoxBA2xcmVqZ
OJo6OY4YG5iOJoK3ocA99Yd4p8g4chvKB3MtShS0DXbDzYvA9Ysi+7qGI+49pYMPx4aff5EHiAr9
m/bbGfJPO6uupZEKQONmWF03/vR6t3NgAjSo5Ah0Oi2d3vg89zZv0lSfvFEdvqo0hWhD+wshPXCj
o7uNysf8NPMZb/1Tpjvn5zN5/9lxmq9IM7nzKl9TSio81uzIs8aeoF2srjhBmqBKjdSUN5DQLIR5
u3xZ5HN3tcMBZfEJeBbMhu32bsA712tO8tA6sM316kco8TC8I3dDj2aFNNl3SXVWWBmgip4YP/m/
vPTEk94PYXy4f+OZUO+jxPVAMIweZvSqu5P4A4KRWC8ZJ3c5UFEMZyrJN1q2EbCrbkuof/iNZK+A
zOMRmaNUU4Fm9hgAHJHmlc5itcPTA5XXHZz1gF54lWFDk2vF2qkv8f30nz7W0+zp46U9FtCwybt5
FOAwjaSRK+xdoXNAwtCp9l2X6bsOqPR9a+KMI0FghacdKe0gE3LIp6HgJWV/vWA3jnJkBJiZ2dM/
GLJSTq1nLvjd+fbWFdGnCIv7jqvtiXJ3OvebQtb37jpmurx+gzdKT1RWP+IasfEtEjaHfz9TrdBY
ttQiMOgDp4Ka7Qhp5xXS+6ObbJ2THt94NIAZg3iL/XvBvfGjVXWrz6fdmgRoxbm3K2YpFl9fHeGk
+MaundmoaMpKmm4ritbl8eRLT3dgiDfjU/kXGbSqGAahiLD3NClhAXujQTAsE9IdzAm8PESyQcGO
LqEx3gf+rGqHOvnEa4L5pNEDQ1pCAZkHhllvkT7bjmZoalR/g+K6TTWV50r321ftUkkggBFNDueQ
lVgvDkljM2m+I/VOKPKGjd/R2qtHFR8aF+5uD2gusi3otp3ca0J0AAbW9Vs6VISAjcHr2wBPdtqy
4SDH8059p4/qZLqAnkeAlqN9Kqfn7MGhGEbhKTeOV3LUehuB2DQObiJQ4iBYBoRGAmliB87t6YYO
rQjtby6BKs+pi47GdzpGR4CGhqIPkJaTjg/fgh08YF4+a++FnNMTEiIg3ScaQUB0OaFL9h2HessX
BTdjrdM5xSxEh5gBVeGiQ52mN04H/f03LY/AIT5X7iQBI54thdhGB0RxdwZ50AclZveoM3mdPYAH
3I9f7wDZvS4x11v1cjZoIOu6QffQB14DuoqYEpQEKPpU1gHNpEufV4EF5wN/gcgczQy1BgrqBSZx
/ho44nRSF0dons3m4Dj385xv1z0H2zwulKfZkOO6BGYcp8VHmZqTbCs90Zs5YMKBN46w6o1E6zJ0
ppvplJu5AsLA4dSYKfE7C7f0+yOOY8XuxA/8zW/ZMXQXtVbTOuAYrfjxYCTPZyAMizz1ROcwS7R/
WAvqF+JL2nimEtlHic3r1Zm6lHIt1tp3lPuYiP8/Dl63PIa+Vj7aM3NuCgUCEVQJYlFs9IvwgD1l
3PBDnkRuAd/k2W9JJ8RtK2G800TCOAnpCv4oLSRGwy5sOUs38UwE8vAHjR/M/SOMo7c5J+CpxJhM
pEZ5hBHsF+t2B8tQ2xKde9ThVQ6ol8nJ+PU/T5Xq8C6bAkMOpkt4AHSLM5AFrGzutkiN8vgDrbTk
suD0/I++kVaasvlU7gcXODRCcFS0b2meWAT+VIkARCN7BTpdx4wTEP1FBsYYfVU4SjzQY4QcFMd1
wXh5jtZZCLGEJrmdp2rwsvvw5C6qkTSvMuoNqBJwdU3zCLE703Ixex13NQ+OUIplx0jisNy1T4Np
j5O00X31xVre0eL8sJImduGCo58j0nhxK2jrNiJxJEQYZryy2iJxFRJxZPr6GZRPCoewr0gGsrTB
4bX8W7v3QNYfDHNAYd2cXW1VQJW3ZA6GG2HZd6gNcP560yhKdHwciA9fAH33a1nH+AJkbpsFc90D
+DyO2ECEH8qew6KFacWOvYOEpYjvCMe8WAeSpeY8dUm56ElFNCVQoq7buxn47axxVd9oE0WP8aYw
hzyuQLOP8Yw/TTC63IokAUSqttoWFtHsny7Yp/Z0mTajVJAlgL9c7Fq+YddHOheA3mCKF3/d0SwD
NMUgDkfAyyT/FI0SiQXTg9O3nSU3Cs172EKMWT5OEaA/WrlizJdMxpPaFTwBoFxjqHCPunTBbMgB
2JgYog2YRQw4MjetLI9hRWp72Gp63Xrp0qbjYI1g5x8fxsqBEbFOdIiTDZWNTFWPl0mECnEMVkXB
/zKWPg1SDpFZ5pKZnJvdWyuEwnYiwne7DvpLNbpNUg0lgKzv7hsebQK9vdmDT/k5+8jYkExrH8lG
vOPpoW5sxOv9CdDeLlE62wRu5ugDc+m9K1jFfEXShYn8q0mZATmkAKfyAJL4WprrLVBl3SmX34Y1
a0Ojs6CHQJ+/o4/9jMObg121ZestmcTWekrTv8UIa24cEmSHSg3W16AcH6tuiQt0NCfexClK4ZhU
Sz/9BBY0IM5Q6OPzXHNbsEMbqt5H40xneBlDXO4TBMKtEnky74MVkqyP0LO9FcrX3cevRjZ2NKIo
/Yhpy7fYZVfVOwvVBylWO0NYrFZqOX0LDBYrDMWuhYsFWEVV/mAADhSpv2G51paNQ0v9Rt7F/Vga
xDkPmSbU5i8W5MwoFRVekJco2iXateQbZ+8a9NKtUnumGM62IEArpIlYRdgc+WOyRX1gEzYuJjqL
Tdi161bgnYV2T48UAq97Ly4nv9bLvzxZI/t5j/YIM9JMFJrl69eUuvep1hxcm1ZAXrvoLxspWh/i
j4OUukg6P+Hx0/Y+k/lBQLJc/RtEovPUYbnyQopx9UPfs5uySEr6B6Otj1sTE9uLXHSw6OcGEQLG
mMCeMaxbWrLx5k8Q+Qaq8172/nNwBARit73Kq6xieAyDCXksZ+v5n3a+hD2FZa+u9/kE/O13n+3x
9Wn3GifU+LSqGLDLlU4+tRU8isRK7YoP0Y+Ucx/UZwFO12NR3MZrO1spbjSm8ZNFUHj3WXId7K//
9jOWXRQBNhHW6UNpd/ZR3dkiTYJwqAd8FsIJo/3bwXkzHYlCMCeDtv56OIHkfKKyFOv5h4IkWro8
C2bGDeO4BMm2ErefJe9AmzLbwDM9g9yTTPn/el3B4Ek2I/vA6+OXfxarIWqDebrklGZa98uZ4L/F
xSnM6hw/g33DbMwCvm3tn1XkgKl63pnEbd4UcJXmFEu/wg32QFJxg+wtT0t2RByFHpPSZx7SlnZr
qEhu1MwuSA/hk0UnRqpBrBqFLjTuEHFB5/p77qU8HKIC3hSvqyWC5+ug+jP6V1O6rgjzLwB0ULLI
dYf7URZIcQsVInEKrL+4wTxctKeFx+dMtLT8j+VC3s577hmCv3c3rpDpa4URKZpFHReF1MKpeB2+
K7yQMO0acd2XoK6RvyYcDn9aGRMpZqbnDLLy1NYVj7LoovIv1tzRPrcOOZOEOYB0RVKB8KTNSj6X
DogHWFZWMDzla0hKcxmdV/isE5Pljl+xQ21JK7jOjMvJQqnjbnrH1rFck30T/z09/bu2soNJxtic
/xixKCiUwPeZ+RiIrAVhgppkh20TCEY1bRQf2N3AYfiSvWlE6mWasSd52pbOqLcVrrsAzdrEnVze
vfPLn9Db4rZNFzo99n0UxBmj8ZClN1jXsagYCOt5g+VNEFiqOSOL4Aqh4HpQrBHLhUk6eWizy8wY
6eK4ecAQ/Dqwx4v1Eg6bYdOSLXbbdeAVfKjhSrvlyKm1pWWToyN0OVy7EwkGExgqLskG1Go9RECM
i4/uzwJA6nYTno9kR1NmoezFYpECxnG3hQUuSD1VNCfJtxooaqiZmgS9yCsZsX+DqTGn/5cjPliR
J7RLBartKc3C72hDWHTHQTJ4mP6hinqevg0orWfpKV8+K09KxmPEFps/Hqmg7VlfwH75l02FqEtY
WjNPQ26m8oC0FunZVi2XfPeEzosfnWB51mmbZAOhh7n9UAmpaQIdC/rU503zhG278tS05BRfpcJG
4lN7TyF1V2DlK7e69442zySjS2sf1Z6JEVc6j3tj+loWxhJ4yP3qaPEmqnc8LZO+9djM7VMk2aNZ
ccpn8qnlRxaizTyymJI9DE4r1bMQm0RY2bA8srlrn8sELGEtaZUIOKKh6h1hUV6vPO+yIZKU++2A
x/Q44DgL6fHs4vYtpZ51zxtUFD+RqnbJvumc2aciiSTdcsyDVcGspZFShCEFwysIGN4V0sqi3mhU
pwJ8UvL6gSvSWmkXtUKwXws1XqIiwCeroP8EQgGdSFBsyN3ectwQgcPTvj2ICMOdQ2DrouO7Shxv
obDZMQvQnh8yCkzhZkKf1pJVkRvCC5AFNtd4Jl75SSE5rHt/ard+oRuQBNcyye0H/xmgqIEEas3D
WL5VBMNnz0fX0gGNetLKfQj5hZ6VsCleRcrl45WG8eu+1baN0+nWKqf4a1xj0lXhsR6wJvoVHHc8
Lhj/rn6+TFhymOxP4sJRCUOK8WkEV7AhBpoPS3zIjGCNIM/eN8fkBia1rhJjyZ+w2V2nKMtLMcUL
gqpMM9XsHz/DBoKEdZHa48cwkFGSAQEgjyvA+NFqaOCdPIk+qPb/CsqfZ31aLDI1ag0ZbBT+Bspq
1QMcTWNmwKPqToa/NIEt+jfdUWYyOjS//Ss2JJ+v/Al01p/2gFoAnCKQ6Hb4OIwb4X980sAyUwbA
FgCOe1vXHu9o+NgEbg+gBFn0bUIA1mxMefO8BaX+Fhd5k8GfKieUfEPwk7ZeMx3LdbJ6WI4ih7iX
jw+X9UWMG7sewLfmO4QUxArFhYmbF3xwqgGRzs1pQzTpggFTDAKjySPWigGawcREbHyCargeq74w
JG3Po/8gFkQf69DI4OtR5Vm6nsrtOfDKK6IFetYnzaiuK7Rd9MURxjgZ8ez+u/OitkU9GdoCaKPY
IbO93PyJ6tdAigwzZKB8VPsQ8Gh9x3hyv22VZ+716UvrsvbzlB147pFjGIbyyTa89kOM8az/rNYd
Bt9IQrol+9jXQv9YBJzfgFhENYcE1MtKnuKuxKivQMkpLkrkYgr/9/AjtQ5krsa3FhMcdxbq4K9A
DV2QnQIngj1ZM6c3SXgexYw5vFQ7/W9fyPXy8IJqyQ45GuQ9BsUTw+e9qripeJ5R/H+sFdDcSVce
3FUZx1JOeFu9gBg3z28KmpcQa7Q9smKrLUNACrS/4olFbucmL99Y3AeZMdqcR7udqN9I9lllyAjx
3k6SPskeZawI9EQJRMSy8YjXsx26/oacrmiwqr5GaiaXPZrlygVc6U7W3WGGa2LTuF8BDPQzAzwT
veQM/9EBg7Kz8Foht5fz3nCL+y96nVTl9vy42bw2SBCuX8BnSbBLl+WLEQx3JS0CmKYPNfRt4wng
495Od+rJWBrgd4ICAUm1BWsuSoJRLkECA1em8HnKxiGeXXICljjFSj/quFUGAYZhc3W/6g5/DmOj
UIJ6g38VUHB+An4dtnqOkIlpK4RzUcoAXv32XfcV8BgpHe/ELrKbyJAZTDfYhKqukrfx/15mPYMy
+oC/LCfE4HSzg7C7dAH2NPkxKymMUVb9gzlcpS3mtmMYvf2KnQe3Ri7jW2mkN+oaynruVF5qQ3vZ
sSW8KAjhHYm8vUGoh6VH+dtjAxxiy9lC+fZGW7r7KRMcdTzhNHSQCVUUZrduJYbhPeA9nnmcHmXj
oJRxRSmjpcdK60VZxJEJURB7A3YWTyo0IrR0sLYrnr644PHyyOnwXcRhtm39vrF0sHnr2grWduX0
Juw4FkIbvoRi0jCPRp0fsr/XrpYeCkBkJL3Zg74YXjbE8NMPCk7nNU4naEP5XqWCpLyRNWwR6Gd2
+ygaN+61peh+DSePBvvf1FkONs7SeL6gUDYLYxtibf9plZHLbVcpbht2t7w0vCCokkqNtDc9zdC7
MtIzfEgr5pJ2ZPe+WXHF+f2CZ7f/6dFX5ZjO4DTeY6szP0jFnToPtn7ESisdZIlMjsbfdA8nkrl4
NZaSZpx1MtG1IBA1U5hrJDNMlfP3jUlXyCevSESak2wTulqSKBuXct7IewT36IlGaduXhBzmJeO2
Vh9HCs0YmkjsaKySq/qB4oxorqZThAGZusC+3F5ds63XHoJA7Nss8uk0w7CinqxboB6qOhPHgdH7
keHJIlWry/J+NsomBFlsfHyfsU9gF0YH8Xp83wSoznrE8xXASQZrYd7rN2YnbuLzz8iHgoyfHUqW
GqWts8n/gyZxH9ruvrS6lEVqwsMkek1keaK5D/dG4m7oSUEe9gP1+t8NliEgW9vTvCHqWXm4e8rc
p1W08xsEasDPz20Px4SsnaQrmngiP1kBtNcXMXQCNOiPPOBbztUr1dCDOpPUzHzHszWyl9PJTqDE
hlC7CWujHLLtFcUGWYs5vwYu9GmG6aHUlzGAmNRvq7bpWvJKTrSx0tAGXRHH26EVCOOwJALykT3x
r0+CVEd2lz2MG3Ey7iiZGkJYI0cXhDfgxaHAT0LI+M3ESq1gkzScWClstRhqWD2neeE3tf30X7t+
jU97mR93GmpvGgvYgoyfbyG4LnoJJ0spHQqT0Wbby5FssznvenS1ImC912AclRo+WzMzBcdwyYDO
Mo+lJhzKaHdyzYdPNzFlu/FHpawSzBFjffLmD9cFpJ5VqZo3MCczu76TaOlUicUwAsX/vA/Yq0dF
SnGCrXri5+Esl7lXb/zjbnHArxIvB6faMOzBeg1h6Qo10zXZCCIA/JYla6BbRvLXTSxbWSl2ZjpM
qj9E1NumfNYQpJQCD12HES4y/wGFwkzXjQqv8zuv+HBDx7bzZSAFv028vMXPnWVq50QZ6KOeGV+q
jAfG/W15UCW117/kppsChZ4qJIG1jougvfuzo6jGF1i0anhh01lxLw/HLEXl4A51iIrsEy4ATjea
4UOVtYhTDqrUXnnBWWT1MiJrqTSQcx7BG7EFO9qvZma4HM2ngXxrU0ARwdh83OGE3TTJKW1fjyNe
NcgFcZtgGbzu9oku3UAVrFLE/qKXSJYHE6qTUJoAcmcgvfIA2hY0A0jqCy9he09Spj+q3zz37OQw
zivTrB7kxvrBJvf4hnmMiaCXSh4xM1ON8n0jQpa2Hbr54w+uRjIoEiMUspEbU21e08wVOhsGg7I1
VTltK2j36nukOxQ2KkX2QX5OEWoYv+vRYyJYaFFBBlsqhLPEy2SEUGizLcSX2toFVIysrzR5rsE1
btqjgdApuB6nF7cN1lYYjFakMfCwNfhuHnNYmZ+SMZ3hgSr8KE/NpqbSXiVd1oomH6VAg37yovuD
IZiAY+ADoP5g/S6P4JXR3KPfMUnfcRGl5acCGZfcbHZUDxpE6xIlVGYy2+miONJ9EbuZCrruk2GL
7udUXARL0oY+KW/Re2HsXAHBPihCh3NnraLTysI9BsWEtQwJXTO/TcwQtEtXqo+g7etFMeygNZTJ
RQ==
`protect end_protected
