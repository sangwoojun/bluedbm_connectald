`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TBx8e4baXZaeSZSFCIO1Sb0+aDuKp2/MUi8BltcYoRGvNKUGl8aVVuEOAPjtujA8+Gdkyl4NBXhB
UPJJ0pkRkA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
O8dD0PdugNMcpy8LpOPVQdZ5kI+QpDhx689zSk9XVBsxh3EDssGgi4d59GnTsB1kY2c4cHC2Iq0s
7VsTCCGQAxJtedNWVuYVnUFa5XaHncAbkev4pluaRAi4qr2dxYx6WUIXxjaR5Z+5R/ejNrEq0LBK
oadAJ26kA3zaJi92hSE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KNvGy0ncjIEwan6o/WJAx84Xr7vmnV/wpPcZEhXoTxM0b8eEdi0UnKG/n1zzjwxoAdP78A/mKCpV
SbNn7I/10Z9ENpas+Lrsm7JagiV0+kZEBWq6htSEhkAY51AUL/wGsJSc4In8ec/50Xtb6C5SpuJ9
3HVWVVBz9e4LjBCCHldKrePHpEkRanVfsgxodJ4X2/b6HUFy/08ejAqpAW8tYxz+fE5JZpogUV9z
lpn3YWod/+1b3rk7Phgavz4trRGSa0DKA6SXA11yKo1dXVW5j3N5SZsMzGzXkL34BeVgXR74H0bi
dXB7bp+3d9FZXv7ZJUCFlec2BxuNMJa3Z1g9XA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ztA2K2xemdfgqC78C27PeSMrMBxcfh8lDciXtedT6ICmhicyvCEmaJlU0KsPmQCiqZRlDMteNW4R
wD501TilA5Et5mEOD4tclX/xTuizKFKDksqrtZ1WBdeKW4DAXJqojGJpga+qcSdwoT1Zne3OzWnu
vAGd2tLnseQnpQSrcpk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GZYmEutPkA2XDyFhv5Z30eQ/TDtmDLoI2HsI6/bt5y7ztcMXuQB8d26bJ6n8hhOL+j+yRVkxQULv
nH1dtEEZUyH0lEJn2Tgb/oSgTrLItQMA/Xn2K4/7kMZOZajo2fxnScJUThdLGnOLtXtN1aFRRpvj
7cJEIN8bIyaJBavPEtabhgzyHgzlxTAc/hXlCMu0uw9g6gKKHvkARnCzQU1aAxR9ZG0ydha42yzD
eti9Gj8bFzMqXH57xu2DGzzDbS/4Y9ciMt7yAI++Udm7FqtdOkLDHI9P520o2ZWnCLGj4IZL5EQT
1Trbg1nKsjm5mZJf0MV3qyeLCOtUOix0J11/WQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22384)
`protect data_block
zqeBd0f2abJBkcUA2mtN7cXteNQ9zkm8/TuTq7FNeQYDLmEbOTO83n9ExbZJGJAxXDfs6i1eHXpe
3LXDWhfPFKBRI/7eXiveulooigeb0aJGyiFBNP4tNeRXgyYJOyPMac5P8mc1olBTiVHZmHxCR4+y
UX/ugZ6SpA3/lB8Y+KBy6DYDFSPYQbLmuYmXr3dpwrmMLoPG5VefXEy3HnYPtXH67UxwsVDEntEB
6Izg6qUoxLUh4+9bpbjNR7wwd8PgL69jqkAwOkI6vWvNfOLXyZ6HL/0Oks59oO1UeGQHZ6xowMmo
/9EYOm3E7jxePJPlS/EuV8Anje9DZ2rke7yD4HBYIpQ3rMFF+T/PW9GXpnJAarKNZGv215sFL5ny
j5eYEJIy9qA4vF8KokuvecEcHxPHKsUYGC5IMulBoXAFpdKoqS05nvuEvR2pTK9jFbSdcZlT/CGZ
gsfBXUMqXin1EKmW3iOrZiJ9KPpYE3CCZLSq6uatE1nd+ex+pzjC2CwZ0RA8TVkTBD9xqspfBwbC
+jJKaAvFlCZ+Cngt4TLtUwSNey61X/C5V/Z7iXDnav/HF93vdbaX9naVkWCTKgtRHwLRCptlERWf
WB/CHnElVwX211ETZ9BpKk18uJ3xlX0xwqrgm24zdyrCaSQ9wcsm2tZOjUf9Kvo/cYnwq8Ti7tZa
B2QjixGNwrAXXmd45wRWdPCATzq/Od5RszppvuChbM5pXmrFyZskSXNoBKIUPC2u6SNruwM3KRbQ
Luc8Newid+iRTWVNxz6/FoLjfm5DlF+tpbBSpaCreYSKfwAIiZYX65hqoofrnVkWJQKAn+6Z5yqs
fqYS7BkbE8jju6pBxecbI/0tfCj2lQLV7YwW/ATnk8s9Y7GASbGyPpQ2llwW/1PDu85hAGWhshb5
3eq9bGHMmWAQz4DcvkPp5SacdeNY5FxCaLJZrTW+bIRiiFyXG0j2SxYluyum8VbP5m0S0evbMBuT
7XR8w2PLELR4Yfeve3g9YENY4U3ayuMEv5P5Rj8k3Gaa2jGPQMf8z5PUUSPIMR3JOVsVEpmNzJ57
OuSicCGGMncPj0EFMlDYoNKebLP5Xac6VGwQTMK7H0gYTEEQr/8HVXnTgsEGRDDV81VaiseOLwfT
iUzVlywNX511benP4dIF7b5o1p9ZYT517sKzcAD7iW4Zms15IcKi/YUBJWp8CLcSqkYsIP9mCMir
L/m8K3okNGPf8/XGjSsbLdOGbVifhyMU+thIsAz+QwSER7Wt2B/qUguyNM7cOD+4KhHyLCZjDteW
DmdXI2Ls6qCVL/B6XelA8ZIDgc9C76nHSvMO9zsHKkeQd80jwnTuuzfff+6/BsGmRWNBfpTn5G0P
5Nd+RG4fYDzK9CX+UYTLnxMGGdB1/zK0tZRaQrsa0c0hDyhn9AFzaW7zikv8Z+HfuilQwXdC2Jwq
S9Y7l7y7G9WYgRBvOcVLkntvevO9FJwp5kcCYKhhN1Bp0HsFJJY1z7So1aJg7w5VM5lAmKF9pmH5
S4/74zKy+4FySBgKuC8m/foqeqNXGRTxH2a6DszhDya7N9HTSXz8RiR5usk4fY3uXC3WSgDwM14r
AyDs32ZkKzqVSnC1b6viX+EFMKEW4XQPLUrVpv73sdBD2cP93449g5WEmcdCLOrWzhN1hrkTcC9G
M4KLPbPtXuDvhBoTZL3iLbDtCk4noKYlIUYVzLCa181dGZAvQay7zDeHvh8RFshR9a+JZIrCT8tY
5D1bOmJfKffMN96UwCg0PHhwPJKrYrfKFGaC/MTtgRi0gER6RKSn3D34D0mdfGhiUSE3jTs06Gn6
nA5/9f6JXbhEj/qSyYIXY3HlyETb0ANRmJ41O+T8iW2ESL6vde4rSsDEkxV+/g/VWwoD41GJ941k
RrGbnPyhpwggw5VTO1R9kEjW9VTdAq6Wi3IlL/p+sqTrMZOA8CX6Ve1lmh93ktmFrcYG9beHepN+
Xeqy39h6Yh7qYlDbnF1QV358CT/J91zAEwEEImieNRcIYTG2ztc5b4x40oT2H4BUMTkbD/iqgUrV
3BgTvyJsxh3En+5yiSNd4aQ0a8j2tsQASEt1vI5oYlHkV/urIZeKFam8tXuUm1tNpDBASXMQbwDC
TF6xoRIbLd5LdSUA1IDCW6O5ddjK7UUShoftVeNNrMPsRrcFyMgkEZoh2vsnwBNS/DZnJydOVF+e
AaNTatjRkUOdZNsynZjciK/3eFIQIownz6JfFao4aVuyGXXPVQE6XDlp3b7lE2B5Y95zqGm0rP6v
RulGHttQGAgyU0yHqQfxODMNJQsOvkQ1U5WCjjuB5wPMYUexIToaW59Ov955Es/bFdYs2SFPmBFH
4qebE5V7bYrNYwSMcMR5hp/HR4qMGGOpLdXP7RVncmvYKZuTairtIsahgsSowb6MW1gyzW6J/Q2t
ZXCDtAxyLkv7uhJ/Gi5bE/6EoqdBfJ19PbWu97R6+bvjo7QI4NCGMFZKCuoTClUyZvwVkdfvOXcE
+MQORZ3MyTzB5JWBHqj7XCp4nVGkAX8IC4I4P6irzOIHHVs4uH53ganmaUrB2rswMJRUjlaqNcTw
0lOQQ85F18Ir/Ys9NIzhvQp+6b6YTysc6Bld2bfaXbJSVWKqE8yBVOufwRwigmFa6liUF3IbtEOA
7w5hHFxqERu275Uc29tdW2Q1EhuZ56FUY+cbsKrSHUEnwLdeNUb+a5+RtwAxXszb30nF4v9zWzkB
LDE0uVr6iNiM5QWl8Ytgw5p87IpHbvpishmMJg2vVBMP4dojiR9X1v/jbEfS+jAeO/fgbl7f+3uW
GmNPH0dBE2dtd5sAfnUIOu4wrEfJwfWekkXTZz3dAPjPvotXS5W+faEaJ59pWnqs70WyGUShKZ93
J4Ha65fLZLqAVivoVWeTDBMD7ORlLu7lYcSZWdZk4fp4FTaLI+YkHoUzG7d4DUd62QV3wH8o9ReF
SmiS87lXmxc02RS/D132fzJPr3Phd0bSs9zIo01hrsF4B2XboulkFDDkeBeJaXkGt0NCQlqVU4WK
T5wDobU1DEBFS4vdBBob6RvlAxkiIJRfjjLBDKn12XJVbBpt1/hcPMeqEdgEhP2EJuhXzlhRdlzZ
ixWOknOyRF5MmyIg9fVNvTt9rfdNjfYGpuY2NWKCelzmp/V7IzHl4sPO8UlYticgh9xrcgIpNcEe
KoSAtlIyXR1UdQJWb7i4P8k1wKyrMc8g8GH+/8KkaUPrUFz2sW/3q4HIY5fLGCzj5IlhApzZaoqL
Hw3ZauDWi5awYmCXjmhinTgwwkU+X4IvhdK6mN8zuaK6neK4WrvxREFYCZabE+s2Scf06Z6uyn5g
1YkhPxD3QTEFeguHnQO6EGDBQBuRAyX6ZEHcRrDe5q8lqBnIqKnK6bRTPV828gxdz/6Il1ngaLJt
DgPSWGaB4fHvNj0wu5SbWJ7jhoRKiFTZjcTrljhwtLVY/ztEiFEZvZd0a3V5MQhU8LIL7KzL7vn6
Yk9Baaci+NCH/2PgabuwYZ7c6JtTRRtV2THVHlM88ZAlizG1YTrBZZR6fFEScgDLVk6W0kr7+dvU
p56UFz/C7z0M1OXL1UKGaEivEK/ZmkfJa+0I/4ZM37UtixLmnAbx+k23tFAECoRnTaL7mKUmG4Z9
7ehzl6KOBvZUa7++dqyiCA+yVoZeLCNHhwahs52expQszQTuvGW80ZxLQdNrGK9Hp4q6DwVVHvyq
mNHG6Dv+Kz1iqdOWCLnygH/us0VnYbbTA1w9GGz6PrQ7ExpXBbmt+fsJYoNb6VW0P7dn7VYJEDWf
sZ+wJTEofxj6KHEZ/UlDN+H99cf315Zu7FBwx/ZKQbh1jRxBia9mwahbtRuJKOTPVU/BAAalxZqM
q3aYBHGYnz30kKVjwoAZ/6OcP+npzuHp+TNjuzYpWcAkc0HhWWxEef2xEWcivt200B/qg+Ju78ld
FmZ4GjYycm243mZ6ul8VDQ2gZ7UWikXrXGr/mwNz9tlUvensongxQ5PqCODaqb/WRj+zbfa4qo8M
G/NddZaCL4p3Zy7iVSyuw4IEvIuKDjF46Oh8fNySj452owgf+m8cCqO3ijl0k06BwlyTvPcc1WQ4
1280AXa3aFdd0SEHJgzraUrqoorUQgH9PSoS4W6ypk4FFXspNihcGl5eiTaW2NQu0T3bZorsBIRM
yqjbYsNApfB5fQYBFVkIvzQQaLMvEzH733rI5BhzRaE9ZYl91oS4b0FxrxFIDHV295TdJ7xpCaRW
R/Ea5KnsTgXIKXbn/4uJSkpAvcWUh8XJkMupCHC5Y5HQ3Dk649IuxIT0m58FUccbC9PT0GKqldRG
TQN/Jn17WE5zn0xlPPZygGMF/78Gc25F7lu8gRcUZ0MymwWaTQfibb3IOB+qPXpU/LRNAIEJItnw
6tqvTzkKcylAX3kWXVH457AgZwl4NRMN9ZbKp5YBZreStjvht4hnywK9+VO5ngUGXmZk3gx1Bz03
Os9w85AGnt3D0DsC7p7Nv3CGSHFS+IIcT/El8V3L6kV3+pIUi3Gd+a/vaPw8sjblE5DFqpDg9emX
Qs6bAHwPzmqfhz8kW0gzNEkNMc23DTuQkHosami/VkJQNCFPyquV99dNlYFgZmvxsXPEDQ3TOKjw
KhL3v6v8S4sV+jBK8DpudRdPboo+0+eCBdrhiXV41C4qKsbCbPkk3aWVbdteG9uHzsHI78i4YvPt
846dax5VD22531vjjpi5tD2CyJib/UZGj+6EXSNFJ5uLRbLPqQDf//kwwyqy8ilCzvY8CDcavk9s
2UXeWpvZE8KHoun7WkIsLSqDGQDwJ+fecYWOPpigTdhGePzAFBrhJlR865oIlSsi+I+3kstPhKDa
ySRj1E7KrcBxaoYUK0MNWL8kaGJIMgHTovKQqNMF7x+qjOEAzxZsqlM8IOJ2cWS4vXiGJnZhIF/S
9/2qy1tIOhLAg5m1SZYeCfLIlDI5ntOD06wKLfwMgH12V5oS0brcPUatXsQVMwbHUC03+89CQtaS
wESq87j8yi2me/87coFee4a8JbUb//RdjFypS7niru9vOpeqi7ByiuzdcUeuk6UaYTveqwAlX7vS
ff9Gn/GZhMLx3GP9Dhj3dRyx3V4mlRgZJKVsHtA93zpHSpxgDnJOsXUNyyQxf7Hs8uYQHPYqyHny
v4TU+waHlTkdnOPrEUT4Hqx77SopWwBNL21ETYrC5PpJimtdgePnPSqtoZCTt1GTarVRu8nmYL2r
DiZRKBwy+zLCjQlMWgXnSxZJ/6sjPw2dcrzf4gg+0t3iyXWA156CS1FTmetLPHbKKSYokggIqBno
W0xtW9ptfVMMZ+eLPvMf8OIvaefiHNK0Skg5JGTXdEG/QX8Ew4eGDeOLzFMQ4k/NP2YeHLqs7kWx
IP6h8Xc0a4LLZOgwKpDWsNFdWKZNRwUY7ZT79Q2K8KRsgElF8t18mDa9Wd5hxMu03QLqK5dONOHH
ycBgGKfMrHoqpedsS9pSUW4tZiKmRTYKMDOABIMZkRnh8hD+HrgPjL7s9mUPhytgHYxZXds2El+5
XvsFpAR8v5t3prgEz+DPAzha9/gEgI5nW8UJovLL6sZxf02+k6dBGmx9ghGcxqFDPIXvsn7idpTQ
Fvx5mFJx3G8xrzp21XrdnrcXPx4KHcHVSStQ8BRNXPVlGYvyFd4qhpb0lLnUq3QTm9fn66Fnclu1
XhBF5Zl/chC21//CdsgVyWtIOZJEZXPjPPzgv/ojr92UBh4tid8fNBdJVhGhlpz88Tz2/s+CIGPQ
ilghQIfRmSlQXrvPRP+DT+VcJ58CB2wTT4FysXuP823IZbNKcMUSgp1h9DvGARdDaIihZthDa/uC
QVA/oAQB+cNi0/+X3tmBmGwVKD6xPHUjWWyJ6aakXefAzEupi6lgpKuJ9iT1yvWmEGyXf+mi66qt
WP82LVQufqMjl5PYus4CY5PjOlhvXhKSzEFA2lKb3Ulhkfthxh5s3bWhH1YnxKYgh0IeOC/XQkck
H/a/oi6ilnqzO5YxJ6s3AJ16ZmHwr0VhGHsRlNbCkkmzYbS4qGS9FmoEWGJTqOsxuINsiaXCz5m9
kSKOmXTQHPhYz1uT8yiViOaNBuE5CejONTyiEaxb+Ouc5ZZF+LmKJsbWS1KeO6Ms1MnLmp1THZ7t
bc/Dc0joCNt38OXCFYuX5npC4mc3cEZ9TSyv1REbjPDXYQQpDVCVtdBba06Z1ywBf2N5P4gTXcMu
pKDAHCfPLdtq6wQk0/6WdjBNFmsLbRZiK5/qjKneWEdgQEkEMiTKm+EpCCWhPKAwTRUUO8xNmzhn
frU/zuk2iciUnXPzNDfRd2axcPlN7Kbo2phQ6x0RmN8ewPjJ2uwvtrmXa4EcMgUaCk4UN1qaznWJ
Z8BiKw+ILlv5BmPuHYEKtBhr8XM9p+nX3cEAXTuKqexcBcTvAYqinNNVeZosfSeDmIkQSIG7twdC
AHTYKXCJKvwwm84Ep4J40XhcVUDxv5MKPd4fBoaCvwgK99QwlJUddRKQEGXaPyEGbBno0aLIcR71
BAbzh3EVIP3fgfzCiIbWL1QmXqw27B1uslItVQei6FFyy9MAk5cb3ApgGoMi4XPJqpLeGevo4DpX
YAVpp1ma0iiWogEi5HJX3bYPS0SPRfymNNkDWaZibyuIHDQouvZWIonJk7kbyKcvI+CoFdtGVZGP
swR3zbtiBInintmmz/etVmSlw0GJkkyzf60uUM1Js45/ffU3X1mYSn/2MysAnkpRzU6bbZr1J+TP
jvZvOkxsu5AVwsYJdYFl4esQ73+Pw46iFvMPqXGrGqO8/4oymqS7pdpD9Ws0mbuyWnwiopx6L1vP
dFJQfw0fZOG9TGhNPrXAZMuZuYglpgkqUa4IUyKaw7rAIKzEuq+AuvYki2ZKbjDdg1M48u375+0k
hHReQ5iQhFLc+v1FFfIYWLloQi/d7nNcY6G3JuLnqaS6K3LnT/x307cdxC6hPcptAUScfnxzFX7D
zAUAiYTbCNrGDDZVWaNWc7neyDdC1jhkMN4xmVmYl2keTVu+1Z3knRSlPUjtE0gIoAakE5IMoqvA
hIVPk85yaGgeh4L1CAFd/Fqq8pKM04+nlZrJ8juv2RajXxj6k8IL8UY1ykTbePrtU84MvZ2tovNO
TCT3pYIgImUKTIRQ9QbFqwoGJhm9P1Gt5etdonSeU9vQ3fyCnvy52vEhiQjDUrD8Ob6IIXTsMqIZ
ZryqKPFYJoA6x6y8Lyn8iq25RU5jZ/13sw2a94sWmDJ57xyA447yIFv0XAhhbKSC4repxqZm3Aih
qqEPmXYAOBZ//XWNb5XZ9FNZ3+9Gn6O6ufvxbu2JGSSkadoZ2LcigluLaN2Ow4Agjnf8L4Uvht4t
6hswIRgHn/H3QIM2J+d+/0pRB/vn9AmcM4Rv/TwtlBh01yuACIB+8/jyHj0Bi8EVrgnjvKIUe9n1
uFJD6Q9C53CAy51gO3cD3xw9eYv7OIGUzEBb8oHqr7Rz34eYBXFBPLWL5WI6kINq00BbG8jbeqwE
7CbQG/a86LLLH4TuzyL7hEgLXX3jmC3iCoNzRX/GQCnowvoXrAEi7RfUTuvVksuiuSvLMnyDZiXz
nWE44mRYizTXYxgycO1H3jLxPfVW4D2U+spG9AqhywtLRYybCXz56q6dDA+PqsnASbUUO32Er5h5
TDYspLWUet8XaP2eQUo6au1tu3WYA65G1HHimFxro4nOc1IZV3JBG+k1a/NAYOgUzW9Sc/N99TFZ
ESmagOvSN/BI/KWNwnNIqJ6iJdxrh7/0tGre9a2rTOvZbEcs+RZ/Rf9UBB1es04+WaAHj0M04ZHw
ceYQpkWbkT0i0TmRokTzvTeOz0Q+1R8gzRfrhQeR8lTNW+YmGohvHmwgbKxhr8zZAnASvVTpcFiz
41RhPj0YiE5lMXbOCf1s71fKF1YIxOnxp0MRtNyCKmHTHV1/Tg/2S9oroRk1rkvt2jmkEyktP4fO
mrfZpY2yHCmR2duRmzTLgLhKSVHVLQNgx/Hg/iJ0nl43ShxQp41MipTPCKBQPX+dsH5lw42yQKXe
JCSCxMILjvuZtSJGanYfRCrm8pczjAApw6/YXU1Upi8bALkkzXC0or+TWnBpvtigZ9R0UyDodid5
LqdFQKbeJ7MUF8qvR8agXMsS6s1YVUSVSeKD03EzOxfkEa2FlYKGq2fkzkm1VT8MWQVCBS7P/r4d
c4MxWPKPvqy+/wBDyTDzzs0ZirtPFMNNqid9uDLMkdUXKqYw8s0ZjLx6CgFnTwqMHKcX1gK1rZGL
jnKMBdfVL91LEyW4eqt150NCsFB9FBRNOQo8tAl/UWElTN3BlTOHMsYLjtzAHfboVCDKTKeVr/IF
xrApHUkPoTbCKhMeom9jvbLxZYnQ8j2UHYK5MTl2dYx7Qozpib5izR/mF0WsRc47TWm0K6oTRplV
6ukwzEnxzvx0J/JxdAG64jB4RL1rT/AWMPhf486gKJUGqS6jHBU9Rnu2qhj3rn6swq/XXQPBz6RG
e+bDDg5dPKXjrf/UlTKV2XMnTdGkkn/nPEMuufvSgGXTtRTOrgBWL0fB61SNR6hhi6buiqIUCmT8
I+yPPZ2lAn0rLO9pNLYwifC/BgfPeS2qE0n1xcDAuv25r7go6CVpWstwsT2SD1ZJSs4NjullTfAc
YYP3dbe/6IgSA3jlzEPB4ZbJqqB0aMu8i17abyskbPM5AXWy1Te9y9ImIDPF5Xps7EFPNabBKy9N
6oJ+XmbF2a19c71PYuJLeBlxQaDFP14tLgpPlYGeA/vGAujB4HZUYjzRXJK/J8DmS1+Ni0e5T9Ix
lnifcIYYduWzpYLIDbvZa/EXxw02ZsNJt1vCscD0DzpsNRAvSt6IAhbcm0TCxlP5RiV91THa5DtR
foSxo+zAeRzB2pWrtZ41Xx5nkRqORYZo41kEHi2PM68P89yMu/IdwEEiw+rn14v/1XWQ/0rksSGb
bA6CTQ4K6R38J4piBGKbI9CVyewVoDVPgSzMt0Ud7ditTpBA9peH9hOTmYElJ6w4LK6oZ9iSmZF3
YCIxqvw9AseQdF7rWs31FN0OXwRlpGMTE1LCJLfaUTFJ+p3yV71YWFcsyEyhqxrvlIlwfkvTbeYX
37uxjEY2J/op6jew6nQGbQXYE6N2CHLoxNfP11PtNQrlCwtsjtYXM/bRtATMeJoy54vZWGoxzGsC
XrPuPT7R1HVjb7t//iD8HvufnImAJUhIUksvNh7in143hjIusfENP3VuqVdptlnksiYgQSEcNhhE
Cw1d/C4vBh7NtXOsjQ/5SWyjCCGdJDJq39q/hC7v1g1NzXf0lcu4frSQTE4A2reZu0B+5+5vRBTw
Av0VVfkwvQ4tbs4SEx+d9dY1f3bxOqvgWK7hmi28KMIef9FcwlvUebBFMmAW8I0ewfAUL4hpQjBO
2EnNs61xdpC3tBQQiTGJbi3GDBSEjl/Ahrzip4Th9QFfgadrWN9YDaRRBVHy2m9J3+glEXI2vuuQ
LqW7PKOQDFVPGV37entzH042f0nYg6uZvn+1g9wEzka7w09VwCSiYTwKoLIlNV4nzINnnTYe6gHP
ogs6C40cdDHTH8Fef8CyIqy2j+eehwILmEasB6Jqgk+5ODiF2wwxcxNtdL1YS1IHmeIuLc28yG9X
iEmVkxl5wjW87k92DfBfYzzslnPNJwjmtDkbc+JtWeuJJDsGzTHEToXQQ1+zqiEk/u/5ax5Is0VS
hgvTaS4MzQDy8SvC5EypxSDas7hw7vNufE45IwQx57XpPhWSiyYD7JEEZqg2ucry8sf+I5Tab15P
vBwX4wVJJSux7daTLmQONCkusgQFI7ReFI70fCvZCk5eFf9sXYp53ksZ5sZamd2XOHEq6LOB7VyS
h9iMgzk/EpePwSf2DKIQEdNXzcIOiOp5q7gxKEQyRCdHBzY7VjH643vJfG/A4Ka3qCF/Lfq8EF0+
46PPd4idHTGJ4dZFnkiluG6HJJJFZ/Q93vhwVuAaU+qRpevE5ngUTADe2JIy6gyn/YybhwtnuAWp
wDCDtMyQBlhYjXdWFrTYEQES+emlGVq0Vj7okgi+gIynvLEHAjtPQEuDbZk/mtuyZpP5wDw+qa+s
05eS2xRvPyovBausk7WjEY2QjgSjMHLlgtBi8qTl1FDvMT4p7bHNArZzdCYJK4FLbH4nSyWDNuaG
BztMmWnRCwf2sZBfgDcRGRC0eAaB72fUPeSiPr0y972vpx3J2sEisiC9aeHSJT3qD14E5640MPj5
n66IH4oHMOu/PuEdyKQVWst5QM4edreyb2r+Ze9kn5T0MDiUVMTUU+5RXfxyrAewKVLovimR5jPl
onDDc2ZBWRId1yoC3UxEWeF14Qsa8ZOH5mqWcLdVF4Ye+ezlaQd/BQTCOX/Rf488cvpkPQqCyoSv
grBpR3Qb34rOMcIcaQ6sKAChGoKe9mU0ON40fNoR2Hc3VXosai/JwPkMauzVJmwkbtSgJ6txFSMg
rAEkliO6QEVtSSPPekPrDtnMAo1Cw7ZGeFH+uCCQ++vxciyXw1aQGUrdZoe67gML1TNrerRAyyB3
7Lm9P56x++8978/Ly3XjTu5XKk9D4zKmEzgcRsD7/0y8g+9mkA2jb0YsVAbeXxKPc+0j3IcmxD1o
Cig7kJIdv0jQeeJ8HAlZStxn31hHxcn78XzUTmLPTcMT7cQN4ZWQDZ2xzO0gNK2yIauNaVwcY2v8
Wm8aL8tTi7WvJElaMflqhIFBEcdZcZBjdnDxjg7BAVF382bFHXpshxqlcB/maXR5YQNvqiH2IDVS
nIGmNb7AUOhj55Z1nsF5cp2GV+zJLn8UxI8qq4AvAsVOZleFPHHuMq3M3g3lNbM0s84LNbIonxyR
fpu66nx+pgD88dgF2ZO8o71PU9kkJEI78Xq6/aX/9bSHSZ20qrOSjjoGOrDW0QxI3z9sv9XrgNkE
viAPINJ9r2RyOrrU1/I5RGT41EP6Lc8cgkH2B2mCqea/CoMBhWo3eEr/WyKeCY3TNzs4K3BSjQUL
7F8RzXfolOoorAfrttOpex52BHeb1kBEICQy1dtsQT/Z6qfmiiw5kSKKW6YleJqnhp8WD0uGkGv4
VI4dBlOli+qMO9pJhDJi1t0WPDb4xE4Gdnu7oIoLllmRPcsl+V7hgFHkIxvUYdBvhZlD8EihWaa7
0Q7IfbdGoEv/20jfuwmmkaacTF9xfD//g7KGDhV6CZwcg0PK4jIIncjdVALcphpfTxaW7fnMDRWr
3VyTdP/ipoEwoHReWjuFvJo/75RXgXokytlvBrgdhL2dy9f+ym13b2Cb5YD3Mzw2a78TV8QZX6bH
D4IEoVeE6fk82Lm1HbIBQEtDUNKW9Z0oAq5kN+OFEN/dRSgGzyg/J58e0mcM9JhLjPrOx8udos//
la5p7ECofAJ74ObTduytkcqyVqLBEQ9Sl+GRwZC2h5m+2KwKquEb0NttW8I1mmfwQZqZxIQdI0Dk
GYIgGw31Q757kQwYr8WzrtLTePHjANs6FUTS+Xs2bduRQljgzrFnDGTfIzaGcw0qnRwnL5tIin5g
IyquyryVB4pNL8pXxOxYzwYQYPFzOxZhHppm1LYB/f2C7rrMYHOhn1REPrn51OQhNZ2VsYyOUogY
snekSA0UDeIsRujjk3hrIyvNc4hnt2oi2T9jMOgN7JKHohnHzeGI32ulUeWTDSVeGaAqfNFk8a9r
c3ukIz3GAsi6N09j0bHDNBMgE7b3BL+0cXPe4G9mil0CfpTxpc1ksVfRYZqWAIwk8bwGMDxVig/V
2qO2BUygEOYutzSEYtxs2Sxoe1cqSsZGXgXaioSzJymY1CFed5HeDNgCnpU3p/JAPo5Fk+2K9jsk
zqyY+75qk3rnWndmPLZS/IWQJETRl/hLwmSTNzs5BxznaJBnZLObXVC6miyD7VVeC64eaPB6Isc4
11++BAVfnBY+2JQbOjAl9jvlxkXMyws2F79PQ/mToUeZo5JnlhdmWzczt7Jdm3mvs+O7/pPIARxx
aPEf8+KOD3UYvOWzAkYO7JOILS2g+dhQbQSBHCzNNwJgh04EwogQdyXEUc7RvIdoYGIvmapZRwGm
Hv7bhlIAfxZmy10hG9DOL8u9ZcstSY8kP1kj5HqBKZk8Ce8NdN6nnU4p7ruMEkLgjkGuH3dWK+UR
/FESMqheMADfD9jsRtagcvMD55bzaCp4AVDcF6eOUraP8XmaPnrFESqxpFqDzbAF/pOcWa/GF+/g
j4xY0v5+FBh3Ogo3ys9ULmcYYiRc57xKi8j3xuPRMS3XFvD5F73hdXMD0wMjSZkHEqymCrjuPIiz
TJQ+2kB8r+55v29J3yi7ZamQiA/2BRkXYOGXOiim2LH947+JlqRkv6oz4mAapD0w1lUz0cCeJxrC
oe8uHpfrBsdfQK5Tvh2fwZ7DJ7U9rgBs7gUeBXrHdFdJDFmMWcKEhgvzHi+7+BM4ciNME4iHGz+v
cBSp9Jd4CEHBU9XNiC+rGXZJGb93GhRoM+0RVa+pOZ2PykvUSY5clDj5/orEBd7T69pRjoSyho71
O3AX075NM2TWSg/qmK6USnUHhe6TIVVmyjDpccZhM+BrWQh1q/PoK9X9sw4+ayWFlvJjLjS+1TfM
BrDCiEFupWcaY+WIYcpBkc2SeLlHbJVtlTHdST0Yf98QioXD5ZUkuMsTERuqz1aGneADTRVcQTgA
j0BI1N6Mibh1Nc5427eFPYBYUC6cAAGTd/wjjdQKvyD9VhyVbCp/MdQx9JbmFiONB3bXlc8pOXEz
fXBDONcUYS7G8kxSBw+VTZCQTQkECSP18fkX1IInIY9eyZWY9h5z4MZPOFn6pgQDPE9AbTgBq7Zs
/xnYqZvnJWDNOD/GBpA2EpYUa4YgDMyHk0Ubt7mehkHUn4g46a+4KIFhv8eL9sYfxk7FRt2Yt3yd
HtYw2al2fS7l6ddL9PCQ6jaeVJjfozb2DiTRspgKBiVSyvLue8dqM9GEkvxa7xTvZJxQz+FL8SBe
nmzK9zaiNTwNPL8at8KgMjpRpp6OfaSUKLG0Zj/h7LpLz8Qk9AlL6RSBk7VdwqaHU21rBujCGJP7
18P1/TJpOlRVruvERBKqaDGflSiZaGQG/6oKn77nLZNqp+xTCSVwWZ6dUnefApT7lz5wJ9nglA4Y
vVXziw1YLDzz+N2ExeyDj0np5ELrB+kJxPChmA/z1WasTX4zAORPIN8P4RthEN6XCVuy4z1y6nk8
lIxC+XgxWVoFOSARGlkKAMenklUUNdefH78biAflYH56akSkBHyJPZgkMVf+T5rrxNDbHKS6KJGP
drI7Scr3D/8wI1iPnMl7rJSfmGSNwJ8DFg6E7a+M63b0VeDykVRPQeXY/U/b+jY5/5k9k01TJUhy
5/DkdmQahfJlUIjMuhwX9/ScTnXY4Z5Z6CnEfeqTRkMJP45EJ+C8X0ocBC0rFyr0KiNyOH8R7ZTL
TvHyfRwD1rt2LvF+3TBsGrXx2RQiJl+KwBd8y7ReYaA3qoe+HuGrR5/MSyAFLPMapu71NgICLvg3
zhFCAC5xvVsF0scFu3CV04TiOFue5OCAEUed6OsHJlCKTpFl80pgSbUubT4hMogreNxv1cU4OaC9
g38rAqglwGF/GSX9EYlopASAz68eP9i1cq4MLRNVMykZv3mi5PruerosEBdXk9SuMZwpdOErY/2y
5gUlaN+jV1KkP1QF1ET6N1lO1qrX7iveElwKIceN6Q8jkeKm5g+mQ02JvLBPyLnOCLG47XsFfdO3
8irOsxkoEft9QOHSAey8nM6z6aMeWYnb1jv+Fi69RI4WdkIIVxMtTmIMwLguxzNC7IodqnGMgMY/
4wGDPqdGxlOjd3+u4ODUt9bEw2kjLupSFUtHA70BImfs9q3gXaRdF74B2uavgHwalTCbHzD7Tolc
01KHJMHJmaBTQCKuO5BDc2Mgj38yQxGTsQuUJs/DS/wbFJ+lUppYBbMBAetYT3VNU8QvAzbny5qe
6dWHKpQMj+47AiGqbECiAr4Xq5/U6USF/1rlcVeiRKVm793v1zLCFSjqS2u9rIyFV+4Xjw0Jmgts
/QCdCIT+ua5lK+bHEZsUyDmhICT09bhrQs5ouQjW+4hWdXOsypzWWNvSAFhBGRz3/+ZtF6Zkreiz
gaHmHfzGksRD8xIQcFaWRIP4QWPE9bNtFZqYialthQHouf5vtT3Z1NKP/76XdoJIxBJxJ1WF4M8h
Qo9AHJ3FFld2B+i75Mar4Lfe01SW4RByZY0yEOdv1Ii9SxHtFZ8IKbmfuwW1PNsSz/FhqWQHxJn0
SDdEgyEFyudNIkWFsMz/uwQAweWcJGHmxssdfUcWhjuOX8TT8F1q3FN+JfqZ0+ZZgmSz8JNKcLCT
NNaCofPKpBYjlnNUexmFMuqgowAc1nGrn5iQCCo8LiWIpsUL8vAyIidiPKdBUYaThbCO7+HVy70a
GDghMPIMUqUEFLEuh+snYdsGQ9LfcRd9B8xHllTgHCUyDlYxpkRCF6hkRcESYkWmp72xhJHgc1Vq
p2A4PaIexQvAwH3R7MUsyXcgS0yyyoWcUW0u/146RP4dXxoflG+KK4dwl0y4qiWPy82DcYVQuPLW
lS1cOf6yj4fGmwsOooZgC4hrvP1nE/pHgOo+yjjZooTkHYGeW0HkAkZpMEO99jgXIojIQY0dIQsc
TBiXHRqoFlk4JpHDFS0NCX0ar2Vx9x7Xdh7IZ/sbCKKydMnbQIq6GuKy6b8x9fWJCniFw+IDMHcg
avs7ExBXOXBGIWe9At5o+YZ1UBU5Gzj5yHAz7+xm57e+VFYGxZRyal6X/DwMjXwikz7La2EUMURR
KkoQ8CtcpXoia16va+VYQ4v+Dj8U/RnHtlS+EswNv8cefswUxk/CWnnoIxELETOekw8QuP/JUMy5
rg3dlW8avqZhNGmxOfmBaL8A7CqfRMshk7FEDiYJwFirkJfnYu3yNW/rl2D9fZjpf+Mq4sfVmUtv
5eEITTWn37O5ByyP124wpY/+7NSEzEoQKyJviE8x7TSZNddO7fVD3YIjqL9PfCTXRRuUp2uh6pg0
NLG9HBqg37bVk0Fv9eYDtX6qVokdbbjNnHe6mddXU4Vyzci9hzhYjzibjr5zamxXaYam5FRtlD8g
BMVIeOnKeKYcdqteu+UpDFkxMT8Z0JVzQ1b8p+H//GkpnCXXwUIIqMuMLA3lOH4FGDYHjheY59Qc
q2DTlWZUzqcFXsxxGm7TrYz4Lsdko0T9S8EeRDSWDf2JElaeVk9udM2o7dhSFM4VYhgJ+j+ungk6
6QpJIWC6JWtL7/0BCmne8JGvEa5uPWPkDYMu+mrROVh/YtsXPrbjLAk+NIlrj/XhENYjggXVDssf
WT9wpfXtOsvpJ3CRocgYzcCD4Y101daYV5vrOt23dY4Z7dgRSy+KRWS3fe/090MSe3Xm3yIzJy5f
pyXJARCfJwQiNgolEkLe2wFx5KD9eYTbUBWTpBcYm0ljmyU+AWbkYSLaHw08iWReVUQQoPwZx6+G
SVIib6v8KCnUOun/pTfIBGpBGTlXQUnbeRNR2f6Y0LWb+6t21/MXkN4KgbRLbm2ABmu7yyYNRgk5
UWJOuHiZMM6hKpDF5lFm48PXiFBJ72v/s8iO62lYZb08hs0rvNEk6PYomKdP9xsvWYKHDczIvDlS
PDRGZUpUQNw0qxK9vOszYyhgsocgBv1XpD+e5fzshaAAVZ9qFdAfRj7+fFg3CeTAQa1lH9C7yEqH
s99FpNGfxUh22br7ItqvQaGd0G2+EGolI2jJvAH3FlOoL2ZB6ShMi1CIlaM0Uz+L7DbuEXPIfZTr
lmucjyqygOzBUTQD+gngp5HtaFGMQlN+7BkFRLHUQat+T29GTpzjfMMRwLZ8a2S7UdKWXJImYzhM
a/Efu40qG3VXZ05hARLGSWbRDrxquwCKRrHwB6Uq8Ftr9NtmVcJgdHwLHiNz1U7TcEJwWUr+1zvs
2g8KnO/mgVufgnKS8if0U/hZOVv2c7oj5Zr23/qzeOBY8NhNArSPmPilogbULDQ11v9qd63qARHC
ok6+0FAnczu0zpHlWke3bLmIp4uCqmDug9OM3zUiTJeLLxsO3io6+qjiZYYwaF4ns4VypqMpi0m8
sS/ZU9J0P0UaPLxpbLpxMjP1Q/tG9fEmInh8R9YfqPM0BYP1zEhY6cojDrlry6bh6BR4Ts4kwhqF
IF8JwPgQOIuPnwx++GDz48SnBfTW1kLn5JG7K1DVoQ+GzE9bdA5WbPg/a3lEwjyZoNu5TL9b8O4G
xf4tTAt0wZGkKapSVsOxaVcePR3PylqkzmbxNm3aBy5oSfR/7MpQ8YvvGMPr73r0o2GpMILV3jaM
z3p4KCZTFDx89yWS2PN2eTzzdvGSVcAIaoMe1ASzzAvN7VJ3Qg1tQrpQXl4/ClJcR+xh5mi4aYHF
Y4NPp91Gl49PEma3PdfDLmR9EHqxHlTeoJy1Ux8Ou6XdKVTWaopBck5LqLpyyapaSlr8M8CfkqlC
MQ0+RuYFWfVFXi+Ig3FWksKXj6vVHNK3PAcoL1M6sVQW0ElkxhCWOzlO0d/6ouGIGsDAbBTgFlj+
UibemAas/ZXUAPfQDv+Jux9pASSp8BzrRl1+GHZcdNUHvlFjNG1JhTP+4+A1ptVxTVMp0/AWdec3
w0V3xT+n4Bv8AJSUx8VoHNW0AVlc8T6+58iy+yhn7veFgIbQ0GE6uINUb+M8zds52NoWMxdaj1oZ
0UzDdnDsZt0qaRtLalss1j/BnTZhOjNGZhBbUhkXVnx/kk2uPGG2Ua5NqAhbwZdzVbReHBvUYuc5
aU+z27Nhw3q+bGvnx7g+K6LGls8OhA/My+RcqFyK+5fQeRpI28zFyrP+7lt+l4nUmAPJe0tU3x7t
Vyi9uJPFmLBnfnQQ9bVT+ngLwjfNjf/SGl8bf+7xhKtmLrq2zusz0gvIg6e6OllTMhdfRKJL8GWb
u7fm/Zpe/e2qfaAIJT5jkfmTOgsNMJxsbS27Jv70gjbI1FnFjYLypQlI+pyWemb3UFRzb3VQl/15
HDPxQTREXvv0OOQB3mXqnAz2NUD8rNxFzbLI2veQsiDPbpntXJHBUBST/dvPe5l1gs2TBdRiHmNq
hUDus9lhlGDi7PGpJItSSOkCf0bfXva2JPUjFf9xWAOXCsKEIisxoLSHYqDS8phrHwok961PvI7f
TOHDPu9kGy8j2ywsCmKbASPO/7F6bTYVDOkL98+U8WmqJmRsexjHiRDc+guMzuSRAAZL+pCr44yI
hoUPPbgroN1DOBUoD3LdqJwLOEaA+7k59Fwyz7IuwWrjp09Zb5MQ0uRz2adf/O39Uyn7acjcDaVS
syoG52hjR8cjkt8iyNKOQ9EBJodLtqOVv3xnL2EH3WJ7S9bQh+782bv1AoCfMNkA0HkRi/q34otD
defZIs7iWSGy/9SnmwA39ungHhRqVjgU9Puz26RnvklddeEJf3JYx3k1iETYoi4JHvScoCidstXO
/8rXtTaiqfQR1QWOj5XKiegb6ddWnhujUCoGt31+YwHtcxLygkJqpJkvdB5YQkUeHtoJfouQyG1b
fwZ7H6rVC8iTbfUyGvigdkmyWPUeRwSy9b6762ysmE9566igdTR8PdDHy72ZJ4effHO22qdkSOEB
wV5ILcpE3a91sZ2HesIMq6017RMmke/eEgDPa1xx3HpSmYx8ytbvdk5FthICZVUug3S3cr7uadQL
HW48OjCydOb5pswTgkeFz0QiETRTLcgIKQnD8lPY0v5uBYKfofURi9GE3NXvVLPnJIO3w191zwYH
1YLMEDEaijwCfE0FQEcrEOwgMOkSkFCUpWmDXV4YWj+FG3M0AdxqBetQb34XGNVnBnHSpLJcNSe5
zM5PJFzoeojEvStLATYRZGnW7KXwr9Tih1YJLuYnUV0WPSfFB6G//De+tHeNq10b71DcviqKHMtc
OEnVwjKQjEMOlEP0p/0Khld0Zs7BTpd2iAAI7WJfua+W8GZXBnB07NXrxL2ZP6E0xhocS16a3lN8
OcYhj9RSCWLYBF2nMhECQmSHafrCEHKt4IgRjer7kSyJ7RRTL4lbpR8/Pf99+O7rkj/uvnnT2uu6
5cUArgx+OB8wq6bsth/qQJ0PbpdN0Kkn+U8ilvqBQN7wab4QKwvO55iKP8TljjpAcRd5Y6HqOHly
Ci0ace6vvqh9T8kvdZxe70QXl3A4KGgVXjtekM1JhqcM3qrzCHjVWU4rbWBtQajCVilaycUxMNdF
NpI5JszH7CSFxxj6roCpxJDqmOJ3qqX8TeeJpwKNengcwz10CiOniwTgIgViT8TLoHP38+lFR8WE
VRUrBrSSfx6YBX6ogMhdDMNqWAUHGh7Eugx9QQMi8GHlucWAvUtZdidtQPPNhjB9nBGA2BAjYe0N
MDYznpOIyswq1kB+7DxbFEf73Muxw7reqYtuMEraWFu+VDefwPVaFDOIH5u5VV5tyaLioWbhMBFa
7/EG6R2eX0kOXUw7Ket86u/SADfZIKOmgY/dlfxFMDp9pJhtEF9DSkK5rC/4GL230d1xw8c/s5HR
Ui1lMGXX/Xge+EPq+fBv+rwGQIcSa7aQ0iBX5QPfGQs5BNKvCKSTcEK9CBiokveHW7OibHffAvh+
FCcgQwHkZYGSVa5M+ZCBESYjocps8TkIOmLhTzBKRsbPiybC4/BBlkVZUURrJ6gX6QwTE2u8ifJi
Ahc2lp2nNFDr4NUUIqL2ZtHoJqypehonDwOuxp90GenNe+mHVtAbBJWS7HorsFRMrFTuKOGvB5/O
d/EQ4Fk/Ryoaqlg6y0ow/KWP1yP3y5FFhVrvL3G0j/IbX2gN5+nUpxeVZQm1hZ1B/ekP7j4V2sLe
CdN0SdXiGhPKH6y7U7U27ipmeMAUrzvaPoeO1kEfg+NRe/MUl0c2l5IWQCRnpAmDU1RRvln6/RVU
iWgO56SLaKYKamcw75E7Q5I3CKJ+J+MkHia7YIp02y/szf2P2VeuM+3mwFDi8myI0U9qA/IqGxtk
YMA2doAXJTrrOVSJReUv4iHxRF9NO2UJuLvS5Vcc8F5VM+H4DbBWe9JttA4a48iNi5WIM7UlO8sx
jJw/TTfMppb3ivhc/Ariq4DHEjG8r8EzYua5MGd66becuXYKqYoMQf+roIrXakVpZZa6SDCIJJDK
FWTlG/vtxWLX9+a0Hk679aKjEP5Ey6hfVlcyizojiuZLEwgJUYeQqJAEki1Nfgtjk4MzIVbtb2wa
YpW5ktx8Mc7U+Wzga3/dnMNk5QYeBl3iX6VwwuGz0pHl/jc85k1YUxHq5pk3+b2f6okaK1tn2xZ6
iEcHtt6hplmuRKZqvafU+YQphUOgGLx73uxlTHyR6ISD48SGeovhQj4nlyk5vtagvYvIa2MZBjtw
FmkMVnzHKzJzA8TVOriHG/Os3hnlrII4uDTrF8K1/KrDH99J8g8siyr/13yoCfBNX7DdlRCHv+/Y
VbVQXWfQnASF8DJpu+fGiijjXWZs0AEYihB3Nqu1W4kHL41qDhaACb1dXLoMbBKZpRBY64jpdBJc
sDuSXt/0STv774Y5TeBFHDy9OPdxoDlXn3AalDBf1hl37E+ZpkBHm1evZjDpRAH5T9bTs1MyUAEn
G7Oit8uy3qKTWUSFj1D2PNKoTrlEPMPT40KX+mxwdFS/NoSLCie/Ex3aTD67Q4qBh9xbRhYrXZUK
YXuBVOV7PG6S0sDcq+cwu90eVDkZ7EZIlOlkrNijZTNzPrL8r+rcOSn9UGF6polosgXmF4GWbqDL
WOlYCec//r5g2SByLTBdJj6P5DvRVMN8VzcYHBMLbAjPm0jLnrRtXM+63wRKBFG2zCUYkOuwO5SX
W6Kin5pnBQCGHJJ8Xw+3Ezns6Zq7WQJvBtAlHaztqZOU5Je7qdtC5nxHjmjDL/j6+SV+O3yTrfx1
8BELq44J+VWUWgYWJEb0a1/wIeIno31JX8d/HWK75sVFss7xmYgT28ZSCZbyZpGBKaH0saI+u1Bw
eXYtLgnZeCnk8LkCGTiEOF7ufidww7Gn6tk5iApfphNqWexhtzVafBNC73IryZcAoxM6kNtpprf+
XdgFX9GwA8+bcbmyBpj7qEDLqBeNZLVVxHc0EVTtXTYo78Lf5SddTp5X/0fu+Sa4vn0dd9K8iF2U
6j/G19vDFXhv4JjF13bSPYUOe9JoVAaqnojLrrKRwdZIMZCkvfL5x98dRZcDgqLmfdh2kE2qLsoj
wRPSj55zu1UOIJmd7InBz/MvF0y1mAZ1n1obh+hUj2hKgbbXJ6qB4RA9ZOW698APc8Mvr+uXT4c1
2EJSHqzTDhxYG3rKZ4BgCf5940Z1DTmufPkRwugtgaX5+H4+lg4bnhRQZ2nKrX58oDwnB2UA7Ya0
id530TEhfnlQ9I4VW5ZGVPq0uX7GJcSHOTyfebnZMbdh6rDMblbvtNAoVcoOFLgqmSpT4B0602An
LOqpFTIOqAzVOBga5PfEt37I89Ap1hXihqQd/zCa6BgZKBa45Uvyz1LKCbvegJAu6NuYkbYSz4wl
Ar0PobUeTfI/ahLYpDZKqNra9L0WyQsWLq0popVvKCUtfoOgvfS/Bb73cdLj06caLdJ6cw5aqghV
sP+ZdhSqvzIvIBnhE1CM4vNLT+zrhbKETqqNQWUXOEBWoyRpuxeX9SIrnQSu+P1mI+8F7Ha8Bv9r
GTcBdgxEgvY5l4XIkJHYNOvfmyJlTIw/xwtH6WEa9eyb4p5AeT6PakPe8tKiN7oiybCMLswafkKe
t+52rO0Crtvb4RDE8A5iTc7pRGyEqDVy47h7GZrd2pr1oG+YAUfGl3zjVKEoM3DTZhlTw9JDaf2d
me0Oeqv9HkrWRy2zYKOPb2cNNaHDK4LQ8MJV7aDy9whqKge7hQz/jOGEJ29orlrgkCjYtUC23SIF
YizbGGlHXWhpEhd+UrwjDApAon/Q1fGhrLu/qh3fdYciFf6TTzEz80e3tUunl0c6OmoCDDAEJDIU
x0/tVhkiTgb84HZtdlvQU1X10x9XWAeVtzSnkkvKuRMQGxdo1b3uPkrpNw2DGyZxhx7O8KwmXYve
bDKNzhaAswHpEmca17F8OHYj/yJ5pGc/ZaGPLKeCIDG/oRySoM9S0tAkgJ6hRdbnafZwJq5Wdkov
IW7skSgu7O4OgvkxIEqnjwVPw9m+s4suF62Dm14+B5M5OqRfgFDxrLKzXdKdKN03aJmtCRJsmaj1
I0WC7P47Sq7e8CEVfHAhpdnIHZcZROlNVnZEy44pWz6ryXjPj3BBpixa3C5m+iV6mGBxovLV+zu6
ksvekM0HoLU7OsZQe6YTh7DRh47E3xrVROqku6EWPPaKcG2FYKozqtwoHjtWQnm3TsVcTuWQiEOD
1VKksdVqEH5iMKkI5tuNZ1a1hl6agPFuMy2a9BsMdHtgNXQRf2Udr6oocCCAsUMKBq1N6aGRZv4W
Ha9H0Np9EDpPvX89VC+VDqFZoXMqldj0R/E9q9wcuozwh7Jcd0OkjJJzK+gfZoj74UX6xVMWljYW
AW1ifAPiEvMKhbCqGOlsLKX/iH3osF/c7Zt8pUWes8Y5iLPn/ym+N389VsPldHAPP2BmvlHLsZbh
D+7TOjaCnoutr8akDpBTdx9oFA8iwDYfJ7lXxFfTsj1Gspev3NfPQrWKI2v+tRw8Z4TWyeG8mQ/Y
Jq7EZZfjZOTkT9oWrKlZtGSCZmJ87t0YEdxe7vZGC1BEZXillUw8R9P51s5cqotxaMXufDu9+tLL
omErbhTrH22Cov4RLb2T5IOyDI0Zj+T9UeSCzBosCSeSAfaFbLX4Wk9G4Sjp9Pim8YHh7hcYMSr7
AoCO7/0fkV3tuVPArGTq/yS/srY7b1fsns5nL00WGvRzT8Y8QutB40twZoQQktbESJXM+Wo1yydl
t8fM/hFrKKBEeOinSE3GHfohQ09+/TnLAmhhyoDmXIUg8kleeVf/RnstTxvGn4YrxzraUjZ2eFIU
DmrOrTfVwUQIufaBpxH+G1oxfvSdutRD3Xl3IUHAIqUDZD7/sm08ccnlDVLj105ENpWqm/huwJyJ
ebwkd9gJiBnkmcyYi4HRsp4U3aV3spaEMx2z6fAH2WSmw/Hyam7k1/VYrQ05Fu/uUsTYdAolz6Am
KnaUkxI4c66I+1CRCXs8ZtPfGgyeiPFzuy6tbtZRc4zjavQNDLcyEFF49p/Ewjt6fyLYfls36wzM
nZOnIDAZElCZjl1QiI+0s/9Nl/a6ml3OOtlSNtGAnUhf7SMrjoY2s8DqtImDhKH6ErXZMuPVB08e
r39T5ztZ2sUKMnIBlnNTo2ZlU37ajI0lEgTCelBAxgqDIj6530mGNN1W7DIvRVJb9GEd2JKVU6zq
prhBRuYzQNVVebbXf7lWis4XJRhHFQ6zTrNNEUUVyn3W3RflXL3cGKq+s1h4CMd4KKbCnMw8jNVe
TmmWHf3Jnc18K01rRNLvWwCmkAKkE02eNrzaxO4V7E4U3zcwsMHpd6BIs0dRxPAScWVQZKB8G8qf
JPKQLTpBof5G0Wy7VL9/qeg4oNYu8+sL/sgVpaxO+m84QOnoWZUR58TyrQZ6cUrrwlX6i7gXakJP
H6Uq0Bs1IG4xtb/mC076y9ZHu7dE419TQI2EsaCko1jB6w6xbzRT4EQyBd3gphGICF/II0O/zm41
448Q9vK1w7dRX/tgdQgYsP3KhUnQYniTVnpfe9R0hVYaDNO17YYP9/+JQIU6lyp8OBDiZvmpz5Xk
hgIxUJWfP8oGy24hG84lIEeFxEGaXuA8AfY6y5q2i8LPa5rDty4VNaeBBX9naHVK9NsBpyQ1ASXc
hrhRXL40+TyviobfBGKZu3IVJ+q2uteK6yxQLbKS5YI6U3Ivs4UpLa3+469bfNTw2pTsJcmdkHT8
U0w5naPWIDjXNq5YG1/wKmquusdLLO7Pf6YKJ4PUwPCelPtb40DWoyXNv4LAwYM6L4yGrPiCTFR8
C2Qgvnl8MeCl27B0VTngv9Z0hh2SLQs6iR6jFLdRY5vx26K5nPXLbQY3gZQVuY3ap5Oalkytsj4B
WRDfyeUb3XG9n5DjMeETvu+V9sRoPz3NeSm6puvDFoujxJ5TjDFgPV28wFCzGkVSDxlkQEg011kh
ww0jbH9Z0qXFlnCDSY+l9XglCR5JzLJn+kh38vD8FGmqgKQSVraakbJbDRIjdKD5JtL3KbBvXlHe
cpbMN3lj2MPQfqEHcWIyRt59dvVHVOmFKQvipGIZJAgtpozofmEa0i81KhXlVbq4eQz7o2ggJ8Yh
NgbAfiz4Ojb9OgYtimcUO1QJsopEKIKZLKQIJumVkeD9Ce6DLaftOj4G9V7Z+JLozWYn5NUbGKqw
igZ45OsBbz6Zt7YxiTSmeG0DtL/2mUttrI3QWV4Srk7S4WHw4tqzxlcqTQgUJQ3BPf9igvNxHriA
Mr+7/6ijWhf6bCq/Hn7ADKg95KpnmBv/Ei6wkTBdUat07YkAwteVYdXolUe0EsZCwE+kpmd2QSBM
nxv7FvqoSon+ILkc8JKm3CklZ1+pkJpH1Xtxd8hWDiA1wnLHEsXNmELkJYxf+KA9s/2qKiELicun
hBWURiXGmkFSdk+5FwCjXdOavoNFzcRPjBV1CmRQopRsLu8FN7G7GvsFZgDJoT60+CSPoq7yLsvF
DaeeO5fyfiUJ8XQFcJ9oOMwx0tQARON1HCQ1Tkc8I1UA0IwGuDNG9imu8mJxexnJ6TaGcx9FiDiR
hEj4oYrhILJd9qoGkJel6rRRGHQD+VivulNQyWbF2rrjDbMvbIaFs3soEv3YuZhl1K3fKFqcrRr3
MQmZ5ka1oApwW5GMtSNNlPRGG/ZD0RPgHEL/94YdaBv48so+9RR2KdbARw/swrAVqV0z8iNd/s0w
cq4k8mw1cBhjrlDJkdOI1pHyAhQKPaLB+by6d1n5vijmYjitxVEOMqrce+pMaP/QtEHNpa9MT9uj
CQ0EKUv37qjKyp7fdCl5DMNmJo3nEoCrGW2lO9Og52PBCNT2GBPrcnHUBm7k0gx5J1t5qS8BX6zk
dbeMWTJUDM7Z8qiVZrCR2NooiRrrGI9Ca0BG6IKA40LGWKE0U8G374WXS0ofIhU9yTi5A6SnMcPz
WU1z+1dlJ/LVgFnMoIyhdeOAr+aWAiyfSxL1nyig07kwMm5EQUai0jclAmm7W6N4uAhlKR8tjMqz
9Ln16KuOItjo+yePnJpMiGnkRyyygNkzXAqY2jG6TWN3sVAAoo01gsCboEBDprWRg53BnF++7OGl
69rnMK0zkdJ08dso8DmNnwQfJvIXHPvvp9yZrnl/M4uxcb32t4/h8g0jcqVz8ySOFbcH1cwgM+MY
WF6U0tREE1wEDjX1AydE0SvMCyBwQ4yfjLy/mN4FW19rxXlQ6I2vzKncLdRldcpF+yUak5yuYLCq
VEqWuFzqRr4c0hd7fvdSGWHo1v/TFY7uTITtFsGscm5DVypnug5XVvPRRwtDRl6sqzTHjeu7cHFH
52CNbEEEtyLnFaLa+hzxLD5hY90wX5DoPwWkFHzFzJdEpBjjVwItZx9Qaj+KzDe6/F2igjezB2Hg
NGa6o2phRn7Eekik2KDnZavLKePFviCc8pSCzeZH+0I7xhFBmcbSjj/d+zCI5GhvKc8Yzz6ZuTBb
KyETJHXFcEeBvMBkyAl93LyylWPsQRM7ID/ff2xfg6/dbQIUgnYVcHv5KiG8EpRC6g8FR0u4sejR
jDdV0zLBT2Lq2UjTnaEnHjq7qAXnS2CJW/9TIahco9tKiyZT12drYbxabedYFg2+k+hD8dTDgf3r
6Ml+OPA6qkc5QsQGcneOSwaSsjA5rtLllzPTpHK8TF2jtYXZ6eCLOQIqL6w3gG6q5XtESFZqQpkV
UbpFDnQN8yHrm4/jhIMnFKhkU5KRF5dA6SEPgmJAGGtsauwktgsb4jCU5yScobJoxarugwjj2WXU
LfDy6+jJ3tgb9FvBOzRGdWXpczZWX1SAeedQk2lbfwaa3R9dr1SkcV3v8S0WTmKgN9rs/rlPRunJ
ixQxoG2C4Jldn5X/aZfsF9wVR6tTfjgsuyXtu+184WdhopPHm4YhzLlEL7bpvpAoRf5BO7XPs/wi
DIwh0iV/jRJr4RMlzQG+B2fyb7cPXuHIEm8bQ0coAGCJc/JJrP8fmBfNWKvIZFIA/RII5rd5bZ/U
gDXtmMeVnXWFlfkBE0EPt7yg+JmErs+VtiXCRSyZiF2RqR26VRSpvkoSevhw1i0gJFVJj/2pXIMb
JYcff9G/uZdQF8EwkWaCJ0HM3NNqh8X6lRzGWnaQn6YK7qSJeskOpmZ2EomVhAixxq5hp6BYNDMB
9nFAdctXb1Gy9sq0tUvh827aCo1/YqS1Lr5Kj+5mcKW1ZK4mqF+ZXlSMDHtR5hyPN5QFhQut+0/0
JmVadSwFyGchwHI10DgjLk1bwkhOfhpEO35VYKAlCqkpe//vsNZsYDWURBrJ+6UJOL3J1Zby164W
26UfKJu7YnfY3n2n65PUPc9+z3iRUn/r2ggQ7xo1E3iRWPdQHJvLlv3ibalXR2V/lWpw8J2t3tLK
wgkb/s0SttZt87vC8utO8K2umGwKKFrhZBarqwmGlcn4RTYQWoN15g+idqmGKGgFMPAq4nMC0770
ScQNai216U7Ak5OAPpLwUZrEe4YPwU+zaFRMQjg44pYgMYAzZOEbgg/6SP0wpRBFIRRN6Mgv4dfG
z6c6zjEDfIaid8O7ahYoqtgP04D0tpwHD4K3QTLojbc+zulqpxRRnE/uWtQ5fOng29xeIiKYEo63
nZ396ZcKxs+/RQSMIjM7nXMxqDvT6ayfpqEGUkzU4X2i+MwIGii5lvSTea/3tlLpP8noMGl+mweJ
p45SIRdQ+ag6rlRsHfYBOQc22p1Rds6S7fGsqzJX3Fx5MqAWgO5KXn/UQi8Ywj35kL7nF6Q7vx7y
ytjVv11f4yP9prbgRdYsch2RFs3LrsZ1+Pkch6fhuxbD0THWH1MT8kF+GXiPZSy393nnbfRgCcua
Qsg288cNfokZah8uPeNOQeowBrjhMRoTQfUW5qV2+Dm+LvaGah3NOB1V/mjDynywq3FAMGGFSXbD
C42ostu7wxvv37qp6wMhF4OKCq3Z0yCc4NBeN4QQctAfiMToXlxC8PUR1LfzLINkdrQKICNEsaBD
K0C1KwzLgTioiI26wAuOpbt25sKNmJfmk9y5W1DRSQoDg904SKXSXGiqqCvrXY6Q9Un/x/Hzk6DX
aF2riyTElH1n1IsQEoVf3jDRfWuthyA7jfPUq47L1T+AzxbljB8Ly4dm0fWjqyGtmUnyM+D3B189
k0WZpT/4KZwFSkSG78uwgNQpCWO2tmVR7AmEb+GS6qND2BtT3bSpi5++cVmQolnB4jiKlInq6Gsu
JPo4mUzIiLi9k9JL8kBbT/p+/+lIM/deaBBAYTcEfJkPpVTi8GiyzL179NmF/KXUxUN/I5FmC0s1
ILeHKpO3rrHGSyPtJh+dI82vN5pgBWqjeqgBknTv36ITinjr8ivOi+XnYoxlQdzFjlslt+5akdfd
tpLYbtM4IblmTz5a46dT9dSCEYJB++bqyt/SMaENSXKkd0ugtyZB2t4pP9sc7GfB6dGczXIsQWSe
C5rnN4ohktgEUUn4svXPUPVOSzQ7CLQAjT+6WXgfPZ6xn8JDBXt36ohrml/DzEblHI+d+s594Zew
DeyFewtmXjWr8Pf/1awbMd4khqGkGOsszlTITV/DzfqqrhCqt2US8LuUER5bM6/ggCA+/h3OxCgT
CneSh3dNk7flo5heJMpr/NzrRQu9K+hejUwhPYyhx8GTEJ7wj1u3X43GBN1ELTU6V/qsmIprzpWl
zYFv+SfdGJRPuxeWNbFe0Mmrks1fXuKmgsBLu9p3AsfxBcURvPpVkpU5r/jgEJuaZIUV1garxT4U
gH22Jb6ySmQBclEv03uyRCLEhnTHjVYaYAeODLeaLriLYT7K93PeLs67B/+mfpyEapvmYQXqPhV4
HejJAEhpFn7xzne1rHOvcZffTgNjSW9EaUbZgSCcsvCGjSQLHFayqyV5XRAcDeSIvBlh0W9qoxzX
ev95nWBU/HF4ISvo70K2aLP0v4dT6CWoy8IrFwi3UWUXD/yo2cc4e+KSxX3z9vhjieU6DrjwLlG0
D3tHFPZMqdx49TOx3iZC5sqeFEEG+7zJJ4de04URv9vi9zAyc+Vl9BUl35uv3BiYSEXZxaa9DkV2
DAsG6ev+ly1BCJfJKzme0tGsvMTKeUuM97eILffkatS4EdtK2xC6jaKR+XBY4eJUBwnJGXuKslHH
P6hHndk6nG+kCgdF4rX8N+ZdLOFNGNe1nDuRRSRDjclyljadWHbktNIxBTd8Uqfk3KM8B1h7oOSi
GRmg5TfXJugzbnrW+3kJmOI/p54YfgfAxyQtXmtMJnXJ9z3OXCGNrR6aWVWN3ptJ6Tm9PVM0MoCn
ULbQIFwVDI7rDOZU0AAzV2jSgz927B2GxERita8umsOwfebG5+lVdLjlHNLYUzmTe0lRsgCpYdK2
LsoZ7Gag2FpDeM7C+9+9ekMQ/yjnM9v9HxGF0W4odb6ACGxhX9HvI2TPbYesXiGWDsAHJVCRmZoe
9WHcp3Dxtp60dIQoZRMG91NTawjlAoJ2on3ES1l6CiMRekXirrdDmSiBACp36Qppef6KuONWknHC
P7tUBmV/TPCnbalq1UIazabmFBMzKxNsMlpDJKvWDhbbRwUakfR76jwu6i+iK4TZQn8/3nYLRFjB
MLOMYPnZhx5TL0s7e4ULKvhzZE83qm0gyLHQjnCjUncuki8mDnexmWefGt85B5p0sg3F31VNA57q
IKILVIbmEiRgdD+dqzaJiGnezDZLAFSWzkSQeHv+d8FPn8A6uflJUma04qoI+vzjrITNzZuLemsv
T+zuOAH/9Bzw2DTjNrEpMBzV+inraejJUUOcDwkL8ZQeQUj0VaGQqNf9NYutMCtBCWK1ZsQ0mI8Z
CC70/KJq6BfUdOkhsrCFj6eWYJYS35KN2wuWSYCuiEYpWj2y9OKi7vPRp+XL0SEnErj3dsxaP6E7
sK0D04oPQfmInxCZabaTewd2to2jBP3NIQtTbyahJ387E8x1MCakouUt48Ot3UF+pihkV+1b7B6R
kTspEdzpRrQTvj0NJ4toheB0JOGUZwx3OKOpa9Uod15IHYYGuZI0uew3KtGOX81QJHAIXOfN6AxC
TH+yd6QcpMBiEmt9U66C0Gty7W79FuPxi38nRIB/NkdQGO8oKrvj1PLu9b+IoKg33mZZrgS5ktgI
PvpfkvqaGdSmP+ZKGva90iXy/+7AwlkNHhVDJTpNTPtKofKOH4g/zSb+kfDaw3dxh8NoiTTOSrTn
jpvqfKYQjfNKMkY9nQ58em9piJ0g1mLnCEalyIGvEB2gjLEbO1oFy2awF6bpHdcZ4IfB+pW29U/e
koapOxPSiLDzBGdnWiWlB3wLWXq/Fgs2Xc61nl3QRR7Cuo9Xc/HtOPA2o2vDbZ0Rth3cmUySFEtl
tQulq+EsQOszR7jKxRv21iA7LbClK80/Yo784mfMxLbw/uxzrSh9mPPZXpwQbXWV2RXGN3UzXuLc
EuCEq218sXMfne6xvMq8E2LUIuLyoOBM2Uw0rs1sXuk1fYR6Chn93RcWSdw3SOmD4DJkqAJsaDDm
ANu+5ab5OzdrZbRtlNastbgkBcjwE0rl7MOJazNFhhDb6gUAdYkycMtPqnCTbAndEIooni+AtwSG
ez4ne/iVvxMZsgyCwygkd7rJDp3BWjLPLH+o+3DHBQzUtimaYGmWCJPSN8ssG7rQuoDcgEvjqPu9
kc+Rmhp+Nm1D0r33CKyL36r/72TDW2LDX5qlVCvAw/Es26bQ5C8Jg1OTntQ6g6DQhSD9DiuMaHaC
52zmB+hLe1qZQgRsQe+yAYt42Si5QgCngIGcDIQvpyazDeWLWo3IWJKhMyLRNkQMA4m65ccGJOqP
wdMI4N481XPaaJAh6WGqfRg6KuZVwGijRCurs1juN+OSzkETyAKs2cyWnoT9716q6XX5nu3icV3z
sXM+frCLj1Y+qQt/iKP1pd/RTcwf1qAZv/TlPgqAJBILZ/e1l7nGRVQPQog0ehgLexcihRWTpFt3
Z2Tp5ayT5EJ91x1ViPKACZ23uNPVgQX8WiT+2NjzWEFSFsGM1qNu5N6rELexmkcI3cT+hNai+6q5
149eihoYM2yAnyZseLP5s1qk6x6qUsU90/YQnlDdbJmQWejvZibU45LIe0OySfwDaet6lCyTLXF1
/XoM6kUKjg6gwyol6JmAcKEtecdKHIhZgxC5QM9Xcl/FAnKcHTNTKqw4oSN27RYJW2bEQMEzXkI+
I8KFbvVZzbqdJES8N98mtCFk4u6uiYuBcgjRra45pZgo7QIC1i6xgptCZvhSO8/FwNS8QaHzGCbx
Ub9y8mx/IsbjTK/7kebW6KTnGyh2/Mg8dZG1e31cSpyRQTrjI1Ruiho0rcYeYvywChvC/rQQT1ga
t/uJUkAtOK5w/+LTy97ZR/lBFbtT1gn13WbatJ9XqS4MagJhLlqem/SFWhND0hw1S43M1Flm7bm+
IdCJQYbX67pdDd4V7Yax4C7OCVVqtfl2ogzsv3Pgb+vUxnXIB3f+HeS6R8Vppa9qMkkXXz8vFajO
XbS83Wc5+psxNuQjGkcJvQUVEUW/CJbfiDXfz04TXpGlepE6zPmBJoF5s0XhQrhkRtGPiomP1fUS
gtr0vFbbmtA+fuYIvk+cwP5ygCDNhPcrOCic87oFPzwOAxn1V96BbNG/ViQiYsegFJhsgt6g/CUL
VxzoqUifmSHQGHleGqAPTRNWQrO0vf6k+UDVU6bf4MCDrX7juQ8/3Q==
`protect end_protected
