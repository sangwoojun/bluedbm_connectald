`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
o/H5BY4mPfAgmxiAgIGg8X0cy5qY+k2+uSjBTcBKt+JDOsjd7zA/Zx5IEBN3APghBzCqErDzWJ98
BHAr9ChzDA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F5iGFCiFmAgG0CX2bxqSTjkViY0B6qayy3QDMLw5wYyecrVrpLvxVlQE9/KOuB7KNPARwGqF1ANU
K3DHxFybZ4cxlLtUQV3+SOkxAjnnGkJcRRueqz+m6R/Fvqe2Fy2znkTfUjA0dFEHY9bakt4n7l3o
xFkJQb9/yCuD5wPx5YE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HTv7veARJ78cKEwNn09gdpP0OrT+zg8d+L94gNPcrG/knJXytcaTZxQmq8GIgwLXWUMgC9RCgx3e
I9CJ7QPWE046nVSvAP/NtuNFYFhSINbK/vcOL5E43yVeeHUREk0lByynP8NOgxDivhKw1CorDb0v
nKzprqHpUpYS0JEGx/gPRf32YzEkQlEX/JhdLZz6KxP74t+JIee527VFB+Mpn6rcahZDbtup9h97
eELwtwdnSsOMfCNueau0j6U6M1sS/+v/bBanIcgQ+BH+FfxoGIzYUPtzdjO505ArdQZi5iw+937n
kaLilL6MDJxQGPXyFg/tMIc+V63RZfkHH0nmmw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UiTI9zCmhmnij2k44+QM9SiB04yZdxbSvuiA7hGd6Mf/cnPebeQsrSwdqAcsvE99hp6dKkAwniyJ
2mBJwHkM0XNfQ6QMZ+oZcfg1cIC0RpYM+xfOJqZQGW5aEC5I7gJCxo90dX7wx2t80FPYcSmYuimq
E7APy0zvKu7UbrcucRg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tAdgQ6j3IaKi+3D2ogyvBqe4an0N8QGhgfCJ02DexVNY70Se2vl8zyUSgSes62Hmr9GK8FAf2xjo
f96pYrgVojqbaTqdBjp7UgMCs/bL6oZ7T/qE2ucfHTsAdqI1buRQNEGUas1MUVUTlzs1g2wM2sw5
i8ibyYk87je2HzGKdx0Xo9g1qRpcpGlIz7sT0KpKEOLbsW2RD7voEQbv17MztQkNnEglDNFwfwru
aQ30hXhSefotN5qvQnqeHROGGk9NvXiU2VgN1lTz+oTOFMUfi2vnArYvL8jeKyvOUdn86K2fjHby
1vR4aPPT2/ai1AG6zcipLfX5NiYRUm3bB0PtmQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 43760)
`protect data_block
iYuQvx1VOZPrLM2uPxIZCEXCmE9pJxZRZIXVjJnhhquJN5Z0U5aFh+FYA9NMz/9DOgpHmkocWkBp
lvnSwagKcGMTdQzJPrAN8RksBiMBxnbHkBDoJjbeMeut1b38fK0wRrBQhGEzW9PAy0Q/neDlx+LQ
ryhMmEjYjgY60FdXb1oKt6yG+qCb/tI8FiAJupxK3X6LKQFDsb9XqTZSSkZY4CZw00MlJrI5S0ep
0bGwQIn4LlfoX7SeA/Aw1FikjgcXLZBzAzj1VvMvJI6BoxXjaJpCzP99lXUD84xe6wZZck4Gu3Wu
3Mc9/06fcYU1ENdXtyJ6o11KTJhitVZkLOQHBdLnNpdaRl0KOiFvFAM5hT0OfNRJT4akfAnWeSbS
iuUsSurJ5Pvy7yFLzHF7vtvkiWsVVPvCDjh6+6XUWqlys6QD3eCYlTuljsLQ+ZT+vxYUSH7XfXDR
Ju+F2kdKBxzezJUWf98M61f3J/il/ysTjNIBFUELEtH0MYzqpW/E0wnq/neqC30KQY6CgaDAabB2
7rnMSB30Ij8jNbLhyTV354KqXtZEmukCb1MF1M/5W3JfOAic6Ijp1lMIL2FmbHl4HD17ch0CeJAk
hYFnJQZ8cxVz4H0p4HmDBRB7IoSRBaQSBJRud15LuxUluqGxUBMkSScQurU6TFF5JAQUhGJtcEGa
AvdeVX9JXZizcbFAXV0h4DYhOyESL3TF/e8hgr/2BENG/9/GNrV1UwNu53R/JcnIWAEQ4/AUqhw8
ed1oi10Lr1xOsh2lgI7PEDdZUdyikZBbtxPSnM0QnoA42bOwSM+LNhGWh/vcUkIlxhsibOF+ncZo
nuzVec3o8S+OzStTogJXu2ZTBjavjJLseoSHP9gd7QFUAovj0BmD9MOR+ZW9MmWowEWNGH1/aHtQ
Ad3hFX3gxy4Shi2bIea9e91Y16wp7qMA3Nas8M1/uY2vOtzEz+IjWJ/JwC/qgejoyK6qszO+ErnU
rEnbgczna26MJE09kNaKTkm3IQ5+Le17PF2tMcXe48uh0cUxBsWYLwetzLtLtfv5Dx4Q6TCYupuS
mNZ0bsDvO9LSaZA/wYhoBvNe6bfdesYY9TFBb4h1CFa2qFDA7fgrvd5oOf+v0IPq3Wtsy60fBAK8
87jBgyu7PyGjOmRcRKSLYUtigDWiJkXEAkRFts0kDA7ehWIn0tYE6sn4/Y3rAakyzDwqC0ia6jFw
d3m6KV3mBdKLcA6XJVssywzq5xAinMSUdkXx/NsXQEikHSQRlgf0BqQepKmqYb9FbMetvlWN8429
5HRDGFft0VdeSpbrRpJRVSkRAtJ7BS3exZA3Sf9lYJh/oQ3cNM4alt/LgFGooYceaXhXgH/p4gIL
LAK1ovisTKp0FjMFVRNUIqAkBIon4R0AzhYO6ScXTAOhk/bsUx1xtkKaQbUBJhTQ7afn62ULYgnX
a6kiyL78d8nDNrCyTTD1IYaRRjj3oQ52K5ddS561Br7xjvK7+CYbIFbFL21rSBkp6D4wnkShpSsN
vV6xTPCRaN3c0NqdJ/RjHpD2KpLuTf6BLjI4DkZz49x+93USNJy7xEdMNUf3Lxf35aKsDh/KiGbq
4cC0etmy2DXnwWvGlR818BOcZAfcgtyJGN/vST+Jj1ymOKSWWXCZG6NoswIGz1LcbA8aajl7ON0q
gciGGeCA+WtCp5wgKDT9Yq5tG8Y+uL2qfVhPcMGnbPch8TXEytUF5eS4ojMMcsTXsPfAStccw+2l
8G6L5TIDLoTZSH/9jDvrie1eTYHvaqtZ9/t1Kj9Ig63c1yzJQv9mUNIwvuEbw8CFhfTM3roYRbAk
oNHInAu4mjsOk6ClgSy3HO8S6zGMSCLDrJjBDC7IEOwu6Y3jv6B1KtkvJYLSDTKPSRUL2thCjzvE
B8oqVByt33K4f2g8HHzJ3E9pwbbfd6NKW8dXHWTvugh2McZr8jOv9xxnLsdCZ7LTZZ67huNwrBFl
km9jl9E8IwfLomSIWVV9yK40m/xiflnjYs4c84YECx+rEPscCdLoSmSHErzRD7X1rtp41wJCQlfz
iNz99vA6Mayp67iThyaokEOguji1MZQOc66tQj242S9Syx4B7dCBQih8ySQW5A/5FmHMQvHIykCT
0K47LkVo0WbXpdbAtND3J1YGfC8cKuoxLRaomVSngX1M3g/eOIapgtEECQ/K+bixEvcrD1oMSf7A
u2MH/eJN8MaBvQ3aeSNuARuNfc0dYBnAu+YBDO2qSPgu06boRdWeJOLdnz5KLOSp71rmPBMxYyIE
J6djeG3aQp9Ghj2i9p9yWRA8EIEcjMUj9Ue1/DGps26F2HsuBbECJphfbW8L9LR5H3fnknZqZ2Ws
UXB705OFecIhYxXaVho73Ad5lKVE02F7nIQCkBG8XOXfWn4F5ATex2iheyobmpHEgEgGlSLH8VRH
rI5xJUHp3uipthfStpQpTfaOwbb7pxCwDaxYp1C4m10CgQWkVoGAzeb0XX5q6/F+6siFYKBibMMS
bEc8MNend0FuvSUhjzdipaU3qqeI0t91WOWFpFh3w8a01qyK4qTQRqAcOXDrBCM3DPbMU6yfXPni
uQNLS9w2AcHsXspwUbltM7fwzDpe8mfgnNlOB8jotslfYk1eYQx+WgmLeB/7GwX2CsJj2XGUTHqb
NIE1R1BE/4raiAAE+FF3DpNJsBvP8JOymjxZ5APmzvztFylRu1FKjgeuSKnRvpXTr8/FWsMJ9ygg
d9PUQdIV/TM+p2AWTqj2Gl+qSFv0iDv+MB45XpAlDT3TWozhuYE+zckfw/NpwYiKbXfjmbWl2LmB
CjvUa+1j9MPywYNunWr0cH2Qh7oZp4ikrQMTr5JCIhMvfQ6GF6yIQm1WyE/mpZQdQlq00bGxBfy4
h0QuhoMxCK+S84EZ8t89k85cL4CGU8/qBIj961A5KtMcroupuhzvQ9HjF2eNjjk7C/Me/iPopezO
alZU8M6jNp/QRXWhPwTI+UtikBjxaFefbHu3M2tXfYFXjhoN19XF0SSLhjjG0CeIpcevtp1/yGh4
5HEbHZ8hWkP/2blN8k6KixfLNvLUx25hnBqC9awsMwfl88jT8fe59zrydDlqyRsiIglMGb8ZOv+r
2suOLih2RRFQ0TOqbOES72psT+i0i7j0lB+kMlnZrBboPcxzBOs4BaQUw+J7oJcQBue/J6Xt3Lr1
iW/c2/K6EkD3Y/0J52VEUb2zf7MzCIpHwn066WT4HLjNtiD0l7mK+1fkKWgB+TD5ypilQYJF/dQU
Xpj2cf/Qvt2Dm6h0cCdfKvqmXY+wMBbWKaovWFs6eKUKNHHLVTI4UYeIJRFzFefXHu9SzWPnj0kj
hCIJ35dXrWAnIq1GJXUB9kjNkDmjGzQjIl2IT/q2kVvuk86ykHiHos0cypIdkOJa4QS4gWhs3ovt
s4MrbwjKJib3Rn+RQXwII4E53tR3GbNSSaAFDA3GBZ++hq1E0cS5gDw0MYoiT569LaLslIbPduly
VDZ4J2XZMjQZiZ3krRJu8Kr8msubdfa0LWrw5okRrDsJv5d+fPU0Nre/zVhL+cqP3NPJtHrfmD9h
1gUNa/G6+FeskhhxyW2wJSUGe+jmSPY0wWH4tEvfZNhNtj6VSuywUoYeQ64T3H8Txvxqewu7RP9y
uJ/q4KqZQGrQ0/S+hWATS2GMcE5sdOao9F9F2vwVv2jyA086dwOqyA7yi5frm5Pj/WW3HcLTApa5
4LeRVz2eZqTTmLZF3VyKM8yFqfSBvCn63c39bMTVxW76LrbY/BN1eoGub0K+UyRjnJU3rNWRKBg2
r6oQTmMU+3jQ+icgB5VKVeBlO2WZkRe+3uZXSZRxtL/dfnUC6oyvponsjirUvKXuDR8xn/ovRVrQ
MnTxiUn0Zhtug2TqxdBufNLw4MxwJHKnIVGo4gKBnQALyHzGOvSHb9G7rj+LFSGZ+qXYtUgYTmUN
OaLaMolvgxf4+1CmSfouiYUTaWzeyvMENv0oGmVThSaaGtwVzOvQbyRhQ25+769hiXlaBR/lnMa+
LraiZgWfjRSA6Wr5VQkYo1pfL65twTYSb2G0mibxq0AsbDqftK9oN+4O5F45SS41XhQXBFrH02lM
GMrXyGuVgwdmMsBAdRB5yB4stMWII/6H9dKCO7o0fN7q8INF3vRIqwn/MaUeygwRIB1lFZL12jTz
2nr1lXmuuW8bUA/vbA68VaWxIdIhzA5KwFgU6djsA0C6q+j+myZe8L4Cu464KhPkxgpVNlyPh3xN
7+KRWpgIX05iSTBc+2TgU+2UhBKzRSAvJ6Kj0n4jfcNNh4QwhWDN5KIiJGgew4x+VS4vr0jXeOWP
yDk+CPvtTamL+jHFPQNiI0StfUFpsJ1QS3s7Vk6JkSdpaG/M5uRVmBz0+OR9kp6zIvodo9xrKQE3
Kq8Go6enB0WYRsQA92DY34nwaEBtc5+WVqXbykVXqhSOHlGSzEkBvLn5fqvG7y5orBBFW+WJnK8Z
3Ag8CZdofWSctsSnLoOjE2ct7sQATphy//yzWvZnT8gCFC4c5eyWVUpr0WYFpmN3H3droQK/KBco
6nJaEpxT1qOoCge0JOhTlsr1rEVnE7XOdn+Nfac6TLX3aNjMrXj+p/A2Ocws+6hkHvu2cR2KMVJL
u7b/hx8Vup3cUEfWrr4K7gBZWx3kcZWxe8vWsDMC+12rBUkMHHLe0zkktoxTf6e50K0FcHZ9DLuq
4zBQWjUs35LMlQaxcggx//qVY51eU1qU0ZnbHPb9IbN6u0B3GshNWZdbYVrjRooTOp59tNee0CVR
/RW/VYxD4Sbs17l0VGrwufQXGYXs1IQFrGRxjxO20Xnsm2sefgP2cQCt9159brRBYARIIYVBAxNC
LygVboxxY5/OA6YWHLSee5+MzMmTSTGyWOxi/eM5cmc+syQWJRivyYP36SgMIsWcvRon8pK/ExzD
H2jMjbkHJ3t/DZngcrUzIfwLqtGBWXtcZ82Oqoxr2ip1dxGNqbhfjx8feI7LC3YuZu2zTcOt5s2L
l1ZWah4aF9EcHLP22xxwzblnodWscGWz5kEf8A2QWozHgZVRLlBO+J5pvBXmbncEiLDeARjxbSug
M8vpOkDKHwUnQx6JnuU+UPOL7nyKudiBN/p+x/jVa5C1c8Hmch4iJ7/pc4f0WZQt16yqAgqK6ARb
poX8BcsPoDARL78YswusWB1NQXlmXFlvQH9eWvgHQuLp0zGZMgmfCKxkQOBzhk1CvGuLp9bzfI6u
ShEgG5drUfN29A+kXUoA6eJENKo5lzT0QzD7U1lJ3gqW2cT0LYXWqzda2h7bXmuQprLX5tXDDWC6
0lLhaR73cMBPkZ66E43yELGslBRj/hUqjinxHzafBF4huu92fZPKk8peOsTXwMY30O6fK0wzPybD
uc9Qo5oqAHJkJxBYvEfn2OEWEBuUlhAldOwOJ1rCYQqncF8me9beNRx0e8kt2bMSZ8HtFYZuUIOd
dkqg14p2HgpNyzdnXYKGg8Njcdmbmjc1UrkV1UiTn5QopoUBGv0DJNuWlz1UwHWfYwQDWE7yzTmy
niU5Rfk5f2AvfoxPA2E9UPH94NsLtcTDzXXfHo0YxeUju0DnYesjRjkET5DrkokqdK4oMfRCBFN8
Cb/wbPlpfrx+85Uruu43gJ6tIZckleck/YNfXoiGEx+aIH6CSuQAahKws2hA+NeGIZtRmAcfl+Di
x7tOOhrWXISqxSpUdV4momdCbQR8tGK19/F9VO6gRchd9vSzhdWOU+Gq60DAF+zxAvrxRYZRXDmi
ScW8EQIss3sHOxrU+edj6CLQovFVenSGC/ynpkWM5MnblKg5xp+V/sHCdl2JJo6c7VaZNSCq1R/w
TaTn+Ec8YQlsBSCVp8/oHujJt3t+1HGgT7nm1Z9Mab2pxTn8zWD8TPj1ipwVHalXRp9arjJYO2ME
Za2XGMXsVlo9LsS4z0rWtHyQsAvWlO3Q1ZiehcPk3XbagY/fL/DyIJMI9rSrbASShD8bXdfx9zGm
faQVK2lxVMdO7Tus0zgozVuzdGvCpvtKofKa8EDjTAofaKZ/XY5rxtDsj+LR/o13ggIzaUsGO4pH
EGdg+qSRnXnOqIjE/kC59r2w2M55YD2vaeSs5yEOTpLyGR1SLzLUjgXWrZ1cTB77oswyZR5fJLm2
v4A+A6oEDBMY2RWo//jZmGoxFbN97n4sZ5BwdyvgfWFPfxUvYa/RU7XyufeYldv9/QBikM0DIDO6
jL8cWN+AUhPAAg6/DoZEq6eB0D2sf0ZbE+nVQ//5ZiqLf/73AACJelZmB3qUm0hvh7aaANivE879
w5vSNGad3prZ5MPJxwq6NDnr54Y4FZ1as9pHtAFs1oKTXLqvwWCaEF9GdxJfDBQ3h0RjpmwMGWr3
wKey4uTJRed1FD4OI/TzzrbWWdXMcKbFLEa4CbX+GtJpsMX8TvqpwiXVl2cP6HPf+KCEfsqoOlKJ
AAuNNWzg/ZGwObxEF35HWSz1gMMdp49NoyTERLS3CNIsl8m23FaN6y+txzKF2zRhoSC8742kaU3q
MtO0q81J3EA4VclivcQMgtffp2Fu1MOprAsoQayJnCrsehNxUOqkw6jy/xrzP2ldsj1ZQPAPLOAX
Zm0Y/KVPsCzEkW0cIIdaubxpPJCbTstbC5DUw4vF62z++5Mj4Bd+kHXCNDbROB7c3pg+sQxEuOe3
IL4a49xeVsE3ShZsfoN9n2pfhDPIFYH3+TRJYNg2MMU/JZN8yXqoE0yJrsN2tcHH+piCTLqtouAn
WUBuURxyS44WxkmjC/YUsAuTfbzyyaIobT7//cSB3mzCbsWpwjOzLs3hZgGs+wCmB6c8+JyrVeZQ
+QPgH3nUsjwaVsP2nxMnBmChWSg9A42eJ8zIBzsFZhjcNi2XMjI2S5sxhsqivANOGEAYGVofPenl
6Ndu5CipItC7h3nG3vU6nXmMMgm+Cgw3v+lBIV22Lqju7fo2T0aCpVZj5DPOF3PLcQqzr8gi6f7X
f1VbZeN3DX56wNyk7Ncln/b72iFVP2Sr91VuzGsWTeFww+7BCtMYcdq7A4H8DFH2Zxkdw7E6Urtz
LnSvk4WeCf1hYLcdQMqZt6TRxVcec8RHy3s3TM24pvEcqTgFBw2ac39cmpTTKkGnXt7g4u68NhY9
/Ncu9rdKj/BbxrAwPuhngFSNA4rlwkqZlWpITgQdmjQ7Y/GMM4MssevoQW1xtEkKkoV6fFJfeSXB
JQ2Ip1kwgP/nzP0x5Ao02LP4uCAycRDceBf7pAvKziPo42KhW59BkD+G45II2rK7DH83o0r02MXU
LDtXUMIECcUXIZ3TA3QVns8IQthO/to1Qe1tgNEcruJ4SxgFRVJwNk2FuQW90AV8KIydhDphzKUT
/weTL4Ha6E3IJ6dOwAeYhJQ/FuqpQ+lUdEFt2RCXgZLdYnsLmDuYh2H7JedOaCuL7yU/z8Blad2Y
NhdBCq35exhVlY07r/aMOZcO2PJZBBNRuwzG+g7zVOVHEUYekkj+l0kyaptElFHMbsyCBcFehTBU
QBeYMdoaKlpCzayUxtxImxbJlxp0gNCg/twTLVHk7Uy9NrtNrtnfCn6OaGR4YIzNyrVaIqt1yT0F
dcU/UAK4FJ0UPasPaL4wFcUBnJ8Sjh+RdxEa8ij61TcCaPrEDalqQEfcgDfIN1pgte9uQ2ljynhj
HBRpQ+wz24upfbqQsSRP3V9uILG725aHc+UfLbIZqLULpRD1b24PG1bojI2fhr4EtGHNm4E2iB9S
yAnade4moyjJZKVjvgXRTXlErFQkMNelDPUirIVtjQp9RrVb6tKFUOZinrJ718O/gQ6TNkN2Fbct
nZkR86ZA6spiITM/Ou78Sj9gh6U5Yh7wV4NaIMwfo703JICJ2xfdjdrwBCXl5l/QVNilT1zVU5++
xzMcNdhGAV37sjPeSfvbrUDnBh1uEpj3l5sRqkFOtz0Wj2Lvf9HLmzetOn+341X31OSlIdG579MB
h71LeGmM1VmhERtx3rm6G/XEtKhxjj83lkzpR4nVLIK7+NcKQstAOWjkYRiz7qqykPEkZrTn5Z7w
2FH1o1sNZuxQp8sdI+dM9JPAFOOsMJIyJMugm3RW/uMz3eZWmWYqqgDWgCU6EuKTzIx8mEPrXSpn
5wzta2iuS5eDutZxpD7//ZzwWyroe1jyQ7SpMRzogK0BvHnuO2J9fMB4bnIOQ+BYY1gmydC3u2Y3
k34LfBGp4WSB5HzFTCpXgW9vGP9b+peKH4A2w5RLNFdOk3GRhsUtJ4hja56v8nTjwOnn+1l+I+ju
yp9uMX2pl5qwVEb/ouGFfuQkmbgQD31VmP5ABtrc4SCpKYRz4ozKv3MooyW7yq+/WWNoCt96sovR
zXsqRhpd7FO8TLvuY/Cng3DeibnWgM6tAxU0DeEbt6bQeRQNj+R+eEGHR89iJnw1PmAk4FjNT2vT
TaeanrRi+p3hI9A5TWfal0z9wNrfqT17PXVNTrcJmEylXWLOUbiSvDWSqwOGDn/aRnTz0ZNmarvZ
XVcQuln4P/NBX42Jt5g0TM4R2LIfXK+4qh+Rk1lFp07NsL2dWh/x8/EfXsv/HRtVZTH9tbxVwqmX
UuKwSuW5wLkRQhPWBwfpDI/BZ4zMNH2bRjOPLBtxZZyqkvm0BBHWNuMbcLfX8gyf4urQc/bMuI8D
x/rPQwwj8d+toOoiBznbqhSA2vYpka7TnAbnWlN5ap4qZdK8oFjI8GMEXRD8IjFN7vYtJZ9QzFPO
kPQUFPQygSELUHCQxFDTdJaFwpsnev1E8OPc3Sply8VCGV3cPf0xrLKWrH3cxvRSHev8qlwiLJY0
Xbo5djGbvJk5CXtVLLcHrzHyTEWwYRP5L3FHpq+RUajkodV52o3qIFPDecy7qQ4ugVOBu8ZHlG7n
fuYrggLmcDR1la1DVv4U44Qx2MYWeG+LZtnSvZ/M9kdNfP0yKS3iC6cNcxUL88pav9ADY7dbdKTB
jbhRWAwQd7LdSoR5+gIiHgZ/pVNtLZYXLJoyqE4t8jT3zGi2lSuQMnVUYQh1O37PCVwP7z5PLyYb
vW0l039So1pJpmKuqt1VJML7CNGAByJ9aHA7lGsy/tMfqsNJ2jaex6+npMXQvcwBn1zu+o7LqvzS
tZHS8PoCjOQd+5jQ6aI1ac7tTydmy1QHn8NjJC4yvd/MkZjdbPdw0lHcYiw1m5wWeiqbeqTMUBNT
mf4PQyken9ABD01upWA+iOUZhfW8D0RbwmLwacNgdGbYo4kdwoGev2UOONzGkAj4Ue+o7/IOVH1o
L6gE4vHFCzcAvWPvymXMeUtc5AA9hi4aHcdQnVM8KTXh0MbP1GD778ZKUQ49rTeNO2h59tlr/1vP
i8Zs+H97Yqx0vJ3N53oZgqcGyZi5hD3bpbSxT5QFVhbKJbWWqWU51bw6B65Uilz5yLl6hKPVWu2L
3dmzDcM2Zw8X4UTej+YO8L6JXbpCNLeX9DeWLkRGjINyMtrtBF9yAPBPnx1+UAAV+vRlVTHl+b3A
JwUvruaY3m+YkJXXrRcm8BP7ZICHObL6ycjR3qvi9XpHSY0BFz6/g/1mm+OWvJFwAbDNFxPn9+xh
EmuI7ospI+IuCebR+bNm1npIARjAcv+w4hydFctTrEwLKex9Kn6R1rDJ7EXHTHpfNzcvy1hnIQNN
VQy9KW4ObFPDeytZimruA/7MB9KmfEDpUxHPlXNUNKXHfy0Z9Q8M5nPikByb+qGynz4RXBLnD9aL
96rVzSjFXJur3DdZh9q7dK5m9lhsOg/3+AhmQsQTuFR+nxbZhrS+3vJUZoI71kZn3tAUVM2Ue704
QxR6vGuydx8M6smbPVCwo/fuZZdjMAOWmSWgXxT5zon6f1qTNO5QsN64Dxnz1FsES1/IQe6//Z/k
X/tb+f4WAGb6cAUXmJEt7dxGekYn80+iGeUkPnfKu8bP5MK5TU0tpIH6gD+VqPG8/tIWS/vqAUMU
t/VmvGN7Fx1Lq6K6dmNSh0+MvOwxEKMG3d9+F7xHsKUSYYlzz0COOiRhuJedI7JUvlteHiiyR5j+
kloZ0R5RILRkkX2D2FLNcdgxOo/KIcCw2kG5RWnVv2ptvmnBOCi8v7MnkCEY+lycsceniHyGRXrF
Xwj9SSn9+4/6PNo7feqpay/HbZy23+IavBkWwJOr5LsBXw3ygUnreoHcoe7KRq+aXfKHif/TcRii
EYxnjcYNwDPh8ZRGTBHH6uTT6NjRh1MtuHMcIZmszOXb3LUmZx8hv+qZBUYfEzHKI5jfaP1aOQ8o
TXhLtOlSoz+yFwlEK2WKXCEzZdoWNkTZmYygRyxpnHVtHEWkj0mtNafZ5l/klrxcgy+q5vFJAV/L
1sWiPZaEI+z8iL2iphmJN78671B/rL90/uhjH6sVbM2JpiDxYqcsv5wU/Hvo4njVH5qp1t/V3Ijl
hRYVrfPHYkwyU+csUKfsuqKG/6cJkga/C2eZ9bFS7cYK0wbjmhWuN7XCO2YIGug2rV5sLMtwFFAE
qqf4HzYOMXbKFap/NypvK5guzpn9LtYjE6qOPR4G8MfdDqfdMJm7AS1gpfVxyVuM5TmgBh3yc6dG
jt1QoJXYewSL1bs6InoJC2SPEZk3muECUE9FnJVmfBGygXIZBKe4/VYH65TeDNtPjZOuQM+oURPw
25KtGlAwmTGv87kvI+a7wuPjMpv2Mzpx4b8cUBLEz2O/fPPVzwx3DTItuw4+giNN4Zkpm+ivLE7s
PHmkjJIPNw8rMv6XyfI8tdcOnzSKmNC+Vggznkf8Nd8y+AZ/gr+/8XX2r167KO0+r8O0KMBQ4MJZ
7mHMEAOS54PgiN1H7nNwYCIMiT/Z+DO4hkZivmYIOGBCh/chdxDpZ0glfgKeewFq6EXMXaDFPGYL
tEAwdX5xZdsIFZPi2FwlhWE9KRmQpBK70klUbtDs00batDrs7UqeFYHJJOHsV+VKa3NEzCRl5I/O
5AAVe67XsJRcJ2stOyk6quPj5RqrBOgs8Q7Kqd7M3EWjujtfWaG+kWmgpUu/1nvpIWV9PVq9XzoM
ErgYUs8x/btTE5iJtSpfj84/oG5AspH030GpV0zXdVsXl3ZUPLgl+yTBlBtxgPd/sxJ6x76hVUGR
xiWI1XtL+5CP4t9G71pGzMPyfTFH9UwNM7EX/J5uaCpCU2Ba6/VZBD83jG1y0+V342G28Ba6TnUd
MPSxcSpAikwquQ0TUiUjED4vzv0eVHF9I8cb3fbWKQObrBMThpCVRnvCPqttE9RWN2WhSqygoKYR
9jhvuORRl4qsHU8CfJLjP2ekFEt1t4VteJrhoh9HMPpv3CRsbEpsEAuK0Eg0RVwyiNMyK7xBy0uX
xnEXJPcFNn4dzAx8tf4+knatAePG8dA+FChDHVTa/1XT7k9DJ7r3Uv5+26Uzuf3RMukKSbLwO+YH
/xUmLVgCTodHrTIV1hrnUhNmiO01MKWvwaLzSHbwvbKPiqLp8kEhrVUmceYep6fQnpt5mTVUBefr
35DECxfyL1za1fvyf7vMmAHBDMF98G2VdR8nmhaOU3N9f/HiOcISvWod1pCOo017Nj+g/ZasaS3M
REmSeQZt6zdIKNZb4fb96lznViOtV9jDc6rB8xlvL1BalTQqhw1FHxHBcZ32IJs8V8CgF3InwPSy
RGpbCy4Yc1jwcKYCZC8H1yhl2WEwGT5AR6X4Ws5kg5OXBVED4NWRdJWGs/yPMX/aw3OOJOlluYPt
6J3H+hii9B0Z1n0UiyC6OawiGSt6cLJr6rjAdTAN6AP7PszUHyw9a2dGeDNmClXBxUSOezA1HDlL
qBA7p4oEiWpkCoUM6C5m0CC8IXTHpcEoq8KHV+uJwUplXNUQfu3z4jsbZdKeYgIBOJ/e1OuBHCFM
6SGa72XA5+w6+ANH9iTMXBV50XvJMZOpUUUntUVZoPxda/jLGU6BPTmQrBJCVUPHYEwke0wrxeVS
cz5hDjPgGNebGZGcWOdR3r/MeIZix0/SYBRJvluONP40/iyA9EUZI0tTu2mOhoaL+O+AelhZqf11
aDNd40rVktE/kERE5MvYAqcLu1uqwVz07H4lEkOWHMzqFB7QLtQr+Vbn/Q1r9Omo0DxgOlzRL1/p
VcKBrVhN6E4oGfZw4SprmJdd7/R4HCBxVfZMl7K5EfG8DTW1z32y4QQXT2dDqiEjfeqlKg7x4nK6
nhsm9h83FI3TeOY3fwVPK3L7Jy185SqgpqGF9/Pv9CNiwrDu94mVAYWY1tnI9CyXOCTllaUn8dmG
k4pSCUkWikZFdJEhb5sOFAG4LBWnj71VAFW1i3LfNXA/+XcS1clNiTE5BGI/Y/+CHCdFOWYfIsFe
ZpohkqtYcxnV0SG6TWtHRB2B18VHKnopUOCUplGJviOH/5q0xSFkWV4+r3zmJvF0zv6ySnUzrUa3
+/BgyoMruFUfMz+fnnCV4Lv34VOMOKXX43nI68mulII59jYCeDAy/X7pCghe6kKHolUOjnJoBbfX
crXz8KokvxyZA80nJ6dVtxAp5mfyDxslKeMM5WbPufgLdRq/vdLSJfOeJfq41HCIwy0Z4Qq/GjJC
S/O9f5JdLX6nnWb6JeWG8FJLkV1/nCjPcCBn9A9ZFzZSygacR0zfZBui6iCHV3F1tTKaPxqqPcDc
kxyvK/sIU5Gp18dcYRwINc5yWCScF9aVpcdV+ijCBZPZw+wmjpthC70baS5a3zH+5jNpNN0X7ZXc
+tEu4lzAw4rBVfl5gKMq7bfZnEJx9PGFPH95lhiAxFmkHdMGRfZcWlMt0X/YxrOghTAdu00At22U
dwaB0RFPhrXSfr/OLi6TbM0aduyioVgnaql0UZlN1HTQ0tZ7F4NkhVQFnO81DvtrV1PTXmhZK3Ui
30dxBISY9cot9JdZd27vgF8tJO4KROWo9AubE+RnAM9tOmHB8sbIm7JKEVqGp+Bdb5pCRAa7wlGH
cP2fqdRVohEamIz58h0qk3b6945DVwi+Aa0Ab24TUS5vNbEfhyhusWVL7klk06USHw1l4GRBism+
eqpVad3Dzfb8/7KenxLfv0X/FKXbZpBiQAol3I/+AqiMZVngVL0nDy62qSAnm2nPgr5ONidn9YPV
wXaY0XiN148ZgsKjIQneSk4KyY+sN++2I3r2sQEd365PnZZOAeTuD+Y/t4aaofXVQihIrZBsxuGc
35eLghX7uVuW6lFii1oo1abm/Y2gjiRabepsNgRkw4iJpb04EacuOUqIpkhvzptPlUosoQvu7bA0
+7wQk84Y9TjJEFowx2tklkDLu7cJ3KrKNz98zjsXTU0BtnC02a5/wckEmA81c6WW3k1tirrTOckm
100IwURj0nXFIAMJmJfiXCfHwYtwwN25ueklmgX9pJ0C5jDVswVU3xxJK/5MARHhoQjzqdeW03vb
/D7xWMkA0jAUlnEJIt6TKN4Q03kU4FBeVYXyYACqskHqLuc+9wi3RhYITXzowdlSYLxB++GP3Dgq
5CUSSmIbyr79XgdABcdqHdixl68mZHd3o6NerhUKN84jdx3jCoHMyBKPWSrPnouecxfu92pdbTQc
dwk+HLQLjvinmhRtMN45bDFNC0pxgDsjrUgSkFP/Yeo67PxFzxuQgS8QxKKCGvGP3yc9AbFM3YU9
zOWY9G1Twl0+DrsDhcPIZm1Uj5eUTkyfz7ccszLmVrOvHq/jcHFNLIflRg0uQ6aY0HL/vZw/ndxE
Mirc2SUzFix+xjmBjLDV4dp8v5oE1frSBbXL+ppSITUgnB5lmXkL6Qh8RI1JL0cewbD37ll/LirM
c0P5dAAXwsL6DM+ZQvn1T/2xFux95aa0GxVHZLfRjiujLt/C4yt1n6xyqG4yoZReAor8go+9u49n
VoTieFgGwHhJoEwMkyXk+J9WPxYnxa4rClWIGiC9QPsNC0bPnIyKMzOHet+/RzErnluWAs1DPvkk
iSQ4lJlea0cyahjLuGg1GGkRVqLQ+hl7V4eJWaAfPmaVpeC7McNrkNIEdg0SPewLPWdmhzuY7rFJ
dubM++ZxbgPFOcux946j329xMuhwQphBq/dEkiTpXvwFAAE26rG4dUdU5jMntD4pnFQ/sc0S/1zp
UYS2suCc4l/zXKRfhw06ei5az9S4ZEtua5gyVSBTfjMnjamcDE3vcLwNoQln3k20bnyJWYDHO+rF
fRe2gmuIvyliyq+0XQVXOsJvEfmMWShgKJDV0wQ78ngWmt/uU4Cjnq1BEur6hkcQUisfcW48OkDe
FlgmYlUEGPnQOXs7IdmT1h2jWx3REc7eqz8K0Ev+QsByTLjHNu0fMzo6PgCwGr4857mLgzoJERsl
szdp4wvBARcWDv2salCaCnHuwNUU/vZlDrUspIKEIiaQo+7qPt7K5r8Lpe7LBRxfQredMHsdgjLI
dtB9vX91Lwzm0W6+O/uo2qzBA7JNT/Q7vqfEWdQM6fH6R6cVxMI0SQZFCdNxDeL12pZVu/FEOAFd
zcEhQB3tdV+RZtrf3fxsNX5cfWlDOK3PwxWRr5rp/y/Hva9qZO9DNdFYB390pj38htbBiIEKKEnC
Q66JnREtZX2+WTlZm+k7LCgAGZ2Vwa15lR+M8UKwU4gPpjTZAA6i7gh5YijeUtwQnsrmuZiGfqKs
IjYLVWYPAkSLmdmqLBBLD2HN7Oe4op+3e3xS6Ea01bnAAIAKip1A35KOptY5f6JemCm95IQGK+PX
2Di0onRS5hNZ0+9/T07rBBZPPFjm701RpcWt1mstp28Rzruw3SU/NwEXYe0sh+6Cu2hdj5flkgzv
taaRzIIKW41Z3nSSqjQEIYsigAp+04CNQ+uyUSiFR+ZbnPUbUM7mvDK1KpQ5diwbl9HiTgRi84uP
DUaydu+CqaiLVv0T7h6JCHi7ZHiqKz+q/I1JiPD2pUcT7MK+I48s8Uxnf8+WrRfCo5Ar9Wc+HR1v
6Xwpz8ay91ISoBQZ3xLMXdeh4g4+tnpFeBZamAcMDRKBmApwwdOzY1W4XhspC78qm/Pqc3BAd/BI
eaPDee3d4CyAXYkQPA479y9RF0GfyGv/HMwDW28o0hWtoHycnh+0Vf6A3p9MpIv23lhEUn30G+Da
wTVTEwKtYjVP8JoOCt6RWMOz+MNTzdF0KazBZzlbHZEuD/P2km8V2XFX7EbwE79JJPzyFZZCohfN
cx/TfKoQ/R6cmaqifNEJ6l3Z2aI8L3prU7oUgRiiNM8AzeD6n4h6OiFicE78dyjaVqJlUEgT/GFG
iUSdVeTLhH7j0atTvuRoH4hH+1EXBXLF8Q7EUVHg0MYQejzcGmAF6UJs2GPTyu4WZ6gSa9JlrtQw
K3H37etlCICfN2Ofk7iAcyKL8Uzw6HNmCYSNCDkwJYHBD9OR/uFjdgR/SvyiTWeCvJLsNk3Svx7U
ndYPS9wUqpHSSkgGJncfx26HF1mOsk3oDDqUx+ejpLltRmtw8+Xqn+aV8CX43+AgbObTIXFEX1j+
W7I7ZGwe4aUIj68jyRqLrmSUk8Fq4TZ1XoToNCdEE60cbSxCnHFe4L5HL+6yEWexAARTldCrriw0
JVDWnh6Y9N8ha9071juBDFdRH6pNqGCQyCxlMaCEV1qZlAKxSYuHYAn/+SzjDL0FbEii5g/xwVKO
vZNRYrFPDxiu9OZVZ7XIIGdVho3Cn+bs7NAH0sXFaBTuyJzNc4rjR0wp5cLWEssOkR8+MszSuu6U
3eq/1dRfvsXZmTBY4VM2zueQWkF43j1K3hyVVW0AwI50YAvJFMzoXzcDneKjaUz0km71i/PhNXun
9retJxBFb/CORLalhHlWzF15+jelUm/z1lEZRfXyHShSEYk9GrLJiRjagIADhKIcIEHSOhmhC6JJ
41e7hm1VFzxMI/yZjTm7StxqwxXVrLINl6o13I1sXKWC/MigqUaEJgFQvr9bau4sAtZ1bhNGOFJk
t6bSi86yfceuP+9RbGCsNc/HmsBkzY+ZqMj60eQyO1LRU2lpgGNhRW7AAD2ERSsJcRiW18qFyb9O
XYezWgVlOPpG00pZ2T3Ra/iip7s2xgNkt5uwOqhXvENl7F9LtYMe24jzRm3dgI7qBh6mn6j5n6cN
CabZD9XDvIc7qhxhR5Wf7mmMF0XHxnN3w9opPjuEUyjyNCjklRcIult6esSN4BmeP0/0kkbimGEE
vXooxwfX9V5qMmK/WkIRq7eedU0xpZtUwgGq97V0WDqg6zi6/tGnD3xFsuyZfo5HHcOvUbei7Kfu
ksCSS3HoBaXMxRvTI6S6rUOa1gJ1adRgaYJBknTjt10ox1ZDgAOTVIt56Zi4oflFEGn7twuXvjxV
+U+qJ9c5gS7Eos/AuvL4impH9HS+TDQV7EvTITQcbkmrIkQjXPTdQdYBZoOgf0cFgsiU6Gu7ROBb
58E2U8Q6aa/jG+1eloK7kcfUmYQBiB4LewEuweGGZclNDhZInetssjR33mUcfkkxXb0CtxnJnmqw
jiAYgES+7IR5WtO5/27oM9j2McgejqxDax0lYSowk1xv2Ce0oW7ewXK9x93qfj+zbsSfDP02/oEL
VAKEK3MgfEZfWbdYw9y6KskUroKSd6rwUsSR5h446tkXCPrZucXPGGwCqIWBe+pSJmuJzdWXvmGx
GSl0FLppPSPbDl8Fs1FgPB4MWQcX5DQRsI6T3n8lp7vYG0LhKvtOir6ytLYBv5gQAezJIbM5pgnZ
gD9p92G9bAFzZwEtn0OGAtwwEHWNpMlXQc2TnDVftU60WaoWpVPiFdTyT3rh4mmDDORZy8hmhKs6
nLzYgcHOCeuM4gD5ajO4C9wAmL4PUkz+0BJruiM4YPnHj7m/AZJ7lIufZr6cC/d1NjqGv4mtPQen
XX/U1MfkvjWIaXFJ0t68KY/7yVg2BMDlo9Otk4NY7bF27vE57B5hMekJeE2SJ37n3RZJqmXLJ7c3
mCs8GGAdt34T8CqswbjvKKa74JJ8Atqb6cvvbJbH1kXeLQfZlhdFZxBWudYR/IdL0LpPygBytXwy
u5bEWO8zIqYAz/jVRhHB/iwSsKn41bU7+vLTovo9WfyvHhzsPHjN8kHv9X5B5yRf4czu4o7miEVy
CX9btW90jvf4hWbTggyCgIJObfuEnjeP1OzqmLDVMkvonSE5mLa0VAge3bkaTVgmlWeqN8qdsihz
cc9dslH60djzdq+QIQwh5K/neywVvrycbrgpPv24M2HoODQy97WlNRw2ngx5lQEBIEUN4/SheJEv
1dmj8FKlThzNdYueiXqrvtP3z8fflbFAy0zdhXPiism8Ftfpkvi0CC5EgnDXDVjYhD6zQ8lXqWjP
eIypaGBELT0TUniY5dKS39JbNpJgqXZBIcT2Nb8hJLNT7xV4I+iGUMd7Ron9+7TrxAHU8yGzB718
8VKrqdPRTS4xtRvIFy1kX8woSeWF9FXV5xRv00Ez/H5ebV9MjmSoenRnwB2+QCG4fkG2mUT0379M
bYK6E9OenbX9KMWBu69PElVP2AnWLkBSSt0yUbLHLgTZK/mbkC8JfQkKzvy4tOCH95chcuV+tcPN
xHRo6oJRXQJ/lWPUyyuHBlYD9lE9PHI0/RZi37HxNXIP6MbWHzNh+iHErnNnhSo9JiN5vYAeNhC/
tBaPNYjGkf6Oi38gOeNlZ5/7zf4YOwDP3paQYKE+7RK0IBFiGwpTjXgJJwZReUidmYOagRjZ13kC
5+lwT3PqkXSpAJNNzrKh9XzZC8wFORYCJ7EAMjmm4FnOUI3Gikwn49FIhTAj9OlF5s0ciw5cUabl
oGkGhJ2Amc2j4/HcsMFNaLBUEJv0Vd9oPZzZ4aUUbXl6aRAxO1Pdq9FQTKkDQMGhd7LzN+sVcmvZ
KPDZRXItsdShfZH0Q7GdGAB/a6+PJPgbVW4Z7082a1dNIS1/W4rvNcAZSptNhLUGT+sQ4e2mLi/d
g3r88oskmiSuWVwA0kqBalfqZgTSVZFLnXnKuTlXiXLZwyhaD4MJLDUOOaUKTNIIpNVPwmUwY2bn
4F8ETIN7i95Z2vpfw+JudXSEnG28fWesylckJJ9JXwRqHvw0z8ZTViyKUb6/Ol1GWcCxDLEGvS2k
uXluGtDKTuX6uKVsJWS9lz8Io5G/HbP3mcNpOAl0dfrseCheo7YWll4/4hSyiBYUcSXziJOPYqWi
EAoTJvjEFWl5G8cOf2ly+L/kgv5lMCKbIQtSUTcPcszxBogWJyOXDJzYRzByf5f5LoeTT6cD+ZWy
u+M7UulxqTYigW8TojCFVDJYjP/iGQV4fSvVwlVEWJnBnwjoyqr4op+t1y1DV2wCCl7o3znOiWLB
K3+GD53V53cSLUCbsdDQOA3ndklXwePHIFUnor8hBYXxcWB5rSizIRqniBZSbu5bCcyaOBpRoNQJ
aglE14u50it0UJK+P52KQ8DABu9O7F8jeDMhgnH40ozxvom4/sMGzZP9IOZ/fjUmoPRomYlz8lr5
61VFIzh1/tvM2Z5q/mZKeqQFNIg6s0C2b9hxhku65KWwJ5QBanUiBYvlYPAPZnpmSgAAPYivVvBN
KHAJoYV7hAvZ//V6/8kO77r4rWEVe7TjIxhiENS6+4ZqgwRAOTYyB+FGRSTS5h6hEppKzuEGOdUT
82jKvaNpUZV5SeLYCEb/q9XsCSuLPgzMxnhISEBD1+H83N+JRbbVfVQMyiyWd7KQ75fJ13CSYplT
Hx5qVwV5xB/cbMnzJCp2PwLtoDEwgWoLtx5XUBvibqMmckh8q06cwr4kHbDyJg8ET1gbbKYxn/Oi
IDIde83ckdBKWsFNxS85sQwYu+tzE8Od5GtwZEHEItQzXbmyxn7Irhh8iLMXe4stMlkzoOgwA8JM
AMDl+AEIWfEbFA/sHGX/njj3VYG7xIk6SmgZKlVQfuNfs2ETNdGPD1RKP08ZgGjxZbXOcZV2STrP
G8a3+9e6hwRcHektq+ZkK2ZvQzx/VmKJQj79e1GJJAEWGsRQOFbtjC9THO1YuSsgQ0g6hN22Spy7
Verrr1Q5gx7kl7qOROgSgu9emXIIHCpWSxhz67pCpGtcTfRM2/Q7pp5SPH/VMagLfYZK8np6DsEt
u+MpGuRiUR19uA+dsFyPklbUoPKs62dleAXaRpYvuQNqpzlOrUYvU/mVZQWLPjmr3FHiYitbCy0W
A+FKgOGonzCuRtpMt7C7Z23jsV9Y6JTccReN5ac4UnGjD9fM8EoeZpFW/rVxUOIGTwXCfupIDk6R
dHwd3RKeFabf9kHSO2wzXqQyXYC8atwE/oAG6xDQE//lh9ETDsY9g/BorSvbZ+gAFkDbr7ZV0qMD
uu/qw2tmIhylK1AkQFCFUtHmrNe3FGLlsYudxk3w9pWPs8GUVzRcCWvBXCfMedBDI782+gNa6lBD
dsy0Bmn1yNbBSq/42CUrj8qhbxuRmeFD3N2AuixvgfIHWVuObTwhRfcDNjC1wmB+39A/EKB0b0Jc
Gf1ctQJAbyjxxcQsgozpsUamL1YOQh3OwI0RHQoEQ/YsTx35bDB32gKK/Y2QXdFmroPEDPrN4oDC
mO/+WlMsyoi+Pn/xm0OmCkL7Cjp3YLN13jEeWfMuOhbKAIZr6jAgX6YFkGWMYp/XccXKylvoM/Ax
o7QU2LGnROXhIoIMJkOxkqVgV6hqaB4JmxEHCRHJSM9OI4iD1jxYaEldKKvNz2mml7DWmScrJibF
P4ftrCNVivEVmhWpDtnkeG4WM62064oiXVRwxwdn5v9kXzGHuLqiaI3WC87UTL+D+sBjpcWN7HAz
vDb/NCuN1fOH+7BlelkhYAHz/HlbX/e0swGDgRHU5+4Exq6X52st1znHCl8LJW6f5aoboV69PRWt
9W9AVYqsnr3wa5Rm/vPeA9bmKbQ81v27Za2syMysqRCJmqW+VlmuDFd+13+lGcOnNffMNT5p4eeC
9dmbdK8Y/V/+JyFVeKYcj6d4eI+8rY9T1d0u94eWmrXg4RzK1JqPmBXm8lPoURgO7aEf5iEeyS2h
mTl8DTT8A0PFEhFJDm5nF6RiYvTow/BB6nRL2RTTyCp9Vvb2JhnEfcQE3fSgDDpzXf6Csxk6jMmb
EZjOBpAJiVGFubZDkz6+z+WRL20cMpV7kTxqHQxMQnRSG0KFLUfpC11R7EO6AzXrhW9y3hmrmTA0
jQigJiB+JbxeIsep5RYNpcVB09YdkXfJ6q98buN7kzb82/QsIjQJuNq9L+wA6gRQ0soCQwtrN6dz
fefNbthCbEKyiTsNKJrzuUuPpCp4gK/aoyFya2h01DfxhguOypnmlid1lntS65HnhXySjtKQFE18
JpHudVDOdCWH8UF2Ck8IgUSn5LDBAA95RcWehUk1AqooXCUqDv8qbgF9ylX1s3PFd+dRR2+fU8Ju
pXlFZxqjXN0mKJZwJzi5cpRCfDkHko1yqydD3tohH6hD0y2770FrVnh/DFBqhcKWXKPvxr6cMcMu
OOD8XZikiZI1raqI7gPW7ayjCGVOatLgM+oTbBPQL+/iO0M0QELMyAT7gCZZBL8XiqC1evEHCdPK
g6kA0E2Q7OydYa7I33cIcP67TcGIdIlwdIrTybGFjSGing2MMp8iEzDjDSyvbu9ZLlB2/3axWpkE
JyGXaDh2WDERvqfs4E9uOwTI1Hju5qAZMw+B2RgUwvtWny6CvWAoMuJX699ZXxXeM2pT26oukYhc
JyZ5okutndWk0ns9gqqOEQ+5SW1b4yIau/dNiPaSL9wDd4KHEBcCrKNqN9Yizp95vH3s3c9hcc1E
VDirgKG8ZrLeyPFNVP3pWa9Fx8IyPPetG1hbOfNsFbRW08TBJTf2kBqN2bSTO20pRXadalKifBRK
iCMC3NU3S0352ex4PBDvBVZbyYyfXABI1cR72DrT/Twt1TUjX1FCZMGgZ8HQQv9MF3Zdx9QMww5L
PfDUiz+ZtcGACZxEwJgysn1tHyRWuk5NFMER3IfctsPqELPIMri8dmqr4fEEH6bdIgWWAl61UX2l
6fj5FHx7jC1W1EMd9AkDkl8HP0BgBmDurlpHlm8WOROF98OtJDfWQQpf1skZwEvCszCdUydpwFXF
KmyNgWHD5y4QPh3n/r3OR7Jwlo3x3u+oRphzoScLOERrNaskFPDjssOnqq513WqJCPWbyUAWcaB1
DWaJHkFZNvtxje1vciB2kQsv9olDsFOHu6oiZ6c7M+Nos6UDc82wfVAMHQaFB0f1REPfgh2jkIs0
uAafbe3vL7YjnTaEdtbnAgoR9gsAvDl/EEumQJqAoXAqjHUVmmBQ8eV7aD6sZQbQFnYo/kpXKpP9
dnaIZBWOJOvUprcemvEONY2UInpwnv1783wwRlb1hyRLQtEpui7N4bgywwcOGA6ZQh/TN6+W+BeC
AFtF755p25R3WPQRJ4296EdLke4mMfB8Pix8l9gxiEKIi+yW3TrvCIdoSUM2xWXYPHyDNIEMpEV5
qsNiIgSkAjpe3Xcf2vmZBB+WWUuRGOq77oQByjb7xEGHSRhR5LRFawTi6bCUuL3fpY8gWIK4ibNR
tYpXhjBneBI7wuGrKWUarzoJ4POjHMMvc5I/HScd6wvQLXNcCPWb/wvko9HL+L6Jl+pVfamuEu9U
IVqyOx3NKT2cZk7UGZiT6GNMgzExv/82DONRwzFbVK1cn7ijA7tc5Gx+LgNr7iZi6mlFkhe7tNrY
nOqm9+RsthG2EOxh36TXGFNZ/z+HD1UokRlKlFzF3xKquIz76FjtifJn+2HWG7JTuoYvZWn9wee1
rgGMYqjBBBlPlLmySZ6Z57+Z+rZ7ENvnk1fSpF0kriktaNs7B2S8qaaIgh3DdTW4vmtqFPJmBw6I
ukaRInPKk+iwa8bJ0F3W5chzpe9D9oBstQyS1UkJ+y2X0oyqAhTM5sJjxOKjsFX2wl9eUobI/srB
Rp7HhaGeUzCfQ1NjJqWeF+nnxZlXzlSfLaOacjj23L4HqnvscD3s7e2Oph8zewofZ56SVhuPDqQ4
u7TjZOzFl9cMuz0pp7fXpSeoEpLNpqT961DkddDN2jS0efWkIT4BHS7n/IbB78+iV3J/a5qx+X5m
gk+vKdjyDc0YO5Pb+Rve5Byd1kwMS1ObRA1TsFPEphD5Wcc+26yCZHNzXaV4FkmxTsdBqfcl+0V6
Z4J2PKk3kfapKOpkaRRQylJKJVUGkNwNWkcT00/kjrlaLi20hB4kYQ/lSf1GXS52hRngOTtaE/vR
OJ7aBvGJ3yiS8m0Skooo9YdgdDl0yuKS1elvFHbHkqqh5xi633HcUjuZYDfUcsgDyfc1OzToaLin
NhdiynMvgwhxdO5SBPMGFYPZHxnQziE81Av/hMLC6bBXzSRDQVb9aXUoR6KTp6gtLNhi2vf9Yg3l
0Qmgt+EE9U9Kufk0DPI1tlSyVj/F6X8LhFIPRW3ec98j/EvF8P6e9tAMqNDGykJoPhtxxdWvOoTw
46/+sahJwOKXA0sO1xWz+Jjo5u3W8kzws9kJHR6xZ41qJoDuP5W8zF2X5jLZy+jN/1P6pLe53ZL9
nW+vErDPXTIkQG3vizVaaLflW8m4nccHE2RbZdJHjxtf6DgtcVA0lxbvhd6FXDtana/MTsJMZZhZ
te/LAg+cmXFzlajmb1rs1cv1GFr+1234/sMvFUEjw6q7kJpmHd7U0b11YbdnZnq34zbtJMR8/8Q1
TbI7v/Aum05Za+C/OYnjQiiNYM8utpkYesFKe/Xl30dBHfSE0TO9s5SNJwwhvWH7TIxwCsUqcKTY
cLfIa1VikIaE7xhUU+ugSXWOG+kRzSI8vyaMxV98pFaB1P2WMmiIHaYJtJ3TsYGpb7Bk+lOK/eVp
M8zSZSqY5otuKTFvVMRO3J0c4OEa0QwO4L2O3zmNmNEUBw2tdLdt9PdnEBZuJrXg4o5sgS7c8wYE
1Ws/MjkyLSNS36PwdFKwOhaiJG+E0MFQS2TN/SIaEwipvdH0IMUlhinMRVrfRvjZ1NHWYA+EnuW5
eXFj9dI4LxEYvAWUfyzCDSB+OaDLoha122c5ivZHYgcZFEtaH1rL9oiskZ6VDXnVfjV/HD1iiAa9
qHXoWNSDZs3w/W0d7SzHeH7/nEydJjGKuDLBJoueT2nXsrFI6aHOROIHnP+KDN2gPPpwIoEu+XaQ
l10wUwYDa2mwix41MDqiEfQ3/1w5vp7ewQ1qMScJiCTmwon2NMp4GgOdL+hMk+2hLu2E92EX0pqu
USpXRkazfyHQTKV2gQKlWbbT4/evbwhM7zxwc75ZqeRkMQLSVRf3Ddkb0lSDBxgrxqNZa6B2Epdj
acrdSoIu6knkwOVPJVc67OgwLQFPF+6cUrlFbzDnl+B6XhUj55qrE0etemAs7ZJefMLfM/Q2rhP9
wDb8v/stkb3qf3CpE13wDofbGV1fd/gFaoXV+gq2GQNnHB5q4ZW9kuTm/iILDK4Z+FY9aBXohFS9
fkrrYOlC2Us2RyTLbNQMXBDecodhh2f5xydS8SaNuEpeGkrfNaFZDJ045AKXL+MqkX6b0OoY8ee3
N0M5yb494IdgqUPTjwHmt3bNgNBGXU/v5epkns18eb139+2xyKo7DJVE5uEeZVGEFXeZMY3f2MLC
JhntvV7WkAEPLXQkX2cwyAUyWj0d01LfdZ1krug0UvLiWTC/U2GVzYM/jZYVAsXZmj7GC3wuvd8g
e+fFKKSJvJVu0C6Z7ph0M9v9lHO4Y4YbQlbE+g8XvVzsmwFEywqugygbsz0IUu1k3Z2axODCsUgP
iMI0bcHdQd0fNZfmAtsC9l+dL7CDedf93pa+SnMweswiidGEpC3GswEVmsARSPs0Qawnmc6L4aOQ
vejuYIlp7gdmuyVJ/GG/WzHV9wjyXyEGiYDm1HFnHYT3it5nPG6TupO4m/9jCMZ9iPt/IMTOWfBA
dnt71wVCLjwy2fTKZEyRljyqhNgMaL6JKsT6PQ5pXf840DoTPrsxeThPNt9wWEs536cJOs3kgMok
TPA6qbRwCor1toO4Lahkn2KVEaYRmWP1ME73Sq8DYKIyiTtRePrmm1PsiqwqQNaifHHGnoCpuLk9
C43tRc8WEomvLc5RO77gdDnw/LkmNtEQQQMCZyN2lBdEstw+NG7SXFO4OhUbLdjQCbVDhjKPP7IB
F7tf7f50LNCD98QBx/xcgmG13XnkZiAawbUyVCcjy5/Aup2NO3pN/EqG74OZUrJd1xFfdpZCtBTu
HEUmqpVecYfIfqe/YegnaaXf2nlqW/ALYvLP96sVEz/YOg/PivNM6PwZC5/7h9tz/eVa6FaAuT0Z
Nk553aT9T1AKLFq4tWr1lwOUObuXPRCyb4w+hkQBoh0OWwUsK7NNF5oCBA2Mz6nrC3jjZPzLAdiy
FDZvEgX3Dt9LKRDx/5EeKXIf3BLzPiQoKiwn+GZMpalMKn0b2ck4rhnT8JqzzCIxPq03LqaJ4HHl
9aT1GQO0smZa5ZaaJnKiN1rsqG1hy2CCpohRgowtfh2i2rg7Ww1JJEScNZhClfzDWksc0KhFj9dW
e2aK5ssuMA+HKtt1DLHBHpX1mZMc6PGXfILpPGO9LLIKlYRaQtKGeReE/SEbFMTdpGTy0TXQm0z0
QAC5lg+05a4AeN9eAs5OkU7t8lmj2pu1z9PPzr+oXy4m8eDy5rUFbXf/ZqB9c38eyoBqD8WamsqE
1rG+Y6DVRPvC1cv65kDtF897HwkKAxUbq51UtUy/l0wiIQOhkoJ/LGmx4x3CC/yGduT/iHnpOT9q
baN40gY96vboFDmipYtNdrzgOO3Pzt4HvGvVXL8ilIU+7ltpt777CsmE4AI1YY0sL7RRE7mtAg5W
wVlX6/4ey9ZSXtfsL1PeuseC/QZYnpjQvcAE8i7FSrDYuoW4PHakWoYqYODAb07HfXEg1EEyxbfu
nf21Kdz8KXUXHm9YuRpEyk7UxoWO50/E2rnbQ212bS4zYSFhX6v9ZoQPyHzZwRMh0zM18ES1yaa/
PeSeudefOVBCNp8RfPT7wKOGUr4OPtfKDUh3ZAa1/dEjqKG/RuZuhZnoSMkrQnEDnzwjxvh5+9ID
O3Fa++zOXuxUgr53k7jSTFFG4LjWKDOgR6H2O7XR7PBNce6S8MBczYdfWNGiDpNpFOiCPSO6HCg9
wGHbxR4YS8M4zHFHHKI4pvAPmEXAUdHT8mNuAycUH29ZYO3UlFQKt0B+7RbSpvW5Dfj9Nh4X5PSa
vEpotnYsVs6qB1Ya8DM7Rfusqiuske+J5XAxlEViGkPcgOS02X4OMrs+1kaD2g/U+7A61XtpDGm0
lTOp54DqYC2BOkSp6MShSdvyew6wbj82BRfWTDrc9p4qx4N8kuODia9tZiuGdnFF9u5MZYie8PC7
S0DP9luHLsqtOj37LqwujnTZLVJfEp4DjMx1Y1dO4F07S+cweGakynaj39EN1HMFxeWXE3MCIYiX
8PYzcaMlS3OzApqu+gu+25KoKQxfbjerKCUHGKUlxP2r8nDriSvHHYTtaIOiLXaNaAFWRdrseBbi
yt8Z7NpTFXtV4nqzx2dOvspXz5r8pCZtjRGJ6L9eajtvJvKLHBdrE/z5FR7gxmd8YKxumgsqiuPJ
SbrOS0HWc9zJtVURx6AgimYwXx7a6r2q9cDB0xTHeD5bvibwrYPATWe46c+35KQ8+tRZR5Br381F
FcFuwru2C8E4gPg7U8mCkruB93Z2KANVv71/Njfw4CZSOzNeIkvPeUf0CJncOHRABS9wUSP5qinf
Nipi3nQYskJd7Phm/ULA1oDpfwmAmAJLiLuasembCZV2tz/eWD2qxss2yA5cmUDthIjbqoT/Qnzd
6gJy2uvST20rsW+sMnxgZAjSaL0BVg+YkWlJXApctES6yEdI/YvgjhdXvUETgPzXnFNpLeMW6oL+
Q+gcmLTyGZGHGFAAVANjdyhYXx/9DnwI5sXiFSt57VtMj/zp1j8m0uwQkcEcp8ffAJWL09TIoQE/
rLtPqSH1StwhQhS5Iz6aVKXb/1Ykq+Z/SVk9tDdWoE7VOKNSgzJHw0BEr/xAsx2uexc6irj5/M1E
5XafClrKEr+1dJZ6AyPIV9BDqV6P1R0ADCRv87DYYKuTYqOfV5aUUkQb7xJKr28tzKuQSaLhgm4W
GAsSBPfh98/KlPsU9KQPSr1b2XgNQKbHw8jUijow8DIntSi7mKtgCYv2RgTaGXsru8GcCb2Ru33R
/pwJJD/QT5oL0Ftpf4GkJZAGO/y53pXaD6tlG5k2n9TIHVXzkfMNLm+9ETQ14T8Z4GfQEX/ZNasL
pmGL0E/BvEN3qTIedFKjF6Ww/nyYsOyXLp03wlfkssABUhgZGZQjT1qlQZ3CYc1D+6pI8qPhMiGN
YKB5CxgoUN3DuNERq82uG1C2BiTfvn8+X0qzJfFYY536/Ch5Bq00nBJN+94lu+7f0A4ijJRK2ksr
wEbVgYfuQbBhPhYO0/mJvOJkfP3YLQigSAgO+H3/ka+t02YY8hbU4D2fNYaoM3tta2MEa9orjT/Z
CYExJGKxe13RsIlENywc20nqX3q3psH4r+Q5uF1aAYNNi6FugkWFNaEWtufeS9cAWDYx54Kwy0ja
ko7WdiWAnOFOfiocVdNZVAX4i6/gsCleWh3ZPIhtEsIdxIHfuRzwsKhzt14Maf14Lb74F2QBhRDU
qtyMmeU2ujy2qQ8tOvVP/HHDyYbwIWo2+dQrKPsTTqRcpoYMyYomgynmRg840CAHcTCl7slfz/Xn
nccskWDamOXMwNZyzh4F4/kM+xcjeup0vvXwM4o3EqnPqlGd8+5rJWHD933Wzh1EuRB/byNeKQAU
nI/Rvaa/3Hv36VqNCbTo9SwHz/5McD8QxRn5uOOOlaWUV7l1Df4lKox9esTm5EXqXizKwS6yVGD1
SpPOcwoO2OgHolTq/5stEb9IRRULTdSmldEGJSgWeAcY1pp44zki1AyCy1AF/rRaSLBiWOi51Y5z
qb6k5Ksap8Qur10F5XmdOFjhVzyNB8AJNQ8Aw5Aq32woogsqoJlCKF4EDiFEtvRlgI/E3AdKbkjO
dXozgUHESQuKWRtdnU/VP215fyHtlu5LQ1XzTJbkn7ubOJAHZZmuxMnMUXLDNh0xHSZPmiTXBfrI
qSRkYjPMc576t83ymE7R4dL9LOah72jioC6mq/thye/mbZeye5juG3fqioHbLZb7TP7vsuVsHwDy
FhQ2nR/k+G3vw5HtBxVVO5d72UosVeRYrzdogQPD1rJj4boElQ7q3noK6yJRGDq4dGLtdpGsuUan
sOAu1dLARILna3QU3X5DwD8Cm2GlHNWwkkz5VvkNk+fI/k+ih7dUfgkT6jXv7kaONH0q9WzWgNdd
y47DvZ1BtcLzYS5/HubOQJjfs9C5Yj89sQlIt8be/d81I4tMuIk8in15gME7UFwssKCssSTdjTIt
a3qU28EFzUMMZQuX867PjYiO5YM0FfsoIjFM3HZ+UR1HZUHaTck6Jpi8QNlegYpDBGKRF1k8obOt
d4fvVB9KODpuDU6GAgReagbWhS1eePTWyPZkl2otmJOTQw3xyNkgeZLBTse++s0mIFPduOamfE9y
4RC4/F9N8yild0FZOOuPfU7rjwUIIjTSwonWAk9/N+CsjwCLhG4+1lTxFDrp2y9+kOBUdru4BdZK
NAeg+cuE3PSL+FaY8fCMxrmKwLMuO6AaQIf7Ps5fukh9Sj3MQGW44PQgo8BLWQmyXFS6xeaWxWzw
FtOeHe+fmPsybRt+yvAjqlpshUXpMbQrBVAYuQiotEdWzbn5z24ly4t2KPQlnSK7RF/vlwZRe+0T
xkI4bu+/jXTpt/MxapTRe6LcSLT9c2E9hzXTwjB+FKU3k0+jHZMdsaufjtvnzCoclk0zhu3hebnx
1MJOKKEzBontIwRqqFSKLuoF6yMQ83+P0e1VyK1TRDfy5X1S3xypVEQ3XicjA0RT0l9gbw96lYNR
x7I91Y4jm4V26CI4F9FplXfTvK5N6nqBGATzoQfoE3su9I3DDVouzIpP1VvffNjRGCFUePuF3oUQ
kGYjoKGHjRGSf9kux3A0mRDI0GaJHwqU2iujkwa+eOiiocfi3xJxQKTWjN9iYUjLQcmLGxwCx4DI
J3+0JG/srvm12BGsJaK5OxCDb0wHfDIV86k5NPhV+HcR8iK9Pv90FLks31mqjDhWEb60qkBEnXuV
pzXUFJRoix3GHOQPMg0VvP1OywAjrwGOURBy2P9WbW8eyGQpsTXmNfVKhJbtRAcHoNBU6XxhCfI3
Z8/E85JLcYRtHEcaW8W1q4ECJOWPR5EtCfZWDIbytbHRHK1q6UDMgnL0GfEmyCHoUTR+ypAs3XRT
wP/tAVlP5sERrlEYeGXc1lmilJ2RJl9ic1kG2c5yKKBi+ypNRiDvALdLdxCUCa+mPeJl149XUsjr
zyaYYUeOiASG7pm+LR3o1JWVye/W5V2vg1w39s/eqb8vD/sYUi0q4XBUFCUrjR21aKtvltZhc0jP
g1/9Kyc9pI6E6ecgQJyfegdmvJbaY45CDR1j3Jk9FYWqhAS4QV7utx1v1yPx2FRuvUoFjzkeesQ/
rGZdVUNxA1rxPNUUyQ3kyiqs86hIpcLLqA9sp2554ysvJRuLQg9XBqH2B+VBw3yvJdIQkdho3eSf
+YrEyw4PaCpfKl3c4qudBwj0JyfRVUVnMV5RwosWMoyWNzaxPCd83pUa1wiPG+C8klV+8ad3qOcv
gP0nfDXDoCLCO5ms8TqSX7KJJdaiIMTVE7ggRwliQUXqT8VJZQsKNV9iT6TaodS4X1icBinmUo1b
MT91LZD8nC3E8dUHuF5WiFNIkzQzMBfRAewh8Cd7NwcJPqQ8o7NLEj9TNc3yju5kqGToXB1xn6dt
JQe0QGC6FQJCs/b2RpGxc7+yoWYLl493h+HKxDlwIpOTjCFbkW9kvKPv7zfOZ4FjPe5aUMSpjHgp
l0p2yDHcWVezmBF0aKmP9FVSxN6wIcibKLuadJJRI75/tLkfArQXJbmfJcu+BDCdnyPETdDFU5mI
8ynmPqtoVGCdFPRz4jIOMYcAKGOsgN4vNmzCwb2NVI9G4lALobNv2mibb5ZLkCek79YpVrwXf4r4
pdLx5ePsfngUSh7t8Elch4Y3cfeh6cvXJn/44QbskQM+EA2K32DfIviicvd4da1BH5VUCfWFnmA/
wSgI0wZUIxEEhBIPHFIXxF/c5jbI+6nr6Zn9JtGbs7e0ocTAa24pTbsBYXcmcRSYXzEdavVMEAEz
OPb0PPZMDDtCVSQk5rj3htGOTM+wyUMbsyan2jSUwbj2RZVqz2d+kbrOmr3PeSxwK+qiCTZB0T0F
f0pNQCK1ZNhgiBW0I4O1HEFIlYCln4BY0kv7lkvnieFA1EKcPnrufbxGwIdXUWR4But2MwqSg+IO
YDF9h1Aij59UaY0lFwbl8D9WXB543Fah9NPQolWTiF/dtmKRBIvW6RE7wlZlqaYSRelj6s4z/T+3
mqPnJ91BmfZ6bP5+7dRVFPfPWE1zoBImjheJzP3oX7+juyqhAzYwiq9X5kKY31aBZLFTZONhF7Uu
pwG1pMbHl2bjcP7eVoqbHNseI6EklhJERfqyMk/+PCan2lkVVU9+lq34ja1QNvoYZjzo0mUABqA5
Mq/zh1OFe6ARlCJ6rjDA5fUlMG3uvhuGp46+3P+tJqAAb+S7uQl7Nw6WbR2U2FDeuNMKLRQXfG1M
P0GKvv2ClmGRJxYgjjIFh4MLQK5+e9v3Z3U/OGExuNr7JfgJ3YUhuEf7bl/MJ8rmtMP05uD/xB2N
RLbzzeDRGZs4tWUQGsoN/4b6zCKGjlNaOZ/mM12oX9aOfng10H/nadZ98i7PzCGlzJTTozD/HuVn
b4+YDYCrSL/TS5brF/oRSH/TR17E95m+9dDAV++/hZVrnx6pjClOrVbuw4irjKKLbjFdWoRYk3t7
rkAhTwiFWrWzH+aMzR7z7dkBy/upqSnuH59s7qUQk0vfnmMS/2r6ZiAoSj96iCz50WjyJ04wFZ9n
sJZRJXJeycvRdp5sGUQEzc2ique0p47qMBPNUOcFtDr9qCeLl6KBb7IBT0vpKw7COobFcfUjk7QZ
r9fQXKJ+NPog39mArHCaF0QkhH9NhsLhOVFceOWS3GrSY3qvhHYokodBv8T4uZYBa3mz18BXtPIv
6qEFKsqlLvAaar8jf/uAtSN79dXySMVkl14GVKE5QVNrKr/uP378ji/KC/ykH422r8Aj9oWhJcAy
YrZ16VQrFbOxfiEQqdGCnXRX2vEPuh7cDy04MaPxlUjlwk/XdmMfTTdLhy3HwJ54Csu+PDeXTxgp
d71rMqxrMH3/OxgFwESo/dBdAE15LSeYaDAMCPna5hI+hFtegz55pJ9rBp1AesILqDlocM7FNhVB
HIXhIguvPnVdp+lSJIDupDVpxcME5LgpYvLBpdJ4gjYul3vVWMBDXR3cWkbx4pgjOCvMcChmiq4K
eM1tAFezVPDgYfNsAkZI6zM9iMng3GSp7RA4/84oiz1eI9yRNgir3aisrygW+gyFl57DujHT0ngq
snMwvb7aeRPhDpuHi+NYREpnBCTpgM8B7yMVPWHhtGRVJnyGEhEygpBFB9yd+WJD3swR0PQTYBwD
boI0UD24yo7BEnXCniUDllckNWjgqnP0M3ruaYFxIzXYZjKSzu5+6WuGh5GrpGjD06o7aboL7/zd
5fVZsGYPQPJ569QGt0iLqr/JTuGtcIbkKHUD/m5YJ5YavCU7FfQZ8cCXI5F5IYpRes07Yolo+dNQ
QTrGuaSkT04iDSK8/Njecrs+L12DCZ2aGifhhbP1jYFJBaKvnP0CcJ/u/QkXhjz2rljX1tA/xxxX
5vRMBzePcDoHYDE6zYWJ8ukDZZjW4e4uG6wMLYK9ADz/gD6AXgx8bLjXhhFA4QtVmwGT6M4V3adz
d6fyDO7YFomqyR8GgdoA5qCrpX9HN7vYwDdOmRdJyIgqVn8gaH4OdHt9xqjLftIUZRBUzm0iN3Z7
tmOT1iiN0cZC584YOPyqyqVgdrEsyNeLKMhCAG1IqQ4BS9KlA7fGCXm0z22g277a7f/FqubUYLht
LpUPhztVIZCREhyzj0fZPV519A/dR9w7NvlswlZ3coRqAKPaw3TGtNKnb57S2emgrbuDx2byvAfF
96mpk2fNA50r+kKXbnQr64QzWbUMOz1HbwfKbBrrINyZtj4KH1WUVCLSVG0kfjwDQBkUmaMH+XTH
ejbzI/kpUZY/OUIk//4MF3/4QrRc/WhYPNG0vAs/SFx7gfPI9GAAyP5zJLEek52lMk16xsz2MeNm
Fbdh0AWAlNqtGgIwvSYKnANfjFP1E3Ykz9lHbxmEqmxXTeJxjY0RaxvQvYn/oOVIKsEh6KSlyNif
dRJspRJOGBsLR+NlDKOz0RySvENNeQ7PxyK+Zo7+k5Nc70XtxyJN/sYIZDuagK6acJqxqDlb+de8
9AzlpRkhXTvjzOPfZn0IUwWnxMNfPOrqJ4EAy31Iur3MXLIHdmzuqulF3ZCTFzvI3rzeREXFPnoW
UTgCa3WO5qHMcsGPG+pM8gb3y7ruAT7HzIIMYxOplc98G8q6WvdQ7Q1Yis4AJ4gF6vAUc6zhyhNk
R8iwvCDDcoFDTqYA5lz6GtIAWQy7s/gflij3/0+zjTPUtkEYchlVAah8CF0xsaldeD0lnI68onQW
NVzxw5EnmMzlLmT98kcQ8ADSFYO+KgRSgIYUgIjboQMRfZDbKePkBcArxbKmOn8QXdKnv6eaBZSt
3bXs9zjOWpfXKuFSutX2gsIoGL7/F3lgrhVZ6L4lyMEZ3xdL4lmVCVwQYrNcKq8uBxSG+OXhzZ9Z
uqNiKtSOkoUuihvX2NCuJnPQ8f77/wQq+xFjmF5fpuYRUU2lXhW9mx1tYavGjzOOxUrLjMsXQxO+
sdzZZs5pJvgjyaJuIuxWjg1KtJI0cW6mEqYkwer1apUT1IxobZHerRtz0wI5fMhdWWnafwxJ8UUB
T1nJ5E3U+tlOFLcVA5yTjAYI82t4Gz3QgglJBlvpBhTga1gvz8k8EpOoZAOTe/+aGpW4nboKUWXx
N1fRUuw1HueS058Fq95gouYhdE1OpL/5noVFH0+huo7IYXxxMRy1QNXpDWczI7aU7LDBKmnjtwe3
CJ+ihtyosyygOgRUgLlKaJ80K/ooZpP9mEp+i1094LYaaPIh2AAdjf32CBEhGXxAC68V2/5JRKZ2
ZB0RAtECkoXbxPdaZjNZmnz95WDrkVPmlQKecrTszEHyivyslv5n0TnI5CEWJyC3bM5MVVl7D3I3
g2mRiOvaFbco20WNLhptrYRPxTDi5uxv66MTvrplqNMr/dCSmtC7/nYdT+RMe4jZIMXvcO5thgsl
C2znkDRNTh/Otsv8sN9erYgYbBvml6/UJUfmRuO+FWwGuly49Xv44nTfJEtB+1e6h6eW2RUQ/pRr
iSXpTU6ZuTkfRq40/bsaSWqycFpc9hbXC3TAoSu1LDUhEMQUK73UYUzGMnjqd10L7HZgLhXJRD2H
v4SS1QkwCbOsrGrM4IomTh/4uj3OjtSXOAmwVsl0vjPGZ2hifFw/PJzkW22z3BPHlpsSARYsxIJR
arqqexXzhqDT0oBSa0h5UH8m1IjfWNsjkUKEcEBOylyPfrkkP18HTCpfDDWHQ3pU/6X3oHosStJ9
MI9aVuqNVKeL9k9Sq3C8Ioy+qudjWDBhlQjuN071EVSNfW3K10bb/HxAC2FIMhQ5yZpskQPOvz5A
ct2Z2k9PDJ626jUg9eP6d9b+QfXwMADjDt6EIn/olVbfFxDbwUlLUc8dYwzjb/MuYEeVsGj4dfcA
xSFUgP1jPu45C44GgIVxjK5fC6YPt9n1yeH/dfyTYZ5FiXTdnH3gg64n6vNPgz311atDfrqYcCuc
7NQsYlaDVmrYSGd0yl0DW2ajFB0p8PZh3L8zMyZmXBfP0cWl21DR7jXDZRzQnGVLYksGhGVZVsto
E8obL6qgy9dOzW+CR8Dd+aseCVV+wBzTqwOGQbxVYoN0dtXKKu6aXWgHImf4s2HiRyJHTJ7I4PLU
HJGE7CttgXePD0kZCfkGl1+x8oGJYVrqESqyRxdfz/UPX1qqmp+7N74causAL/Rv/jkqJn8BMPSw
Tw1NToO5UNEyzit4FTa9RRgUa5B/Y/PbC0LyOAU0OLQ+3MXuyHgFn6FRti/UX+wIIZBBQ5dxbTzR
ffiJqCpx6/A5LiNTFkQjJ+02MD5VhaVXM+aI7jq1jQDJNV5WaMSw6sbcvyd8OWSkoofpGi2eb9x8
Wv/QZq6RP+cVIxPDdneBy7VpXGfz7P01d469H9F/dtRpB6qH/Qeuh20cx/7nvfbHASmXVPxmv6NA
MS24csOH0Tvh18koBXXDJBbSFMzOsBXbpvkQmo2c0H0s7vH/lVO1Zw6oleFEpX9qv8pbNW4vtqBS
/wD6+LGdCoF91d9sLWAirekeOdLcHqhUnzK6yjthTPRxU3zgffe7konD4AyPwvZ0WEQOhb/9RAp+
YlUklyrOKJPOKvxjFndRVDY5saTfaVV86nk4jJ1vne+OUzBdMqnE6EipAZQIGVqwJG2kpo1LBWqo
LT3n1Ne633IG4hrpEFty2QPRBRYQYXzvO4mzCPSLATYcN+e2csQgq0XR4Py62+2R+VqXnoOFIFAS
aT7UcdcrixmveqfM3UtHwy2J1JcjEkTyHnp2/+aDee/yUrwblRfrU9Tv0GnbTiMcmWuIai7VmoI+
JBKq9YJVJn/73gJ7rDUJ+xPysK3GIsQoEW1/GUhsK5MKhk6aioiUkSaLgrqUgVwdxjM3dlm13M1a
xG1xeKhVub4ixayR2oxQ5iz+jBS5gCa6z6s1FR2NsLHx8K41ATXKADyxwp1wdJnV7GbxWjWqWvHR
O0TSM0kOQZFni53ZKi319DvJMuHOp8x3ty7kIUCJXIRCtZWeyFo/LObHS3qNl0G6p6OSzvMzjpcd
/IuivnrOsMBfBWLCLrH6lnh22c2chuYceapSRGvu84qbLT/ZjBuU3TESn6E8R+pMeyUKfkYolCR3
J61tBX8LeUpIKg9bbjOTzJNXFMJKC2lCrzE58LvO0TJZ73bFCS6akj/4qesdTZmgb6+/yH70pQG1
BRXtKb0zDO1duDp9IsxAON1mGtzfvs2HRskrlQGHhMTy3UZS4HS9W91t0R4kCNtFKfLoRb1RfIyD
uLVe+LonC86FGsKip2Q2yWBsqLZUBJNV9kW5altydIV7VDZ10DZ3YS8u3gwCsBbjP8io/Z7vKPUP
W9LnQxut/Te2Vjbg3YyNz53mX2u5BAuy5AZibDTHrSyunEPCwuWHkjcgDCdYX/MhLIQVDKD2qEcn
b9pXYa+W6WFe3DL4QS9DrjYUDmXxU41O37tcUxDhKRiqHdc9UnCYLCmRJdGv1wP7vAWZi2bOFDtb
ReKyJfmZviZw3usGbY1Mdl1FuVtAUB9DDT4dBo/rPB6U7smpTPMVXJGNp9DcF5vYij/Q/AOQAF7q
qIYxmoCYhZ2zTjQByNzNYBzIp49+OdaUp8vh3YQcAPkSFZ64Iom82p0kBKnzi5tG0QHmAXwlyaH5
F9qJmCrfWbZ7kcqK0Oewx3c8VQILREjazHNI5ahlVK+yTwIRMobdtTWpTreNgOBxqOLcDEhjbwoN
054t2Pz3kA+uoFtyvQaqp3CqMbugWFALTySROl+cofiN3XWHT98Xxa8IJTQYhmzbactdzzfmJA/b
qEx8zH9h+L956DCrVIGHXtun9hZ1P43DCaYNsa8MkBjJB3qSlxlqalX/lMpPmSORUnbZfPhkhpUA
BO9tJ46tsGdC2bcKiGTJFM+4vitz3BKhNn5xyNrWS1ah9TY/4fQvsAxUc2ZwhKeoBSA4Ek8w508F
yfHq5BP0XdWj67QLgEX7IcUNcy4WAjR144jyX7RYEnOtf1BRCsqf8cGUC+DhwCc1Vya1ROBkNB1v
Cr8X8ykhYSlxJCyjj4oGldw6p81gTkLCd0jofVfrwuiJXkWh7ghbQtAWNllmmG1kXbA26rOp+IHv
b1H/RUjOuF2EclzYf9sYo+Z78rws2AN4KLHgMRPgD9rYy8aaWN+F+qjv7HagJpNCEpTekIKM4TKm
QTA5TPwpO4fvXAY5EOjMgHQix7jTteP2PwowTH9V+XzLMZb1gu0tW5ZoGjPGL3K+oRkcpZMZaHxc
bKfaLnqC4dQQbzAAX65tG3GWEIqQiGcdKtz07ZUipozBodL1B9asSV8Lr8XZoHz0Pr5LIdVNL97a
YB6f8QWaB5N9keTxxzKuiQ67NQxhE/JuhSfRwo0YiFFMpzUafeZCkg3+U0lopKjO/QDBRZi0QlVz
baVBVjRkpLOoaZNcH42yhTqbqc7GRHb8/1Skg16men8+mSdF1wTYqn2QJIToH2SaxdwtuvHm9Gbf
ioF5Ou9+1CbH3Bo8ebdrD9UrfqkcZ1ZzeZWxY4JGmXGaRA64NANcYVj/s/+GDtUAmK2tGZerAoP5
Q35+ufrlhnwkQZNZk012V6IcDvpK2K1vb8OwGRlwsZDx08X+AD0xAfUF/7DV7tkYNjDvXzQI39+O
Bgv6Tr+w3Hy+uuvMrUVtmij8h5EkkRU7iqNJ0bcwDRYPtEz5RQhMXndchonjyQEoJvb0lb3qLPrH
BqFoG4JpZgbQp3OS2yRtAD14PId6QUYZxtmy1D2Vf+iOvZoUOMBZ7BFMT+BeuOUW6uPfzG3lXxdL
4oAAPIZMfcCNwps4LCONwsrrbf5g28Sqvpi6WFsAR647Kai/FrQH+7j1VEsVaiKIBGuyxu9zrOAq
Dan2w15Q8mDmCqQK91/87XjkInlHg8PzYAuUVHgR4/9WEd9W9lY6vrePaYzx3+0G2Zo4B4G/yhGT
DtB0IPImULptUJV6vu9wxSkHXpGd/IHI+EUJXQbkG6gIaJFe3sEi03wDar1wbUm7nIQyIUaV5QBe
VqDpoXY6746AzwKMN53K4bWrSV1C6FemTU8SJufULlIkknW4D7LDBPZIOLcDqEo0+b+WLUfNVMi9
23v0U0ElcX5Ft+8yApqsdEqzj3EdoxJ5qT/Ecj+cxRSPyX6p2QP+M9NQpK71JkgP4ICajU7Qn0zN
RqfptMWpR0PpipdFFwjGSB3G5aKNYM7wCbTBSZeL6Ru5isbF6M0w7XyL08FWKBoBFFIoLX+cN6NB
PdtRtJPkUV03Picky13HQ9owiU5wsm+Kv/3XvpALMFk4t+xwgTGLHSJCf1Ny/8nMXWyvbhjvULm9
CywMybFhR2HGYcKNbbrJI/erAO/Qha0SYF50JKv3q/BkjLOzQZAgiCCACICdClg01Sgmu22GBkNC
2QqcBtkQKf3gg7Sj6YuXjHO4Z8yeWPWSoJCCryXRnSjg+y2qRtaWaKtTgXqjvZLqpY5nYJg8s7n8
58pUoQjmIZSxw+fN73a8gIKSqwqBpWww35AKqvQ+g8rd7xBbZnZEY/ghXeXC2X2DTRGsiVFZLHae
ZaEzsC+oJzi6tnIrzEcK6VAeUmzQ5JkREt86zfmOf+lfW3hywX8ssSIo1YL1KC7emE17SpkcAE5E
qO8OpXCPHb+PK6MQI5RBTapuTcsp9McaPdqHZuMVPi+88pftvyPdk6jzFJfk0myhtLslPoDOcDAg
kBn6FVWdjjBLZGq9eCk4e/6okaxPTGInhFVSLoBz8U6QC0ma5g/duJJfYKAtgKTWjKTbTdgmmBY4
D45gKsJ+MwUWobH13yH8lu14/HzPyCJSjLmBXuwUBehdJTQgHmitgKZSqumyBFNJ1E1ZlVci/TQb
wQLnC07zjv/yE6RZS5AKp2rUbMS80ir8Ph7bXEADdBlL5HmQEidKQpJADoZErZoSa5d8OpfHHDPQ
MkgaC2GhFLMWxCaZRTTNTYRFsZ1k3pf3maCFHVhaL5DH10IweT1IDqlmJrU9RUljeoI5p8FH4BoA
vYUvBNqAOfXqmPy7017Ou3JcZFj1spdlSOBj1TdZ1C+ziBlJjnWqbkh3xrcDm8LBzauzeDfVjNmb
eqSA180E1dwUD9vRz780XuyVneW9ldQSwVPY2mmKxan+UaYuH9GlMRE2Bree2qvmzKsn6pkInNSb
6bfvZeUYToijmFwEyhPDNFdx4UBhyLZRfWQp0tiRU4NOd2/7DSoeb1p2NTXUEi2T3GRBuaMuwBk/
NHXcd6Qp+eZOViGZL0ZF7AbblSIEDYrowDfen47q9fKop9+jdOtN2CmCClk+f9gknTeCj+Q5zWLm
Rz+TAeR4KmhQT3+BPRKo07bT9bl26WBk7bpPRVqtanEN+7rNwcwCgX+lP7su9cqc0Z7hsYmhlNY0
9gDO+g9lL+pNuWkpY7Jz6HkAe/JCid5Ml/Dk44EeTLerXYX7NEpIV57rksmJw6uhsI4jy5GZMY3/
nYb5WAoHwnxZQaBXwRhzGQ3BntW8OQTbbvoruFONNt15MYUCmBSruDjAe+dDojJLjACsiPb22MOd
ITXKBf+gT8SXmlNrORAOx+aYvVzw1nhBxgjOrhqUwmF28XkITxtZDhULERLetffLo42npRP+Be7h
X0zn97/2QVu7uiIQCnhlIElO9DpRT/rQ+i1G8AQKyQcGNmiHlFBuAcAZhF+WE02Rro6RV6wkRPh6
SUHIvWFtSd/yOBbmKNlwByXa8jYo6GGEtr5eQSq9s+Gc6vasrSFWzh2SSOaR4caGpwXrY2XaOhy7
8tw7YVyYHcOuCe7XG0o08maiHmVmwJi1zs9A9pLKESfMt2IuRmyxcV+QW5MYpJCRvQPtWoKBWhWa
9ogGt/+iy6ArNuFqmKTn3aAZQpZLdqluXQ74ObwESJYI1wZlN0nfyma38XA+3iqPMyzlr8Q3VPrN
/dtozPsATtv2Zl7zKE9DYPXW+m1kgyfiq9qyOKjAIDK1lVgqTp2B6CQoy11Kht+yT+VpNTAk5JyH
/tM6IItaWC3VPcE/gzrc4G0e0k3kRqcQHM900/hNJarY+XSUMW2adofoqlxoPey+SR6sxQ2w3jJT
rU38uwQE7dKvwIM35KnKlIwE/FRXWEnqGTzmXWSCp/qU+MQszcmvo8bB3WbVdYqqVPdChjTirqIa
pfWprONqF/Dkykqnnk57J0BCplORlTcLkud+EbLGUDnBo/v5RCOdkCIBTpanmVJtmH83BlL+ZcDv
z4MOOR595dVRLXSpdNyRcuAhF4jUoJ5L03MFMw7k7nB4ibjGs+bmcyjTHDBBCFr66Y5nfGyzhV+b
gbPyWiL0STXu272sceoKvsxMecRTG0+KSbcXPsF2+k8WnjwsSc0CWrbwO78HtV14av+FFscMbcU6
7+ueDpd79d7uMkPBh98WKSsjueXQGXxzf78kHj6PbUkXwK6ZMHAAWwoXMDanb0NfmOlpUflw6iQz
YFIqtjDQI5tHyuHK/P6xuJT6iDfA3/yyWFZtFb9YiF1G8jGeQFHSwJpNSlQ8P64dDTG/EdZ3vHwa
NE5xuld1o8fgpxvtM3pSne2uHMjLoPw5qTDbiP6L1Jp5tKGwBCSFTOe3xUfcBpUOMsGqWHyF8Iyb
WAkRTL1X+2F990oLHXqFkZpBbXqyymRIeHQTqNw7HihJokxVOY3N33bPaI07rqbtZJLlajdpQiXy
rZMcg0Qxn5nFlz1/kYqCSI80j2qAZ83JMw/tvq4jTr7mbrnatQJFIT2qj8TfQbycCweJPUX+Y3H+
q3+JFFmpki5LNaI+bszOFtAi6QA+wLZgdnVx2BqoCj6CBo/e3HGTCsXyBS2esmE6JK2ClV/wngFK
BXI2XGDGpRMGkVsnmEzhBAp+WLufj9ytWmrgkyKF7J5ADBibC9iTUvUx2cYDy0CXDEXqdcq09wNV
LHMfSVSHw4uUCqYq44tRNR202Q9FvsmEaSFMzkne6YGYebtkSEAYYlaGuuufi28ly8n99PWvlJWL
6+hoNKumDZMERuQPBYGklsW3kRCQ/aLpbd1mX3Aeq7RXa2rMfZcfNVpMLRtlC1VVjFCdp9GFs1Ol
ZIIU9B8HLSQP+ciE/HnKPKlBYgUBOCXaukVPltTAgBuvn8BpJu5lEbj04RICUuZJJJnPDEv3lfgw
C6T/uDWoDwCUxmbS6r4hIfHOCCVIzo92cDAPd2Xxh4au6PeExEyuPzM820kbMVtzYH6nXjvx5IPB
Kr4H53kh5W2CkE1KWlF2p03n1SBY/JqxrzpcYEyjRnj+xwS+rLmyCM3g82euKgF6UvUvUoaJX7af
I7dK+2QmKvxyCMKuRE9zkkwvOTvfeWTgbhf/h5pDcVIh0YWfisjSoptqZQ5Yttjagq2FsFhjYoUW
ogDyQ4ackBz6T32fCp5JV6ZMYR7bjBOTYgxQnBeLNOEJ2b7gAGzduJFOWNR1AEPN7HjAmVoCbkUR
6BJUPJR0joltjWFcfrvGTyd0ApTI3ak7UXBGDSF8hlu/4YLUS4Fc776bPuJYopl+j8ADQ1eKUNFn
5jsMa4Wjt9p29jLBcaEn0s4KLcSWJYhyOg33BBylY24qXz2wZtxZed+AyFxuMpXmmcBeD0uXXYcG
az9Tb2973/9gssILeThb0KXc3nxfJQ+RtT3YZFGsHF7GZ0RjWTGKdDF2/u1zHlC/g09Eubwu0l7+
eEc+PPG205G8p/SEJm9L1Efh72zMDN0SP9jOgOPUD9g3o9hKaJVyobhQkatZ7AkhG8FKtF6J/Nl1
ZdM6Av7h4tFFLxRPuOqZNGYgdQMnKB/enJuIaDX4df3rBYTB3zES5Ell8VzR2VfwN1UBNib9ncZm
llNYDesx+qTbYWUguhp87sW/CEiEAatwoWxkiX/Pg57V/jd3cu0fS7xH3Pd2mBDafoEy5bBE0Myh
t5zOLHJemp7rDHKLKs4rkdeVi53wXYi4vEaU65rSDTF7lzmmz4K1IUoMq5QbOwbDTssL+tzV/iei
2Dxs4uEW7vhVnJAc0FSuAQkfbvuiYL9RrXCpG/fhk5ExlLSTt2P9L7t7RVzCnP6VCoL3ukm0VgOl
Qmu6h+8QA+GT3IlfqYhvmn8O+zCPzOuLJf6EMxjeyLRcYDF03pWex0OxdkI1HLvDW/BV2LjaCRF9
6sZm/QZII/4dgiGys1SenCAcC2IQLwvj8lf94A9i1a5QkBiCmMSaA238iZuAI6DXsiZNACUEQ0NZ
EL7NLTXPhR0Pjuw8P+qZSlWbK48X2y+o0H9FQ+2zhcDQesRxmofmVZIno1rUp+DOcIfA0A1xlNW1
qcqR3yVJV73Wjz5KynXXGxgtPGhKI2sQYhIN317RtJm6MdrVohoKOFEONJGO1pJvMTC2TYoigoXA
PdFuexiB6pILLLFkWPLPM+sHYMRNR+6unIKp9Fbur1bQw/HB/k1BMIlZTO3JapCXWkAJrnLN3PaN
zFctSZs5IhtISq+Tl9aYirsLsZWlZ+EQwnfvgogiPe3l2AEKbRW2SYaKVPJaOZy0ZR+fKauqBCD4
+Vm504dkfCQ6sFCEYRwFIP6n31OWF1XFIG9aLxxakiGK/iObdTp9npLPCk5FL9NXMdJ01nJrimjc
/dyw8EC1f2sUEfgaxGcevZjsYUTedpfeV9KfShZyGn/n13WOSauVSKYRoUPl/VKJhp3hmY7eL6N6
FMHuz3s3aTKXHIHj+F+vYxjsNB4feRuQI3Lz8e1Q+3dtYcyCilu2tDE46FdV4kbw1JqXZfTrt09A
GTrgEctd7d0bN9dH0f/UXS4xWdKPB/86Nx8pE2WcEmCRC3QX/KHIZXAi+UcP8Coq/AjsPRwt7pAc
Q5EgZgyJkPWE2UBgbzTq166DT9Lkp92slHAhmNh/70o/jR/b8/hK3U1JI4bQjbNHUlM2F5sz9rY6
I+00GZupeb+MI2d+0Rr7BlGpic1PcpYanF9nktWDtxOuoE6yjw2bgFXxZjAN3o5Vf6UbkrliW73H
u0mpCVoCN/oAovIeue/JEFcSLirnkoW8p32XcG+Fjs1mC232I+Y5w+SnfJ+465jLNdokTS/AHuZZ
yOe8s5GtZ5Qv5VSe5L77mLHCeoIfVarxzFLBEQ94KhsdTTMWCeTtcl8zsUDQmPALeNK9HnNMTQ8k
awZZ8bT6QfjF5DjXsNrgw4nOTv6sWFdPpVzLvXLaSoXR6x/SIp68h7ea/sJapNRZzYzTGi/nAe8t
XvKVTVZWvpmPoVNehsxvV1P5nzHVfNL3+A9GGWtofDvdT6TzCEDxw/Ukw2WFvhW9hcfemjgbTXhs
5LJ8OIBVv4775ntKHxU7yv/Q9jvsQ2zEwLO+r2GEuXmecoPrL/0ANgBjT62b8D95SQqcJTGa2rUJ
GcUBaVSaIcb5X93+O/bWx2xUTPG0hLdK5cG/RHEG7LqAY2ZBeHt1wCf4v1ASswnXpAD/nqaSIJjP
d5iT6VvEwtw6+jOjAmSVYo4S5mZrwuw3J0aR5z1dDXDj82+atZG+MREI5F8fEb2q2ylvIz40f3BT
Ho8KKn6cXaDrDuYueAIR8FKD0hObztvKoK+6jrwl/qkKjMqBGfOgFi+Z9mf+u8zY181XtgVV2rNn
rRvqVoUgEfLg/iEMPaLe5ngLRNQQCsa7Zan8zpEucXRSJznVLFyMG3DcSIuYqBriO5bezBhhdVez
6SXm/hy2h3GRf2B5Dr4nZ+/Xi2rshMPrNbW169WDUvUqxxbi0HrYdBymbOHQUfH/ttKoXrhejNiU
F0ymXRfnYSccfoCvI/p+epzeBWnt2p06JZJpwaqeXJfLPsbgMtQDQWjsmLN00o/y7BZCqmcfKkEl
IQ/oDn5HGUFibvhBkGyfuB2lE/XR7MLZrBUCUzO5vWBBVHALPvuP3GeFs1HOUkr9mScZgELYCjXy
+m5C4FMCcqMDcg92J32kkR/mU6266MbKDDAwboxAiekWtULHGlFZjvqlmnxiae2tFGvI65bMJEek
Ftf1WI0VUWEiNXad/ZbNsIE3h/5mz8Od+987y+twt6AQj/fwGnc89Xej5XOdhS4e2L/a2qOBlfOW
auqiNh5EY9NEfk4/P+f4tTH/7l51w6KvlCt0nxNVX39IbQVpSweQrkoJJDlzNWktmOnstQc+6V4w
qG3gbcn8MK4JyceVjl1GjKNVynBv2fatPyRrDO/HDeO9svo5+PKevFQpPgAj+AgR0oVmQPdqQnSb
4VZG4w0If4JJubWjo3nkYMTm+x2xH5dsg+msr4aTIrfU3GyUBoJpKZvG2Ci1P9MAOpAHutVpnErB
MIgdbkMBTzEe6CQ/r5XUlluIy7AwbRhABOdw8oQXLY642N4GHT/1HhwYpvcQe+kZpqC5sWNeTpTp
dz08hNNBBbnJIh6tkW+BI7c7QnpgPL9PVTyx8vB4MVJanambqVv3E30ceOolJrc9uIPuamuujUG3
7o+4suLdfh8iyJzVhJsbUcD4Z9GbqqacHpMZCCuhWhPU84rzatB/ca7qixdHLqVdOD+v6mmlmqJV
fuukoieYxNEo6pIVLpfP3fKuCYuEIh6LBLzhjyTWUC5Na1wKjlTS4Z/GauUfb4a8Oec9B5hAQgOV
qvLwB7id+ERAZKphnY6tgHsBv7tew0apCPyYqVhMPm9wPK23u9DeZ2urS2Azbtk5nSTs6jqYJOPf
/zm+2O9fhNKpumjo6o9CuIL1OJ6NOWksZBi4d+ZqG+alL5GmwSiKPVEF0NEgtv9zF9IUZbYK6mVn
6qR9d9tl2AYXXEC8G4PGmyHTZRQK3lzt5WIZzPtyLG383QyFNyz5wpLhWRLFFwlZuQvYjnw72hAv
THoXB1LVcPKWpwV6f+VKJZ47EQ3xZliictwajZW9fymfhdVgU5xsacZPLd3T4PBJ9ARS3Gee+tQ0
LDB0KAt6HHIoPnG1NlKjV0lI+Q8EWnLReyk1v1BWvjyQ7ma7ATqaJEo7az2qdMfCP7stjLODgWnM
Hmk7ylgVbeDNzbAX2SXgy7wwWzZQcXCe6cB57FtRiy4vMlzUs9zMyQnB9PEOc6pkb0usB4DqqlAm
oJq/ELk6JPMt5YjULqKDVM4dLqvjXponsQIoE+muVTAXoctbxFWOs1P4PeZ1H7d53reeZbrw6RKJ
H2xIL8EQKXD2XXax9RJ13hqSfJYytJYcXedduetIZbqqHirS4KAHZpSYSEBWAF8oExHaWXuItzw4
XYuE07wriNZI1rn0vL4Q/mwhG4C3rlSUVIS6Lh1XFLg4sgDv2p7Z378Y07tfK5mwzlilQmudTe2X
HBTI/VbWnB4MzIDw1oE9GMSBzC3y4GGNR/lMV5Zc2K03tYqbxirsDzbBmAYlr1LXe65tEJH2Fl3e
7s17uprdPry0HE+ct0ZmESgQ150D6tkuFgPjTgSK+R81C/OHnkT5fJSFwGVAbLFxeWA35L68waAh
ub1hNQdN8US+JkPkZUdZA9CIzexZgOxjZQlmxmZKZw6ZCn7nu1IUrUggqqDWgraAph1bg81anLz5
8RPJ+ppMyhJJ2IXw6rryCRqBNjfvAg9UF8Gem3ta3rvnmKu80JMhFBcqd+bGyf8hqHP0jPtNw47Q
4HWl5gb+LXwnyZ8c/xJQ31vT4pLCxeOi0lmwJQTUI6GuIuiu9ODvg/r61YJbgbad2VdCSgSRLuwm
mLkyemIJtLjmIUOFuqcH3cQYOK4DFkIRQ1Q5qQ3nF7tyXFwtN8kxgGL81UvzI1coBEJ5kaR3yXbQ
64KvCZDjvR56TRbQ34ndCArN26hazlWbC1Y8BLPcXHir1Yu0p9E88ISsuQjsnhPCC6AsMyiUF4RB
somI34/9GZy2LeJtLIHYmHACXjD+zF+eae3VUV7Y8Kcxa+sEApc3SBfsOYVizgCSrhgpIXdw21hp
kesd5KnSDIbrlU3zn5YVh15YIMIpPU9w3BbgOIonCFQ18KJg4kKG0vi2simOM9Zuq9Oyi3k2AgT2
kXD+qx4wdm0sswzZZJlMannSUHhsxE17t9jsvM56i0Hs2g2CQltd+lc6VbnXwiDXhzZH3IcFudFe
WoB04CgHRTkTvZG213bDmuTmnrc2s8VPpgTlfMwTRjuUaKH+tKHVymGOF88dIYXcoOIA07eibV6j
jPeZRYGjYk5S0JfS2EbFbfO/3cCjstSNSIl36Jdo/Lj096Bcx631hTk5ZFlgoVdIuW4sPtpQFkow
H4UEiTLiT6IY05uLutHOJDprk2epcqVtHB3F1NPyzZlr/ybqJKC+bkL+CiBCs7SadphBZ8h4S/va
g2Qwh0WAEtBymjdITZleXw+Okpnivu3qRWB0FCiO8VscJwcHvqEX6yUYMVaJesyyWgVWY8B6ThD0
punk9AS5i0fZPYM4Hkr9tRts5dn3bno2ugNiEcItcJAbgg628zyBNdn4dU+noaJGh6VbBDjQSl7f
Ca0mDeIXciLHjYC10CeEF0omnp38hBDR8aDwzTbLrerkJUpf0rMDlGjhMapy7IBAbIzPrJ+MR/+3
iYfkZDKGjzhoaY/2szDHQFmEkBzw7p2hZQi4eAOOXLJaMyepQDbWdQzQ9QGZYS4XLG1PQv7LJoqE
JEsG0vvsox7A0ffyARpGLibYBCsSMyPJth/NBF92l2pfHC3KyynY8S0Vmwjyd4dj/GSPyArpaSND
c44/jpVsy7nKzzr3Vio+TwQ0YUi1AcVcOK9fm0vkKmtnonZpLZrNskJKIo9UO+gz47wODy/Os3Hk
ULuvfb5y924PWxfT67wZTyQrYV8ImiR+yrd5srqsR9z3WAyckTRkn/qqKl9i5KK27hjDM0NdVXJR
P5FJdral+3og5g3w3YiejD+O9x8Ztv34r7gsvQxCA6o+0LCpH1TlddgXSXV9gwmxXgSAJoNh952+
dzDmNRgOqh4xc/0LvFe5LACWcFfbfV7Zxg2ZUFvp7vskNADcSuljNSy2w4xUpEWQmZ4BuOwmgqxJ
9MfaE0kUouU2MjDsj1eAjLhno1T0lI3kaCFQA7HvK2w5UdvrO6v2yoc7Hx6BzQKu4FO+TqzAsLvY
+5DYkDKhr25IRzUzrghnbZDaZyNKMcQXhnmps6OfK3LPCc7lPqSBMsA4lSPuOQYcOx/qy1fpi+Mx
O6o2tFE8peb46dT0smmm6EwXdJu4JTEYcxvyasPJeFmdYSW3YFcXvb+6QN0HT8UV5uYq9eCSyY9K
/43SaKpbzckNY0Hn757i0BDlKF4tvX8mAwNZuIT49izFoTMFcKZ9gwKxAMu8MAS+FsaestKEaidE
NNtriWiCHzzwy+BWgPWB0aucZeTgjZKEdjItJAmZSNbHAkRvJRkqcDdc6Z4o4s0Jre8+eou30k7v
zp/zeUxVWOKtMy2P+grSgJUT4nO6SXU+gBu6ahzKj4FsLxCNrUq3ytIzJZB3oV0xO2+dIuxxrs03
aKsjzOfugt+ipO5YtGFxH36YXNYqMQpBBdtbPHRN2yNcAXQLfwW9SD3AL06P9tvSggjZ6gt9OmQ4
PEz8fsajuFhFiFwjmhG3+hn3neJWoMj3UIZgSG6BGLz/GJalhlK/JEisdButus833b8LzgS1+pgs
fvr6U2k8n2d09ULsMQPLKtFKHtnUtnEwIzmHpSWTQaos+oiXP/6kp3y0RE8/njqsDOenJle1XWov
pIhHTZrSVImjijkOHOumuIsbFDO659we7ufdqNgt4tQXzvIdyZ4vtAvJ8LLdShrRfbY6lZ+qcp9F
M+ZVeNaILgymgPx1EiNmyZYhfW1ueaPmZeC1rG4Sn52hwUymNdxWFLb0c3MvyJJ3a3BfS/bGEgDb
olaTI9JQrlgI/ZIhe4lvNT/2xTai3ScqBpA0tEtSR6rCZpBVBUPsGtxSJ+RST3jfkp6Zc+uQQV+D
q7tWWdlveHpE3jKUQmCfwKzQ3f7I2y5B8zhmmn2wlzoIvopQdNSCNOLd3/LR8eN46ySZm6rZNPBl
cApE9jQRoaE1bCdeaOErmRBb9JK0eaE0YonBbzF0NSHPRklAHWuJfDavSENcO8cZwUu+STCNM7uJ
+geCyaBsPZKyvS7X6FjDbjMvjJwPebHDP9D3uEVvchpIfFhgKYbACkee2YJTNRNlIp/c/4q6YlqT
pOO/aELmrNwoldAu46Z3oAcTHGw5NP7DscvufZS468N+9cClNquiSy9HX9mPSwnwDEarGM1WYUKK
+9ABDO93oODToh7nZjmrDXiJV+dtB2jqZspDDc7rYtHqOoe1g2eH8gETCV/v0tydWVklZDruiJeP
AZrYsYfxuEB+Uz7pLv44s67nzACd7pNrSvDGOpJ4Vkeam4ot03ii1Oh6vFoWX3n+z9LeirSt1/FW
eWUyhEeOJKKAUzimuExp7qQj79HYAHvNvurF8MfNQG+QxksSwrLPYd1BF0T/sUoj2Xct6R1u0BmS
TbDw0SWIDRp2EENImdoJx9uuKtZ6X4yPql9YI9wHqqACPJAJLPrs6mW+P8PRILI9cZqSrpADlMop
Y30WipOstYTY+vhEaYbgTlBqAcr+ZSScszqE9M9E3nQ/DK3uRcffPoD7OYntFcjUuMZ/v6NMZbK7
4ZFCGwPs99DoSBbm9fDvf6TvjhY6wmlQlEYunbOko3L6Xe3V+f8K4VjX8R5r+HWPCIiiYhCsu/4l
92Mae98pkWZav23p8Z/OUs5myNBqgiDmdMFUO0dhwqYTLlzdATG8Uk3SI/sb18QMb2af9SeqhHyZ
ERiZYI8zdJoblIX/MgkhJX2VEmvoIOt/R+Q6rLqlCwzyf7S2vGGqlBmnr0mnlAdf+dCjL9diIx+E
UV7u6xqzaJoYDzXP0Y2ga32a9y4yIRFlSzOQp9CrSQXBCwHOEkcq64pIPyyol9v/P5Rs5cQqA/x8
EQ4s9ZpmQTAKGmz+F/6lXTTxTJ703OYcXLis99WxWx7g94j+LNuSpmHIQTiSd0uWFxDp6Wu0nT2c
KXLA029QD0DxLAVHiJ7U6kp3LiU3env0ZTJxj9oux4fqs+PxChi/YETo9PsBIlk5ktd/HtSNkf+J
n6HSdhFDSHY8h83T8KvyN3GXLMh1C5n6vobb6RRNIZ3kCB8jV0Y2F26+QJVFuDt0iLP5cWkDyr84
LgtERsEQrX2WH1HAyr803e01KDK5NTII6NPYJZ3AJqabGgld+GQD4n4FZ8DtqLaoFJ13hxQ65eku
tyMqflUXXSl6g8aZHaraJ0/TCl9c37mgSGmAO9m0x5pMwX1zKaQb2roLz6NgV/Li+Qpl/Hky8Hwc
LU1T/5YzNMY/rOPxEj2JNCvEDkDNoIvTJF4YBuadqz+KBXJcsyaGngXj0+NPP10pXCRHUsCFb0QB
YWJTcNsb1JTQFDI80MPdmqNwoJhsfWC72Q2lAy6jGSFWL+vGrvEuR2O7HFx0HQg/vKMbowwsVWY5
icW+qi57zAPSDinsGtz2b6UCj1bUS40jZlQOcqTMjiFZoNeOeQdirY8Kr9FW2lRFBxv9XrgOwPRi
m/8Wkj20so1jmKrO9NZkodf78X2zdmRmMDS6ebJHMeUg7Q+v1MiErECKgvv+1GJd11BOPoR1dSGZ
v83qTnD97vtKPQrs3JUNfm3IN8teWmyveTsQp/ANbg1BuGsh0N1sWYqNsR1R5CZeesVU8qItnRj/
xhb3HVl16XhVySbAItx7aEqlHugFuoaF/LNpk5+p+5P98r45Gt/g3ksr9Sx3ja87UoQYMt7JDdg0
naWBAIGtsBmjPq2G+wFzEJOKF2HKyTqji4lNQ/cOHvaTy9+IkV2JICbt9B2ldbempnTbIDIYbXE3
051rjocdUstTburGlftVJIS2mC8k9WJSnQGTk6QIgqSwTukL6Tn75KsV4cojiXlm+NSnkuccLlCG
D5SvLDcd0SHu0Y7Vaxr3apcowMBp7khAuthcb8Yd/cg3nNjTpQarRfEHBWOB75oBUkTAEdB/kZgP
UfhDgDXR7YHAH2fRvzqPbkOxuzP4oKHfv/L+ZQiBuFGjI+8OVjg3QmcMf1EliCyDbMYX+0PpmNrS
4xqN0tlKwW+hrWdgOYsojsnw7pscl21cMntGrqQIeOtlptFW2DnAHKYpdE9s/qU43+MSUR15j09W
6AUqVu74Ii4pv6eZe8xD4qdisx+jxw64sZbeofZkzDtLK2w5xa2Sz4ogT7PalA6nRlU+50VekRy5
5DpiKAWEh+CxneFuQHvCeAOOgDggK2g8WFsEBjf0UrxYdcpPsWbaVBOhRLKTIE98srpKh+LZsrXj
AXKTb/OSpdL85ziBPhz+87YUs1Xv6X9ITHg1OtDzwxoSy8VmurPiUTZlWE5qIgygXn/V7ZZMwUhX
CrIPCJOU45IXJADDsOoU2osxLj+LuYBDHJngd8PAm9Uk6cROpg5Or5PS+XHZ+bNcI7blUT9hsXkV
2KydoyY4FUkDGiWJautaTU1Qflcl7aXr7smqMpSEjNk/5XKePUZ+aUtDt0k9I26Mthdb8Ffvn8Iv
iIeWFxpgmp+MoFh5odETV1DNdgG+G7K3I7k3Gcozmz/sqLr/p4SG4ajKiw7ApSbYKUI/BkwJY9h9
ylyoexc8JBV7oAKKTu/NCcgcGmRtUoHcZ1gMJb9nbnkIPlVfx480DiKhWNe6yHCu6grNgRAhppgZ
KqDza+kV/9g8eYfGqsEOFNnKP0Dy6r6j4KGjH1m52nni0g61/1zxpPyCOYsSvxN5+2ANAWMJOoHg
8ZfTwheAw0aKnY6CV5iBZZr3K9sOcaeqkgJtXWIArH1N4619iWz+YT3b6UezodvTyWtpliwJciRc
xuN7c3dWQiY7I3glHH+xSTUsXnATXapMR1SRBHL6clyucgZ/h4zH89rGsvOcgF38QjX6B72v2hdE
bBKMOUXCKbihK7WMSsKwHq7NSgT4YDJFYIORu51Gg1EfqRDkGTTZOXIX9vGiDPyeNA7hwXsqAujT
KJyDCWsc2IQbxCsp3XiE7KQ3yMq2yiLgzpNt0SSXh/fIlpA5Y2og+AJqO2GmppR7+P5ItzBI4OmY
rKNTdJ2FJFEX7myuU/5DrcszvnD91u687yts9XPHaVl3b2PbBnl8NdOnNDql6Bm9HjNX2CSamoJ4
zrmUHgU40Pst7adM6jWeYWJHkU8SciLSUaDi3YPDRDzkhCXOwlAeHRsAQ7usYvi0KIjUk+C9MxzB
rMptVZ/J+6cXC78K/YnTiO7v/gaNGM14xc3iNeN4qhzOOW6YH5THjhIkN2uKqxBLj+WMtpmq8xSo
GvFLqHEqTSA35UdQq5bOKgw7CclzAWLQacU5tsBfezNm1jpNxPj4WU84MfA6XZTjnQ7izq0rW+/m
ueTHwljxPZHY/FYkG4RaZxIPJD2iAgEDwG2GBNlAXSluCr+yHttbjeBm7XgauMU7InfV3rfImQ29
9UMfsU0tVvqNonWH/ZGgKqdKhvHX0T/+2iJltijLdsTGxnidvW3MPNkGuuHqkFODtYm6UUVD3Ki3
6WZjGwSLPDIqqcNK02XluNo23+c6eemkOooz0YjEO7Av82TOeV93Jnj5cCXe0krXqgAxoj1WaQ+6
dfvB1nJuqRX7q4aYwkpMozENMqnOuPreNZpuOeq35TkFftiWXC3TUruThpNazMcIgAfKgSSn+SYI
k4mWCVfo9TTPUebPBYq1VNi5OoO8UfQKLHt/Ff2y/+/PzafWVM+xyzk6RxxWn/1I1DgDsMKDpDS4
Pmi+Oq5suE5ljL5EblLZ0iisRl+C+lca0cf0efcqCqKEJXh+EFV404PahH+hyPbtrVezDWDlKlss
YvtiSW4Y9Y9j6tTEMlbXin2fAOMASY1OoPz2030W/OxbnyTo7KCu49MpeN7PFHevhUmWldfWqnRy
/0d2T97IPcr040AribbN/iHrcZsRQSA6sUB2xTZAnHCoSmxKAWNd8pSSbWacOqJK7NgbffxHGUdk
R1V9DcsX/bD4J54JH0OEOoYwQMTiXnugRMhNT8NZ5wEnHXaiWIDJ5tsUnZqYRlyoegX/0f2FsbAj
UlZntP7umGi14xyCojty8dMKe1E3WshvyoByPv6o45XV2pv74RaiXnTXgeMCZ/e/cJqZy0hSBKTA
No+RdlkRXWrpbgyoLjM9LcOUFs1ZWeStcQtX0C12wRPWAByiTZ7FKCVi4tiDZT97SWHFAcQ1eR7u
b9JttXEmB4JFTQ2VXyH1PcfX/40u83tmZVCkaE0emjyHIAqever/M6alIel7G0H4gnLFH1xHuKMm
cmcqxdoDyRV+KkzDLjsBOWbVOMBmhgHD66NJerPAoe4b/hdJcEyvpHX6oGfjuSO1vXrYpiPPbKO5
6bqOBLm4Iyc2SA2NP0LebYeRjV5UZ6ITvIbQ1ednhE4lLgSHNZfa3ri1SdTO8m1w0LpGO5uSVzSR
wGDDIlyNOuCwWAj3m/Szd9VXgGsJkNedFF2F/5i23Bh4C1LQBJILGC4nHiOjqNqKlkALEkvvM8X/
2s6myU2t91jHr9cORKdzcG21kyGqNInv9hqyoVVT4+QHBxLN9ufG8rmFrgQGxayGkuU4bi7UeZpH
rk8qL5rKstLHDP7wDbRlfL+OtwjybyRGdcyUrrq0JF2cdZupwWoGBwFX3zEFuuPqmdb3H4RptmNX
jmYFWjdRxF3bBUwwTQqnOAEjOp4s3EkrdEHaL0hMfdb1qy1AVTwuhrTXZa1ixVtk+jHQMT8dUjSJ
nf5UZYduX24x4G8ummfGVkqQ0S+LVKHO7xQAJTDKrgOqOawnGYNzUVtRTjjZADXurzqAykGRjqgC
yoHJpn0r5IcZ3XRcUiBbcExuNezRpPu5kbKN8elhT1wy4bw/jWLmjQx4H3yhpZcNtQTFZ8HIFK45
rL2sUZ1/q2WNOsYWHqpp19oBkY+QiVFS9Bpg7WjmfieHZQPc/9hw0313rUnPAvocbfYNqyKg0D9t
Q0QsFGE5ugE5Awq/LVbW+hxpgBy+ofMmTdx2c3JH7S/TW14kS4dT1y2N2fCl1YuPhZ12GT9dyOwh
r/mDH99G04r2bQ6ho+MrpfCV+WFuK+qf4W3jRq0iEYD0BIpyyOgOO54FpLw9lenfPtWrajreYQ8k
PTrpDRUVYlNQdurMQ3xGxHL2ZYfZkyRSYfHEth7UjrEk5a+IZDTsBp8hf5ge6tbjZ4zRbjJ0YjrN
9jURmAE3eZy2LGb0zfJbKRsMwbnvdf56JI0CuVIOVvlqPWLxAmRq5snoNlqLPkNi/eu3rO/GjQJo
eqkciqPFznAob7lXC7GtsT0/90SQa6V9eLBp0/ohCnIB1/QlnBdXn1isEQq7pu+3LHqSACBKWLn2
AKe0CPUL2ZBvi7z/gTtBvLP6a9notB3ox4dUNo6td95xs9R7G0Ntne7WyDV54hjy3JRtNjo55nq1
3QFGGZS5nKMdYqSTvFJ60m7pzpCm95jhLx/5s1wCtggFhLCCL2ea9Atjd8h7FQ46kbblMuAgxljr
mPX3yEQ3E2qWL5XIeFG9wFCP26p8qXP/kR0Agwx+cR5Gf1MOWsWlpITxLpBMDudLh56k4FEXoHsA
VTevH7TgcRvFji+CtXevVn3zwLiMuiUwiwXg1EYt5d4CADqTpcD1BfboSOTxmocDAbL9q4nWqpJT
lVm7JF/SVQ9aTj3LsMKy1UqCCqNry88pz3P6a6P2Nh1mnwcmSC8+TzEVwd5NM/BDwRCsNggsuB5I
tdzod5WsmXySC/9cn1l3q58YOMrVftkqokvOVZObHQZa4nUSVUWloDW9vEGeIptWCasQIB+WFWk1
t3Kk4Crs8owTtJM6+JpdiCZOvoDfkEJQNNxx2wzJ2bKxaNN72bBPeQc/tKxNpGKHTo3sqd684HG6
I5+xAx3+vDY4ugWx5ZUZVy5RUe7/iVc9ObQzmP9S51ydrWKidIYSWTG1w7pGtFWCB8aRp4hc8FkB
e3rwFaC7koS6KNKzihMwUo6VHt6GEuMaq0RhQTxwHibKs+gEXquWtRMkaECeQ34MC5hMZE2k7hAp
YyXYFPy7SkJPRQu3G1PO9/jVF8iGiefY75CzEmvoQXwfQegkm+98rlXRZqxPBPnklHVRD7l37DdG
8UvuOLhoFFcyMek1HYO9rIt9G72JhEwV7OsoMXoGtO643cCTU8UuCUvPDue5mJnbcSUbVPXQzjWP
n1yLHgo7sX576jSOcjn31JAVzSvrnDKqAuI1s4rCQ9I0869ITtpu4LyGKKZghagpqoYbb+5cbS+9
ESavjOg/W1Y6yRy5f8Wsk+RhQevY8dHhFnOxDqDNHo0TgI3gk3zrrt7DHOQp6echcNTNrjCE+Zk9
p7ZV8QQR5XbPbh1ljMAoVBE+FTfbeQyhc1rdFkCXveIQK6Iv1rWlr/HEshx2KP6METwSWg+8eqGu
13gzY3olg3VdmpWLCklAWNk4g0SQafSjyS7Sh6HGLtVL3KvvXyTFvHB+FWztlq6jx1gtiJzxapOn
tJ6hfZ46dcI1CxlOUe3PpcK64i6VXCgfcYu/vcQS2AQggSXO3mvn59PG4eRwa9hDvISgFX/Y3DWO
1Fm+ymTfMYS1mxv2PQ+NRcQTjFboLu7S4mtmBIVq4qf08zwW0lr8b63rGpbfcB0sD2JAXDfkY6mE
dRob2b7KIy0PbpNOUvqPmkJVJvIwDuUksIKAhGrrLibaQtVrrj+Jv+gGEJmyliJJkiJBOu6r5JrV
U8RU9Cg3xDrATFQMjKGJzommvSgUwUftzZBaTa37nwqWI7hEtoC66p2UGRqQCkwUQZ3QStCuu7Ga
9dM2P8LF3sTeAAYK5PUrVHYShglNk28QgnE2kXjjSYdn0U7ARlKikLN7CK6x2rcRTkvuPh7Sut/F
lrOUk/g7vpdN+Bj8VtltNTiSuDI0fyOFLrzyThGTCmnmtkXmNJqMcJhN5hAuzGAEgDCXrB6z9vvY
rgzjFfjiAN33Bcu+D1Dmh9sAHQORcXaE0FdzKvltKfdHYRIRtETgBQ21cY179ASgHwvXMSR8HjpN
GnzHN1CZhR+YCXJr1ldk+vHdiZ/oV5mu0BsYYIDFsuf/i3VCR9WhxOzHqCZWmRsPyRc01DNwgJ1z
aVNuKSpGwYNE1H17l6lgpgqMAfA4kTZbHC952uEEfb/xeeBKvoLwXvnJmiHR3lCcIGbWW6YI/q6l
AHCCdA36X7c1AwfI+tMadt6rdeco/mwq1dwgVZEBpM2bD92F8aoJIxGd2QilAxnLxwNCng0gqtVG
j37fN6nneXN+gXwi8RmqDVMgiZiCCP1frGci3WcMfyT/eDkXC/4LqPRh29fKmXQ0A2VxomRYMikt
O//25TfqJAtflQYZT/FNiIf9jJV7edIJQQiGZCdNC3hfPDlbhJ3BOSDB6aC4X4YzLN8amFs8D6pL
cs+EHCPz+xUUbC23oWJClypfW0WH9v18VUz7zeIK64uzseIvTRcW41RsJIiRpQIYgIjjfEhmqQgd
4FKMe6X1MWxcCTx0/UdGqyAorqz9sZBD0LCHim7chpzqiPFXMHhiPFkLD3LUtJitfmQOjw/21VBn
t/7maiIIw2YDyLxZJHh4XlvkkIevLSLTV1AQ28Mie5MPRck0qlp2vfHEfP/R+42g9w63UfMuxCWt
fmTL80t0Hv+ztDLbwvyS5jrGj7BBHnOEzPMINwDDyh0qyjl5PT/allqrPf9PPUsCH+mbzmFheYY3
oGi1kZhhEMG6yQU1b63dnxKgqBhuFZPIiTCbZabOxGkpHFGKHUXlmMKLycQJdFV9DmxG6HNqdyng
2bBNvYY5W6xI8EuApt/iRq/7cBXVRTTBj8FUxuMo5tumg5d9qEBmDgPUYDbPBqGqOt/nB3zGAofs
2tih87H2spN6FvF7WgRycyCGLw75AyjoWz2oHjwXV6t2nsNzePHECSFsJfBFCRlAQVUYMU89ae5l
DChHDq4jD8NpgRzBaacW0hEFvntVMLepP5LLVXecnGesTsXnD5zGRhwoZTKUlLtNoh6QuZJYXq9s
JH4Lg7e1RigvEBlm9TOKmyQ6tPWk+iGFM80vFurnuvTrhERxembcp+KvGuvhhW/oyigfkr4uIBJ2
QA1Q1CQiiflu3OXQx6tDXE5gIYrYEyuPUyqQB/J7no6TifpvVkoZ7nxgbqWZFL8CPDEqEfhTYT1a
v7mdnTLg7NyJ3qBHjOLUU6oquW/yaZzPskYuTTS8/Ob/q8irzvxzG5zNeIEdXEhc7ZupsVkK+yGg
T/VQhSvWrGJiInjgzbmnBZa25bJFRKkeGyjmcU5O1UBG7Ow5923Fquji+yCJ8a/iORcjspjjJhrB
oncdFlRSxoom9vzuuKKHP6WhqABXHsTyRIREnZj0+PZbA6nEHYecVuuR41OYNKHrOAIB2L6a6nSa
ryHw40qLY1PZRkuItwCofrw8anK25UEunE3GdsYgxK3Pm/V7ehgzNzRzqYNLMMkqGO3oo++EME0/
NMUe3TyyhBjMWcqHCZ9yjFFKLVSeGagB6mIeex4u7BQAsfYnEhh52BnTNno0zJ73TcvFFym0YJlO
WwGpm/68FcAimVE6z9V39L2QpERKSyHUQ/v3Thi40KR3xSv4BmfxEZ3iOdX7NlEvyGzp0tVf1P4s
b+Rc65+9MUbdzSs8d+7R2qVwOGaEa77ta1UgTj9/uYFuvVmUbqLbA53KyUFIni5YRWl4RSKiQP5i
fkhPrRml5OCrf4DHRx7MSrXT727iEA0R0Uac9kZTRIUQSZWqgWajzmgG9ALGq3bEgaXkDmj+EotN
gPKRf6LGOLAauSfNBJg+rQ1/VJ4Ai0Io6nUHH9HDxNP0a7+lbUuuuY8S5HhNhAYdn3sarljHV3Zo
Th6IiGKibBZSf6u+r8gRve4P5BHzpDHSCHxZG5lLb88Xj+zgkESsrLcbZpO6TBJwJtjek3OQEAay
X1n0gDgFSwlwVUJ49oCz9MTkLq9DIo9kY/cZ8IDqAewHf2uBs/DEkY2YXUJm9DBx39vtC0qB3vHg
X48nb4m1hQ/CtkoLmaB6eEF8BapAdZVIaYbT5fxGCJh7erlAeyTP8kJoIIATP+1tLKvN8ZlwBpK1
ssict/pWdbzrAKh9tG2hJgq960M8fH0ZjadVo1JTeGEwN18Wpk5T6VmON22FzhlUWcymLljSeDof
egHTjrmksk3u7E+si1p1O7RHhSfpW1YDAh25jHuNaopSnkinsMTwjkEI+2hTWn3mgt4nDPtJeYS0
hopNjHbC9kF0/HnTG38xKflIjKSI2sBxubywKYXuXQc8bF59OX6MAx4r3oelPgHMTH9xnKeoOPAN
kxervah5ZWQrkVSLd75hmR8Smr3bkZ3mEQkATsjyA9M7qgifhrEVF6uR8kRkQNFWE6aTNC+A7e6S
eWuqZWW21tzqfu2XZtQQnYh4oLSuMseJzDNwUCNKLA73l8cduFvlZoDlj2jBFz7uJ6TF2c58MiU5
Jy0baiNYhFWjJWVwb4bLAb8MnQxMcCNFztKzWfW/5myoR67YwqT47mCWW1JeWRGKXHZedc/Zjdbd
hRLCdUvktZsBEZaOTCWGHuSzhwlLI37g/znMwPNGjv9NgqMknobvRkm+Jw227LFKHnH7cw5+cgUt
gFGEY9+2uWB7n+QszGnu2Xhha2btt2u+UqOS52YXtDn8enBjl9tPInBfoSOGzHGTVrVvh73NFSUl
PnwCkY6GL6g5UQPRR4a06fHIk0F5LUNr/uhbUaxJMLUAmviUrnnvONpZ0NskA0qfxnpOe7GFU+zv
XtfnCosV420SgINEx47AD3hovD4ny68dzw1iUHLp3Pl3b/kLxApEA54ieO+c6LG/AEl9f+pkCQET
TxDu1ysqfeUMSxEUdAr5iQh8OCJYtChtx9SoFw9pjEuo66O+dRYFkM01JqewOT29ofKscRszm91D
e1jqeqXRNRNQBkKKRq+ceicFAoLRwnRZ65IMbq7RZyZnVyLxJs2uJF+UqQYrPFGXFzINeVwQXHYi
U2jCV+BEARtRNHPuXHbJvQ1MkIHiCR+GHDfLeFfLe8f4yO/MR/PA5jkfWXPNUf+ERa9O/MDdV1Em
qOXpWpMSFM8Xv2oMeZpiMZJJyroQfACTFSRDy2ms+eQhj0UkHanTWxdZJirsjaenazUHiTm2RPjS
5JleEhbHKE104oTg6BZwh09i0V9GptLfiJ0qB7BQHbq8KAGvuZC9k3R3sbhaIu4Ycm1NCemtm3JP
n2ubOZ0BG6cssvpfNU8PiSxmxa3bLHSUJf/gDcptuYcJNNrTbSd7DyCCKI6/qS3SSXewxarw/CBs
BgPlB0qIaQQHBpVMaqGrcLVZSONIdIv/OnOMourpK2reFvl3uDAifrDJuwEd37P3JRykTFPxjbjW
vE1tKlOiWCiM+4eGwr/n0oG5QWEprEXK/l+h+NlVlFL73L2hS00BfLpVmlvHwL9OM6RX6r7TmmWn
VTjt7mxivzcJ49fSM06CJglJceTCOn9s2pxeswGCwkop9LG06rSIYSDly/vpHs9NqDt/bMx96qDy
yHVnl3/10jTUraRtD84bWQxd9gAb4DWiGPIcNwy7dySerJDweNC6MHv6qpf00D/12kDiWxHIc8mC
GNy1OaV48HcOqEYtTFYTcRodlYcXqCYkxD0zR/4Lkkq28SNedSppVEBV5sFJ0TskK00SG4gZ0kJ5
ODa7194pttN2nyTebQr5LZXPk/tZIi/M02QtPArr4IAPUl8PVjngjjIiVULjMw3Hl3St4Nz/u9Ij
/XQ6l/BRZsDlzsBZ3wy5A0dHuGvstgYAsCfVlkw7b+zDbg6s19GGZMbqylQmJsu+DrheTlErbDLn
MwEzMk/tCmtQhmZcU+PrYUKrraJUd5znWOxYQQB/x3ukGh2JeqKaSOdOuKxFRiUZJUYxe85/V0/H
qoMMjPLh1/7+FI26BzWJ9qhF2vr46G7IG2r+sn6UlljuUbt6OGS8XZQbZQ+CaYUhxcUza+J/6Txw
lWMmkoqUo8KmaRyBl7q1Tq0N/U4EqH4C2zWsc1VlzLOhcRJqcdfT3j0ORvGhY+v2WCx0fqKSCkCM
sJwkUJBgitgx1Sh809Y4RQGbNGY6U/eDxf+NHxWFPcBfklXHHDJ9EUGBj9G3C14tR+6yTaK7u14P
HQfAjTGICFaj33zMgpihCcuef66LeUzvKw/+MrMA/gsDLyJ5lHQSu/OECwwP5YwZmdW68MQSE6c/
PF8srONnDbKMT0kiRkbbPJAlzG4HqSsPzx4Es9MxTVHITN2/Du1EBFRUz8Ls24bT1Mn21KRGkVUq
+7dQCjwQDv5RJOpfEIS60wsk5sSQ9Wiy/uCnuvMk5ex4Vl9t4dty5FZPLkp3qxyPwX4RE48U2rw3
/BhRTcFxyUK2H+9GGjACYFfT6nQMCn0juT32wlgIzgOU/FKYHUbtAbCtiAl6VF+9uCpXtmo8TzdC
qe1SvSQ2LMgNdjKmIGzp9/c5b5Kc/f/TXg2OLYYqG9H70pA+Ujson3X8IufSCOERYxFGFU06g4IY
W9weTcyEmioDCRJI4siyxm39w+zP6xZXGNnibkQvYBy12uZyVhmJMOgECnNy6TGntLTXDQvz2CFA
pfWP7yS+5e0IrQyv40NwfhIJGFKXduIQeMZ7aENqawgAYRPE4Q3F/WnOKLdRzPWE/4UQ1uZblxkj
N5f1LB+pMIvsZJ90GcUvTkkCzYxSJLKw8axd9mWCCQbJTjyaEn/ZaqkMwlVzvWLeNDH0wBMejFae
QsDc31nAY7ydCJkwlr7cbyCsFFxKr3lGZCYJidL+TaAgoxUvWz7pCs9ljD4S4ckj0R9jwxLE7PpH
Do02E1w5/9KsXlBq4zkHSM78kCOlygvGa6uqDh03xA9oWIfIkp/A4wi3u3gVaJHn2+0GZBZj5LVZ
MmPahSqo8VZCsuNrwo4PsKJdSG/aqaad++uJkpraABHik1Z3dr6tmb2+6JuHsSS2nvy/lDF6Vvqj
OZeD9oSst5iCJMt66w6xQcunIykc4nBBY6HxCunHuxrJ+3EP/AK3Ffccw9ti5uvg4sIzpWdrR/QN
oBPnG9NmzSbg2ADMW9hyRiWAqVS5vrTmyeFSIMsti+BtCSSfE9DrRHrcQhiSS4zmamJpc55DgrJx
C2MHG38qJGWwa71s2ygKt0+jQsgFVKI01tOTZFG+NHqjfhe2bsZXm9hx2aB6Ks0FNkzbsv9J1Mr6
XGawGeaYh0Ng+ijKJjHJY7qV3uk3hsTC0n6f7CUDqItmxLsy8e5yNX/UXdy6wZTkL+nWO9xM3hep
t/27c7rwCthL3XZvz2YJdsiOdBGHTRYq3Ym9nX8/iF6KInCg/UaK7tCRDanviqKKgGUD8NmGr+0N
mByNpFMNY6kYx0wXw3y5LQpnVAOS7KnI0BfmEzGfvWC7GwX7T+DCcVxfTEulBVS9gvjM5+YFaz2O
E1TJeQw9hrZeb/m4UpXnGzvDyh5/+BF5Ow+dEZes4XvMOgRtmR6xF9pItNsrjN+dzdtgbLFM8Civ
VP9tHzANwSAGxcS3MeQLvtdjHtJ9wPKy9AlMq0HIQ52MK5OWxcbOOzn3Vk7MRH6uCqRSlJ0Y9NFH
c3MbonWook1miFOcDJ2BW+vewq1lR4bydqMVlS7FxyWO0EFmWhkOu7+8IIzLz7tSByJqaLPdRaO1
I0oMsnSfie4SRHiEvsJdDofaZCX1qLRRxnZa4a+SZ168BtjCprYxkzY=
`protect end_protected
