`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UdbgCs3cOKfXGxwnGiks0foSAFvwu9ROCUdMQ+AbMfhiX/lZ/Hu4YqR2htbQ9SD4/f/Tdh5V4hGM
Afm9uEwtbA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LIDtf7KxUZv/HGcq00SIH+MDkmEUf5uow2hx1fhg8jCi6Ll8OSHG2wGKqJTBVbw5JikkNc1a/TPu
uP7oBo1KiFG9M0j6eATOp06ZCJeHMJlkzMK+wiQHVfPW3GnvVyjAj8gyVrz+Uo966warOCINo5j4
m4SUmVESN4CDRKnPtGY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TzVRF/JHDw+ctQ3dOwuk/u9gMPVo/gR2oTfB/4EjD2w2WR13GDHdieVc06VMCx+lv1PedAGTfDtH
rwyLfSYBP724mmzIwqa3Qra03YFj5Dej/ZrpxSnMZVr73Br4qAEgj13cSeeQnpJ3s5fBPNyevQlc
WK2dw/80GgcdwGGSvnZV99RQOCYgYy6RDWXHtbArF3Db3+QCWRlSbHXh0f/CEnjpbSW/mVrQHXa/
gMGEQ1Tjl5xjKZHVUsytdhBZeqYnVHiIMVkpPviB/405OnWPT6Ltx+SIn4QI2IPOndaMJHePGzho
s/eYvJ6bdrWV4kVtvsmvS8ci2isaJhPhctHZLg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
v9mghB9fJKxWdc5G+f1Nqy5bvIICdfk0wHqMBSIOv1adS3vnD1rqW2JHTMpFwWcxo29gUodj9p8e
rN9/sk5+GNaNaGOoapP881u0Rdp8CN7mCR/ehSEN9VqsVfXAFjfCWMCRNY239M+2hT/Mh/l9gNJN
qrKrgihakPaPycx8VS0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jxxhSPb7ZmgXcgFeGop8SDvbtRv3TNH5EBhJ1uEJKtXm+dWbCWoDy36uIk7sUtnAvp82nNgUi45z
Mp4HWtKKcQkS9afRKgbvYPvqNVtpO+2jUTU9TkWvMXrUy3SDvGpXvV9KXTYOccgu1yepsIKD28zu
icuUbsOOGMiDgSKe2wZ9YeykmR9Ln+3OOo7Ik94XB34MteuqoTOrfCpooA8Z3vzEA7/QLKHCoX1c
yZAB9AdLiY3Ehw2tGMPNB95ditpsIBzq0XThpsnJZuM+e2Fq4DZ/VPLFz5wraKg1svQMnX30HY45
yAippTNn881HYuRTryLu8/QnmWk4EcA4oY9cSA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11008)
`protect data_block
BQ7/u6I5CkNnpMDyDyz7h53LT8nrlV2SL5kVGvwZ0k8KGCPWrTVQs/SFbJcWuKat/tjKn+AsyqYM
Yt2cK98ha5gppETLVSiibou+GXejIAKczaFUE8jBAVyJyy6WBp4P/SLb6Aqrfp4aJMXf2PgPCN2P
ojL+umR4SAoBFqqMnya0Bwjg5DQicEUvu0wKCt6gxBw8AYhcZwSwrCClZyfGvSLcHZ3sQWAEx9mH
/6AqcHRqailToytoATQT6uqCUYZf5wVU+ejpkBi4vJUb7q95H9K11z7Ycc32pQeB2cE5k4R3Cl2j
XBHidbQ6DMu19YcKLFqL0MnNlJNmWymYq9EDmzpld1xtR3kAubA78NNW7lN6jBrD3sYTCyDMeX82
X6NxTEaYS/G99V+zLaWc6D1JrrRs8QpXkzwN5P0clefwxnc7wNRfecMakPaokWcfwWi0serS7iz+
TuEXphjtZ9+D4uTX+wYSSXP6pAg/D8OvJ8VNXF+gNhdYYMdjctzspwU5afyqImu1Hkk2vwYZH3no
RdtWO3pLPccfukqBtc5Jr31wzDLxqY85cIjG/PCg3rqLK2+TLGWLINDvVzx/CDljoNzVpDXH/443
96OaHFwwwsrTC2x2WczL01Hnhv3QKaOvTVdBsO99yo3pJd/Iy0LJN/Ct5eFUd8e33CTsTCwGwIna
Fznx8sjQFRLbIS0XMQKYErmF0BmAaIB3rFX5XfnPIRYCZ8XDHSC/0718yfgL8vZ+x9H56RXhV3W9
YEK4wzWMXlF//D0sx5jL43H79hYDiijx+TIiedNpZ5fqLD3JpYE/Iw4+fhGmj3d7YQ2hltrUMd34
FO0lT14G6/kePXQGtfQGUmD34PkXVGnssaMB7EWAHp2MPOQXZv5aKiPGOWYFh8cAFMpF/hhBaWm3
jRGkYhxIfxv0noYJHvp2MU+++bYGumhykcw5qM2DsX1tDFU4/hLUHLIMrnRatb5pb/+gzf7UZEoX
GYw9RaPGa+Gtvh3p0o861p/Z0d4x9GeiPgFIV311pwzXjmjtVxvwM3fkPZil9tT7i+O6RPwT0Kye
J5AL1SHj1nXdIGLG6GF7cIgvCDnUrIl6vvclhLIvMjKUFBE6pAoMdIZQf89DgAI1fnP4iKxiez0u
Stlnu/TzP0Nn0lWgKrfQKcHQW0l8qtRBguwFRwbHrV46qelmj9hmieBBNH5hw/Q1hojRG/Z4wANA
jUInRQ9/JpYYVAfC6V6+4sPpYhd5jKIxDX/Me92kLIR8W1CShOGVbXywEBg5YA9TVlnCZx+vCuyR
6YeilGVpO3i2QtybNREdSuY4n3lYlV5gLau6ByIz90wclNR1AS1OHRH3ZUTJBMdzhdC8gSB0gFRR
V37J+YGJXZZjRs6XiAOyqR7mIyceG+8DBfry7rnBKD98ReKRysI6L9QxxyDQbQUHwGRVlwmDdoNq
bcDBcWNWuWORr4ytUvCh89nb8jf0Ry/LJqaWIhRkMg//l8uCLlL6P6a8z/7d7UaCcQ9qDWXOLgVG
FSFxNtRMcM2ErUoaeJwWEAsE/jbza40uv4TcdqI1aYcA+r5dHONT0wy+7YroZgxOMM7E0REswCR9
kGK025cJwAHJCsKqPP+OFgUn1LccnF365k6jJztds3aFQ/4QYY+RBPqEtXNajwm53MPQkoHRlwi1
yXNdcKaDUVYGJdvmJJIzXOLijPsOJtICXDtBH5dKAV8cgb5sNaSChA7atRmwVnNNhf1tBeo4PD/W
lqa0x675I9LAynto4KzVmyh3MLpsfSgdtvMMoHIQfhB+nWkBmQni4dGbkgX32rtZPt2DcQN/pFam
qxiwbsbG0acR8AFuNWsEqKgT/l5RkqEJrS05r2g+VCRGDXUxOVhC6ThR83/iP6+58IlmidfdHF3R
LhMuRAbm17MVDOJ5P60ootqrvFkM2mFNfCfbVGjeSzuE0ErAEXBJq+/hqnfx4MP8n2KyG/xly1Iz
0xB+VWKRiEIat2vt7bL6uBt7xPWYFGEeqWyEhafYGFi8jpa+Elg128QD5W2+0KCN5sTliTtm5NoY
BFDZ8a8EaCRG7vRFpcNW9KvD4D9Oc4vnT+zqHOSdf/czOWm/d5jqlZJCxjGa/2cqb2ZNqdsYo/Jc
4c6UxTxD0o8nPctOsOrug+2Ub5HyYVJkwrnrO6q8p+Qqa/JpOHF0YEkEjIkslQvZ4ZezCaiX3v6/
Iq1yqJp6lR1zHhpwM20PWQBP0P1/WrSjUJPUBWLaWv61f4S9cK0LclXya40/wqMVZAPzuOTisakW
Naw9AUjcTScSwQzJIIZ3nbvZWR7KcjrNs6rCRx4pLX7tZMd9QMaegeQLgX9YqilIxibZhE66R0mL
JoxnmRuOmrgKI8b7DwjxV5LBA361gClxDZJcRj/rreWN44WgYpDPAN7j/W5Xxj5/ksLjUPhuYBo9
HtB974AVEtUuW4njJgqdfS9JPcWQGY+fuK8sfiqTxYoSayWJKUZYBv+bEtl6gDx39LTHW/+qj+nL
GT4QcBmUZ5SRcwMoDTt2+RJrP/P0uflZPYHVjYLlYbsK2rtoxf6i2MVijUPgoUyIMHFPejr2SKA9
jcm7w+IxPZf+DUCWY/MYC4K6M6ng+VYv+n7L0Z/Bc7c7BFac/pMpLT7Id7vr3XBIvCRC6kHqE4To
T/OI2NmIFUe+9ENoV//cCAPya7hOEkVC5km+3kWZbdLCJHqJO4Y5W3P2atKEvS15KGwmpolayywV
v/IOz967quNx/6j2OY0qjiyyZ86tarYv0uuECPySVgs2PTm3Q7f5H5oVAqKEKFYIqIgYt09qJKoq
tZL0/PdghflE7EAi5hwCt3fgkaslYarPyP0zSmCYU9XBFhhsnYBXsaiB/Te9LC51mv5BIno4I3vi
UrR7FLU/nm1UBTmuonf0Anc4WA3GbhKS23wsD9V6L++tpBE6xnYR9QfrZC4l24GSHxlCNAye++g8
+nvzoP9JaojtCv2TAoGF4yrDlLTOhYfBjpsgQ1ENzN0oWvhOwGlGX+Ut9chVnP1bI6o8366hPIj0
/pSGiYZW4FGahNaMXKHaprHJISQF+EbTd6QlQGfUuYHhaar6aqpeWeEZZBfTV+gS5pz5beoLIrjo
24uIuNZu/zjF/rOpM1lYdHhRVmsTH8V7yFykdFOObUYgO3Y/YPpYuNbtjAXXSjCKHjQiSWAdt2EF
xvFmo85vWdsYlb/1OApgrPE8NjmzOV7qCz4nRGTz6b1IeTqnPuWRyETxpNm7lU2Vt2x4XuqF7riP
w+bdXffgYvu+M8LaB/SzboK3AizjvRHNjgpkRMSRZmOZhobqlCZ7Ce1W0TA9kl22xnCfJtJzfx9O
FD/3xeyyqyNq74jZbjf9iYl0mKWMeG3IKsAorYzixMeNXGWFKvB49yiROLa0avSJhmaXANMKnhhI
9EzcUwDJdv4EbDUaDGTMNgQ5bXDmu/zS9gf5Aaxd3OaPwqtxgajl9ZPOAWxqkj8uNC4cQblBNZbJ
kuN20rmy0vR7hWoKMdhsxSdZ6kpgcSCSQ7YZ9C4PaPpcS2GGsA3xEmDXgYC4id64N0AdAxNvglyG
vQ/JkQgKqOdIBdnTy8oOKjcZDp5mt89dfaakHa6hkNyUPCoplMdI/F1tyecIoV35TcT7udg/Q7ZM
rC27D4fsmz6ENeOHKEAomrdAgnYU9ZQUEsCEcXWkTu2zu4j+2nBwnS/Nd3nchdN/c/9bu2JxIn8d
SdT8eKuT+JZpy5ej0l8pSXaCdGaWZR6FEAGEPWKAU8WeNZJnJH5Z6g2G39oiIfK1cWysqtMVhN9W
NvARkalE8bWRzLkD3BucrLLslO1piKgl5+RkvLaKvYIE8pmw+z8cDXRuS+SThSCZDgWw6xG0XDLR
rsmsMaRgxJB7HfAlXMxm6BHr2B8KEBk26vGnZw1u3tuM4ZBseIn3LtzN8hUBZox1tgsDyzGFRBRj
OcCvjrxc+bbK2cqLERzq4iyRmFO+vvCkvzrhnAohWT9RKaXM13F2GQ8zFEqBvPzdwPWDntfCqbDP
672KtnCVqinsueWPcFDQsecpmNvDrfSwl8/0STDBj71b3Rl64HJ4rE0ry9JxQ8l6qU9uVLRygekh
izB3OFJqYHgQF28haq9liIOy6LgS+Ftpdm1jgGw9IoPREXwYJJ4c1sM3/yuC2t9a4wpXW10FCPuq
3Ld8rjkoe/M6VuLxHI95r2s3tFj9Hi8mArLgvZiXM1KPQHAFYUK8l1NXfvgCaCVUTTyVuBVC9rmU
zp2Z4wPKGaf5QJpHecyMRCeZVXrFzemNx+bwtnSXYKEOQZc+sG7AysGtkijfRFbJfUYsMtTWZqnt
A9bE7TPVHMdE8oCFgDaitca5gw1dZxEiq5GM9UsUt/jhQ501UGvY1Tgq6bgfKacBI7C9Ski7uNjb
UYcT9D+zg1gO/chZkv5pwqm6/3eACSSdY0OLX8fZdJAZzj5xGJqImdGvxNpxei23l/dIw7/U8j3O
BRHLny8F8bXOArPoew6q8RVvyXxW/DxdxhZvjb3T2tJdtCbDJXe9eyHMiabadZN4GVdNRfjPuT8E
ceNK2ikltFianWjWKgr2feo2SAXZuvb89+dGbMqZajZ4Nul0+hg0hmmIirDdOFU1/RjJcrPNb3Hy
9pQvzqNNaZBDKfFvqwp+X4DNOkWaeSqc2Jw64KuEECv4fGFT7TXwat/JszGMrcSPIy05tszuhNiJ
43YxAm3BNjVt87i+1rfn+l6ewuK7nVkvAi8kGSzmhPfUD3ZPh7j7zLobSpHiSkH5D9iTMEOmzhSz
HxNgzjNS5YDzavBYi+X8c/mW2A60HZDXnZ9Uf6mwfepOAs7MEDrIV3YK+8nqw8Yk6bQ5wyhV2JRn
kpe8ZuBGP5Itg8XEOWxbU0ugeyQPtrpoy6sN0V4w0E1K1kWf+CeSWctruXHM34kh7wpc9yf+4xUf
9TbIFZfjGudGsOuq7v3MWPojUFoxGDCflsEcsDo4L6NpfCkRFLKrGUldC3clzRKQAyjnYevny8HH
Dd4AZ+o79wf8/WoCFtymRGxXwpgDLv8YVDE1PtEvSbSjpQipiH/cPmSqu9Q60krkmANcZ3R16YG0
1RnCvwp0lABB+HNvu5/xSuAbKMt65MHKMLVwcTUU6wJkJBTxSk9gWzCs+f29XMKJLafzKnZ934g9
Xkm6Bc21FvRiCJ4naBM+tiYNR8Npl2mC1xx24cSFzdRtsUPCu1KQchAjYIvzauVM17sJ7I0Kvjex
6ZUGzsFfsi+EvsrFifB4DUjyCuKao0NegVSKEFzyHLQ3OOszYZR7Q+RlTp33XCdE1LcsmbDAptKR
n8pyxMeYxrKv64IpwilYKP23bRPfg6+fuMv2z+kIbuHrGVh6W7FqaHm6hvaQmNV0wpoF4lPrWUoH
blvvrjYsS+bUe44szawxl1ujhFrfLDFSw2VAgSfb0QgPwSxjtFb/uIvvHRMpIVProk+P1s/t9JkU
E8O5TAe/jaR++nHQXuOGPpNl/4SCKb/r0grjSVF9kXYw6oBnylccd7L89qs0gG9lZZc7KabkCCyL
HBcGnqCnnmeflvg6WXPomUiMi0pyVswzqc23jaScZusLntfaDf24oLl8OB/tID7Q30ZPyfZAYVy1
U+VgWOzV86TeET0hnXDI7LPYQTCK/6VuZOcOy8d8GDKLOEcY9t7K1tFVBcPOYtXEKAuCMB9U/u37
Q/n0YGL/FD6BBsKLtLTtJ+fkr0scL13naOzrMabU/SoUdeVo18M2uAAbwZ0Iibon+d9m0VEu/rva
njM6JHvdw5eJqpSRXj/M9/u4RVInn4yw7X6qk+u5elnIXnR2euj4Q0pjjD7uqCG0CKzVGSHIxaDJ
GEO7hUFZRZn93qZTactyv+9YbAhcQcKdE8H9I96+ncXPLMbpe9bq4uDkqUI+IMmUv1XPqH2/4ssf
kIOaXuUDjCntTwUg02h+3SKyRcDlHCr6cqdTheDYO54JT3Jl5xKDWQMVA9ppEJnQMVcRvoC+L8r5
TSyvbSYlebGrbUhj8u37UX/k5x3bLQUmp8f9VtQAwiY5gpd1bWNBT0tbTfgiZSqBMByfZfXp9zsA
AfZqniMQGF5Qx4q4tM9bX3nAau7eEZ7F9bJsuaPaCP8ezneqfd/rq82UCO5y7SrCCmiUmOx/ich/
uFr3SyFAYSXF85RZIQtLl6HEL9W47pLmOAnrG+Zl4V+4wblhTx0i2c59xLA6oGUXd+hDERFFXKdF
j11Iujq8QMfzimqXUP1VKRajdDak/zbctNiX3LtphF09Rzfvn6RgFNfOlG1ss+Dc4DVDtZ7g3gpK
eUcaPIpIgKxuRjz93R6EeEO7Nl5lNJNdMDBAMm1/ElHUUfSRFn5CPrRoT1y7DLUjdO9kD2w33Qh5
b3CZAiisfeyDkuVeQLcaUD1EKhfIgmRGt+7bEolBzJmT9r9K9lCWV5hP3qT0x064uEUYqf2DSuj/
mhF9dkmR3XXDCbp8/Tn27jBgq9oUqNT5ay+g+KwfE0n+PqOOf8f0atY0HtXzMNFs7Y0tIYdakWRT
ubeW7PnFUV54BGJhy3cvRDU0e7LSzqNTbhJotfgT6w+mOCaDxVl+JFV2F7hnNwejVCqWtIhHdaY4
LHXY+WTzasHm8b+eTQ6xdAe+FJ5Co53GTNmCKonZcZHWNQzFx2Yqi0aWzjaXEYUVehfgVoTkAh5S
F1sswtD9fLtKvnAbe9AcQTbnhjQRuh/XdTymWjJzvz4snLVCks2fjUUQtkBicmYwk73z/45DveK3
d1Ek5A7hBMo5es36tpVgGhjDKtaEMyhEiW0b0GOrFlm7aYCVBSiXKAYZjg5RLJSDhXx+mGmsHe2F
hwVmX5yraQAcwgVhWpHEagx4HtK15T2nA2n3ngrsW8OPyPdBDj8fvO3sKG4D0qOqGo8Go5siLVx6
oUX2mmeVSJeqEqgbwF79jEwEI8gY+EtiYZBu1voQ+76IW2wjxcKcqpe65c7BbkI9hxu7GPkY3QVw
yy4S0+Ya7yUpWWWXMX28/cy6QPQyTy704hpbpvp3xuBS68ksrdnIbUo9TsTiHDWRT+ORao3SQiHD
DuMoqXYLZ+Duqf5ysCum+vzOccQXDwoScDw6VUCfzvc8FOQvk30uBpcxYy0bRI6GatoL0LU5I/za
rS5xn0mBkYmzF4uWQYej3XCEH/z1MMeaWc40jX3fdXDM7tb/L11Azlb+U3VaiZfYqj+R7YVIYQA4
uL0Pht9/HK8DfUeKnRt2nlrN+OLKPFTRbIvABDtt8mrbcTNmhVUcXoqxVXiBJcWY2a4XX0F5o+7C
WL4vqRUagXEn8qU+Btij5M8Q7R2GnqXllqDVBiiiVg2HfvqX0WHxHOMecEk+7gYiUC8PbE3KGuGM
ya9QEyDX/n4YxpwJTbhx3EfJ05gJMDIXHih8ma5olqfMKYZs2pg8yu+LcSBNmWVwCLr8TwsRmsSR
FrrzD8vXk0Qo6F3I7UuqYW/yxdAhyoDX4lTF3j2g6FgaPB3DxGBw4K/a3COD+EJjd/qNGDsEryIR
Ju2h1CBLEbyZNIpkPmb52ikPaHFcqP51/ABt4pkmXvjeJkYmjNs/x4JyigmosuRQ2+MjDxjaSOta
N5ukk5vTmzuLGaLJCkgtyd55jb+/auWyY1LDH0Pvb3VClsuet8D6rgpA57stjSxYJqLzC9uLYkQ1
kLi7X4uof6xDr2DNcyOonTg6M1S45xlaKO3mt+BAi+xGfNOMj0LmpI5u5W6aiArK106I1LNQnkdm
7mmcU6A2ARA4h2rEvxep0872NQRfIU3U7pbfyAtxZMgNu4jx9Pt7yiFuxjaHNszvxy+mjeWYiT1d
JtUW6OvkXLXj5cRATnt+BgDsRIOyq/gZUzUpnEjE+NmQtYmCmuuWtT+X3gqSYhG32N1SRHs18Q4y
KVgUEZr/m+iA6sosj+iu8cbGDjhu5UPkgPuvixbPCkZjFGxa1Ca8yhthL+X0wOKDD3rsjqUgPks3
HvNu64OpXK0Pom0m4gqtfD25UOvVyuYEqy8JKGs4xI3Zx5Qwhefpc6OhZ4njxtbtybjvnjJBBcSl
birLdYfreTpc0TAlkSvcbTK4hmcYJ3d3rMUfkCrOISLQp8MmJe40EvTiGVDPppjLrCsFtxr1istO
AqFfhSmO/oW7yUQRsd7J9KW6dQHlknzuGl1xb8+EKH/i1aW1KbBdF2kpIG7uYDMILvFfQ2v/AXba
nH7noCKT8TA8kIAG94JPI2wiHTwutPfPMnb57MBImH2RQD/koZrbXWFL/L8Ziw735ZOM6VFiULQn
7qFtpeYzgxibaADvDtejIe/n1Rd8GdWNzkf2NFO9eBWI9oxSbNILdavpsdo1BntvoLh7f/xmjZHg
P/bPajPc/rxgo7JfSqjDJNFgtiPGboA5E91Z2PpeBclT+dTL1XnFRlAB19OAGGlxabh72Dnz90Nt
1wqpxuCqYJ1XClKD8bXN531DeO/NKeG7cu1kQdrI/d55xXQIHI1QPYHtOjUTkLB91IWv0xo8Gxp8
gPpJE3AQkrmmaFJHaz0BpBblWyjD5PmIEjmnjBmUYHaS32fHdT7Sp2iGEL0MahvJmGbTjSLyW99g
9eTZ/kPSaE/IGeyrtcrhCS9tv438FwFv0+Wj0yVaPVlhQERezConTEMPlsCnnzZf90uaH/S0KYcO
MYIlcdtuUiZ2wZHGKPzZqGMKr2B/IA3x6XgkMu20wQbQYmkcB70AlQFc7WNBVMTFTJJsKiqYJgsI
EGkXG7CRnNoG/w3IHwnW2/G/SqpaZPhFFf/PBnSNkH0ZXHmshK4QjzRQYDwy7WXWOXg3wRQJW4Uc
ejbOfFHyvsuXvs5eZVFfM281oAjdhT+sXU+mZxtsAs9YyFGsNQ5kUlsVqgWpN6peSWaUStjEMewk
Y3RQ5mvuC/1He71XUwzNx11cnzzk4rSaXIRyW7ij0CP/32SaBSPbty50n43SruhGwoaEOYm/1fy9
5MzQLYgg2tECIkhHGmeILxIgDQdOqSVbETyeG6HUK8GIc21N2cMS9mpljwvL+EWjXYMqz6Hym3M1
Ii9O4nqPBNqoELdNmICsJKjIHl3PqQtsn9cNPnu7GviZGz8MdM//lKv5XSEdKcjhtERrkrpVzZfp
ovh3bZJsYVgLBna9k/026GLdplMek5Emd2eIShg3nHjPSLgGe+vrCBqIX8xl8s83ifeqS9vk1eaa
/MWKm24gh8i8Q3nWcKp45Ts8GqL8Zc2Nxelzo3mnmLGBO6gcjLHCEsqUHJj3rPzJYDgtdiwZ+Qm3
AbrXgj6AFmhC9SHGu8n8jpyX0ES35L2HkUV2gJTpQKKelljTio4ENMOxVx+ZBpJaTif+k5WoxzIG
NXcnevJeD4LA2dOZ8LE49NCywyx54+/q6gmopYerMDd5NM66PM/yKTs8ACDjWKxMpLo3TuojMaiz
4/jG5Hn2ev5zycET9my9ZA+l2oE/oh/S5BUGoHeH6U7NltQa8GqXSBhSK0aflK6RTS39AgFteQZV
AoU+K4wd/mCEBukdc0cG6VazakwsttdSIbVHWvzN7/4uAXsxrdIdlZb707mqwaKtbx4FVbS9FRs5
QRwM+HSgGACT2Wdq1KRCYq8WF1v8WLcvQRo3d1oGZCM0W/4WdEWPaJWN1AgSg6IC27lBFdBsOdkv
fx9sL3FcWlbUBcG1qfsg+6LfA+9qwtn2Mga9jOoiJhZbGAIWDzmnCH4c2+KXENTPKwhGJtiUNnwz
3u5DbF7KBLMPU5zJTV1FO74i1Gs/epaYetiau0Ro4JPKVYMI8DYOqMLUnxaUybEiBqL9OJCTSImX
gNlATUa+yQZ9vhPY/xbm4KPDMgQJvCKk12jB0AnzN7jQlUF0XDPCO+rZ0cU+sFboEiSTXG4S7a0X
dtdlSKhgvJON73UrCZY5GJzF58ggwWWiqVp+JUUqtLGSxQ0mn+7jqNXMYSb359KsXOZUFEJGCmxd
EHb9Y/DKpOpXmHpqPiuJjchBJ0y2PsNFLFQqbBaAmjzw+6P8J5L3kih10o9C+Ecfhw/LCmfBb19p
MLTRJm9T6lDn02Sdbx4P8+yXQa9N91DHoqUntQA3zcfsRf101jNTeof2rXEQJq2goK3qurmSVO/8
bHHI88XngHpW9XLmHFUGKF+oOVgcJa05UbIHZN2OsWpupurn7y0b8tdYaFPqSAyb/f1kz6btK4yK
eqOtaW8sooGZfdciWQXrOwZW5wbpit+Taih/KhxfeitfGIunfZcbiSQerfxU6A/O4hV09wNUJcIW
9NIsXYtCZvHOcCtGnbS3NXyYaOXYTC570THy0n875k4S1suoLDhVoJQbXAY2zvw9lO9KUoM0dOOy
1uoTnhYzp+PM5MVMPnz+o8+Sj6QTnuXb7Fdmvs/Pw0BzpjLYCxDiakDA+hjdeMxrr3xWH9dan/6s
K/3tlYnvrx0mf6DFXo2e7R180S63uD+CzzyLCqIfL9lsa140VQx4923GVfXihMoBX/PkF3MkSj5X
yTGMvVwHMyqjTb6M73u5ZJ8pyihvkrAm2BMACgQASq/Wh+YqHpDVc6ptCZQdF6dJj8GSshtixun4
MJBX0RMCKEpeocD7QeVtJ5EiqyB4NNXeAoxvVJvtdD8CJqjtPJW3ECkTJMCBxpnmGxoHbDwc7I+o
eN+Y0FL6qnPQnxZ9KWCWR9Jyru81XFjhVahg7ULxVWqS9iSAa8QIWmuTx6rCmnttoFOWJqE7Oj1O
tdxptewaDg5CTiAMxijAlSO2Y8o0LcxoCHjPCDiIfXR7kc82vNPwilWFJBDIwYJhA50putR0Z612
IefIdF7kPfDa9lnDFjKSLBOp5j2gBoufpU+hsxr9TPu7gY61TiOSpD/LmnJYkqShfzDdwUSyyT2c
8yoh1ONZ6S8hGvD7toCnb4oG/ZvUcVk3N4NUO6fa3FHtpzSDxoBYIeX2jodLFAab9yy1y85mWdre
FquFVg5SKWI6JaIkAz6/yamYXR6x19vDJZs6ZomIo5SwPoEADS93y5uo4QKqEhiOCDeoIYBBom37
h2DghwXZzd6YOfutNRNQj5n/Ht2Eh8FYkgjFPg6w1H2GB5BgJwE2p4D/iXzK5voSyKbnWOx/vsBU
IKqYiD6ozU3X5nmBSe8jge+ZiVsTHTiRQ7Arw87Yyq85HsQ/Y4s0PizvqsizirmeDHzG5FB0GNBp
OFr2Is5Bd9PX8RureGEKd9oQA9CAQjVUnNvMkXj8b2gaOBCWQdkh6ZjptzDyh1bDV5U7go3KYKvm
+bBbAoU7h9l9z77wpdGV1ONJdD1YpWVP3PB8Crx646fQ3M5dWp0m8KgmZFn5FYRUkPq7yUVOk0Lr
sAMTLfiFJ5D0Uyf4fL0fXPU/CI99umud1NKq+j94NguzLtMCntlYerTZL9C4FEVvwjSJGhUAES5O
QJ2c3NXWO/5JYxBnqguBIaawKoX1kKNFMjEfhh2Nrh+brofK9Z0Q3w3o+YIromYfmHDA6vkbPKeE
Z4sxQyfd1rKkptm9nhNiXFPcas92FON/mYezvP22qDH5QISgZFywEpGp6P5u9gu/bq+6hmwwx5MU
RJc/VaboKA4cnXXGRv+2xHSqTUIb35oWgZ1wQkLEHiOwjNPTlH1Y6P3Lq/RG28E1Aj7+dNEb5XJ+
VpAZ9S95fvpr2duow8oActlei8g4e7dGYeKcjgoVHvCsFvRIOI0QK4Cz1zQ9Zt6bujHgZ+xT5rik
fVOLmXT+/H8hAo0eMmBquU2cxNZ92ll1P+ejyeGKrAYy7n6FTHJbmQTBXdmkMIXZYRlBY9ASn0IW
4dgjsxGZMh6wwmOZWQFYVaRgGne7jADn3PRPbmhvAeLL9nAfgi6tlvq39BKk9T+diHuOF58RYi51
1ZqMU7ehQg7SOuoB16fYlkNlfxja2uOBg8QRBWXf+euUjOgB7gabOExePOuBp2eSTnY4U+GbxEaN
aDxETHffS94mHmmU+3VvBGzGX878KyD7q835tubDDZ6ivItHm6ogAR630IBkYPQ55isi+ayfcfXz
3Cmp7aIlXYMjGse+g/TPyDo7aO253ttB7hJ3mNa2/teQhpAwN0I7U6a/j9C3eCohEkzL+IEzqHLN
XrSbbFxDCTbV45J+TkgGgdF8SFTZtzjnDkCC/pnrScN4LSxKifyacCnM+tIY406GNQB3oUBNJCxl
1l6L7iMNPKUZIP9Lblk6BgnH+hUxKQiBe0SumZpeOVO8IGJtql71sO1Ecn904U43ixiV0n/noVye
6xVad5zv0Iav/oyBqdNz7WUKQNemmI1BuucO+9D/f6Uvd2sXeNu7fSNlddaBzIa3am3FJOS277Sg
CfiS9Zd3dBghpZ2oM/1LSGFH4sb5PlM3ixdfgTWhPm3GASrqWSqEmjxOMFwC93cRtortxQqCic1A
p9nPTa6U7bginheGpkwS1gKhucBNh+qTJIbBKMuKkDXWcNJiYjWt+769KMLI7Vf/wJpiaHT2sxqF
iPhIecIWCeAMUwFLhLpP6Uvdhl/RO6IQNysr3CITUhYRiG1JDSPRqAypALbVZjeUGm0caC3JU+g1
URwX8zSWiSdxeRygj4HwK+rJKp2m9i3k0nRl0h6Zpr31d8zHfPt1L1Qe1N5jqfE06gbg9b03gMUR
x/SqIj1aEDIoV1tf5kopkr60OWAqKDpIa5KonAcvLmPxzocaqRDoibxwhHxOCPy2RO+1cbflULKm
SK87r9LHrQMX1jkBtenW6VNq5AE8RJvJBu/0bYpLnHVoqORjBUKvz97bcS5l+jvmE3GMmzSxI6bY
/mlEiVcJUfCRo/kqs4UuX1hv9rZgm13NFs5J9dOVUtyEZvbxXcswVrnmJryCHdAfYBVK53/tMsOH
nOhDQscqXxV8QsNxfmixbEFzqg0oDH6H4dGKqaOr5J85524TlnEKllsK8ZTHmByr7tVXvzVtNoBy
+o8Co9uxACvqW0AzvX8P//R7TmwlHfZ/ihqxz83BkOL7uhzJxbhVjljcy0oe/oagI8q6CnNWdUQz
wOUq5yoCWhClX9udH2fk9ymCtLkLyJQvUCIWVQH4VIeAmllmrZ/5crY8RNekHkyC98lwkM3wSDw8
ZxuCxvTjuOGBwePGAkpSPoRhEjGBAmY37m9uUjIPduaAwmKAjHTxCVQYl6N80CG14j7j/WnQ1hph
GXmS4N7QD9T4WVJ/zFTbDn5fOU9nu5TWP2xIZU74dSkRvcAH7JU2IOj470/Efz9kAU0jeDgkn51H
TCgZPbFyv9tBauWn8ZyD9t0m02/n94NtqroqSLGXMXgMaxevZeufVmoe0/bHZuq8H9P3x2u3l3YB
L6LOsOFAUGZBn5K8evNIUcDIn9ydFJKVCTRaMST2n26v2hTMhwvOxe2Eytn5cA/IX65ySsH8WDoX
+Q7uDkKVHlqBjxdGnylHKM/iLF92vHvrDUwiBM14GCXho8vsqdqfttYdT4NQALo0TbyHhWw6LL2w
yhlsWb7jD4zMCsQtbe4H/iHnsWkA5KvGI0kBD0Wk9nrH5TgbgaCzpzEIXtfmBI3TItPeVSACaMM/
1uCi3OBiluwenWiZoah8H9QDg/cmFVfTKhx4nWtluS0viPbNWPHEJvd67OgXnDEPeZCNvXtFgJ3i
7r3GoSBlTP39K2OFpwfLdZ5cuNxkTlh04GsHA4JhAFp948ckQ+knuIb1oPNa3iS3qLm7Kd/5eLaa
T22ObJ1v2x2a3rYb3ukJy4FKAYJJi8wGq1VRgxbut35JbrQkh/8kzUQQznfsgPLdmc3Q2/W0cDFU
cSlMLS413VH5L9ksUJJ1Gck9VrtFj5PsRG+s7D5hBJ+qDA2HHxUhyBHJVzK0v7RE6UlLNE0VG4XO
/JuvcxqjueTlINt7Npm5NG/UJnfuWb9unmnQ3Rq5DB8pVCUCZizbCMCMywslw6isndCEA6agwTVn
Q/X9Oq9ygI8Z0kWFyFJMY88N/Ro59B4BC/7F5zLpYFeHAJg+xQvtZ6flIbrfdzlYnGE/vr7a/1Fa
4GeglEpUn+nSVhePtu/ZjGYCdIXA3BuVjHDAHXTDBO94flu+9xjBoiCOV8dEQyAAiCaazaFUTQEG
pY0X99048qq1ao1Kjg0IKjLqt7jnIUMztOSuBJ1xigIYhT2FknguOsQJZgB+D1g5oyYyXV3ZWw6G
uDkv49jhhbXdCMc6Lp2nPh1Z9H0yq/5g7EnLF71wVcurz9wtlnkzXL8p35oY39hXJhbfRH7+v3Bi
/xkixlwLmyyXSs034ScWd033kssopjC45HTSCyTY2MzlKK8eiLz6k0dUyXzzMa7QWhF0cEJjW1yk
85DJS9i5/TU4ylDs0QyISJrmRxMxxNOpqcaY2zDvTM/D17hgwpCUytSU+N2HoHeA0h9im9GpQrmP
0rDWViKfjbJ6JtfdLRirIPaRY0gzKRqtmADm6YWChNiVO3cEj8EF4Jv1AIforjBLRXsrxa6R08yl
L7uXICxc4l6Q8VZSgkHFOgpTE6CsqViKxBxmqhfrc1UC41PfA69KNv0d7AbIQ4hWnSS7/BgFwtMJ
vJL4sJ1/QAtOxxPIcQk/1TP8Pqhc3QxUWXP5S/G8k5vm6TGGkhk/yYUmtSwOSVrSibVPo9sCUmIQ
UgtqTN/V5QvRYRxwW/3Y1uoSbVgORaOTamIlTVTENCUIoEicBYvzIrwJ1klSb7ed0vFLNugCjdFZ
APRqoJeCXA==
`protect end_protected
